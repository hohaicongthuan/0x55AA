module layer_10_featuremap_268(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398db2b4),
	.w1(32'hbba8ebe0),
	.w2(32'hbb917f2d),
	.w3(32'hbb4802c2),
	.w4(32'hbbadb42a),
	.w5(32'hbb64366e),
	.w6(32'hbad2b9da),
	.w7(32'hbbdf2711),
	.w8(32'hbbdc397c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8041),
	.w1(32'h3aaeab85),
	.w2(32'h3b1dbc8a),
	.w3(32'hba905958),
	.w4(32'h3b80e583),
	.w5(32'h3becdd2c),
	.w6(32'h3b4074b2),
	.w7(32'h3b165fce),
	.w8(32'h3aeb3938),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf68b61),
	.w1(32'hbbad8c46),
	.w2(32'h3bfae04b),
	.w3(32'h3a9ce34f),
	.w4(32'h3b9395bf),
	.w5(32'hbb8cccd5),
	.w6(32'h3c8ffb30),
	.w7(32'h398db31e),
	.w8(32'hbaf36adc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba378520),
	.w1(32'h3bd66f02),
	.w2(32'h3c88ddae),
	.w3(32'h3b31e8aa),
	.w4(32'h3c216b87),
	.w5(32'h3bef042a),
	.w6(32'hbb746dbc),
	.w7(32'h3c690b43),
	.w8(32'hbb64a386),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8edd5c),
	.w1(32'hbb918454),
	.w2(32'h3c0e0166),
	.w3(32'h3b48265e),
	.w4(32'h3c006aa6),
	.w5(32'hbbd48477),
	.w6(32'hbcbac1e8),
	.w7(32'hbc99657b),
	.w8(32'hbb87f05c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840b60),
	.w1(32'hbb23292f),
	.w2(32'h3badc16d),
	.w3(32'hbb9df885),
	.w4(32'hbbade8c8),
	.w5(32'hbb803ccd),
	.w6(32'hbc0daf68),
	.w7(32'hbadfe513),
	.w8(32'hbbaeba77),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5970e4),
	.w1(32'hbae3445e),
	.w2(32'h3b4ad57e),
	.w3(32'hbac1ac84),
	.w4(32'hbbd7a54d),
	.w5(32'hbc2a1f9c),
	.w6(32'hbb7f8d21),
	.w7(32'hba3e0d83),
	.w8(32'hbc3d5385),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75e17a),
	.w1(32'h3bcffc89),
	.w2(32'h3b589cee),
	.w3(32'hbb9abe15),
	.w4(32'h3b8ad99a),
	.w5(32'hbb6912bf),
	.w6(32'h3b72df29),
	.w7(32'h3b985f89),
	.w8(32'hbc2b8b82),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1fad1),
	.w1(32'hbb83ea10),
	.w2(32'hbbc09c6e),
	.w3(32'hbc067307),
	.w4(32'hbc19fd95),
	.w5(32'hbba779c4),
	.w6(32'hbc0091c4),
	.w7(32'hbb97d07c),
	.w8(32'hbb82051e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01bfdb),
	.w1(32'hbbf63876),
	.w2(32'hbac5ab3e),
	.w3(32'hbb44ca8c),
	.w4(32'hbbd270e5),
	.w5(32'hbc41f050),
	.w6(32'hbc1ec3a4),
	.w7(32'hbb8fee29),
	.w8(32'hbc0fd4da),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe20e80),
	.w1(32'hbb81a149),
	.w2(32'h3c0374cf),
	.w3(32'hbba3258c),
	.w4(32'hbaa3f89f),
	.w5(32'h3bf7565b),
	.w6(32'hbc638264),
	.w7(32'h3a8545b3),
	.w8(32'hbafd731c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ec0a8),
	.w1(32'h3b37035a),
	.w2(32'hbb9b64ce),
	.w3(32'h3c6f3855),
	.w4(32'h3b8bac36),
	.w5(32'h3c0a8b23),
	.w6(32'h3c7468c4),
	.w7(32'h3c37a3c1),
	.w8(32'h3bf14b7c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babe287),
	.w1(32'hbc6ccde2),
	.w2(32'hbd213913),
	.w3(32'h3c81e55a),
	.w4(32'hb9eaac1e),
	.w5(32'hbc0c54e6),
	.w6(32'h3c8481a3),
	.w7(32'hbc4c011c),
	.w8(32'hbb516110),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8e1f),
	.w1(32'hbc2be8d2),
	.w2(32'hbc0b87b0),
	.w3(32'hbbac5171),
	.w4(32'hba59ebaa),
	.w5(32'hbab2973e),
	.w6(32'h3bd6c1ec),
	.w7(32'hbc6c303e),
	.w8(32'hbc1f3a14),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4015d),
	.w1(32'h3c0c3d0c),
	.w2(32'h3a8c5ec9),
	.w3(32'hbc0127c8),
	.w4(32'h3c0a042a),
	.w5(32'h3aa1be0b),
	.w6(32'hbb7b6ee1),
	.w7(32'h3c13f1bd),
	.w8(32'h3baf4b6b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff7375),
	.w1(32'hbbe53f43),
	.w2(32'hbbdf627b),
	.w3(32'hbba5471e),
	.w4(32'hbb7eb80f),
	.w5(32'hbc690bf2),
	.w6(32'hbb5a59d1),
	.w7(32'h3abf4e26),
	.w8(32'hbc8481f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac9ac),
	.w1(32'h3bc564d2),
	.w2(32'h3c2e6ee2),
	.w3(32'hbb40a232),
	.w4(32'h3b87bdf1),
	.w5(32'h3b9e275b),
	.w6(32'hbb9cc613),
	.w7(32'h3c1ab1ed),
	.w8(32'h3b081227),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a160d7),
	.w1(32'hbae6716f),
	.w2(32'hbc83d192),
	.w3(32'h3b30c086),
	.w4(32'hbbcee4e4),
	.w5(32'hbc0ade32),
	.w6(32'h3b937c8b),
	.w7(32'hbbdcb93d),
	.w8(32'hbc8518cd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8a8f),
	.w1(32'hbb809097),
	.w2(32'hbbcf207d),
	.w3(32'hbbd00559),
	.w4(32'hbc0f1a39),
	.w5(32'hbbe4dce1),
	.w6(32'h3adc194d),
	.w7(32'h3bda4d77),
	.w8(32'hbc3f1e83),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fb42a),
	.w1(32'h3be098eb),
	.w2(32'h3c42b643),
	.w3(32'hb818d9dd),
	.w4(32'h3a55cc63),
	.w5(32'h3b8b6676),
	.w6(32'hbb388ef5),
	.w7(32'h3b1b4a62),
	.w8(32'hba464b91),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60629a),
	.w1(32'hbc0b46f9),
	.w2(32'h3b613128),
	.w3(32'hbaa53bf2),
	.w4(32'hbb765def),
	.w5(32'hbc0b3c9b),
	.w6(32'hbc1e0dd2),
	.w7(32'hbbbf0066),
	.w8(32'hbb49c9b4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985c536),
	.w1(32'h3c0700ea),
	.w2(32'h3c35be08),
	.w3(32'hbb136cf2),
	.w4(32'h3c10b972),
	.w5(32'h394f6696),
	.w6(32'hba28d31d),
	.w7(32'h3c381d15),
	.w8(32'hbb44ac1d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53f2ea),
	.w1(32'hbb242055),
	.w2(32'hbcccb227),
	.w3(32'h3bacbf98),
	.w4(32'h3b6d0eb7),
	.w5(32'hbb8dec51),
	.w6(32'h3cef2812),
	.w7(32'h3adb10a9),
	.w8(32'hb9fed919),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb448458),
	.w1(32'h3bc9958a),
	.w2(32'h3c1025e4),
	.w3(32'h3b69d609),
	.w4(32'h3be663fc),
	.w5(32'hbbe20609),
	.w6(32'hbae1273b),
	.w7(32'h3c6deb11),
	.w8(32'hba2a9d88),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a3b0),
	.w1(32'hba641005),
	.w2(32'h3ae83c60),
	.w3(32'hbbc7534b),
	.w4(32'h3babbf61),
	.w5(32'hbade2d7c),
	.w6(32'h3c2fac89),
	.w7(32'h3c76c1d4),
	.w8(32'hbbecbc94),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c95b3),
	.w1(32'h3c08d9c5),
	.w2(32'h3bfc4577),
	.w3(32'hbc659121),
	.w4(32'h3b89d777),
	.w5(32'hbc6a0998),
	.w6(32'hbb9862a9),
	.w7(32'h3c42651f),
	.w8(32'hbc10a1d2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88d19e),
	.w1(32'h3c2d2746),
	.w2(32'h3c7f6e6b),
	.w3(32'hbc3fbf9a),
	.w4(32'h3ab9c1b8),
	.w5(32'h3abe5779),
	.w6(32'hb8669fd3),
	.w7(32'h3c98d0cd),
	.w8(32'h3a5b5445),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e3449),
	.w1(32'hba90e91e),
	.w2(32'hbbcaa585),
	.w3(32'hbba63434),
	.w4(32'hbb35d4bc),
	.w5(32'h3b3ce20a),
	.w6(32'hbb2b9538),
	.w7(32'hbba171a8),
	.w8(32'h3ac197e9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29bf9d),
	.w1(32'h398abec7),
	.w2(32'hbb874a16),
	.w3(32'h3befda5a),
	.w4(32'h3b8ef717),
	.w5(32'h3b863495),
	.w6(32'h3a26add0),
	.w7(32'h3b015c4f),
	.w8(32'h3b1ed584),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a73bf),
	.w1(32'h3b5535f6),
	.w2(32'h3c4ee779),
	.w3(32'hbbb4b3c8),
	.w4(32'h3b32b4e4),
	.w5(32'h3be73fe1),
	.w6(32'hbb9e3ba5),
	.w7(32'h3b19502d),
	.w8(32'hbb63626b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87e06f),
	.w1(32'hbc3d04c6),
	.w2(32'h382d018f),
	.w3(32'hbc0fef27),
	.w4(32'hbc29cd90),
	.w5(32'h3b148d84),
	.w6(32'hbbcd1b4a),
	.w7(32'hbbc51381),
	.w8(32'h3b537e6d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b9961),
	.w1(32'hbbc78137),
	.w2(32'h3b7a1766),
	.w3(32'h3bcaf593),
	.w4(32'h3b7f4e40),
	.w5(32'hbbb619aa),
	.w6(32'h3bceb182),
	.w7(32'h39a52d2a),
	.w8(32'hbb4ece1e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32bf9a),
	.w1(32'hbc5693e9),
	.w2(32'hbb2d1702),
	.w3(32'hbc10251d),
	.w4(32'hbbbaada1),
	.w5(32'h3b85cfef),
	.w6(32'hbb235e50),
	.w7(32'hbb876d2e),
	.w8(32'h3bbd0e37),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84685f),
	.w1(32'h3ba37e8d),
	.w2(32'hbc41aabb),
	.w3(32'h3ac86b53),
	.w4(32'h39fa14fd),
	.w5(32'hbc4ca0b4),
	.w6(32'h3ae73b05),
	.w7(32'hbb48cafb),
	.w8(32'h3b49b012),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3289),
	.w1(32'hbc0d7390),
	.w2(32'hbbbee097),
	.w3(32'hbc255cda),
	.w4(32'hbc1e1664),
	.w5(32'hbb74488a),
	.w6(32'hbc2e3485),
	.w7(32'h3b196454),
	.w8(32'hbc628ec1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae5559),
	.w1(32'h3c1a03f7),
	.w2(32'h3b98555b),
	.w3(32'hbbb0aadf),
	.w4(32'hbbbde2ef),
	.w5(32'hbc4b7213),
	.w6(32'h3b6b5934),
	.w7(32'h3b926f39),
	.w8(32'hbbb7c5e8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69c501),
	.w1(32'h3bed52cf),
	.w2(32'hbbfe21c1),
	.w3(32'h3a400e25),
	.w4(32'h3bffb1e3),
	.w5(32'hbc646f55),
	.w6(32'hbbd9caf1),
	.w7(32'h3c89acbc),
	.w8(32'hbade2f9c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1df8),
	.w1(32'h3cad4398),
	.w2(32'h3cb9ba42),
	.w3(32'hbc2e2682),
	.w4(32'h3a3cbc58),
	.w5(32'h3c258088),
	.w6(32'hbb0ebff3),
	.w7(32'h3c620e27),
	.w8(32'h3c6d33d0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ea2b),
	.w1(32'h3bea69e1),
	.w2(32'h3bf6cf83),
	.w3(32'hbb181ea9),
	.w4(32'hbace8cd5),
	.w5(32'h3c086fad),
	.w6(32'hbb2c305c),
	.w7(32'h3b3a6777),
	.w8(32'h3c78aa64),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdf1dc),
	.w1(32'hbb964a3f),
	.w2(32'h3c052db2),
	.w3(32'h3bbe5849),
	.w4(32'h3c40a068),
	.w5(32'h3bb9fb02),
	.w6(32'h3a972a3f),
	.w7(32'hb9e1be5b),
	.w8(32'h3badd987),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f931b7),
	.w1(32'hbb06881d),
	.w2(32'hbbc6c32b),
	.w3(32'h3b0e465e),
	.w4(32'hba94905e),
	.w5(32'hbc162138),
	.w6(32'h3c880542),
	.w7(32'hbb5c960e),
	.w8(32'hbc24c346),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cfe76),
	.w1(32'h3bce39fa),
	.w2(32'h3c44501d),
	.w3(32'hbbbcd0ec),
	.w4(32'h3bd6eaeb),
	.w5(32'hbc43cbe0),
	.w6(32'hbb8b13f6),
	.w7(32'h3c158ce2),
	.w8(32'hbaef8402),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e0c09),
	.w1(32'h3c7d4a42),
	.w2(32'h3c53c10b),
	.w3(32'hbb9232d2),
	.w4(32'h3bd27a4b),
	.w5(32'hbccf7ffe),
	.w6(32'h3bbd45f3),
	.w7(32'h3be7f3d6),
	.w8(32'hbcd869d6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b70fe),
	.w1(32'h3bc93d49),
	.w2(32'h3a1e4358),
	.w3(32'hbcf95ed6),
	.w4(32'hbb847394),
	.w5(32'hbbc9f6ce),
	.w6(32'hbb315c6a),
	.w7(32'h3cba9c04),
	.w8(32'hbc333fd2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5be6ed),
	.w1(32'h3afef728),
	.w2(32'h3b9e120d),
	.w3(32'hbc33db70),
	.w4(32'hbbf7e250),
	.w5(32'h394de537),
	.w6(32'hbc863e30),
	.w7(32'hba962730),
	.w8(32'h3ab70aad),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3d7e9),
	.w1(32'hba138a0a),
	.w2(32'h3b7869f0),
	.w3(32'hbbaf3dd6),
	.w4(32'h3c1f8128),
	.w5(32'hbba70002),
	.w6(32'h3ab90a36),
	.w7(32'h3c80dcf9),
	.w8(32'hbc3fd9e1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8760ed),
	.w1(32'h3bec98e9),
	.w2(32'h3c0d4b5e),
	.w3(32'hbc1aedf4),
	.w4(32'h3afc3048),
	.w5(32'hbb5a4238),
	.w6(32'hbb57b3e8),
	.w7(32'h3c4d6b0c),
	.w8(32'h3b87aa70),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becf8a1),
	.w1(32'hbb13e8eb),
	.w2(32'hbc4793d1),
	.w3(32'h3c3a5f9e),
	.w4(32'h3b1979b0),
	.w5(32'h3bf234f5),
	.w6(32'h3c63af66),
	.w7(32'h3aaef682),
	.w8(32'hb91b9cba),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefb126),
	.w1(32'hbbb10175),
	.w2(32'hbcac0ada),
	.w3(32'h3c381888),
	.w4(32'hbb3cfee1),
	.w5(32'hbc2f328f),
	.w6(32'h3a8c24cf),
	.w7(32'hbc3229c3),
	.w8(32'hbb54a517),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384aa75a),
	.w1(32'h3c140484),
	.w2(32'h3c2db698),
	.w3(32'hbbc9b36d),
	.w4(32'h3b2e6ca6),
	.w5(32'h3bc414f8),
	.w6(32'hbab86bef),
	.w7(32'h3c1c278b),
	.w8(32'h3a5b2dd9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61fdc0),
	.w1(32'hba99fe39),
	.w2(32'h3b73d149),
	.w3(32'hbbb32f58),
	.w4(32'h3a84874a),
	.w5(32'hbc49df12),
	.w6(32'hbb025e4f),
	.w7(32'h3b7518bc),
	.w8(32'hbbb921ef),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991fd9),
	.w1(32'h3bf5adcd),
	.w2(32'h3b94de7c),
	.w3(32'hbba758a4),
	.w4(32'h3a892ac5),
	.w5(32'hbbcc615c),
	.w6(32'hbb1de81d),
	.w7(32'h3bb005f3),
	.w8(32'hbb96be72),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba861e78),
	.w1(32'hbbdddb6a),
	.w2(32'hbc461781),
	.w3(32'hbc11834a),
	.w4(32'hbb002e92),
	.w5(32'h3b9bb4ac),
	.w6(32'h3ce75f21),
	.w7(32'hbbefdafa),
	.w8(32'h3b38b494),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9641),
	.w1(32'h3b840c6b),
	.w2(32'hbbb09296),
	.w3(32'hb943e53a),
	.w4(32'h3c148b4a),
	.w5(32'hbc035911),
	.w6(32'h3c43a9f3),
	.w7(32'h3bdec8fd),
	.w8(32'hbb7b9165),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c25d3),
	.w1(32'h3ae5b678),
	.w2(32'h3ba60ab4),
	.w3(32'hbb34f28e),
	.w4(32'h3b3a8961),
	.w5(32'hbbc9aa46),
	.w6(32'hb9a3c4e1),
	.w7(32'h3b7ae86a),
	.w8(32'hbabcc143),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacecef),
	.w1(32'h3c11aefd),
	.w2(32'h3c217cf1),
	.w3(32'hbb3ba179),
	.w4(32'hbab77853),
	.w5(32'h3bbf570b),
	.w6(32'hbb99e817),
	.w7(32'h3baa46cc),
	.w8(32'hbb6ce3a9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a35be),
	.w1(32'hba541a90),
	.w2(32'hbb56e2f3),
	.w3(32'hbb5df878),
	.w4(32'hbb80c413),
	.w5(32'hbbb43937),
	.w6(32'hbbe6b06f),
	.w7(32'hbb843a58),
	.w8(32'hbb9623ee),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4985c2),
	.w1(32'hbb8ccb6d),
	.w2(32'h3ba4ccbe),
	.w3(32'hbb62a8a9),
	.w4(32'hba4462e2),
	.w5(32'hbbec54b1),
	.w6(32'h3a119f56),
	.w7(32'hbc11f35b),
	.w8(32'hbb856c55),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749080),
	.w1(32'h3be9f1b1),
	.w2(32'h3c276b9b),
	.w3(32'hbc429fa4),
	.w4(32'hbb0b4c01),
	.w5(32'hbb3e3562),
	.w6(32'hbbd2d8a1),
	.w7(32'h3b9b3933),
	.w8(32'h3b7628c6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf84266),
	.w1(32'hbb3d6fcc),
	.w2(32'hbbaf682f),
	.w3(32'h3a97b4a2),
	.w4(32'hbb091856),
	.w5(32'hbbf60660),
	.w6(32'h3b95474a),
	.w7(32'h3b0c7689),
	.w8(32'hbba023ce),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb473fa7),
	.w1(32'hbac8c178),
	.w2(32'hbbbc9813),
	.w3(32'hbbc2f5a6),
	.w4(32'hbb6bda37),
	.w5(32'hbc5e6cf6),
	.w6(32'h3ad5b12e),
	.w7(32'h3aba43eb),
	.w8(32'hbc8fa645),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc319c79),
	.w1(32'h3bb2ccbb),
	.w2(32'h3b9468b8),
	.w3(32'hbc4b6fa0),
	.w4(32'h3baaae66),
	.w5(32'hbc498364),
	.w6(32'hbb475551),
	.w7(32'h3c5317ee),
	.w8(32'hbc7194b1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba587608),
	.w1(32'hbc0396b6),
	.w2(32'hbacfa73e),
	.w3(32'hbbf6cf46),
	.w4(32'h3acc38b1),
	.w5(32'h39c6af89),
	.w6(32'h3af208fc),
	.w7(32'h3bbf099f),
	.w8(32'hba24728c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b0d71),
	.w1(32'hbb2e2578),
	.w2(32'hbb86c3c3),
	.w3(32'h3a071657),
	.w4(32'hbb1df92c),
	.w5(32'hbbad7af6),
	.w6(32'hba03e867),
	.w7(32'hbc0171ca),
	.w8(32'hba4d5e3f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ddb9d),
	.w1(32'hbb12bc12),
	.w2(32'h3b0a284a),
	.w3(32'hbb45a6e0),
	.w4(32'hbaa291b8),
	.w5(32'hbba6393d),
	.w6(32'hbc266570),
	.w7(32'hbbe7bc9a),
	.w8(32'hbab58f96),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab756),
	.w1(32'hbc0ccc42),
	.w2(32'h3b5aab56),
	.w3(32'hbbad33fb),
	.w4(32'h3b764fd9),
	.w5(32'h3a418655),
	.w6(32'h3c0cd254),
	.w7(32'hbbeaf12c),
	.w8(32'hbb34746e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53e347),
	.w1(32'h3932983e),
	.w2(32'hbc7d2ba5),
	.w3(32'hbb92d7bb),
	.w4(32'hbb6f8417),
	.w5(32'hbc28d61d),
	.w6(32'h3b90b617),
	.w7(32'hbbceaf81),
	.w8(32'hbc4a3a9a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fc596),
	.w1(32'hbb264258),
	.w2(32'hb92308b1),
	.w3(32'hba2760c7),
	.w4(32'h3b9d8c79),
	.w5(32'hbbab96c4),
	.w6(32'h3b4bbe74),
	.w7(32'h3bd55dab),
	.w8(32'hbc48d3e3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10c15c),
	.w1(32'hbc2de8d1),
	.w2(32'hbb5984b2),
	.w3(32'hbc8d4eba),
	.w4(32'hbbacd1a0),
	.w5(32'hbc8c43ac),
	.w6(32'hbc78ac8d),
	.w7(32'hbb22c660),
	.w8(32'hbd07f884),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf5429),
	.w1(32'h3cd15dbf),
	.w2(32'h3cc23ced),
	.w3(32'hbcc1eb31),
	.w4(32'h3c053f21),
	.w5(32'hbb1dd737),
	.w6(32'hbc06063a),
	.w7(32'h3d1b0342),
	.w8(32'hbbc6d008),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0086d),
	.w1(32'h3c5bb92d),
	.w2(32'h3c4c1e49),
	.w3(32'hbc21e442),
	.w4(32'hbafed2a7),
	.w5(32'h3c50c557),
	.w6(32'hbb9ff43a),
	.w7(32'h3c0d768e),
	.w8(32'h3bc6b94a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b820484),
	.w1(32'hbb8dd21f),
	.w2(32'h3c28e35b),
	.w3(32'h3ab9397f),
	.w4(32'h3bb01519),
	.w5(32'h3bfec4d0),
	.w6(32'h3bbd67f7),
	.w7(32'hbb55f1c3),
	.w8(32'h3b92e989),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7fc2a),
	.w1(32'hbb427ef8),
	.w2(32'h39d46598),
	.w3(32'h3b55bd3d),
	.w4(32'h39f5cdec),
	.w5(32'h3c36b083),
	.w6(32'h3aace41b),
	.w7(32'hbc0e715d),
	.w8(32'h3c10554d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54b1d3),
	.w1(32'hbc3673c3),
	.w2(32'hbc939c73),
	.w3(32'h3c479340),
	.w4(32'h3b3f1ed7),
	.w5(32'hba64639e),
	.w6(32'h3bdc4eff),
	.w7(32'hbbab4558),
	.w8(32'hbbce4a69),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9819476),
	.w1(32'h3aae5f22),
	.w2(32'hbb4d0a1d),
	.w3(32'hbbb2f261),
	.w4(32'hbba068fa),
	.w5(32'h3cc572c5),
	.w6(32'hbaea4337),
	.w7(32'h3af8ba77),
	.w8(32'h3c9cc96a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762a7d),
	.w1(32'hbcb0b129),
	.w2(32'hbd12eb0f),
	.w3(32'h3cb8b1b7),
	.w4(32'h3b22e224),
	.w5(32'hbbd32309),
	.w6(32'h3c029781),
	.w7(32'hbcd1f108),
	.w8(32'hbba9801f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9f365),
	.w1(32'hbc0708b2),
	.w2(32'hbc0f44cc),
	.w3(32'h3b66dbc0),
	.w4(32'h3b05e863),
	.w5(32'hbbf6ad54),
	.w6(32'h3cba86b3),
	.w7(32'hbaff0d36),
	.w8(32'hbc44107f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26084b),
	.w1(32'h3c14d9d8),
	.w2(32'h3c52dd24),
	.w3(32'hbb4a2aae),
	.w4(32'h3b488bd9),
	.w5(32'h3cadcf07),
	.w6(32'hbba01a7e),
	.w7(32'h3b928c15),
	.w8(32'h3c8729e4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956c97),
	.w1(32'hbcafa0dc),
	.w2(32'hbccf6c7d),
	.w3(32'h3c8c49d0),
	.w4(32'h3a21ab0c),
	.w5(32'hbbc9ee84),
	.w6(32'h3b895701),
	.w7(32'hbcaa00f1),
	.w8(32'hbbed33fc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485681),
	.w1(32'h3995f1f9),
	.w2(32'hbaf75f13),
	.w3(32'hbb0f9b68),
	.w4(32'h3a46e56c),
	.w5(32'h3c48c09b),
	.w6(32'hbbdc5af9),
	.w7(32'hbb3290eb),
	.w8(32'h3b70f289),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f391),
	.w1(32'hbc5b6d97),
	.w2(32'hbc77262c),
	.w3(32'h3c7d8753),
	.w4(32'h3b998ffc),
	.w5(32'h3c06ed4f),
	.w6(32'hbb55e8bc),
	.w7(32'hbca5d007),
	.w8(32'h3b1573f2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036a1e),
	.w1(32'hbc0e56b0),
	.w2(32'hbc90de65),
	.w3(32'h3b949f47),
	.w4(32'hbbb23f7f),
	.w5(32'hbc0c41f1),
	.w6(32'hbb2a1efc),
	.w7(32'hbc1838d2),
	.w8(32'hbc277675),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdca88b),
	.w1(32'h3b3e495a),
	.w2(32'h3b810e06),
	.w3(32'hbc44c844),
	.w4(32'hbb4be265),
	.w5(32'hbbd7ebbc),
	.w6(32'h3ca2ef1c),
	.w7(32'h3a2883e3),
	.w8(32'h3ba40769),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0750ef),
	.w1(32'h3bc1001d),
	.w2(32'h3c628340),
	.w3(32'hbb254731),
	.w4(32'hbb0f7347),
	.w5(32'hbb552ba6),
	.w6(32'h3add905d),
	.w7(32'h3ab34a5b),
	.w8(32'hbb2164fb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16cca2),
	.w1(32'h3c1aabaf),
	.w2(32'h3bac377f),
	.w3(32'hbb072d0d),
	.w4(32'h3a519de0),
	.w5(32'hbc06e131),
	.w6(32'h3d037310),
	.w7(32'h3c3160aa),
	.w8(32'hbba76112),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23cb27),
	.w1(32'hbbbe4409),
	.w2(32'h3c110992),
	.w3(32'hbc178743),
	.w4(32'h3bf55773),
	.w5(32'hbb4234eb),
	.w6(32'hbbae4c7e),
	.w7(32'h3b0c4155),
	.w8(32'hbc1eada4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dc3ec),
	.w1(32'h3cdc1ee1),
	.w2(32'h3c979a0b),
	.w3(32'hbc86316c),
	.w4(32'h3c24d5b0),
	.w5(32'hbb769053),
	.w6(32'h3bf1bb7c),
	.w7(32'h3c85e4d0),
	.w8(32'hba8ada5e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2efbd),
	.w1(32'hbbbb6a4d),
	.w2(32'hba2d4f66),
	.w3(32'hbb1d349e),
	.w4(32'hbbb54e3b),
	.w5(32'hbba93d63),
	.w6(32'h3a5a6da1),
	.w7(32'hbb77ef0f),
	.w8(32'hbba19701),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba75db1),
	.w1(32'h3bc5be30),
	.w2(32'h3ba08f4e),
	.w3(32'hbbec5d27),
	.w4(32'hba17893f),
	.w5(32'h3b9cdb0a),
	.w6(32'hbba44d90),
	.w7(32'h3c1793c3),
	.w8(32'hba247fe0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5aaa0),
	.w1(32'hbb3b65b4),
	.w2(32'hbbb61af3),
	.w3(32'h3b86c0dc),
	.w4(32'h3bdde12b),
	.w5(32'hbbd5d68f),
	.w6(32'h3bb1580e),
	.w7(32'h3a630f9e),
	.w8(32'hbbba42e8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68b8e7),
	.w1(32'hbb755eac),
	.w2(32'hbbd0eb98),
	.w3(32'hbab7bb20),
	.w4(32'h3a42e625),
	.w5(32'hbb98df98),
	.w6(32'hbbd3edae),
	.w7(32'hbbbfdf12),
	.w8(32'hbaf17dfa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca58c),
	.w1(32'hba5c7aec),
	.w2(32'hbc60f3a5),
	.w3(32'hbbb1ac62),
	.w4(32'hbbf2ba5f),
	.w5(32'hbc85c6b5),
	.w6(32'hbc555afc),
	.w7(32'hbbc5e1c7),
	.w8(32'hbcca99ae),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa178),
	.w1(32'h3c47c098),
	.w2(32'h3c8b11ab),
	.w3(32'hbc800d69),
	.w4(32'h3bbeb31b),
	.w5(32'h3bae2061),
	.w6(32'hbc25c6e3),
	.w7(32'h3ca096ea),
	.w8(32'h3b24bf08),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b222301),
	.w1(32'hbbe8e402),
	.w2(32'hbc47088f),
	.w3(32'hb9502344),
	.w4(32'hbba968df),
	.w5(32'hbc022c4b),
	.w6(32'hb7296e7c),
	.w7(32'hbc67a0c5),
	.w8(32'hbac2ab0e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b0828),
	.w1(32'h3b607a19),
	.w2(32'h3c104efb),
	.w3(32'hbb386ced),
	.w4(32'hbbada2bb),
	.w5(32'hbc3943af),
	.w6(32'h38eb3a86),
	.w7(32'hbb3496d9),
	.w8(32'hbab439f9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd8b84),
	.w1(32'h3c2344a8),
	.w2(32'h3bc470b9),
	.w3(32'hbc590388),
	.w4(32'h3c0e9d3f),
	.w5(32'h3cf2ec0c),
	.w6(32'h3c969447),
	.w7(32'h3ce9e098),
	.w8(32'h3cdf65b5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb51c5),
	.w1(32'hbce8b470),
	.w2(32'hbcd5a12e),
	.w3(32'h3cfd5259),
	.w4(32'h3bb42413),
	.w5(32'hbbcaadd5),
	.w6(32'hb9714c59),
	.w7(32'hbcb4a03c),
	.w8(32'hbb363c83),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc64734),
	.w1(32'hb9cf0051),
	.w2(32'hb978c230),
	.w3(32'hbb009c96),
	.w4(32'hbaec0860),
	.w5(32'hbae402fc),
	.w6(32'h3c5fbaf9),
	.w7(32'h3b9a6ffe),
	.w8(32'hbb098335),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65776b),
	.w1(32'hbb61f2ae),
	.w2(32'hbc090f98),
	.w3(32'h3b5c4805),
	.w4(32'h34ff0d00),
	.w5(32'hbbdd0eaa),
	.w6(32'h3b7a9e8e),
	.w7(32'h3abca062),
	.w8(32'hbb6b7061),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e6571),
	.w1(32'h3bb3d125),
	.w2(32'hbb8d7a9a),
	.w3(32'h3b72a3de),
	.w4(32'h3c08c322),
	.w5(32'hbbe61259),
	.w6(32'hbb1bc94c),
	.w7(32'h3c0b70c8),
	.w8(32'hbb977464),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc244af6),
	.w1(32'h3b57f0ae),
	.w2(32'h3b37999a),
	.w3(32'hbbf4c0ff),
	.w4(32'h3bc3468b),
	.w5(32'h3bb9260d),
	.w6(32'hbbbce4c5),
	.w7(32'h3bc068d0),
	.w8(32'h3c11e4ef),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16479),
	.w1(32'hbb0ce9b9),
	.w2(32'hb8080176),
	.w3(32'hbb36697c),
	.w4(32'h3b649169),
	.w5(32'h3a6cd716),
	.w6(32'h3a00b073),
	.w7(32'h3bfda632),
	.w8(32'hba81b83a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb728cea),
	.w1(32'h38cf9313),
	.w2(32'hbc09c48b),
	.w3(32'h3b203f66),
	.w4(32'h3b2456c2),
	.w5(32'hbc272cd6),
	.w6(32'h3ac2a89b),
	.w7(32'h3ba5df04),
	.w8(32'hbbb6cabf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491c53),
	.w1(32'hb9c97bdf),
	.w2(32'h3a63724d),
	.w3(32'hbac96dc1),
	.w4(32'h3a078177),
	.w5(32'h3a8b5139),
	.w6(32'hbb0dbb6b),
	.w7(32'h3adf9f20),
	.w8(32'h3a8dcca2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2aab),
	.w1(32'h3b4f9b4a),
	.w2(32'hbb93946e),
	.w3(32'h3bbd7943),
	.w4(32'h3c31a066),
	.w5(32'hbc0e8389),
	.w6(32'hb9d3658f),
	.w7(32'hb9a270cd),
	.w8(32'hbbead821),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66bdc2),
	.w1(32'h3aa90b25),
	.w2(32'hba96b5f9),
	.w3(32'h3aed5e08),
	.w4(32'h3b376c12),
	.w5(32'hbb4cbfeb),
	.w6(32'h3b069f7d),
	.w7(32'h3b2a97e7),
	.w8(32'hbaf3a457),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbea8a),
	.w1(32'hbb2310d1),
	.w2(32'hbad51f8d),
	.w3(32'hbad0bfb4),
	.w4(32'hbb0aeb3d),
	.w5(32'h39fbf4c4),
	.w6(32'hbb11dae9),
	.w7(32'hbb4e5eab),
	.w8(32'h3a8ff9f8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50758a),
	.w1(32'h3b9dc3f4),
	.w2(32'h3b5ef3b9),
	.w3(32'h3bb4c4a9),
	.w4(32'h3b670641),
	.w5(32'h3ad118aa),
	.w6(32'h3a99e5d9),
	.w7(32'h3b358fc7),
	.w8(32'h3a54e067),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaec8c8),
	.w1(32'h3a97bd94),
	.w2(32'hbb5eb28d),
	.w3(32'h3b8423eb),
	.w4(32'h3b148ea4),
	.w5(32'h3b1a750a),
	.w6(32'h3ba8d5a9),
	.w7(32'h3b387b90),
	.w8(32'h3a9eb017),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447578),
	.w1(32'h3bf3ac4c),
	.w2(32'h3bbcc052),
	.w3(32'h3b625d5d),
	.w4(32'h3bede459),
	.w5(32'h3b63d614),
	.w6(32'h3b217d1a),
	.w7(32'h3c0328d7),
	.w8(32'h3b49e6a0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbc1e1),
	.w1(32'hbb9cb525),
	.w2(32'hba3b4054),
	.w3(32'hbb60639c),
	.w4(32'hbab2f69f),
	.w5(32'h3b56a784),
	.w6(32'hbb75f603),
	.w7(32'hbafbef13),
	.w8(32'h3b5ca5cc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a0182),
	.w1(32'hbb84426f),
	.w2(32'hbaed72ab),
	.w3(32'hbb57b849),
	.w4(32'hba1c302f),
	.w5(32'h3bbc7d8b),
	.w6(32'hbb8886e3),
	.w7(32'hbb2cbab9),
	.w8(32'h3b3fd1c7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b75cd),
	.w1(32'h3bef7933),
	.w2(32'h3b8ebfd1),
	.w3(32'h3ba3e7b9),
	.w4(32'h3c0e4efe),
	.w5(32'hbabdfc4b),
	.w6(32'h3b1c3d20),
	.w7(32'h3c1176f3),
	.w8(32'hbb64bf0e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81de9d),
	.w1(32'hbbccd9f2),
	.w2(32'hbc41e74a),
	.w3(32'hbb9af3f6),
	.w4(32'hbba5e059),
	.w5(32'hbc0256a2),
	.w6(32'hbbfaf6c1),
	.w7(32'hbc057c85),
	.w8(32'hbbd44f14),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cda4a),
	.w1(32'hba9e5c6b),
	.w2(32'hbb47c278),
	.w3(32'hbb0fdbcc),
	.w4(32'hb9ef1bba),
	.w5(32'hbb0860ea),
	.w6(32'hbb0f1d6a),
	.w7(32'hba41f4cc),
	.w8(32'hba33056a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eac01),
	.w1(32'hbba1f0d0),
	.w2(32'hbb662daf),
	.w3(32'hbb7c3e35),
	.w4(32'hbb8983cf),
	.w5(32'hba0bd50b),
	.w6(32'hbba7309c),
	.w7(32'hbb72bc76),
	.w8(32'h3884e1d6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad14022),
	.w1(32'h3ae5d057),
	.w2(32'hba92909e),
	.w3(32'h38885867),
	.w4(32'hba17f468),
	.w5(32'hba76c0cd),
	.w6(32'hb976b06b),
	.w7(32'hbaf8e68a),
	.w8(32'hba4ab727),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba719c),
	.w1(32'hbb8180bb),
	.w2(32'hbb908f7f),
	.w3(32'hbb736930),
	.w4(32'hbb4d6319),
	.w5(32'h3b5f0142),
	.w6(32'hbb5cb403),
	.w7(32'hbb139ee5),
	.w8(32'h3b1ca933),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d0c9),
	.w1(32'hba351742),
	.w2(32'hba9779e0),
	.w3(32'hbadd7718),
	.w4(32'hba1fead5),
	.w5(32'h3b2433fc),
	.w6(32'hbb3f7262),
	.w7(32'hbaa2eeff),
	.w8(32'h39df13fd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7d1b0),
	.w1(32'h3ad38f3e),
	.w2(32'hba8bbce8),
	.w3(32'hb994880d),
	.w4(32'h3a50635d),
	.w5(32'hbbf8a009),
	.w6(32'h3abee60c),
	.w7(32'h3a755c33),
	.w8(32'hbbcce114),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc09980),
	.w1(32'hbb22eb31),
	.w2(32'h39e527d9),
	.w3(32'hbb4337ed),
	.w4(32'hbae10335),
	.w5(32'h3a315ef6),
	.w6(32'hbb42a152),
	.w7(32'hb986d637),
	.w8(32'h3a98e9cc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086006),
	.w1(32'h3ad285ea),
	.w2(32'hbb8a58eb),
	.w3(32'h3b9602f1),
	.w4(32'h3a40e8d8),
	.w5(32'h3b36b442),
	.w6(32'h3b92e0ed),
	.w7(32'hbb1d9911),
	.w8(32'hbb76e0b4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21297),
	.w1(32'hbb48d32e),
	.w2(32'h3b84acff),
	.w3(32'h3a323e94),
	.w4(32'h3bc7f257),
	.w5(32'h3a89fd17),
	.w6(32'hbb1d40aa),
	.w7(32'h3bbff1f0),
	.w8(32'h3b8dfe5d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a466),
	.w1(32'h3b4cd029),
	.w2(32'h3a95af17),
	.w3(32'hbabffed7),
	.w4(32'h3b3b78e4),
	.w5(32'h3b4e23e7),
	.w6(32'h3a2cbf65),
	.w7(32'h3a6d6c1e),
	.w8(32'hb92f1fc0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8564b0),
	.w1(32'hbaa481d3),
	.w2(32'h3af9f6e6),
	.w3(32'h3ae5d0df),
	.w4(32'h3b3b1f0d),
	.w5(32'h3a237f8d),
	.w6(32'h3ad7b4cc),
	.w7(32'h3b7790f0),
	.w8(32'h395c37d3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad69379),
	.w1(32'h39911e19),
	.w2(32'hbaf9f9fd),
	.w3(32'h3950dc27),
	.w4(32'hb9da7e18),
	.w5(32'h3b34a86d),
	.w6(32'h3aa75bab),
	.w7(32'hb9bd2efb),
	.w8(32'h3b58450a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9ab6),
	.w1(32'h3b4415cc),
	.w2(32'h3a243700),
	.w3(32'hb9e0b0e3),
	.w4(32'h3a5c708a),
	.w5(32'hba905bd0),
	.w6(32'h3a55bea8),
	.w7(32'h396cbbad),
	.w8(32'hbb2ca132),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc99c41),
	.w1(32'hbad33e24),
	.w2(32'hbc12a5f6),
	.w3(32'h39750eeb),
	.w4(32'hbbe0742e),
	.w5(32'h3adbd09b),
	.w6(32'h3b97911c),
	.w7(32'h3b3c7e2e),
	.w8(32'hbb880dbe),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3400),
	.w1(32'h3a9473c9),
	.w2(32'h3b13c225),
	.w3(32'h3c095230),
	.w4(32'h3b1ecbba),
	.w5(32'hbb9a6073),
	.w6(32'h3c2b88e3),
	.w7(32'h3b75fb24),
	.w8(32'hbbbfbe46),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f71f9),
	.w1(32'h3929d0d7),
	.w2(32'hba073b7f),
	.w3(32'hbada3615),
	.w4(32'h39f050c7),
	.w5(32'h3b318e96),
	.w6(32'hb948dd2c),
	.w7(32'h3995fcfc),
	.w8(32'h3bfb17eb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7755e0),
	.w1(32'h39e7c18f),
	.w2(32'hbb00891e),
	.w3(32'h3b535492),
	.w4(32'h382d050b),
	.w5(32'h390a4275),
	.w6(32'h3be3ad46),
	.w7(32'h3af0ab59),
	.w8(32'hbac11cf2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80e75c),
	.w1(32'hb9f15c47),
	.w2(32'hbabe4e47),
	.w3(32'hb9da193f),
	.w4(32'h39eee192),
	.w5(32'hbb38fe2d),
	.w6(32'hbab0e605),
	.w7(32'hb9b1234e),
	.w8(32'hba7eae7d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53ee0f),
	.w1(32'hbbe7d6e9),
	.w2(32'hbc3e82ca),
	.w3(32'hbbff8fbe),
	.w4(32'hbbcfcac1),
	.w5(32'hbade2432),
	.w6(32'hbb9eecc9),
	.w7(32'hbc08752f),
	.w8(32'hbabaa890),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bebf0),
	.w1(32'hbae5e976),
	.w2(32'hbb8adf75),
	.w3(32'hbb5bdb96),
	.w4(32'hbaab3cdb),
	.w5(32'hbb4889e3),
	.w6(32'hbb55357d),
	.w7(32'hba2e45a8),
	.w8(32'hba7bbad0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3a108),
	.w1(32'hbb8e0e91),
	.w2(32'hbc2d8d69),
	.w3(32'h3ac234a8),
	.w4(32'hbbb6dc4e),
	.w5(32'hbb825a4a),
	.w6(32'h3b25a126),
	.w7(32'hbbfcfaa7),
	.w8(32'hbbf3694e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7fbdc),
	.w1(32'hba9f158c),
	.w2(32'h3a62ad1f),
	.w3(32'hbb8419b5),
	.w4(32'hba20f1ea),
	.w5(32'h3b8c56b0),
	.w6(32'hbbe12609),
	.w7(32'hbad14ba3),
	.w8(32'h3b6365ca),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17082c),
	.w1(32'hb6974a3c),
	.w2(32'hbb2657b1),
	.w3(32'h3ae2beba),
	.w4(32'h39927d2f),
	.w5(32'hbb1dc01d),
	.w6(32'h3abd2eb8),
	.w7(32'h3adaa3ef),
	.w8(32'h3940a144),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944b56),
	.w1(32'hba81496c),
	.w2(32'hbbdb7c96),
	.w3(32'h3bcbf9e7),
	.w4(32'hba384f40),
	.w5(32'hbb8e5b9c),
	.w6(32'h3b88ccf9),
	.w7(32'hbb53273f),
	.w8(32'hbb936111),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb114695),
	.w1(32'h391b8846),
	.w2(32'hbb698161),
	.w3(32'hba8bbf5f),
	.w4(32'hb97df90a),
	.w5(32'hbb96ab42),
	.w6(32'hb8f94f63),
	.w7(32'h39f6df2a),
	.w8(32'hbb99e73d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aea99),
	.w1(32'hbbdff2bc),
	.w2(32'hbc2a131e),
	.w3(32'hbb20df8d),
	.w4(32'hbb80d4d7),
	.w5(32'hbb1f5557),
	.w6(32'hbb9eff30),
	.w7(32'hbbdb0031),
	.w8(32'hbbaa7878),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6773a3),
	.w1(32'hbab5f35d),
	.w2(32'h3aeb5d45),
	.w3(32'h3aeb9e82),
	.w4(32'h3b457074),
	.w5(32'h3a9fad8e),
	.w6(32'hbb0f98b8),
	.w7(32'h3b2d5f9b),
	.w8(32'hb897fb02),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b7418),
	.w1(32'h3c4aec65),
	.w2(32'h3c121ed1),
	.w3(32'h3abb6f81),
	.w4(32'h3bc50f0a),
	.w5(32'h3bfdfe41),
	.w6(32'h3ba56f4e),
	.w7(32'h3b921d6a),
	.w8(32'h3b80caea),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d1092),
	.w1(32'hbb2f59c4),
	.w2(32'hbb7189df),
	.w3(32'h39d3c104),
	.w4(32'h393d3854),
	.w5(32'h3b1bd69d),
	.w6(32'hba4761cc),
	.w7(32'hba753b61),
	.w8(32'hb990f4b4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25ffbb),
	.w1(32'h3b252d2f),
	.w2(32'hb997d029),
	.w3(32'h3ac2b95b),
	.w4(32'h3a8709fe),
	.w5(32'h3b861549),
	.w6(32'h3ba6a61a),
	.w7(32'hba069ca9),
	.w8(32'h3b8cb1ef),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8846ee),
	.w1(32'h38661a74),
	.w2(32'h3b71a971),
	.w3(32'h3b0529e4),
	.w4(32'h3b2a8edc),
	.w5(32'hb9dcff0b),
	.w6(32'hba4c7732),
	.w7(32'h3b58ddc3),
	.w8(32'h396409f8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8fab2),
	.w1(32'h39a5d0c3),
	.w2(32'hb992af0e),
	.w3(32'h394e4526),
	.w4(32'h3a9544e3),
	.w5(32'h39f57362),
	.w6(32'hba13a172),
	.w7(32'h39c1d228),
	.w8(32'hb923c330),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0b49c),
	.w1(32'h3ae6c2f8),
	.w2(32'h3aa4861b),
	.w3(32'hba3fce04),
	.w4(32'h3b961bc9),
	.w5(32'h3ba1eb53),
	.w6(32'hbaf9e56e),
	.w7(32'h3ab20488),
	.w8(32'h3b8fa7c9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a71ba),
	.w1(32'hba9a6d7b),
	.w2(32'hbbd0039d),
	.w3(32'hbb4e6474),
	.w4(32'hbab57863),
	.w5(32'h388174d8),
	.w6(32'h3890e58e),
	.w7(32'hbb0dd14f),
	.w8(32'hba3850e1),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d51d6),
	.w1(32'h3a7d1622),
	.w2(32'hba67eb93),
	.w3(32'hba9f4270),
	.w4(32'h38ca43e6),
	.w5(32'h3a987f5b),
	.w6(32'h3aeef156),
	.w7(32'hba987cfa),
	.w8(32'h3aa55b9d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a83859),
	.w1(32'hbb6f339d),
	.w2(32'hbbe7c876),
	.w3(32'hbb3154bc),
	.w4(32'hbb95e5d9),
	.w5(32'hbbf4ec33),
	.w6(32'hba3d8ba1),
	.w7(32'hbb8f72c8),
	.w8(32'hbbf871cd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bda22),
	.w1(32'hbb69c949),
	.w2(32'hbabe7d5e),
	.w3(32'hbaacb009),
	.w4(32'h3a873cc3),
	.w5(32'hbb9a5e1c),
	.w6(32'hbaa46e41),
	.w7(32'h3afe7ddf),
	.w8(32'hbbacd340),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa8e2),
	.w1(32'h3b1fd791),
	.w2(32'hbba03e55),
	.w3(32'h3b9154c3),
	.w4(32'h3a26d837),
	.w5(32'hbc129b13),
	.w6(32'h3ba762f9),
	.w7(32'hbae94403),
	.w8(32'hbb1883f0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe17175),
	.w1(32'h3b66e65e),
	.w2(32'h3b179bef),
	.w3(32'hbba21d4b),
	.w4(32'h3a9fc072),
	.w5(32'h3b5ef1cc),
	.w6(32'h3b17c62d),
	.w7(32'h3adac3bb),
	.w8(32'hbaa63dd6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1756),
	.w1(32'hbb24de9d),
	.w2(32'hbb8e82aa),
	.w3(32'h3aa735a6),
	.w4(32'h390cd268),
	.w5(32'h397a1d3f),
	.w6(32'hbab3fcdb),
	.w7(32'hba58c446),
	.w8(32'h3a895673),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b141127),
	.w1(32'h3b987a0b),
	.w2(32'hb893360d),
	.w3(32'h3bca2a41),
	.w4(32'h3b849d1d),
	.w5(32'h3c2f0fc3),
	.w6(32'h3bd58004),
	.w7(32'h3b92f8c0),
	.w8(32'h3c185fca),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ba0a),
	.w1(32'h3bc8bba6),
	.w2(32'h3bf3d743),
	.w3(32'h3a37e977),
	.w4(32'h3bd02f46),
	.w5(32'h3b1f6a0d),
	.w6(32'h3a36cccf),
	.w7(32'h3bb3b54e),
	.w8(32'hb9102c38),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f31ce),
	.w1(32'h3b826eb6),
	.w2(32'hb91ec7d0),
	.w3(32'h3b74521d),
	.w4(32'h3acdc417),
	.w5(32'h3a341463),
	.w6(32'h3c14798b),
	.w7(32'h3b1b994f),
	.w8(32'h3b35c54a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b522d55),
	.w1(32'h3b75a194),
	.w2(32'hba91dd7d),
	.w3(32'hba4b42fd),
	.w4(32'h3b39f3a2),
	.w5(32'h3b4a586b),
	.w6(32'h3a76a744),
	.w7(32'hb9d0edba),
	.w8(32'h3b2fb873),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44cebc),
	.w1(32'h3bd4063e),
	.w2(32'h39f6eb69),
	.w3(32'h3aee4b25),
	.w4(32'h3ba7ff52),
	.w5(32'h388f5e80),
	.w6(32'h3b03c4de),
	.w7(32'h3b38a634),
	.w8(32'h3af119f5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcf0cd),
	.w1(32'hba25f310),
	.w2(32'hba923c17),
	.w3(32'h3a06f7b2),
	.w4(32'hb9130b17),
	.w5(32'hbba69eff),
	.w6(32'h3ad7bc51),
	.w7(32'h3b27d2e0),
	.w8(32'hbbb7ef04),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2509dc),
	.w1(32'hbc13be17),
	.w2(32'hbc0d75d7),
	.w3(32'hbba923aa),
	.w4(32'hbba66408),
	.w5(32'hbb8d5f9a),
	.w6(32'hbb94ed9a),
	.w7(32'hbba691dd),
	.w8(32'hbadde30e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a792855),
	.w1(32'h3a0c8a54),
	.w2(32'h39c771ee),
	.w3(32'h3a4b7569),
	.w4(32'hbabc2197),
	.w5(32'hbb6a3f98),
	.w6(32'h3a0c6c1f),
	.w7(32'hb9c961fc),
	.w8(32'hbb5e8ac6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944686),
	.w1(32'hbaf1f673),
	.w2(32'h3b0015f9),
	.w3(32'hbb0bce83),
	.w4(32'h3b0bd15d),
	.w5(32'h3a1ca411),
	.w6(32'h3aab37bf),
	.w7(32'h3b3e7f38),
	.w8(32'hba12917d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aa0e1),
	.w1(32'hbb7952fc),
	.w2(32'hbad0f489),
	.w3(32'hbba0780b),
	.w4(32'hbacaab59),
	.w5(32'hbacfcc5a),
	.w6(32'hbbbe7570),
	.w7(32'hbb72d663),
	.w8(32'hb98f8328),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab62bb7),
	.w1(32'hbb26a4ce),
	.w2(32'hbb27fc72),
	.w3(32'h397394af),
	.w4(32'hbb8a8aac),
	.w5(32'hbb03bf14),
	.w6(32'h3ad8703e),
	.w7(32'hbb19f8cc),
	.w8(32'hb9e7acb6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacada7a),
	.w1(32'h3abe5e66),
	.w2(32'hbb5ac282),
	.w3(32'h3aa8dda3),
	.w4(32'hba4598b6),
	.w5(32'hbb0e92f8),
	.w6(32'h3bb7f887),
	.w7(32'h39d65e1f),
	.w8(32'h3a89e90e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e4335),
	.w1(32'h3b1c99f9),
	.w2(32'h3b9fa5be),
	.w3(32'hbb9ba0bd),
	.w4(32'h3b0f2e4e),
	.w5(32'h39d90a5c),
	.w6(32'hb8ad8de9),
	.w7(32'h3a4e21f5),
	.w8(32'h3a372b6d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb550d5a),
	.w1(32'h3926cd58),
	.w2(32'h3b30eeba),
	.w3(32'hbb14b946),
	.w4(32'h3aeec485),
	.w5(32'h3aceba46),
	.w6(32'hbac0f452),
	.w7(32'h3a5a3323),
	.w8(32'h39efc722),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a533f1c),
	.w1(32'h3b945970),
	.w2(32'hbabfc8ba),
	.w3(32'h3b8bd5d5),
	.w4(32'hb9d4858c),
	.w5(32'hbbb5c6bd),
	.w6(32'h3c0e0b96),
	.w7(32'h3ba3fa8f),
	.w8(32'hbbcf48a0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43f342),
	.w1(32'hb9a5f144),
	.w2(32'hbb6387bf),
	.w3(32'h3b1a0f0c),
	.w4(32'hb9ff7e9b),
	.w5(32'hbaa95504),
	.w6(32'hb96346ac),
	.w7(32'hbad8179a),
	.w8(32'hba9c4cd8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22aefc),
	.w1(32'h3ac1bbe3),
	.w2(32'h3abd666b),
	.w3(32'hbb5d20b5),
	.w4(32'h3b11fa87),
	.w5(32'h3aa1e671),
	.w6(32'hb9a478e8),
	.w7(32'h3ae94813),
	.w8(32'h39f2da7b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a15ca),
	.w1(32'h3a31617d),
	.w2(32'hba6e5732),
	.w3(32'hb6df84a8),
	.w4(32'h3b1de997),
	.w5(32'hb9163d3d),
	.w6(32'h3a828e97),
	.w7(32'hb971b1c3),
	.w8(32'hb93d9e4b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823942),
	.w1(32'hbb28341d),
	.w2(32'hbbdbe658),
	.w3(32'hb9f149f6),
	.w4(32'hbb23bff4),
	.w5(32'h3b24b7f0),
	.w6(32'h3b715008),
	.w7(32'h398c1086),
	.w8(32'h3a22468e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971e15),
	.w1(32'h3b55bbb1),
	.w2(32'hba5ce650),
	.w3(32'h3af553da),
	.w4(32'h3ac239ad),
	.w5(32'hbb040f00),
	.w6(32'hb9c30913),
	.w7(32'h3b21bc71),
	.w8(32'hb9f075a9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb598af7),
	.w1(32'hbba41050),
	.w2(32'hbc0893d1),
	.w3(32'hbac9edd0),
	.w4(32'hbbd5150c),
	.w5(32'hbb3b8985),
	.w6(32'h3a564635),
	.w7(32'hbb88873c),
	.w8(32'hbb3c5371),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd6a97),
	.w1(32'h3a220a8e),
	.w2(32'h3b311651),
	.w3(32'h3983a03f),
	.w4(32'h3aeef506),
	.w5(32'h3ac77930),
	.w6(32'h37ee915d),
	.w7(32'h3b2c3324),
	.w8(32'hba61aacd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a241),
	.w1(32'hba123264),
	.w2(32'h3a535e7f),
	.w3(32'hb96231a5),
	.w4(32'h3b7b28b6),
	.w5(32'hbacf51f6),
	.w6(32'h3993b84e),
	.w7(32'h3ab62083),
	.w8(32'hbad02b3d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12839b),
	.w1(32'hb98ade05),
	.w2(32'hbb0efcbf),
	.w3(32'hbab119f4),
	.w4(32'hbb26c0ac),
	.w5(32'hbbe0cb31),
	.w6(32'h3a134312),
	.w7(32'hbb108564),
	.w8(32'hbbd49d69),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb66774),
	.w1(32'hbb6a66f9),
	.w2(32'hbaa8434b),
	.w3(32'hbb580cf1),
	.w4(32'hba74dacd),
	.w5(32'hba73978a),
	.w6(32'hbb8d6d79),
	.w7(32'hba2e996e),
	.w8(32'h399c86cf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e1bc44),
	.w1(32'hb9500b29),
	.w2(32'hba52f3eb),
	.w3(32'hbabd9376),
	.w4(32'h3a72a228),
	.w5(32'hbba37111),
	.w6(32'hbadc0653),
	.w7(32'hba4294c1),
	.w8(32'hbba35cb6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7601c),
	.w1(32'hbb881b63),
	.w2(32'hbc028240),
	.w3(32'hb9c0f94a),
	.w4(32'hbb881d90),
	.w5(32'hbbc599cd),
	.w6(32'hbafb15e3),
	.w7(32'hbb98119b),
	.w8(32'hbbc48e7f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090fdc),
	.w1(32'hb9d22f0c),
	.w2(32'hbb74b054),
	.w3(32'hba39ef08),
	.w4(32'hbb68f494),
	.w5(32'hb7c602cb),
	.w6(32'hbaac1477),
	.w7(32'hbbd37f78),
	.w8(32'h3945543c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09fc3f),
	.w1(32'hba987fae),
	.w2(32'hbaa052bd),
	.w3(32'hbb1e6117),
	.w4(32'hb7bd9ca4),
	.w5(32'h3b03d44d),
	.w6(32'hbb44406d),
	.w7(32'hba97b0ae),
	.w8(32'h3b38384d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa4ea0),
	.w1(32'h3b8d3979),
	.w2(32'h3b688df1),
	.w3(32'h3b39952a),
	.w4(32'h3ae10cef),
	.w5(32'h3ab01add),
	.w6(32'h3c324e45),
	.w7(32'h3b86db39),
	.w8(32'h3877ad92),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee1424),
	.w1(32'h3b530708),
	.w2(32'h3a8291f4),
	.w3(32'h3c1c4f4a),
	.w4(32'h3a5bf551),
	.w5(32'hbaec8b8d),
	.w6(32'h3c3b2f7d),
	.w7(32'h3acffef0),
	.w8(32'hbae1e921),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898004),
	.w1(32'h3bc0fce6),
	.w2(32'hbb92ddf9),
	.w3(32'h3b4cbafe),
	.w4(32'h3b87f0dd),
	.w5(32'hbb55b1c6),
	.w6(32'h3ab7d331),
	.w7(32'hbb50b310),
	.w8(32'hbb01b85a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46826b),
	.w1(32'hba3ec197),
	.w2(32'hbb3fcba5),
	.w3(32'hbad637fb),
	.w4(32'hbb1d64ba),
	.w5(32'hb90c91e2),
	.w6(32'h3a2b653d),
	.w7(32'hbb1cc523),
	.w8(32'h3b0c9c6b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c70e1),
	.w1(32'hbb97ae14),
	.w2(32'hbbeb7544),
	.w3(32'h39a4f53a),
	.w4(32'hbbdba40d),
	.w5(32'hbbbbe611),
	.w6(32'h3b112565),
	.w7(32'hba3b822d),
	.w8(32'hbba9d747),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc94d12),
	.w1(32'h3acab76b),
	.w2(32'hbaca59c5),
	.w3(32'hbc045cbd),
	.w4(32'h3b7cef6f),
	.w5(32'h3b7b5097),
	.w6(32'hbb32e50a),
	.w7(32'hba097d61),
	.w8(32'h3aa46c02),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be800c7),
	.w1(32'h3b57a05c),
	.w2(32'hba812f36),
	.w3(32'h3bcdd769),
	.w4(32'h3b653c5a),
	.w5(32'hbc18be6a),
	.w6(32'h3b804dca),
	.w7(32'h3b3766d3),
	.w8(32'hbbbf5cb7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf1a19),
	.w1(32'hbada5215),
	.w2(32'hb9edb990),
	.w3(32'hbbafc336),
	.w4(32'hbb3b3ce8),
	.w5(32'hb9e2e1d9),
	.w6(32'hbb8ed7c5),
	.w7(32'hbb3a876a),
	.w8(32'hba6e0509),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba578b78),
	.w1(32'h3a91dc34),
	.w2(32'h3b0b6d5e),
	.w3(32'h3b0263fe),
	.w4(32'h3a846623),
	.w5(32'hbb6b0e7d),
	.w6(32'h3b9587fb),
	.w7(32'h3afbdf14),
	.w8(32'hba4a05a1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eb80b),
	.w1(32'hb80865da),
	.w2(32'hba868932),
	.w3(32'hbb5a9bc9),
	.w4(32'hb9a4dcb2),
	.w5(32'hbb643aa6),
	.w6(32'hb90cf2c7),
	.w7(32'hba45c681),
	.w8(32'hba864346),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74e215),
	.w1(32'h3b08fafe),
	.w2(32'hbb370d26),
	.w3(32'h3ace7927),
	.w4(32'h3a31e9b7),
	.w5(32'h3a9d1f27),
	.w6(32'hbb05d157),
	.w7(32'hb9c8f9b4),
	.w8(32'h3a761464),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50c6cf),
	.w1(32'hbbb20f54),
	.w2(32'hbbb7ba1d),
	.w3(32'h3ad643b8),
	.w4(32'hbac78854),
	.w5(32'hbbd89705),
	.w6(32'hbaf50dd3),
	.w7(32'hbaada940),
	.w8(32'hbc02dd5c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2493cf),
	.w1(32'h3a509b07),
	.w2(32'hba2667b4),
	.w3(32'hbb70517d),
	.w4(32'h3b90f2fd),
	.w5(32'hbb6649c0),
	.w6(32'hbb6cde5c),
	.w7(32'h3acd1e60),
	.w8(32'hbb372d86),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fcaf),
	.w1(32'hbbdafcd7),
	.w2(32'hbb8eabd3),
	.w3(32'hbbed18af),
	.w4(32'hbac3f29b),
	.w5(32'h3b2a9a42),
	.w6(32'hbbe3857b),
	.w7(32'hbb1ba38d),
	.w8(32'h3b39e107),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2ade2),
	.w1(32'hbae476c6),
	.w2(32'hbb8dffe3),
	.w3(32'h3b1da5c7),
	.w4(32'hb99dd515),
	.w5(32'hbb6111c4),
	.w6(32'h3b0caa54),
	.w7(32'hb812235c),
	.w8(32'hbb7f49ef),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d7767),
	.w1(32'h3aacc0f2),
	.w2(32'hbb158a1d),
	.w3(32'h3afac946),
	.w4(32'h3a652ab3),
	.w5(32'h3af1d45a),
	.w6(32'h3ae380aa),
	.w7(32'h3a649c7d),
	.w8(32'hbab609d6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5cd49),
	.w1(32'h3ad696b5),
	.w2(32'h392a0617),
	.w3(32'hbb2d4801),
	.w4(32'h39e60092),
	.w5(32'hbb3fb13c),
	.w6(32'h3a2e5419),
	.w7(32'hba409689),
	.w8(32'hbb6b06b1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafd668),
	.w1(32'h3a211f46),
	.w2(32'h3b4030a4),
	.w3(32'hba6a257c),
	.w4(32'h3b6181b3),
	.w5(32'hbad5118b),
	.w6(32'hb98bc1d1),
	.w7(32'h3b109055),
	.w8(32'hbb3f0691),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a763d59),
	.w1(32'hbac4b5dd),
	.w2(32'h39acb546),
	.w3(32'hbb1c8545),
	.w4(32'hba9b5b9b),
	.w5(32'h3b34bd41),
	.w6(32'hbae1d61e),
	.w7(32'hbab12431),
	.w8(32'h3a8e063a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8a067),
	.w1(32'hbb8d684c),
	.w2(32'hbb6bc50d),
	.w3(32'h3b09511a),
	.w4(32'hb953f23b),
	.w5(32'hbb1959c3),
	.w6(32'h3ac9a3f1),
	.w7(32'h39f36afd),
	.w8(32'hbb1dbad8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae189),
	.w1(32'h3b22a29d),
	.w2(32'h3b9aa318),
	.w3(32'hbaaf2260),
	.w4(32'h3baf05ca),
	.w5(32'hbb24f050),
	.w6(32'hbaa215cb),
	.w7(32'h3b93e13c),
	.w8(32'hbb97b298),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298bca),
	.w1(32'h3b420b86),
	.w2(32'h3ac75257),
	.w3(32'hba8f7dc6),
	.w4(32'h3b519291),
	.w5(32'hbaa8bc4f),
	.w6(32'hbacd2c00),
	.w7(32'h3b5e837d),
	.w8(32'hb95fae0c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fccd1),
	.w1(32'hbb0f7c12),
	.w2(32'hbafc7d04),
	.w3(32'hbae4c51e),
	.w4(32'hba803a16),
	.w5(32'h3b0343fa),
	.w6(32'hbb2f18d8),
	.w7(32'hba916f24),
	.w8(32'h3a4f1329),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b555),
	.w1(32'h399883bf),
	.w2(32'h3afc636f),
	.w3(32'hbb656b85),
	.w4(32'h3bb2992f),
	.w5(32'h3bf321e3),
	.w6(32'hbb95af3e),
	.w7(32'h3b8988a1),
	.w8(32'h3bb4abe8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b9505),
	.w1(32'h3b063808),
	.w2(32'h3b15b814),
	.w3(32'h3b9251b7),
	.w4(32'h3b863990),
	.w5(32'hbaadc535),
	.w6(32'h3b007d6d),
	.w7(32'h3ba13dc2),
	.w8(32'hbab1371b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb281baa),
	.w1(32'hbab136f9),
	.w2(32'hbb43d444),
	.w3(32'hbb02df18),
	.w4(32'h38351a11),
	.w5(32'hbac4f3d4),
	.w6(32'h3a18141f),
	.w7(32'h3a2b4e97),
	.w8(32'hbb577797),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da7e9a),
	.w1(32'hba9968e0),
	.w2(32'hb9264b7d),
	.w3(32'hba410ec1),
	.w4(32'hba6aeb73),
	.w5(32'hbb203344),
	.w6(32'hbae03cbc),
	.w7(32'hbac4fe28),
	.w8(32'hbb6273a8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60a98d),
	.w1(32'hbb472f5b),
	.w2(32'hbab0d8ff),
	.w3(32'hbb0cf0e2),
	.w4(32'h39d39591),
	.w5(32'hbac02094),
	.w6(32'hbb110f0e),
	.w7(32'h3a0d903a),
	.w8(32'hba470234),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9d10),
	.w1(32'hbb878c92),
	.w2(32'hbc1cffbb),
	.w3(32'hbb797323),
	.w4(32'hbb1410ff),
	.w5(32'hbb8c33a2),
	.w6(32'h3ab9dc59),
	.w7(32'hb928a24e),
	.w8(32'hbc07a75d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853313),
	.w1(32'hbb9ae05f),
	.w2(32'hbbc4e9dc),
	.w3(32'hbaa57498),
	.w4(32'hba50600b),
	.w5(32'hba1fce39),
	.w6(32'h3b32ebbb),
	.w7(32'h3b85c7e1),
	.w8(32'hba949cef),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9a8fd),
	.w1(32'h3bcec6f0),
	.w2(32'h3baf1fe6),
	.w3(32'h3b63c7c8),
	.w4(32'h3bea29ee),
	.w5(32'hbb3d3760),
	.w6(32'h3b858345),
	.w7(32'h3bf23ada),
	.w8(32'hbaf050ce),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13be72),
	.w1(32'hbb0a3fff),
	.w2(32'hbc3d8dea),
	.w3(32'h3b8a5f52),
	.w4(32'hbaf50ebd),
	.w5(32'hbc10b36b),
	.w6(32'h3aeb371c),
	.w7(32'hbbd2847a),
	.w8(32'hbc08149c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabadb9d),
	.w1(32'hb9c0db0c),
	.w2(32'hb932a5f4),
	.w3(32'hbad29d5b),
	.w4(32'hbacada91),
	.w5(32'h3b581e83),
	.w6(32'hbb1dba27),
	.w7(32'hb999a805),
	.w8(32'h3b417a27),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c900),
	.w1(32'h38d0203c),
	.w2(32'hbaaa6387),
	.w3(32'h3abf5a09),
	.w4(32'hbac5a34a),
	.w5(32'h3b1951f7),
	.w6(32'h3b00310f),
	.w7(32'hbaa3dace),
	.w8(32'hb9c77e64),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c214b82),
	.w1(32'h3c461bd1),
	.w2(32'h397eba40),
	.w3(32'h3c2b972d),
	.w4(32'h3bd5c619),
	.w5(32'hbc0963af),
	.w6(32'h3bca9f64),
	.w7(32'h3c3f9d6f),
	.w8(32'hbb78b46e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad22e69),
	.w1(32'hba365b56),
	.w2(32'hbaf38e04),
	.w3(32'h3b7d5315),
	.w4(32'hb9539722),
	.w5(32'hbba73c8b),
	.w6(32'h3b9cb35c),
	.w7(32'h3922d478),
	.w8(32'hbbd7df1e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d8564),
	.w1(32'hbb42b7b6),
	.w2(32'hbc205743),
	.w3(32'h3b2aec82),
	.w4(32'h38cdd0f8),
	.w5(32'hbb2f6c54),
	.w6(32'h3a89bd52),
	.w7(32'h3b15044f),
	.w8(32'h3ab5f3bf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85a252),
	.w1(32'h3bc89ca2),
	.w2(32'h398a4c5f),
	.w3(32'h3aadac76),
	.w4(32'h3b87f3af),
	.w5(32'h3bc7f590),
	.w6(32'h3c173544),
	.w7(32'h3b94e43f),
	.w8(32'h3bd926da),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b321),
	.w1(32'hba4e4083),
	.w2(32'hba157b4f),
	.w3(32'hbb893cb6),
	.w4(32'h3924b545),
	.w5(32'h3baa89a8),
	.w6(32'hbb3611fc),
	.w7(32'hbab3208f),
	.w8(32'h3a162fa5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf1fcc),
	.w1(32'h3adb4e0c),
	.w2(32'hba7e777c),
	.w3(32'hb99d4fb7),
	.w4(32'h3a4580a0),
	.w5(32'hbb2846a3),
	.w6(32'h3b90a4b1),
	.w7(32'h3a84bcc2),
	.w8(32'hbacc1417),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ad82),
	.w1(32'hbb4626b8),
	.w2(32'hbb7303ed),
	.w3(32'hbb2b3202),
	.w4(32'hbaf4d034),
	.w5(32'h39313fa2),
	.w6(32'hb996004c),
	.w7(32'hbacb1946),
	.w8(32'h39d07888),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84fd6d),
	.w1(32'h3a9efcf7),
	.w2(32'h3b402360),
	.w3(32'h39d14774),
	.w4(32'hba21d99f),
	.w5(32'hb9c9e2a6),
	.w6(32'hba87d335),
	.w7(32'h3a767d5a),
	.w8(32'hbb43ceb9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba621ab),
	.w1(32'h3c4df893),
	.w2(32'h3c08be2b),
	.w3(32'h3c161bd5),
	.w4(32'h3c01ae00),
	.w5(32'hb8576373),
	.w6(32'h3c247c51),
	.w7(32'h3c1baa02),
	.w8(32'hbaca1cf3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175fae),
	.w1(32'hbb8ce52d),
	.w2(32'hbb567e9a),
	.w3(32'h3c049ad8),
	.w4(32'h3b599ce4),
	.w5(32'h3b43610f),
	.w6(32'h3b21866f),
	.w7(32'h3a4eebe5),
	.w8(32'h3a0f76d5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba205981),
	.w1(32'h3aa69942),
	.w2(32'hbbacedb2),
	.w3(32'h3c0a71e9),
	.w4(32'h3aba30bc),
	.w5(32'h393f3a98),
	.w6(32'hbae915d8),
	.w7(32'h39fc49fa),
	.w8(32'h38c59089),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969fc3),
	.w1(32'hba72976a),
	.w2(32'hbb1fe0c4),
	.w3(32'h3aef24e3),
	.w4(32'h3b4064e0),
	.w5(32'hbb73a794),
	.w6(32'h3bd6cc7f),
	.w7(32'h3ac3f0cf),
	.w8(32'hbb206b1c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a5978),
	.w1(32'h3b7e957f),
	.w2(32'h3a75237e),
	.w3(32'hbba2deeb),
	.w4(32'hbbae7fc0),
	.w5(32'hba95a60a),
	.w6(32'hbb89bf52),
	.w7(32'hbb7729c0),
	.w8(32'hbad10ecd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d0a34),
	.w1(32'hba729e06),
	.w2(32'hbc1c3314),
	.w3(32'h3bf11cc2),
	.w4(32'h3a4c8075),
	.w5(32'hbc11488c),
	.w6(32'h3b22353f),
	.w7(32'h3af423a8),
	.w8(32'hbc1388d0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b944),
	.w1(32'hbb7221ce),
	.w2(32'hbaf98bf2),
	.w3(32'h3bb7a204),
	.w4(32'h3adc4524),
	.w5(32'h3ae633eb),
	.w6(32'hbbf2a7a3),
	.w7(32'h3a83bcd8),
	.w8(32'h3a484c53),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa61366),
	.w1(32'hbb07297f),
	.w2(32'h3aa004f7),
	.w3(32'h3beff1e0),
	.w4(32'hb94157e1),
	.w5(32'hba5ed14a),
	.w6(32'h3baa1934),
	.w7(32'h3ab93be1),
	.w8(32'hbb181bd7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba991589),
	.w1(32'h3ad6e954),
	.w2(32'hbb295625),
	.w3(32'h3a568ec3),
	.w4(32'h39f26a29),
	.w5(32'hbb9809bb),
	.w6(32'h3af7baa7),
	.w7(32'h3a304e16),
	.w8(32'h3b1759b5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72192e),
	.w1(32'hbb0705ed),
	.w2(32'h394107f8),
	.w3(32'h3be220e2),
	.w4(32'h3bfef5d0),
	.w5(32'h3b061a74),
	.w6(32'h3c85b4e5),
	.w7(32'h3a53a233),
	.w8(32'h38c1b05c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba426449),
	.w1(32'h3b0a380d),
	.w2(32'h38e4a772),
	.w3(32'h3b699f98),
	.w4(32'h3ba9475e),
	.w5(32'hba872512),
	.w6(32'h3841c292),
	.w7(32'h3a8c15db),
	.w8(32'hb8adcbe0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb633f3a),
	.w1(32'hba33960e),
	.w2(32'hba734b73),
	.w3(32'h3b809bb6),
	.w4(32'h3b7af444),
	.w5(32'h3ae6c102),
	.w6(32'h3b530418),
	.w7(32'h3b8dccf1),
	.w8(32'hbad4bb51),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978f405),
	.w1(32'hba2ad20b),
	.w2(32'hba7067b9),
	.w3(32'h3af1551d),
	.w4(32'h3b0db609),
	.w5(32'h393bf406),
	.w6(32'hba90a651),
	.w7(32'hbac0323c),
	.w8(32'h3b832c2b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45426e),
	.w1(32'h3aa114fc),
	.w2(32'h3b153d1c),
	.w3(32'h3b04d66b),
	.w4(32'h3b518e93),
	.w5(32'h3bd30c5e),
	.w6(32'h39e7a576),
	.w7(32'hbac9e352),
	.w8(32'h3b611ca5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba394a0),
	.w1(32'hbc0cd4ec),
	.w2(32'hbc23bbae),
	.w3(32'h3b3e994c),
	.w4(32'hbb32735f),
	.w5(32'hbc06bfc1),
	.w6(32'hba81b742),
	.w7(32'hbb9773de),
	.w8(32'hbbaadf0c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b90b2),
	.w1(32'hbb467681),
	.w2(32'hbb9052ee),
	.w3(32'hba9d032d),
	.w4(32'hbb56d2cd),
	.w5(32'hbb910c21),
	.w6(32'h3adcb349),
	.w7(32'hba24765d),
	.w8(32'hbac1bc97),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac18ec8),
	.w1(32'hbbad1c9c),
	.w2(32'hbc1a6221),
	.w3(32'hbab8709c),
	.w4(32'hbb9fe354),
	.w5(32'h39a9012a),
	.w6(32'h3bfcebe5),
	.w7(32'hbb8a6674),
	.w8(32'hbbd23097),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b167a0f),
	.w1(32'hbb2f453f),
	.w2(32'hbba30499),
	.w3(32'h3c377eea),
	.w4(32'h3bc9ba9c),
	.w5(32'h3ab17a58),
	.w6(32'h3bccb534),
	.w7(32'h3bbae024),
	.w8(32'h39ef7d64),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f253),
	.w1(32'hba4c005e),
	.w2(32'h3b3fa50e),
	.w3(32'h3b9b8864),
	.w4(32'h3a29c7ba),
	.w5(32'h3a1ba9b2),
	.w6(32'hbab3088b),
	.w7(32'hbb404abc),
	.w8(32'hbafec6db),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9ccac),
	.w1(32'h39caacf8),
	.w2(32'h3a4aef07),
	.w3(32'h3a82535d),
	.w4(32'h3a723831),
	.w5(32'h3b340285),
	.w6(32'hbb58f52a),
	.w7(32'h38431296),
	.w8(32'h3b78e9bf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fd815),
	.w1(32'h3be1ba10),
	.w2(32'h3aa5fefd),
	.w3(32'h3bd8d99d),
	.w4(32'h3b8f3d1d),
	.w5(32'h3bb0d8b9),
	.w6(32'hbadb94f0),
	.w7(32'hb9fd48c8),
	.w8(32'hbbd59ece),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b355),
	.w1(32'hbbd9b196),
	.w2(32'hbbd30560),
	.w3(32'h3bd3c462),
	.w4(32'h3ba1f528),
	.w5(32'h3b4fd83c),
	.w6(32'hbb8fca20),
	.w7(32'hbb3846ec),
	.w8(32'h396249a9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9486f),
	.w1(32'hbac0bf40),
	.w2(32'h3ababd71),
	.w3(32'h3c2c02bb),
	.w4(32'h3c59f13e),
	.w5(32'h3b41ba64),
	.w6(32'h3beea481),
	.w7(32'h3bec719d),
	.w8(32'h3ad3c856),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b366431),
	.w1(32'h3ab48cb2),
	.w2(32'h39cb3c03),
	.w3(32'h3bc608fd),
	.w4(32'h3bed657b),
	.w5(32'h3999a5bd),
	.w6(32'h3bc3984b),
	.w7(32'h3b32742a),
	.w8(32'h3a833e92),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d563b),
	.w1(32'h3b121f3c),
	.w2(32'h3ae788cc),
	.w3(32'h3b1c51a1),
	.w4(32'h3b82e43f),
	.w5(32'hbba5dce7),
	.w6(32'h3a909703),
	.w7(32'h3b38cf53),
	.w8(32'hbb2f7498),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0b8b),
	.w1(32'h3bac607b),
	.w2(32'h3b242d4d),
	.w3(32'hbb895a89),
	.w4(32'hbb803a27),
	.w5(32'hbaa025ef),
	.w6(32'hba5ea8a2),
	.w7(32'hbba1ca3e),
	.w8(32'hba4b4a88),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fcbc92),
	.w1(32'h3a92d902),
	.w2(32'hb837e7f0),
	.w3(32'hbaef1a18),
	.w4(32'hbb253da6),
	.w5(32'hbb984b64),
	.w6(32'h3b016937),
	.w7(32'h3a2971a0),
	.w8(32'hba1841d1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fbe1f),
	.w1(32'hb98a98dd),
	.w2(32'hbb1eb52a),
	.w3(32'hbb294ae5),
	.w4(32'hbaf42b11),
	.w5(32'h3a236c83),
	.w6(32'h3b33fb9d),
	.w7(32'hbb8fed9d),
	.w8(32'h3aab1d4d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54f900),
	.w1(32'hbb64f350),
	.w2(32'hbc1fc146),
	.w3(32'hbb94c4e4),
	.w4(32'hbb30f570),
	.w5(32'hbb78c1af),
	.w6(32'hba227ecd),
	.w7(32'hbb361b9a),
	.w8(32'hbbc3f907),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91de51a),
	.w1(32'hbafba052),
	.w2(32'h3a320971),
	.w3(32'h3b44f4a7),
	.w4(32'h3b577551),
	.w5(32'h39cc6543),
	.w6(32'h3a102b0f),
	.w7(32'h3a920cf0),
	.w8(32'h3a8c0644),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b76799),
	.w1(32'h3b90fd7e),
	.w2(32'h3b10cd17),
	.w3(32'hbb29d699),
	.w4(32'h3b7db7bc),
	.w5(32'h3b02c501),
	.w6(32'h3c05ce96),
	.w7(32'h3b92814e),
	.w8(32'hbb442119),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule