module layer_10_featuremap_109(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940f0cb),
	.w1(32'hb79250c1),
	.w2(32'hb95ae2e4),
	.w3(32'h3921f019),
	.w4(32'h38a6354c),
	.w5(32'hb94cf15d),
	.w6(32'hb8e14250),
	.w7(32'h39870120),
	.w8(32'h39d9931f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6df9c),
	.w1(32'h3867c977),
	.w2(32'hb4d32628),
	.w3(32'hb797985e),
	.w4(32'h392b9a18),
	.w5(32'h38de74cb),
	.w6(32'h38e8e880),
	.w7(32'h38ae2e1d),
	.w8(32'h388954b6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8641518),
	.w1(32'hb97994f8),
	.w2(32'hb92af2f1),
	.w3(32'hb6e305f8),
	.w4(32'hb97204c3),
	.w5(32'hb9801db8),
	.w6(32'hb8b5459f),
	.w7(32'hb8cc0aa0),
	.w8(32'hb8a5e072),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c672e),
	.w1(32'hb9fe8f1f),
	.w2(32'hb9f28c3e),
	.w3(32'hb97fc03e),
	.w4(32'hb8bdd5da),
	.w5(32'hb91d9aa3),
	.w6(32'h37ae8bb0),
	.w7(32'hb8f95cda),
	.w8(32'hb9437243),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a1a3a),
	.w1(32'hb909caf9),
	.w2(32'hb9098948),
	.w3(32'hb859efd0),
	.w4(32'h38696323),
	.w5(32'hb740521a),
	.w6(32'hb8941c68),
	.w7(32'hb9799f34),
	.w8(32'h38959d4b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb879ad6a),
	.w1(32'h395a97fb),
	.w2(32'h39851e87),
	.w3(32'hb88f107b),
	.w4(32'h3946f302),
	.w5(32'h396e1ee7),
	.w6(32'h39520f1d),
	.w7(32'h396bbbc3),
	.w8(32'h39833bc2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945973f),
	.w1(32'hb8cc51e7),
	.w2(32'hb8e717d7),
	.w3(32'h393eb36c),
	.w4(32'h38bd9126),
	.w5(32'h383ebc0c),
	.w6(32'hb7fef6c8),
	.w7(32'hb909730e),
	.w8(32'hb8116995),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f34c6e),
	.w1(32'h397005cf),
	.w2(32'h39cd432b),
	.w3(32'hb923d9e7),
	.w4(32'h3998736a),
	.w5(32'h39af700e),
	.w6(32'h389537e4),
	.w7(32'h393c1fa6),
	.w8(32'h39b04546),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e3133),
	.w1(32'h3829bc59),
	.w2(32'h38cdfc8e),
	.w3(32'h3999141a),
	.w4(32'h3849100a),
	.w5(32'h3945530b),
	.w6(32'h3824cd59),
	.w7(32'h38a4255b),
	.w8(32'h38e6dd28),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8107db2),
	.w1(32'hb98b6475),
	.w2(32'hb9d1b3eb),
	.w3(32'h39105676),
	.w4(32'hb84dd200),
	.w5(32'hb9827caf),
	.w6(32'hb972535c),
	.w7(32'hb95af925),
	.w8(32'hb98e65fc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c23e33),
	.w1(32'hb9971a7d),
	.w2(32'hb89126de),
	.w3(32'hb9710537),
	.w4(32'hb954f757),
	.w5(32'hb94f6ec6),
	.w6(32'h398d83c2),
	.w7(32'h39715b76),
	.w8(32'h39890d64),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9206ba4),
	.w1(32'hb932af76),
	.w2(32'hb905b755),
	.w3(32'hb90a9bb2),
	.w4(32'hb8f27e1f),
	.w5(32'h36874e10),
	.w6(32'h37cf671e),
	.w7(32'hb7157a44),
	.w8(32'hb905d577),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b481d8),
	.w1(32'hb97eb6cf),
	.w2(32'hb73126db),
	.w3(32'hb8f11924),
	.w4(32'hb7ff241f),
	.w5(32'h390dffa9),
	.w6(32'hb9917169),
	.w7(32'hb780df89),
	.w8(32'h382da51b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39057d30),
	.w1(32'h39687f76),
	.w2(32'h39cdec5e),
	.w3(32'h390ce98f),
	.w4(32'h39a13633),
	.w5(32'h39c61134),
	.w6(32'h39b296d1),
	.w7(32'h39ad7c7e),
	.w8(32'h39dd4074),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb3a97),
	.w1(32'hb9d69c26),
	.w2(32'hb891f7be),
	.w3(32'h3a096d21),
	.w4(32'h39627adb),
	.w5(32'hb7871aba),
	.w6(32'hb8c35039),
	.w7(32'h37b5d112),
	.w8(32'hb818625e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9461010),
	.w1(32'h3820817e),
	.w2(32'h37af4349),
	.w3(32'hb8b8296f),
	.w4(32'h3921c94e),
	.w5(32'h39159b67),
	.w6(32'h383485a0),
	.w7(32'h391cf376),
	.w8(32'h38b6f082),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386bcd8c),
	.w1(32'h35f345e2),
	.w2(32'h398f53d6),
	.w3(32'h39456c80),
	.w4(32'hb85c7865),
	.w5(32'h38121677),
	.w6(32'hb8ba1adb),
	.w7(32'h3826dfea),
	.w8(32'hb86a2ba1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8813431),
	.w1(32'hb99104c6),
	.w2(32'hb9927ed8),
	.w3(32'h3887d202),
	.w4(32'hb8903b7b),
	.w5(32'hb971839d),
	.w6(32'hb96c49f0),
	.w7(32'hb983fd0b),
	.w8(32'hb95d9c28),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b42855),
	.w1(32'hb96369cb),
	.w2(32'hb9263436),
	.w3(32'hb94008ca),
	.w4(32'hb8c0d038),
	.w5(32'hb9300f8e),
	.w6(32'hb9087ba8),
	.w7(32'hb901f37b),
	.w8(32'hb9200076),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c80ef4),
	.w1(32'h378cb1fb),
	.w2(32'h38d4959b),
	.w3(32'hb7d4d6a5),
	.w4(32'h3838540d),
	.w5(32'h39204f71),
	.w6(32'h384b8019),
	.w7(32'h38f6a60c),
	.w8(32'h38c12372),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ff0ca),
	.w1(32'h386a634d),
	.w2(32'h395882d6),
	.w3(32'h39484299),
	.w4(32'h39017679),
	.w5(32'h3983eb03),
	.w6(32'h38e858ec),
	.w7(32'h3977573e),
	.w8(32'h39756c2b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39388377),
	.w1(32'hba4f6e33),
	.w2(32'hb92ec925),
	.w3(32'h398358b6),
	.w4(32'h38c7a27d),
	.w5(32'h3794872a),
	.w6(32'h38d95450),
	.w7(32'h395f1566),
	.w8(32'h38862f5f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e91e79),
	.w1(32'hba2046a5),
	.w2(32'hb9f966bc),
	.w3(32'hb9aa472c),
	.w4(32'hba013303),
	.w5(32'hba126346),
	.w6(32'hb9254f35),
	.w7(32'hb9775831),
	.w8(32'hba1ffd4c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df9a2e),
	.w1(32'h39740e80),
	.w2(32'h39975af0),
	.w3(32'hb9b5bd7a),
	.w4(32'h39a5af5a),
	.w5(32'h39929b14),
	.w6(32'h3926efad),
	.w7(32'h39a4294f),
	.w8(32'h39a406e3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964275a),
	.w1(32'hb839c1d3),
	.w2(32'hb9519d36),
	.w3(32'h396845c2),
	.w4(32'h3983a58f),
	.w5(32'h3918fa28),
	.w6(32'hb788563c),
	.w7(32'h38933fcd),
	.w8(32'h38710ca0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce96ba),
	.w1(32'h36f3d1c6),
	.w2(32'h396c99dd),
	.w3(32'h3929690e),
	.w4(32'hb8500cbc),
	.w5(32'hb867cb23),
	.w6(32'hb94e88ef),
	.w7(32'hb909c512),
	.w8(32'hb9672415),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38596aa1),
	.w1(32'h3714e758),
	.w2(32'h38be78ea),
	.w3(32'hb8de423c),
	.w4(32'h3820e1ce),
	.w5(32'h39260bc1),
	.w6(32'h37f29c86),
	.w7(32'h391265fd),
	.w8(32'h39058b77),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39562b9b),
	.w1(32'hb9214467),
	.w2(32'hb9aad84f),
	.w3(32'h398a16bd),
	.w4(32'hb81e9d53),
	.w5(32'hb6fbfc8f),
	.w6(32'hb9066832),
	.w7(32'hb7d67aa7),
	.w8(32'hb7fd654f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e0049),
	.w1(32'hb9bd05cc),
	.w2(32'hb8fb5d65),
	.w3(32'h389dc72b),
	.w4(32'hb9c08eed),
	.w5(32'hb8cd5585),
	.w6(32'hb9549dad),
	.w7(32'h37a6d67f),
	.w8(32'h38b0c191),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986a1e3),
	.w1(32'hb6c4eb4a),
	.w2(32'h3528753b),
	.w3(32'hb8f6a369),
	.w4(32'h37cf71e5),
	.w5(32'hb82aaa8d),
	.w6(32'hb704ba97),
	.w7(32'h38d1fff1),
	.w8(32'hb9161469),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897d2b8),
	.w1(32'h387ddbeb),
	.w2(32'h390cfa43),
	.w3(32'hb8bff3cd),
	.w4(32'h38dd9ef7),
	.w5(32'h394e11f2),
	.w6(32'h388b737d),
	.w7(32'h391b99e2),
	.w8(32'h3932bd48),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39005b37),
	.w1(32'h387c3749),
	.w2(32'h39222cf3),
	.w3(32'h394d08b3),
	.w4(32'h38a15d48),
	.w5(32'h392c542b),
	.w6(32'h37b69aa5),
	.w7(32'h391b7468),
	.w8(32'h39197a26),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f21bfb),
	.w1(32'hb8ca4883),
	.w2(32'h3826932d),
	.w3(32'h391ee9c8),
	.w4(32'hb901cbbf),
	.w5(32'hb821f57a),
	.w6(32'hb8857829),
	.w7(32'hb7ef55ab),
	.w8(32'hb926a803),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fcf5aa),
	.w1(32'hb793e002),
	.w2(32'h391e6618),
	.w3(32'h38b28e96),
	.w4(32'h3847df75),
	.w5(32'h39989920),
	.w6(32'hb95470de),
	.w7(32'h39251352),
	.w8(32'hb921a019),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d78250),
	.w1(32'hb9853f7b),
	.w2(32'hb9ba44b4),
	.w3(32'hb8100d53),
	.w4(32'hb9423fea),
	.w5(32'hb921bf6f),
	.w6(32'hb954fda4),
	.w7(32'hb97784fc),
	.w8(32'hb9606d0b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1a9a3),
	.w1(32'h382fee87),
	.w2(32'h390be16d),
	.w3(32'hb9215a22),
	.w4(32'h38e747eb),
	.w5(32'h394ea4f7),
	.w6(32'h3733f70b),
	.w7(32'h391959d0),
	.w8(32'h3958c7fc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c5592),
	.w1(32'hb910b0de),
	.w2(32'hb972ea05),
	.w3(32'h390c2626),
	.w4(32'h391d226f),
	.w5(32'h388950ab),
	.w6(32'h38a7d688),
	.w7(32'hb6afb104),
	.w8(32'hb81b64f1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b2c9d),
	.w1(32'h3907f229),
	.w2(32'h36a23acf),
	.w3(32'h392f1967),
	.w4(32'h39b29bbc),
	.w5(32'h37cc1d47),
	.w6(32'h3971e2e3),
	.w7(32'h39a5fab7),
	.w8(32'h391f2e5f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932cfa2),
	.w1(32'h39acf353),
	.w2(32'h397e8e49),
	.w3(32'h38cf8f77),
	.w4(32'h39ca7094),
	.w5(32'h39a39f96),
	.w6(32'h39a011cd),
	.w7(32'h39f3cc4c),
	.w8(32'h39d84efd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982d95c),
	.w1(32'h366f04cb),
	.w2(32'hb7c12043),
	.w3(32'h39599f5f),
	.w4(32'h3835a805),
	.w5(32'h38120e69),
	.w6(32'h37b760f8),
	.w7(32'hb5db18a9),
	.w8(32'hb53115ee),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb806dc7f),
	.w1(32'hb93210e0),
	.w2(32'hb8df1ebe),
	.w3(32'hb6e4d5db),
	.w4(32'hb8fd7e5e),
	.w5(32'hb83257d9),
	.w6(32'hb92a2ef5),
	.w7(32'hb801b2c0),
	.w8(32'hb9023189),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8efed92),
	.w1(32'hb828036a),
	.w2(32'hb8ace7e7),
	.w3(32'hb907e81d),
	.w4(32'h3865140c),
	.w5(32'h37e2e682),
	.w6(32'hb8c33b9e),
	.w7(32'hb8f8630f),
	.w8(32'hb9246376),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915b961),
	.w1(32'hb7f2150b),
	.w2(32'h3899ab7f),
	.w3(32'h38054bf6),
	.w4(32'h37008fff),
	.w5(32'h38977779),
	.w6(32'hb7b8f78f),
	.w7(32'h38c5864a),
	.w8(32'h38499026),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38886386),
	.w1(32'hb85f6bab),
	.w2(32'hb9c5d5e2),
	.w3(32'h37fe317a),
	.w4(32'h391b0327),
	.w5(32'hb96e996b),
	.w6(32'hb8b21408),
	.w7(32'hb990d769),
	.w8(32'hb9c10eab),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a52cbc),
	.w1(32'h3724ed0c),
	.w2(32'hb755440f),
	.w3(32'hb91f1eda),
	.w4(32'h39d7a617),
	.w5(32'h39073563),
	.w6(32'h39902de9),
	.w7(32'h393d4aa9),
	.w8(32'h38a9a34f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88446c6),
	.w1(32'hb98ba484),
	.w2(32'hb92a08ed),
	.w3(32'h3887fba8),
	.w4(32'h39292408),
	.w5(32'h37ec490e),
	.w6(32'hb924ac43),
	.w7(32'hb9048188),
	.w8(32'hb97d8af1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5f77a),
	.w1(32'hb991f969),
	.w2(32'hb91296c9),
	.w3(32'hb8e2ea1b),
	.w4(32'hb6b5455d),
	.w5(32'hb914e2c2),
	.w6(32'h3962df72),
	.w7(32'hb772687c),
	.w8(32'hb9874878),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e72cfb),
	.w1(32'hb9bce09a),
	.w2(32'hb949bc6e),
	.w3(32'hb96b07a0),
	.w4(32'hb999fc23),
	.w5(32'hb91487f7),
	.w6(32'hb99cc643),
	.w7(32'hb939e0a2),
	.w8(32'hb953293f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9536e),
	.w1(32'h3851aa69),
	.w2(32'h392bd3d8),
	.w3(32'hb7ce945a),
	.w4(32'h384e7ec9),
	.w5(32'h392f1edc),
	.w6(32'h37c51453),
	.w7(32'h3914a494),
	.w8(32'h3907cc72),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb787c),
	.w1(32'h394613a5),
	.w2(32'h398ce9be),
	.w3(32'h38e4f218),
	.w4(32'h39751810),
	.w5(32'h3997504e),
	.w6(32'h39363bf7),
	.w7(32'h3982a5e6),
	.w8(32'h39b917ce),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3783f),
	.w1(32'h38f42b61),
	.w2(32'h387c00cf),
	.w3(32'h39b007c8),
	.w4(32'h38f35d60),
	.w5(32'h3684c0cd),
	.w6(32'h3904fa31),
	.w7(32'h3820dbc1),
	.w8(32'h388e46f3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8575f6a),
	.w1(32'h3660f660),
	.w2(32'hb95886f9),
	.w3(32'hb8c9a23a),
	.w4(32'h38bd54d5),
	.w5(32'h39a16a5b),
	.w6(32'h388a04dc),
	.w7(32'h394bfb1e),
	.w8(32'h35c195ab),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39280f34),
	.w1(32'h39c081d6),
	.w2(32'h398b25e2),
	.w3(32'h3a3d5004),
	.w4(32'h3a05fa2f),
	.w5(32'h39f66dae),
	.w6(32'h39fb78a7),
	.w7(32'h39f945b7),
	.w8(32'h39eb11c6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f5155),
	.w1(32'hb7387cb1),
	.w2(32'hb9226c90),
	.w3(32'h39b29776),
	.w4(32'h396c7b30),
	.w5(32'hb79f0309),
	.w6(32'h3753b647),
	.w7(32'hb9971eb7),
	.w8(32'hb93909b1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5cdb8),
	.w1(32'hb9630fe1),
	.w2(32'hb919d60e),
	.w3(32'hb8d48247),
	.w4(32'hb9023521),
	.w5(32'hb905a980),
	.w6(32'hb908a758),
	.w7(32'hb8bf10ee),
	.w8(32'hb8bd867e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9067ffd),
	.w1(32'hb8dd8b7f),
	.w2(32'hb94cac59),
	.w3(32'hb93edffb),
	.w4(32'hb7c96ecd),
	.w5(32'hb87e03c7),
	.w6(32'hb8092804),
	.w7(32'hb94f9f90),
	.w8(32'hb907c1f3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94aa57b),
	.w1(32'hb8686385),
	.w2(32'hb8ade5fb),
	.w3(32'hb88eee9d),
	.w4(32'h38bd60ac),
	.w5(32'h38f75b5b),
	.w6(32'h38d2ee0b),
	.w7(32'h38635168),
	.w8(32'hb8ae410f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890e5ee),
	.w1(32'h390e07c7),
	.w2(32'hb8da848a),
	.w3(32'hb6e8f9ff),
	.w4(32'h38e0f6be),
	.w5(32'hb73f77f6),
	.w6(32'hb8f789e6),
	.w7(32'hb9692d0f),
	.w8(32'h38836677),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d45e08),
	.w1(32'hb793ae4b),
	.w2(32'hb7493efb),
	.w3(32'hb878223a),
	.w4(32'h38fe2084),
	.w5(32'h38bec642),
	.w6(32'h3804a867),
	.w7(32'h38ce741c),
	.w8(32'h3922daef),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38549522),
	.w1(32'h3912fd0d),
	.w2(32'h3970d593),
	.w3(32'h38012659),
	.w4(32'h3925868a),
	.w5(32'h3968cbdd),
	.w6(32'h38f941a0),
	.w7(32'h395bdf40),
	.w8(32'h398c243a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922f0cf),
	.w1(32'hb90d186b),
	.w2(32'hb91361b9),
	.w3(32'h392af424),
	.w4(32'hb8a649d3),
	.w5(32'hb84f7b73),
	.w6(32'hb91723c8),
	.w7(32'hb899f9d1),
	.w8(32'hb772766f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9166c84),
	.w1(32'h391fb50c),
	.w2(32'h395a9a2d),
	.w3(32'hb85c4b84),
	.w4(32'h39c2bc6a),
	.w5(32'h39c55a6e),
	.w6(32'h392770e3),
	.w7(32'h399cb54d),
	.w8(32'h399f47ee),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a85e1f),
	.w1(32'hb7b91c14),
	.w2(32'h384baf15),
	.w3(32'h39c36ec3),
	.w4(32'hb98186c6),
	.w5(32'hb81beeef),
	.w6(32'h386ca8f8),
	.w7(32'h38d397f8),
	.w8(32'h387df0f8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcbc76),
	.w1(32'hb8d937be),
	.w2(32'hb992efef),
	.w3(32'h39162770),
	.w4(32'h379c5803),
	.w5(32'hb929d760),
	.w6(32'hb7282238),
	.w7(32'hb94877ed),
	.w8(32'hb933e8bd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9597b11),
	.w1(32'hb93d17f3),
	.w2(32'hb8c569a4),
	.w3(32'hb908cc3e),
	.w4(32'hb8bb6008),
	.w5(32'hb9057a36),
	.w6(32'hb7b3f1cb),
	.w7(32'hb79a37b7),
	.w8(32'h3858b50b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d7dff),
	.w1(32'h37bca5c2),
	.w2(32'h38d54a48),
	.w3(32'hb89cf75c),
	.w4(32'h3911e499),
	.w5(32'h3969d3ea),
	.w6(32'hb8cc240a),
	.w7(32'hb88ada06),
	.w8(32'hb800f3e0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3893d489),
	.w1(32'hb705d2d6),
	.w2(32'hb8468f00),
	.w3(32'hb7063cfc),
	.w4(32'h3952bbfb),
	.w5(32'hb73342ec),
	.w6(32'h37ce1b06),
	.w7(32'h38515259),
	.w8(32'hb8887f7e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7eb14),
	.w1(32'hb9349a34),
	.w2(32'h3858528b),
	.w3(32'hb7750a98),
	.w4(32'hb8fa5dd2),
	.w5(32'h385d3fa7),
	.w6(32'hb9502ba6),
	.w7(32'h38c5593a),
	.w8(32'hb88016ce),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f893dc),
	.w1(32'h38beac52),
	.w2(32'h388e9f7d),
	.w3(32'hb955624a),
	.w4(32'h3964d9b2),
	.w5(32'h397b4c1d),
	.w6(32'h382c542f),
	.w7(32'h39453967),
	.w8(32'h394389c0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397be651),
	.w1(32'h399647d0),
	.w2(32'h3911a0fd),
	.w3(32'h39648443),
	.w4(32'h3986ac9c),
	.w5(32'h38cdc32b),
	.w6(32'hb85fa84e),
	.w7(32'hb863ea0c),
	.w8(32'h3896d7bf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39544471),
	.w1(32'hb8753531),
	.w2(32'hb8909eca),
	.w3(32'h388b647b),
	.w4(32'h384e9835),
	.w5(32'hb762bd67),
	.w6(32'hb7e9bb73),
	.w7(32'hb80813bd),
	.w8(32'hb82c65b4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e3eaa2),
	.w1(32'h390c9724),
	.w2(32'h396254c6),
	.w3(32'hb890186c),
	.w4(32'h39451bb3),
	.w5(32'h39688124),
	.w6(32'h39013a6e),
	.w7(32'h391e8813),
	.w8(32'h39796d86),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964e2d0),
	.w1(32'h38e79f54),
	.w2(32'h3937f1db),
	.w3(32'h394dd893),
	.w4(32'h3908ed00),
	.w5(32'h392e18c4),
	.w6(32'h38dfc362),
	.w7(32'h3921d38e),
	.w8(32'h396d592b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918174d),
	.w1(32'h382ce15c),
	.w2(32'h392cd2e2),
	.w3(32'h390d6e48),
	.w4(32'h38f1d8ab),
	.w5(32'h3973fb53),
	.w6(32'hb79fad83),
	.w7(32'h39313a0d),
	.w8(32'h3951957e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39280495),
	.w1(32'h38104e2a),
	.w2(32'h3791a903),
	.w3(32'h3959c114),
	.w4(32'h392e6dce),
	.w5(32'h39341810),
	.w6(32'h389224e5),
	.w7(32'h38f5f5b7),
	.w8(32'h3942a599),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382b79bd),
	.w1(32'h38a9ab28),
	.w2(32'hb7b1f49d),
	.w3(32'h399a76a4),
	.w4(32'h39a695bc),
	.w5(32'h391f1ef7),
	.w6(32'h39be7d6a),
	.w7(32'hb81f22a5),
	.w8(32'hb9bdc031),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d9b4e),
	.w1(32'h3904a52e),
	.w2(32'h3981940d),
	.w3(32'h38bb52a4),
	.w4(32'h38e6a20b),
	.w5(32'h3973c9d9),
	.w6(32'hb8297598),
	.w7(32'h38e87646),
	.w8(32'h3954f2a9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3752de69),
	.w1(32'hb893e56c),
	.w2(32'h387d8a1b),
	.w3(32'h3923878c),
	.w4(32'h387bad61),
	.w5(32'h3904986b),
	.w6(32'hb8180485),
	.w7(32'h38b8ae7b),
	.w8(32'hb809001a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf9f11),
	.w1(32'hb92a213b),
	.w2(32'h387a08b3),
	.w3(32'h390be380),
	.w4(32'hb8bf6bcb),
	.w5(32'h3623c722),
	.w6(32'hb94a36a6),
	.w7(32'hb8b62525),
	.w8(32'hb96f0e21),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eddf0d),
	.w1(32'hb885081a),
	.w2(32'h38e226c5),
	.w3(32'hb96ee162),
	.w4(32'h3795da68),
	.w5(32'h3919d01e),
	.w6(32'h38bb58ec),
	.w7(32'h393b2b5c),
	.w8(32'h394520e7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b1cb04),
	.w1(32'hb8e63f7b),
	.w2(32'hb739f5eb),
	.w3(32'h39573aff),
	.w4(32'hb80772cf),
	.w5(32'h38ae1b9f),
	.w6(32'hb87b285b),
	.w7(32'h391866f8),
	.w8(32'h380f734e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c78f8),
	.w1(32'hb8023ebd),
	.w2(32'hb6eca850),
	.w3(32'hb8cc625e),
	.w4(32'h3903c036),
	.w5(32'h3915e8db),
	.w6(32'h384a52cb),
	.w7(32'h38a2b81f),
	.w8(32'hb812e8f4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38162fc8),
	.w1(32'hb712f7db),
	.w2(32'hb880a547),
	.w3(32'h38ee6f56),
	.w4(32'h3721b8d9),
	.w5(32'h37e5f424),
	.w6(32'h3814a893),
	.w7(32'h37a76ddd),
	.w8(32'h3822fb46),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b35f42),
	.w1(32'hb8a32bbb),
	.w2(32'hb796a1dd),
	.w3(32'h37cb5c95),
	.w4(32'h381fef84),
	.w5(32'h37a1760d),
	.w6(32'h37f73953),
	.w7(32'h38998c5e),
	.w8(32'h38d0f562),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384eb5c6),
	.w1(32'h3696bed1),
	.w2(32'hb8a4dfa6),
	.w3(32'h35d76329),
	.w4(32'hb90e787d),
	.w5(32'hb8715ee4),
	.w6(32'hb8040652),
	.w7(32'h38dd4b5d),
	.w8(32'h38a9c826),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9510447),
	.w1(32'h3956001e),
	.w2(32'h394cbd82),
	.w3(32'hb8d302df),
	.w4(32'h39a588e2),
	.w5(32'h39a22274),
	.w6(32'h3955c721),
	.w7(32'h391bd983),
	.w8(32'h38985d2f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987e543),
	.w1(32'h398c9e8d),
	.w2(32'h395addbd),
	.w3(32'h392bc436),
	.w4(32'h3843f6fd),
	.w5(32'h388ec0b1),
	.w6(32'h398cd39b),
	.w7(32'h39891486),
	.w8(32'h391a4f0a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b3e8c),
	.w1(32'hb702a111),
	.w2(32'h388deca3),
	.w3(32'h38a2eeb8),
	.w4(32'h384a5352),
	.w5(32'h39101d68),
	.w6(32'h37a3da57),
	.w7(32'h38fab2e5),
	.w8(32'h39170dd6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371fd1f3),
	.w1(32'hb927be61),
	.w2(32'hb9132589),
	.w3(32'h39309e6d),
	.w4(32'hb811afa4),
	.w5(32'hb91d30ae),
	.w6(32'h37bd48ce),
	.w7(32'hb7cad367),
	.w8(32'hb921b58b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932d108),
	.w1(32'h393832cc),
	.w2(32'h395cc076),
	.w3(32'hb9187388),
	.w4(32'h39a0ae89),
	.w5(32'h396e2e19),
	.w6(32'hb84636dc),
	.w7(32'h3937d4db),
	.w8(32'h389ae749),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba0773),
	.w1(32'hb6bbd45f),
	.w2(32'h389c3278),
	.w3(32'h392a273d),
	.w4(32'h384441da),
	.w5(32'h3907bbb9),
	.w6(32'h388e9f08),
	.w7(32'h39510feb),
	.w8(32'h3964546e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb423c798),
	.w1(32'hb92f4209),
	.w2(32'hb9901762),
	.w3(32'h388110c4),
	.w4(32'h35cc7836),
	.w5(32'hb9344a38),
	.w6(32'hb801b8ba),
	.w7(32'hb7cb7d98),
	.w8(32'hb96d3281),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a2b5a),
	.w1(32'hb6fa425d),
	.w2(32'hb8245245),
	.w3(32'hb9009ab6),
	.w4(32'h3906f83e),
	.w5(32'h37f6680b),
	.w6(32'h382118d6),
	.w7(32'h38e5fca6),
	.w8(32'h38c9be6d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382982e7),
	.w1(32'hb8d7e636),
	.w2(32'hb7b63139),
	.w3(32'h389927a1),
	.w4(32'hb8937a2b),
	.w5(32'h365eb748),
	.w6(32'hb793c0d0),
	.w7(32'h39005a43),
	.w8(32'hb918ea3a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b79330),
	.w1(32'hb895ca63),
	.w2(32'hb8d70cb2),
	.w3(32'hb85c0afc),
	.w4(32'hb913d97e),
	.w5(32'hb93ca24d),
	.w6(32'hb6f39e81),
	.w7(32'h37c54f5f),
	.w8(32'h36435f79),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2c8f7),
	.w1(32'h393f3e7c),
	.w2(32'h39a7ee19),
	.w3(32'hb9ab52ba),
	.w4(32'h38c9b93c),
	.w5(32'h37d97bf1),
	.w6(32'h388d140f),
	.w7(32'h37148992),
	.w8(32'h387f775d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5fcec),
	.w1(32'hb94dc458),
	.w2(32'hb91a2c7b),
	.w3(32'hb830cbbc),
	.w4(32'hb92d0502),
	.w5(32'hb91463eb),
	.w6(32'hb992b4a1),
	.w7(32'hb91ff9c6),
	.w8(32'hb99f7e3a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5b94e),
	.w1(32'hb969b8a1),
	.w2(32'hb9bb72af),
	.w3(32'hb9c9e46a),
	.w4(32'hb9864c42),
	.w5(32'hb9b09741),
	.w6(32'hb99d6fc0),
	.w7(32'hb90b726a),
	.w8(32'hb9365c5e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89830c5),
	.w1(32'hb7d06ccb),
	.w2(32'hb744bc23),
	.w3(32'h36cda35d),
	.w4(32'h396db088),
	.w5(32'h39935e83),
	.w6(32'h3957f406),
	.w7(32'h3999544e),
	.w8(32'h398e995c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e7a72),
	.w1(32'h393d7572),
	.w2(32'h37b49a1a),
	.w3(32'h392ebde7),
	.w4(32'h3a1e21ae),
	.w5(32'h39df213e),
	.w6(32'h38ea3233),
	.w7(32'h393d7633),
	.w8(32'h392f544c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d66d8c),
	.w1(32'h398b6ed2),
	.w2(32'hb95b7961),
	.w3(32'h3a256d80),
	.w4(32'h3a20474c),
	.w5(32'h390abeaa),
	.w6(32'h3955a401),
	.w7(32'h3914ef02),
	.w8(32'hb92a530a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfbd4d),
	.w1(32'hb6a71543),
	.w2(32'h399de07b),
	.w3(32'hb9c45e81),
	.w4(32'h39916306),
	.w5(32'h39df029b),
	.w6(32'hb8ca2355),
	.w7(32'hb9a50dda),
	.w8(32'hb9fa1757),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d353b),
	.w1(32'h397be4a4),
	.w2(32'h39bef876),
	.w3(32'h3870820f),
	.w4(32'h39a35ded),
	.w5(32'h39c6708a),
	.w6(32'h39fc6bd7),
	.w7(32'h39bdd1b9),
	.w8(32'h39b4778c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc7bc9),
	.w1(32'h38f300cc),
	.w2(32'h394a9dd3),
	.w3(32'h39f59f8b),
	.w4(32'h39725d6b),
	.w5(32'h39807d51),
	.w6(32'h391b11b3),
	.w7(32'h393ab39e),
	.w8(32'h398b77a8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39875269),
	.w1(32'h39147f56),
	.w2(32'h390c295e),
	.w3(32'h39b69b2a),
	.w4(32'h39b3d747),
	.w5(32'h39326500),
	.w6(32'h39156407),
	.w7(32'h39952a91),
	.w8(32'h390a94fb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a623a5),
	.w1(32'hb7e19f3d),
	.w2(32'hb615bc32),
	.w3(32'h398802ed),
	.w4(32'hb759beb8),
	.w5(32'h39491f82),
	.w6(32'hb9033606),
	.w7(32'h3825cec0),
	.w8(32'h39345ff8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386654bc),
	.w1(32'hb9556818),
	.w2(32'hb8eb5a09),
	.w3(32'h39346904),
	.w4(32'hb941b37e),
	.w5(32'hb95074b8),
	.w6(32'h3852b156),
	.w7(32'h38abb516),
	.w8(32'h37b4786e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937d98f),
	.w1(32'h38d36f60),
	.w2(32'h3941781c),
	.w3(32'hb93f0c77),
	.w4(32'h390b1cea),
	.w5(32'h3987fa38),
	.w6(32'h38e8758d),
	.w7(32'h39726240),
	.w8(32'h39792966),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d4602),
	.w1(32'h38e636ea),
	.w2(32'h394d5dcf),
	.w3(32'h39181bd3),
	.w4(32'h391b0fea),
	.w5(32'h391581ee),
	.w6(32'h384f0ce4),
	.w7(32'h38db68ff),
	.w8(32'h38e8e408),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ba514),
	.w1(32'h3912f7c4),
	.w2(32'h38d2f7d5),
	.w3(32'h398145f9),
	.w4(32'h399218e6),
	.w5(32'h380af6bc),
	.w6(32'h398e5107),
	.w7(32'h3977c5c9),
	.w8(32'h38c940bb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387050e3),
	.w1(32'h37aceee5),
	.w2(32'h37cc3f59),
	.w3(32'hb7c2beb4),
	.w4(32'h3828c137),
	.w5(32'h38854e81),
	.w6(32'h38853a22),
	.w7(32'h3903fd2d),
	.w8(32'h38af166c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d9953a),
	.w1(32'h3876242f),
	.w2(32'hb99556d3),
	.w3(32'h3904705f),
	.w4(32'hb8184166),
	.w5(32'hb9238b3b),
	.w6(32'h397524e4),
	.w7(32'h3919feea),
	.w8(32'h36db945b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a00614),
	.w1(32'hb8b9ce8e),
	.w2(32'hb90aa498),
	.w3(32'h389a9ded),
	.w4(32'h380503b3),
	.w5(32'h37c144e2),
	.w6(32'h382df413),
	.w7(32'h3826597c),
	.w8(32'hb7c25e99),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89940b8),
	.w1(32'h388cf86c),
	.w2(32'h3901f548),
	.w3(32'h38fe03ef),
	.w4(32'h37d01936),
	.w5(32'h37a7de69),
	.w6(32'h373538ed),
	.w7(32'h38737a73),
	.w8(32'hb854a524),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885e1ef),
	.w1(32'h38f8530f),
	.w2(32'h393f2211),
	.w3(32'h37838f24),
	.w4(32'h398a5bc9),
	.w5(32'h399b094c),
	.w6(32'h395bc531),
	.w7(32'h399deaee),
	.w8(32'h39978b10),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39670841),
	.w1(32'h394bd624),
	.w2(32'h3990438e),
	.w3(32'h39bbe7ae),
	.w4(32'h398a4903),
	.w5(32'h39a33d0a),
	.w6(32'h395eac55),
	.w7(32'h3971e123),
	.w8(32'h39b3181d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0398a),
	.w1(32'h394ad9fb),
	.w2(32'h398aec66),
	.w3(32'h39b673ed),
	.w4(32'h3936e532),
	.w5(32'h39583cba),
	.w6(32'h3945b670),
	.w7(32'h39779eaf),
	.w8(32'h398d70f2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f4343),
	.w1(32'h394ce2d6),
	.w2(32'h398cc0e4),
	.w3(32'h396ed001),
	.w4(32'h39386e2e),
	.w5(32'h39687f21),
	.w6(32'h393f0c49),
	.w7(32'h397039d2),
	.w8(32'h3996164b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f7b6f),
	.w1(32'hb99fad1a),
	.w2(32'h36e9778a),
	.w3(32'h3986c938),
	.w4(32'h3910bedb),
	.w5(32'h392d5ecc),
	.w6(32'hb9341b57),
	.w7(32'hb89d86e6),
	.w8(32'hb90d46d1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aacec6),
	.w1(32'hb9486678),
	.w2(32'hb96450bb),
	.w3(32'hb902cb46),
	.w4(32'hb81b319d),
	.w5(32'hb8eea319),
	.w6(32'hb98ccc21),
	.w7(32'hb98b91d2),
	.w8(32'hb917185a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810aa3),
	.w1(32'h398870b8),
	.w2(32'h391d2950),
	.w3(32'hb928964c),
	.w4(32'h3980140b),
	.w5(32'h394d617c),
	.w6(32'h3994b73b),
	.w7(32'h3975f5e6),
	.w8(32'h399949ed),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3832931b),
	.w1(32'h38ff9dd6),
	.w2(32'h38bd601b),
	.w3(32'h39754fba),
	.w4(32'h39307fba),
	.w5(32'h394d2b56),
	.w6(32'h393681b7),
	.w7(32'h397475d2),
	.w8(32'h396b7b13),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385942e7),
	.w1(32'h38cb197d),
	.w2(32'h39abd5e3),
	.w3(32'h38a966d7),
	.w4(32'h3982dfe9),
	.w5(32'h39e5c9e1),
	.w6(32'h39016850),
	.w7(32'h399e5613),
	.w8(32'h39c85dd4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998f4ae),
	.w1(32'hb9b22cba),
	.w2(32'hb7d09e9f),
	.w3(32'h39949bff),
	.w4(32'h3889cd07),
	.w5(32'h37fcc1e6),
	.w6(32'hb881006a),
	.w7(32'hb887c256),
	.w8(32'hb91c9ff9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394488f5),
	.w1(32'h39b80cd1),
	.w2(32'h39a766f9),
	.w3(32'hb92806fa),
	.w4(32'h39c48cfc),
	.w5(32'h39b51cb2),
	.w6(32'h39db905e),
	.w7(32'h39b835f0),
	.w8(32'h39e19852),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e99ae),
	.w1(32'hb6754ebc),
	.w2(32'h390e640b),
	.w3(32'h39958d3b),
	.w4(32'h386e8567),
	.w5(32'h397c0911),
	.w6(32'h382f84fb),
	.w7(32'h393faea5),
	.w8(32'h395d150d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390fcae5),
	.w1(32'h374fe780),
	.w2(32'h3828973e),
	.w3(32'h39869ab2),
	.w4(32'hb7d568a3),
	.w5(32'hb6f3d05b),
	.w6(32'h38427de4),
	.w7(32'h371a54ff),
	.w8(32'hb7ac5086),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94aed2e),
	.w1(32'hb8d391f6),
	.w2(32'hb77e44f9),
	.w3(32'hb9123a3d),
	.w4(32'hb7c4cdc2),
	.w5(32'h379636df),
	.w6(32'hb8ee5bbd),
	.w7(32'hb77f3c86),
	.w8(32'hb87e043b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb775abab),
	.w1(32'h3853efa0),
	.w2(32'h37a0d446),
	.w3(32'h37384867),
	.w4(32'h3869b0f8),
	.w5(32'hb87f60e0),
	.w6(32'hb69e577c),
	.w7(32'h37cee1ba),
	.w8(32'hb87e8308),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3688a8a4),
	.w1(32'hb628ebe6),
	.w2(32'hb6c14270),
	.w3(32'hb7586270),
	.w4(32'hb5d08745),
	.w5(32'hb626cd93),
	.w6(32'h35e268c1),
	.w7(32'h36322eb7),
	.w8(32'hb7527d3e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73e935a),
	.w1(32'h372ec1c3),
	.w2(32'hb5331801),
	.w3(32'hb7cd7863),
	.w4(32'h36ed9a9c),
	.w5(32'hb73adfd9),
	.w6(32'hb63f3809),
	.w7(32'h378a3f9f),
	.w8(32'h3711b0f2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64521df),
	.w1(32'h3852aa91),
	.w2(32'h38094f5c),
	.w3(32'h388c806d),
	.w4(32'h38baaa7c),
	.w5(32'h37f5db20),
	.w6(32'h38806232),
	.w7(32'h388566bc),
	.w8(32'h380a6b6c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fbb9a9),
	.w1(32'hb78198a4),
	.w2(32'hb7a264d6),
	.w3(32'hb7fee699),
	.w4(32'hb79708d4),
	.w5(32'hb81a4e10),
	.w6(32'hb793e715),
	.w7(32'hb663fea5),
	.w8(32'hb769616b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3eaa7),
	.w1(32'h39200ff8),
	.w2(32'h38c44053),
	.w3(32'h38d40d69),
	.w4(32'h391cef57),
	.w5(32'h38a8eea6),
	.w6(32'h391e1983),
	.w7(32'h394f4f80),
	.w8(32'h381ab4e0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949371f),
	.w1(32'hb926c61e),
	.w2(32'hb8d45c2a),
	.w3(32'h3512e743),
	.w4(32'h37409808),
	.w5(32'hb84c8446),
	.w6(32'hb8b06a6b),
	.w7(32'hb8e74ee7),
	.w8(32'hb8da9b58),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c7fc8e),
	.w1(32'hb7192000),
	.w2(32'h36199491),
	.w3(32'h374aba32),
	.w4(32'h3735e1f8),
	.w5(32'hb839b845),
	.w6(32'h38451113),
	.w7(32'h3809f15b),
	.w8(32'hb88c0073),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8325393),
	.w1(32'hb7217b27),
	.w2(32'h38cc1ba7),
	.w3(32'hb90d720e),
	.w4(32'h3839b4b8),
	.w5(32'h391b3f46),
	.w6(32'h384da440),
	.w7(32'h38b0a453),
	.w8(32'h387ef98b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3bb28),
	.w1(32'hb8c5dd84),
	.w2(32'hb8d753ef),
	.w3(32'hb76c2ad3),
	.w4(32'h384d6a79),
	.w5(32'hb80a42ba),
	.w6(32'h3840fbb3),
	.w7(32'hb863628c),
	.w8(32'hb8fb36fb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74ccf8b),
	.w1(32'h37df5521),
	.w2(32'h36c474dd),
	.w3(32'h372acc17),
	.w4(32'h37f95647),
	.w5(32'hb820d98e),
	.w6(32'h3825b8aa),
	.w7(32'h383ed2f4),
	.w8(32'hb8250559),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7269c4d),
	.w1(32'hb7891945),
	.w2(32'hb7670e87),
	.w3(32'hb8105972),
	.w4(32'hb8a4c14b),
	.w5(32'hb8ee82bf),
	.w6(32'h372b073f),
	.w7(32'h3603fbb1),
	.w8(32'hb88027ee),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74f63ea),
	.w1(32'h36f6fec8),
	.w2(32'h36e86ddb),
	.w3(32'h3712eac4),
	.w4(32'h3805ce02),
	.w5(32'h3788c589),
	.w6(32'hb743ba72),
	.w7(32'h379053ed),
	.w8(32'h3746d5c6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d69110),
	.w1(32'hb830c4ce),
	.w2(32'h38333d9f),
	.w3(32'hb8df104f),
	.w4(32'hb7a746f7),
	.w5(32'hb759d225),
	.w6(32'h38c1b3c3),
	.w7(32'h38e452d1),
	.w8(32'hb7f5ecf2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e743c5),
	.w1(32'h38ddf06a),
	.w2(32'h37be971e),
	.w3(32'h38c62d7c),
	.w4(32'h38bbfc49),
	.w5(32'hb794bb3b),
	.w6(32'h38cde822),
	.w7(32'h38b4e4d2),
	.w8(32'hb6db938d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3500e10a),
	.w1(32'h33ad46af),
	.w2(32'h34d607b7),
	.w3(32'h3601712c),
	.w4(32'hb5b78945),
	.w5(32'hb4a4bfd0),
	.w6(32'hb52704cc),
	.w7(32'hb5fc0c5b),
	.w8(32'hb60a1b3b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ad17d8),
	.w1(32'h35eb916b),
	.w2(32'h322bd7ec),
	.w3(32'hb5095e9f),
	.w4(32'h3519ddc7),
	.w5(32'h35393fb3),
	.w6(32'h35a0844b),
	.w7(32'hb489feb7),
	.w8(32'h36924cab),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8fc66),
	.w1(32'h37b64a48),
	.w2(32'hb77f482a),
	.w3(32'h32f60b5e),
	.w4(32'hb79b31cb),
	.w5(32'hb784f49a),
	.w6(32'hb721a11c),
	.w7(32'h36e85a60),
	.w8(32'h381cc67c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ee8aed),
	.w1(32'hb8834618),
	.w2(32'hb8022599),
	.w3(32'h370e9636),
	.w4(32'h3654c39f),
	.w5(32'hb86e1097),
	.w6(32'h38d7d703),
	.w7(32'h38183cae),
	.w8(32'hb902d8af),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fcf4e),
	.w1(32'hb9316e68),
	.w2(32'hb8f97557),
	.w3(32'hb9421dff),
	.w4(32'hb8d8821f),
	.w5(32'hb84dbe11),
	.w6(32'hb997a748),
	.w7(32'hb8f5bd34),
	.w8(32'h3690b7e3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3501e783),
	.w1(32'h3540eda5),
	.w2(32'h358ba3ff),
	.w3(32'h35e7912d),
	.w4(32'h35d82591),
	.w5(32'h3607bfbb),
	.w6(32'h3593f125),
	.w7(32'h350b9e79),
	.w8(32'h35a8c919),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb819da82),
	.w1(32'h3634dcf5),
	.w2(32'h381196e3),
	.w3(32'h370f2d52),
	.w4(32'h383c8b48),
	.w5(32'hb79601d0),
	.w6(32'hb80820f2),
	.w7(32'h369a1778),
	.w8(32'hb7cb4030),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ccd2fc),
	.w1(32'h37386312),
	.w2(32'h37e869f9),
	.w3(32'hb7528842),
	.w4(32'h375cce2e),
	.w5(32'hb82c14c4),
	.w6(32'h353db5fe),
	.w7(32'h3788f527),
	.w8(32'hb8676343),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9899b9d),
	.w1(32'hb97d47b4),
	.w2(32'hb9090786),
	.w3(32'hb986ed18),
	.w4(32'hb922b07a),
	.w5(32'hb87f6bbe),
	.w6(32'h36a6520d),
	.w7(32'hb8295aaa),
	.w8(32'hb9225eba),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a27331),
	.w1(32'h365fb844),
	.w2(32'hb7c31b6e),
	.w3(32'hb625b058),
	.w4(32'h380b9fdb),
	.w5(32'hb754cd10),
	.w6(32'h379c04cf),
	.w7(32'h3706ccca),
	.w8(32'hb800c9b0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4484b),
	.w1(32'h3917f359),
	.w2(32'h38b458f8),
	.w3(32'h38c7500e),
	.w4(32'h3905645b),
	.w5(32'h389c0575),
	.w6(32'h39008185),
	.w7(32'h3914899b),
	.w8(32'h38cca32c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a7d042),
	.w1(32'h3716c98a),
	.w2(32'h378ec85d),
	.w3(32'hb704eac3),
	.w4(32'hb6287e14),
	.w5(32'h372ad066),
	.w6(32'hb6d1fd13),
	.w7(32'hb4e55892),
	.w8(32'h374c8e78),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ecd43),
	.w1(32'hb812c4c3),
	.w2(32'hb884bf01),
	.w3(32'hb8970570),
	.w4(32'hb8893605),
	.w5(32'hb8b8a80c),
	.w6(32'hb6826865),
	.w7(32'hb79bcb77),
	.w8(32'hb89036ee),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39651fd1),
	.w1(32'h39476506),
	.w2(32'h38a2b1e6),
	.w3(32'h3946bcb6),
	.w4(32'h39845bb6),
	.w5(32'h3900aea2),
	.w6(32'h398f2c67),
	.w7(32'h398f9ac5),
	.w8(32'h383c82e5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37918121),
	.w1(32'h37b33bb4),
	.w2(32'h3657c4c6),
	.w3(32'h37c5fbc4),
	.w4(32'h38286054),
	.w5(32'h37c09702),
	.w6(32'h37b8a920),
	.w7(32'h3829a189),
	.w8(32'h37c2c6c3),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb737b3af),
	.w1(32'hb7e96aec),
	.w2(32'hb78e5cf4),
	.w3(32'hb7c24de5),
	.w4(32'h364c0a38),
	.w5(32'h361c6e69),
	.w6(32'hb6bb71dd),
	.w7(32'hb64965ff),
	.w8(32'hb792b3f6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364a1269),
	.w1(32'hb63d52fa),
	.w2(32'hb6d0b7ff),
	.w3(32'hb6c5b5d4),
	.w4(32'hb62f43b8),
	.w5(32'hb7526771),
	.w6(32'h377be01e),
	.w7(32'h36a081eb),
	.w8(32'h34c83c63),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a7881),
	.w1(32'hb68f7ecd),
	.w2(32'h373f69dc),
	.w3(32'hb8ccdfe7),
	.w4(32'hb84f8c84),
	.w5(32'hb8b3c23c),
	.w6(32'hb821d670),
	.w7(32'hb816ddf1),
	.w8(32'hb8fd7704),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37739d45),
	.w1(32'h36630ab6),
	.w2(32'hb649f297),
	.w3(32'h36482d4e),
	.w4(32'hb7436bc2),
	.w5(32'hb4cd2e12),
	.w6(32'hb7165cc6),
	.w7(32'hb64f7b29),
	.w8(32'h361ed233),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869eead),
	.w1(32'hb8028284),
	.w2(32'hb83de004),
	.w3(32'hb80784ba),
	.w4(32'h37a188fd),
	.w5(32'hb7b0fa42),
	.w6(32'hb59522ae),
	.w7(32'h38134022),
	.w8(32'hb7ad6f42),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360c0060),
	.w1(32'hb617b880),
	.w2(32'hb6ca29ef),
	.w3(32'hb39abe58),
	.w4(32'hb64f6ea0),
	.w5(32'hb688d7af),
	.w6(32'h34d4a49a),
	.w7(32'h357043c5),
	.w8(32'hb63f917a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ef221a),
	.w1(32'hb7ed7887),
	.w2(32'h37e1e14c),
	.w3(32'hb87c35dc),
	.w4(32'hb7e50648),
	.w5(32'h38b8008a),
	.w6(32'hb911cca9),
	.w7(32'hb84777ec),
	.w8(32'h38ee81b3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60a877f),
	.w1(32'hb5f52a38),
	.w2(32'h3589f359),
	.w3(32'hb563caad),
	.w4(32'hb4b855ab),
	.w5(32'h361242e1),
	.w6(32'h35aa1f61),
	.w7(32'haf7583cd),
	.w8(32'h3596debe),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71340b7),
	.w1(32'hb6fd491b),
	.w2(32'hb6b87c4f),
	.w3(32'hb62ae157),
	.w4(32'hb5b2979c),
	.w5(32'hb5d0aca6),
	.w6(32'h34eecc0d),
	.w7(32'hb7018bd7),
	.w8(32'hb6c9c9ab),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f3722),
	.w1(32'h38846637),
	.w2(32'h3813d93b),
	.w3(32'h385fda62),
	.w4(32'h37a36afd),
	.w5(32'hb8925fea),
	.w6(32'h38fafbf7),
	.w7(32'h38aab738),
	.w8(32'hb8978275),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927be77),
	.w1(32'hb605be3b),
	.w2(32'h38286380),
	.w3(32'hb810a41e),
	.w4(32'h37e2c834),
	.w5(32'hb6ba9e14),
	.w6(32'hb850726a),
	.w7(32'hb7bf24a8),
	.w8(32'hb90455a8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36835bf9),
	.w1(32'hb7120cf8),
	.w2(32'hb760c44d),
	.w3(32'hb7ac1fb9),
	.w4(32'h35f40d80),
	.w5(32'h3754dd1c),
	.w6(32'hb7c6da40),
	.w7(32'hb7129273),
	.w8(32'h37ce371a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8875d77),
	.w1(32'h34cde99e),
	.w2(32'hb7886ae1),
	.w3(32'hb7128595),
	.w4(32'h37b6e799),
	.w5(32'hb86396ea),
	.w6(32'h36a9060f),
	.w7(32'h3710af64),
	.w8(32'hb8903aae),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783d607),
	.w1(32'h37cdb085),
	.w2(32'h36c26770),
	.w3(32'h381c6b5e),
	.w4(32'h38362803),
	.w5(32'hb76b1960),
	.w6(32'h38225b56),
	.w7(32'h3845bbcc),
	.w8(32'hb668b75d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f812e5),
	.w1(32'hb90d4a64),
	.w2(32'hb898f8c8),
	.w3(32'hb8f05254),
	.w4(32'hb8345650),
	.w5(32'hb7a5c0fb),
	.w6(32'hb90423e7),
	.w7(32'hb70046a0),
	.w8(32'hb8d1b890),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7920189),
	.w1(32'h37104008),
	.w2(32'hb7639ca4),
	.w3(32'hb7afa934),
	.w4(32'h3811e143),
	.w5(32'hb73f3394),
	.w6(32'hb7baf714),
	.w7(32'h38318d26),
	.w8(32'h37244815),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8769454),
	.w1(32'h36baacea),
	.w2(32'h37816a90),
	.w3(32'h38547203),
	.w4(32'h38c3364e),
	.w5(32'h3741cd3a),
	.w6(32'hb83aaeb1),
	.w7(32'hb70eeaab),
	.w8(32'hb80697d5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h339f4e8b),
	.w1(32'hb62976ec),
	.w2(32'h363e7935),
	.w3(32'h362a3cf3),
	.w4(32'hb67253fb),
	.w5(32'h35d2b811),
	.w6(32'hb6755967),
	.w7(32'h3614915c),
	.w8(32'h364e86b0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d3612d),
	.w1(32'hb510a100),
	.w2(32'h37bc954d),
	.w3(32'h380fee58),
	.w4(32'h379e0a38),
	.w5(32'hb82c47b4),
	.w6(32'h38cada9f),
	.w7(32'h386ba335),
	.w8(32'hb85a83ca),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5abc658),
	.w1(32'h357f50a3),
	.w2(32'h360f02a0),
	.w3(32'hb5e2f0d4),
	.w4(32'h34ad5be1),
	.w5(32'h35afe635),
	.w6(32'h3564f6df),
	.w7(32'h3585d73a),
	.w8(32'h35a4d954),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f11767),
	.w1(32'h37cb156f),
	.w2(32'h380a4e52),
	.w3(32'hb778aa3e),
	.w4(32'hb6e055a8),
	.w5(32'h37dc270f),
	.w6(32'hb8118933),
	.w7(32'hb7960497),
	.w8(32'h3746f5a6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb752bbca),
	.w1(32'h375a80f0),
	.w2(32'hb720d2e5),
	.w3(32'hb658e09c),
	.w4(32'hb6f32044),
	.w5(32'hb75e667c),
	.w6(32'h3770aa8f),
	.w7(32'hb4cc2895),
	.w8(32'hb78c0573),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849887e),
	.w1(32'hb84d6d49),
	.w2(32'hb78e91c3),
	.w3(32'hb8a97068),
	.w4(32'hb86da847),
	.w5(32'hb85b5e98),
	.w6(32'hb82049cb),
	.w7(32'h36e83feb),
	.w8(32'hb822161f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a90adf),
	.w1(32'h35b7dad4),
	.w2(32'h35a67083),
	.w3(32'h34841bc3),
	.w4(32'h3616e481),
	.w5(32'h359136be),
	.w6(32'h35627448),
	.w7(32'hb5343198),
	.w8(32'h35a44c3e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e6b624),
	.w1(32'h3456cc82),
	.w2(32'h35eddc37),
	.w3(32'hb5873b59),
	.w4(32'hb642161b),
	.w5(32'hb51fa2b0),
	.w6(32'hb453b7fb),
	.w7(32'hb561e289),
	.w8(32'h3529f454),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b72db5),
	.w1(32'h3542e29a),
	.w2(32'hb788a016),
	.w3(32'hb73217a6),
	.w4(32'h379dfb1c),
	.w5(32'h37a2b4b8),
	.w6(32'h3828f18d),
	.w7(32'h379672fe),
	.w8(32'h37b2cec8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc0d0e),
	.w1(32'hb8bb7e41),
	.w2(32'hb89782ac),
	.w3(32'hb899f8c7),
	.w4(32'hb8874243),
	.w5(32'hb8372625),
	.w6(32'h38cb04a7),
	.w7(32'h38d9803f),
	.w8(32'hb83292f7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37239db1),
	.w1(32'h33fc8f48),
	.w2(32'hb7fa8c9c),
	.w3(32'hb7b6b52a),
	.w4(32'h37f37b0b),
	.w5(32'hb7f2b625),
	.w6(32'h365a5dff),
	.w7(32'h38021595),
	.w8(32'hb84651b2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d8c4ed),
	.w1(32'h36565b2d),
	.w2(32'hb51f0222),
	.w3(32'h379e9c1e),
	.w4(32'h377800ed),
	.w5(32'h36919eb6),
	.w6(32'h37ae18a1),
	.w7(32'h37c04ea4),
	.w8(32'h374ce534),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba445277),
	.w1(32'hb9e3be7a),
	.w2(32'hb94b74d3),
	.w3(32'hba2947e3),
	.w4(32'hb98fa53d),
	.w5(32'hb8bff28b),
	.w6(32'hba097387),
	.w7(32'hb98c4c73),
	.w8(32'hb879f1ee),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39153829),
	.w1(32'h39a17dca),
	.w2(32'h386eead1),
	.w3(32'h38553519),
	.w4(32'h3955f360),
	.w5(32'h381efc55),
	.w6(32'h39a7fa73),
	.w7(32'h39828da6),
	.w8(32'hb8874ad9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3656f896),
	.w1(32'hb66699af),
	.w2(32'hb7a25636),
	.w3(32'hb6f39d66),
	.w4(32'hb6d4cdd6),
	.w5(32'hb725cf1c),
	.w6(32'hb744628a),
	.w7(32'hb785af71),
	.w8(32'hb6eb288c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b9e0b2),
	.w1(32'h3606c006),
	.w2(32'h35b6ee0a),
	.w3(32'hb5911787),
	.w4(32'hb5a3ea7d),
	.w5(32'h348fd80c),
	.w6(32'hb17b5977),
	.w7(32'h35e2ff8e),
	.w8(32'hb5c80681),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351b4501),
	.w1(32'h36236fa9),
	.w2(32'h3676e9c9),
	.w3(32'hb5075ac8),
	.w4(32'h35a1229a),
	.w5(32'h361dcdb7),
	.w6(32'h34791c82),
	.w7(32'h36220f3a),
	.w8(32'h36639072),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4fde373),
	.w1(32'hb38cd8f1),
	.w2(32'h35cc9596),
	.w3(32'h34693c9a),
	.w4(32'h34b6b0c8),
	.w5(32'h3583ec8e),
	.w6(32'h35ddc104),
	.w7(32'h35a4ef24),
	.w8(32'h358c966f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3627ada7),
	.w1(32'hb7435afb),
	.w2(32'hb796a1c4),
	.w3(32'h36c709bf),
	.w4(32'hb80c0038),
	.w5(32'hb7440c2c),
	.w6(32'h383b1de7),
	.w7(32'h370e1126),
	.w8(32'hb7f5b5a3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be3775),
	.w1(32'h38b32b62),
	.w2(32'h37b35588),
	.w3(32'hb7b9ce09),
	.w4(32'h37d93f8f),
	.w5(32'h38290b17),
	.w6(32'h38fda8fc),
	.w7(32'h38809ba2),
	.w8(32'h37422127),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918574c),
	.w1(32'hb88d9ef6),
	.w2(32'hb80ab21d),
	.w3(32'hb8a77453),
	.w4(32'h3744ab41),
	.w5(32'hb85c2705),
	.w6(32'hb8d266b6),
	.w7(32'h38154f36),
	.w8(32'hb7766f96),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb717ec57),
	.w1(32'h360f2072),
	.w2(32'hb68f7ff7),
	.w3(32'hb7a08dab),
	.w4(32'hb794362a),
	.w5(32'hb7b038d9),
	.w6(32'hb76e0224),
	.w7(32'hb6e3ade5),
	.w8(32'hb71e7900),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ac950),
	.w1(32'hb9415ca4),
	.w2(32'hb8a68d42),
	.w3(32'hb95ecd11),
	.w4(32'hb8d6817b),
	.w5(32'hb8e04e2d),
	.w6(32'hb91a14e1),
	.w7(32'hb8e98eda),
	.w8(32'hb94beea0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b9cbf7),
	.w1(32'hb85427fb),
	.w2(32'hb86d43af),
	.w3(32'hb7e98a24),
	.w4(32'hb82b93c0),
	.w5(32'hb7a2316f),
	.w6(32'hb825247f),
	.w7(32'hb54cdc9e),
	.w8(32'h37384cc5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h338c2461),
	.w1(32'h351e41e1),
	.w2(32'h35a6d17a),
	.w3(32'h35968a04),
	.w4(32'h3534b968),
	.w5(32'h358d0d46),
	.w6(32'h3571fd39),
	.w7(32'h3584f308),
	.w8(32'h35970228),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72e74ae),
	.w1(32'hb7933756),
	.w2(32'h35842138),
	.w3(32'h38044a44),
	.w4(32'h38ace834),
	.w5(32'h389d1bcb),
	.w6(32'h380f19f9),
	.w7(32'h3889633c),
	.w8(32'h375fb093),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35939b68),
	.w1(32'h3622d43f),
	.w2(32'h362bd65b),
	.w3(32'h3606d0a1),
	.w4(32'h34dd49f1),
	.w5(32'h35e6c8b0),
	.w6(32'h3683162b),
	.w7(32'h361a95d1),
	.w8(32'h3651b1d0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c9993),
	.w1(32'hb896141b),
	.w2(32'hb7649f89),
	.w3(32'hb904d3b6),
	.w4(32'hb76bec9d),
	.w5(32'h381fa476),
	.w6(32'hb8f8a91b),
	.w7(32'hb78a3e71),
	.w8(32'h3875dd46),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39601284),
	.w1(32'h3974860d),
	.w2(32'h383a2159),
	.w3(32'h392e5345),
	.w4(32'h3960fea9),
	.w5(32'h381d4df5),
	.w6(32'h3935070b),
	.w7(32'h3935b7cf),
	.w8(32'h38a5f266),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376f4ce3),
	.w1(32'h3832b638),
	.w2(32'hb731fb53),
	.w3(32'h379abce6),
	.w4(32'h37b065b5),
	.w5(32'hb89a65e5),
	.w6(32'h385c72a1),
	.w7(32'h380877ef),
	.w8(32'hb8cc7e26),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ec9e7e),
	.w1(32'hb6d114f3),
	.w2(32'h36030329),
	.w3(32'hb6c3641b),
	.w4(32'h33f8d938),
	.w5(32'h3704718e),
	.w6(32'hb561ebc3),
	.w7(32'h3747fcb8),
	.w8(32'hb51b5429),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c2203c),
	.w1(32'hb6f8bfca),
	.w2(32'hb819111e),
	.w3(32'hb43b8bb8),
	.w4(32'hb73cd41e),
	.w5(32'hb8e73634),
	.w6(32'h3877b05b),
	.w7(32'h3865164e),
	.w8(32'hb8bdb0ce),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b01687),
	.w1(32'hb780abd9),
	.w2(32'h36f6337e),
	.w3(32'hb7e20020),
	.w4(32'h37defc72),
	.w5(32'hb59547df),
	.w6(32'hb82f6b14),
	.w7(32'h36a7013b),
	.w8(32'hb76934d0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a45cef),
	.w1(32'hb93a9a0d),
	.w2(32'hb8fb72dd),
	.w3(32'hb9b09598),
	.w4(32'hb88d1dbe),
	.w5(32'h381693bc),
	.w6(32'hb9a8ba06),
	.w7(32'hb9108326),
	.w8(32'h37ae8855),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363cecd0),
	.w1(32'hb5e90030),
	.w2(32'hb5745d90),
	.w3(32'h35ef21d9),
	.w4(32'hb607b0b6),
	.w5(32'hb5e53bfd),
	.w6(32'hb61997ff),
	.w7(32'hb5a0c22f),
	.w8(32'hb5da0967),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h347ee93e),
	.w1(32'hb64f9358),
	.w2(32'hb561c3d6),
	.w3(32'hb6717c8f),
	.w4(32'hb5db5ce3),
	.w5(32'hb70cc9a6),
	.w6(32'h3512385e),
	.w7(32'h362d2926),
	.w8(32'h36ca484a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb820fdbb),
	.w1(32'h370a8a1d),
	.w2(32'h378f35c7),
	.w3(32'hb7eb3163),
	.w4(32'h37554649),
	.w5(32'hb6db25f0),
	.w6(32'hb8bcba10),
	.w7(32'hb77bd8b3),
	.w8(32'hb822136c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917bd00),
	.w1(32'hb8999fc6),
	.w2(32'hb77a711a),
	.w3(32'hb83d23e9),
	.w4(32'h37ca5dc9),
	.w5(32'hb795a4e7),
	.w6(32'hb8973b32),
	.w7(32'hb63c1ef3),
	.w8(32'hb8478746),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b23ae),
	.w1(32'h37e7e542),
	.w2(32'hb799f825),
	.w3(32'h3671b1e5),
	.w4(32'h383ba2ed),
	.w5(32'hb8043ab9),
	.w6(32'h37dbd9bd),
	.w7(32'h382a0c19),
	.w8(32'hb6e9473e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d39d66),
	.w1(32'hb808745d),
	.w2(32'hb88c8089),
	.w3(32'h384e945d),
	.w4(32'h37959d90),
	.w5(32'hb88b3e3c),
	.w6(32'h38a0a2e7),
	.w7(32'hb75c3a05),
	.w8(32'h367a77d1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6836716),
	.w1(32'h362f3498),
	.w2(32'h3726d253),
	.w3(32'hb686e0f3),
	.w4(32'h369c2557),
	.w5(32'h372952dd),
	.w6(32'hb70de6ac),
	.w7(32'h36401696),
	.w8(32'h36cf0ced),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75e2059),
	.w1(32'hb60c483a),
	.w2(32'h370f9722),
	.w3(32'hb7ae0c30),
	.w4(32'h3538dcd8),
	.w5(32'h37860f7e),
	.w6(32'hb6f9d293),
	.w7(32'h364ab17c),
	.w8(32'h371768a3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dbe224),
	.w1(32'hb894b9a5),
	.w2(32'hb8eb90ef),
	.w3(32'hb85161a5),
	.w4(32'hb81cf12f),
	.w5(32'hb85cc53e),
	.w6(32'hb91e6bf2),
	.w7(32'hb89f9091),
	.w8(32'hb90742ba),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9f617),
	.w1(32'hb9214fcc),
	.w2(32'hb913a8ab),
	.w3(32'hb99d348f),
	.w4(32'hb7a54529),
	.w5(32'h37d69c42),
	.w6(32'hb9a68d06),
	.w7(32'hb9321364),
	.w8(32'h3801a441),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a34689),
	.w1(32'hb86a737f),
	.w2(32'hb86daba9),
	.w3(32'hb89b2a62),
	.w4(32'hb87bacf4),
	.w5(32'hb875a35e),
	.w6(32'h360f500d),
	.w7(32'hb884159e),
	.w8(32'hb966b85d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5fac9),
	.w1(32'h37c7cdce),
	.w2(32'hb6c2717b),
	.w3(32'h37f605de),
	.w4(32'h382c9d9a),
	.w5(32'hb81358f6),
	.w6(32'h38226c15),
	.w7(32'h38bd5915),
	.w8(32'h370a1b0d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b42c9),
	.w1(32'hb8696fdb),
	.w2(32'h35d1de75),
	.w3(32'hb8a73206),
	.w4(32'h37cd8859),
	.w5(32'h382b6e5c),
	.w6(32'hb7822d98),
	.w7(32'h38684b6d),
	.w8(32'h38035711),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361e4ddc),
	.w1(32'hb5496022),
	.w2(32'hb51c187e),
	.w3(32'h35e3a506),
	.w4(32'hb59d5be7),
	.w5(32'h3517d023),
	.w6(32'h335fa45d),
	.w7(32'h32ee49a0),
	.w8(32'hb4e38fe0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57a6348),
	.w1(32'hb41b624c),
	.w2(32'h34d4157c),
	.w3(32'hb48ead6f),
	.w4(32'hb53a4088),
	.w5(32'h3405b517),
	.w6(32'h36057c34),
	.w7(32'h36044725),
	.w8(32'h3603d711),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a17226),
	.w1(32'hb715c60d),
	.w2(32'hb6ff4b18),
	.w3(32'h3511572a),
	.w4(32'hb519af17),
	.w5(32'h3719fdb7),
	.w6(32'hb7653c71),
	.w7(32'hb7490470),
	.w8(32'hb756e566),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c31daa),
	.w1(32'hb59b3217),
	.w2(32'hb52e8b4a),
	.w3(32'hb5821bad),
	.w4(32'hb5fd7425),
	.w5(32'h35bb77fe),
	.w6(32'h3525dee4),
	.w7(32'h35d49f6e),
	.w8(32'h35774075),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb4744),
	.w1(32'hb6e861f6),
	.w2(32'hb6040e02),
	.w3(32'h3750a9a4),
	.w4(32'h36bebdce),
	.w5(32'h37154b5d),
	.w6(32'hb5a7a450),
	.w7(32'h37504820),
	.w8(32'h372bb453),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a886c),
	.w1(32'hb8a86f6e),
	.w2(32'hb7b4396a),
	.w3(32'hb8ab234d),
	.w4(32'hb68adf6a),
	.w5(32'hb80cb66b),
	.w6(32'hb856c114),
	.w7(32'hb73df070),
	.w8(32'hb87be955),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77b66c1),
	.w1(32'h37b8bf87),
	.w2(32'h35340813),
	.w3(32'hb80d04c2),
	.w4(32'hb7de2767),
	.w5(32'hb7462b36),
	.w6(32'h361515eb),
	.w7(32'hb7cc0dd7),
	.w8(32'hb8d520f9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3d9354c),
	.w1(32'hb5c33567),
	.w2(32'h3624d2f3),
	.w3(32'h33a7e7a4),
	.w4(32'h35e2fb63),
	.w5(32'h36751a3c),
	.w6(32'hb6863008),
	.w7(32'hb6658cd1),
	.w8(32'h361f9cd0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958f5f8),
	.w1(32'hb916e2b3),
	.w2(32'hb94b25d7),
	.w3(32'hb7b1698c),
	.w4(32'hb84c3f77),
	.w5(32'hb8251f1b),
	.w6(32'hb83d2cdd),
	.w7(32'hb90f1af3),
	.w8(32'hb924f96d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eb2460),
	.w1(32'h373009db),
	.w2(32'h379169c2),
	.w3(32'hb6b2a15a),
	.w4(32'h37e34e16),
	.w5(32'h376f4059),
	.w6(32'hb831e908),
	.w7(32'hb7c50b51),
	.w8(32'hb7992c30),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368c5bdc),
	.w1(32'h36ec385c),
	.w2(32'h3606602f),
	.w3(32'h35f20ca1),
	.w4(32'h361bf746),
	.w5(32'hb40a0cf6),
	.w6(32'h3656185c),
	.w7(32'h36ca3927),
	.w8(32'h36590ba8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df4044),
	.w1(32'hb8aba1eb),
	.w2(32'hb85630a5),
	.w3(32'hb8e184e3),
	.w4(32'hb87c6e5b),
	.w5(32'hb85d90de),
	.w6(32'hb8c6e1f7),
	.w7(32'hb8c83a46),
	.w8(32'hb8cafcf8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61f42e5),
	.w1(32'hb62a0e26),
	.w2(32'hb45f3bd1),
	.w3(32'hb5f33beb),
	.w4(32'hb5a1e5bc),
	.w5(32'h35a3a6e9),
	.w6(32'hb5850414),
	.w7(32'hb5395aa9),
	.w8(32'h35c5cb36),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3620a1a3),
	.w1(32'h35ddf5ef),
	.w2(32'h364a2379),
	.w3(32'h36190d72),
	.w4(32'h36884358),
	.w5(32'h3656f1d2),
	.w6(32'hb5a8d32f),
	.w7(32'hb213cb5f),
	.w8(32'hb6544a47),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e04a05),
	.w1(32'h33c380f7),
	.w2(32'h3545e82d),
	.w3(32'h360916d3),
	.w4(32'h34127dc0),
	.w5(32'hb50deb6c),
	.w6(32'h358cd034),
	.w7(32'h34ba89c4),
	.w8(32'hb4a32f2a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb515ca6b),
	.w1(32'hb59385fc),
	.w2(32'h3593d2b6),
	.w3(32'hb505849d),
	.w4(32'hb5f50d05),
	.w5(32'h34229059),
	.w6(32'hb5b09dff),
	.w7(32'h34f0c23d),
	.w8(32'hb55e971c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370d0eb0),
	.w1(32'h36f4fa2e),
	.w2(32'hb58422f9),
	.w3(32'hb75ce794),
	.w4(32'h379b329c),
	.w5(32'h37cf2974),
	.w6(32'h372d82f3),
	.w7(32'h37f5d2d6),
	.w8(32'h379ab464),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e0b643),
	.w1(32'hb7da3a02),
	.w2(32'h38062986),
	.w3(32'hb5e1c33f),
	.w4(32'h38a98ab7),
	.w5(32'h381adced),
	.w6(32'h374bedb1),
	.w7(32'h38c6b4bd),
	.w8(32'h3763fb2c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce2ecf),
	.w1(32'hb87f1c2c),
	.w2(32'hb7cb5f25),
	.w3(32'hb8a9307f),
	.w4(32'hb81eed80),
	.w5(32'hb888c942),
	.w6(32'hb89e62ba),
	.w7(32'hb81b99db),
	.w8(32'hb882d7b6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92df4ac),
	.w1(32'hb90bea37),
	.w2(32'hb8c83672),
	.w3(32'hb881290a),
	.w4(32'hb79d2943),
	.w5(32'hb85100cb),
	.w6(32'hb89f8e18),
	.w7(32'hb85fddf5),
	.w8(32'hb89ea93c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351c33e8),
	.w1(32'h35663629),
	.w2(32'hb668a3b9),
	.w3(32'h3607176f),
	.w4(32'h35925a40),
	.w5(32'hb65121c3),
	.w6(32'h362a5989),
	.w7(32'h366a1423),
	.w8(32'hb5b3cae9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62ffa64),
	.w1(32'h362b179b),
	.w2(32'h36d95e21),
	.w3(32'hb58216ad),
	.w4(32'h36539e39),
	.w5(32'h36b856cb),
	.w6(32'h3646e237),
	.w7(32'h370ad30b),
	.w8(32'h362d3625),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb513a123),
	.w1(32'hb40ebd2f),
	.w2(32'hb28ce497),
	.w3(32'hb48b57b7),
	.w4(32'hb56a0767),
	.w5(32'hb3a09972),
	.w6(32'h34c43d0e),
	.w7(32'h3419c968),
	.w8(32'h323007b9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4bee10d),
	.w1(32'hb56add62),
	.w2(32'hb58d638c),
	.w3(32'h3354ba94),
	.w4(32'hb483f033),
	.w5(32'hb48956df),
	.w6(32'h35be7686),
	.w7(32'h35b889ad),
	.w8(32'h34de1d51),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8439b17),
	.w1(32'h36d1df45),
	.w2(32'h36fb5ff3),
	.w3(32'hb79743ad),
	.w4(32'h375158db),
	.w5(32'hb882c642),
	.w6(32'h381a275d),
	.w7(32'h382da342),
	.w8(32'hb8905062),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36589c78),
	.w1(32'h36341724),
	.w2(32'h36477d96),
	.w3(32'hb607aefe),
	.w4(32'hb472b456),
	.w5(32'h365012dd),
	.w6(32'h35a704e6),
	.w7(32'h345f9273),
	.w8(32'h35a8b495),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3741cc5f),
	.w1(32'h366d3c06),
	.w2(32'hb738aad3),
	.w3(32'h371d9fe3),
	.w4(32'h375fce39),
	.w5(32'h368bb146),
	.w6(32'h36d00b1d),
	.w7(32'h37166693),
	.w8(32'hb6da9f9a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b6c616),
	.w1(32'h379091df),
	.w2(32'h37323cd3),
	.w3(32'h375352e1),
	.w4(32'h3786e031),
	.w5(32'h375c3f85),
	.w6(32'h37a64689),
	.w7(32'h380c36bf),
	.w8(32'h37ab5bf8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb549b9b5),
	.w1(32'hb52d7a7d),
	.w2(32'h34a58946),
	.w3(32'hb4db04ac),
	.w4(32'hb55e1cbe),
	.w5(32'h35bc92cf),
	.w6(32'h34573df4),
	.w7(32'hb5a079dc),
	.w8(32'hb45408d5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e33fb8),
	.w1(32'hb86888e9),
	.w2(32'hb83214c3),
	.w3(32'hb890ac68),
	.w4(32'hb7ceb64a),
	.w5(32'hb73e42cb),
	.w6(32'hb8711af2),
	.w7(32'hb82b3f5a),
	.w8(32'hb6c952fc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375d5004),
	.w1(32'h36f8e4f2),
	.w2(32'h36c43ca6),
	.w3(32'h36b8b288),
	.w4(32'h36eb56fd),
	.w5(32'h36c07c30),
	.w6(32'h370e60ea),
	.w7(32'h3723080c),
	.w8(32'h36acf726),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890ad3a),
	.w1(32'h3827eb7b),
	.w2(32'h3889dd87),
	.w3(32'hb8f6c87c),
	.w4(32'h37d949a3),
	.w5(32'h38262d34),
	.w6(32'h389efee7),
	.w7(32'h38b5a79a),
	.w8(32'hb82b5808),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4e1a45e),
	.w1(32'h34d5434f),
	.w2(32'h34879f8f),
	.w3(32'h351d27c5),
	.w4(32'hb5107f01),
	.w5(32'h34a254aa),
	.w6(32'h32ddefa7),
	.w7(32'hb4a7a2c5),
	.w8(32'h359f3693),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b397f),
	.w1(32'h38b10e30),
	.w2(32'hb70a8f58),
	.w3(32'h37885b06),
	.w4(32'hb7124fad),
	.w5(32'hb8fd99c5),
	.w6(32'h39139176),
	.w7(32'h3911b14a),
	.w8(32'h375f55c8),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule