module layer_8_featuremap_126(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885c39),
	.w1(32'hbb9bff2f),
	.w2(32'hbb2a3e9e),
	.w3(32'hbc02529a),
	.w4(32'hbb3e35ca),
	.w5(32'h3a287f2f),
	.w6(32'hba07a29b),
	.w7(32'hbbef0328),
	.w8(32'hbb79b930),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac86d60),
	.w1(32'hbaf1daf3),
	.w2(32'hb92d2063),
	.w3(32'h3a934c69),
	.w4(32'h3ade6deb),
	.w5(32'hba1a8c43),
	.w6(32'hbb014514),
	.w7(32'h39a2f7c2),
	.w8(32'hbba2fe0f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d6642),
	.w1(32'hbbbbf3e8),
	.w2(32'hbb138f26),
	.w3(32'hbb464fea),
	.w4(32'h3ade7469),
	.w5(32'hbb881e9a),
	.w6(32'hbb53ab4a),
	.w7(32'h3b1b5f3c),
	.w8(32'hbabd36e1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02002c),
	.w1(32'h3ad6306c),
	.w2(32'hba82f3f9),
	.w3(32'h3b1a0f68),
	.w4(32'hb6f61744),
	.w5(32'hba8b8a73),
	.w6(32'h3c6f80a6),
	.w7(32'hbab38a50),
	.w8(32'hbbe7e9b2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03159e),
	.w1(32'h3948e265),
	.w2(32'h3a762149),
	.w3(32'h3ae36bea),
	.w4(32'hba65ab61),
	.w5(32'h3a5ace19),
	.w6(32'h3a85950c),
	.w7(32'h3b21f168),
	.w8(32'h3b8f6fb9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a446591),
	.w1(32'h37c80e60),
	.w2(32'h3a643d01),
	.w3(32'hba4802ba),
	.w4(32'h3b1e161a),
	.w5(32'h3a3c796d),
	.w6(32'h3b9014b1),
	.w7(32'h3a39bfe2),
	.w8(32'hbba85d3c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46d48e),
	.w1(32'h3b60a20d),
	.w2(32'hba786eda),
	.w3(32'h3a8714ab),
	.w4(32'hbb0a1bbe),
	.w5(32'h3a48bf02),
	.w6(32'h3b5fe8e2),
	.w7(32'hbae86cbf),
	.w8(32'hbb7bb3c8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78d611),
	.w1(32'h3a9b6d6d),
	.w2(32'h3b99cec8),
	.w3(32'hbb17fd49),
	.w4(32'h3b6a5d90),
	.w5(32'h3acac63d),
	.w6(32'hbb359756),
	.w7(32'h3be307bd),
	.w8(32'h3acffecb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29c557),
	.w1(32'hbc2b0950),
	.w2(32'h3b3988d9),
	.w3(32'hba5c4578),
	.w4(32'h3a92672b),
	.w5(32'h3ba04b8d),
	.w6(32'hbbc0a082),
	.w7(32'hbb647815),
	.w8(32'hbb652132),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7d470),
	.w1(32'h3b48e730),
	.w2(32'hb97e1d04),
	.w3(32'h3b598d23),
	.w4(32'hba3f58a4),
	.w5(32'h3af3f594),
	.w6(32'hbb1def6a),
	.w7(32'h398f3da1),
	.w8(32'h3b5cf803),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf5f9),
	.w1(32'h3ae4ebc5),
	.w2(32'h3b0c254f),
	.w3(32'h3b41e6ed),
	.w4(32'h3a82253c),
	.w5(32'h3a655f8c),
	.w6(32'hbad1c736),
	.w7(32'hb7cbb0b6),
	.w8(32'hba9e3106),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e8a98),
	.w1(32'h3a837f79),
	.w2(32'hbaeab57a),
	.w3(32'h3b38348c),
	.w4(32'hbb55bf7e),
	.w5(32'hbbbec664),
	.w6(32'hbb0429d5),
	.w7(32'hbb0913e7),
	.w8(32'hbb7fe649),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad09cd1),
	.w1(32'h3b1c49c4),
	.w2(32'h3b00a903),
	.w3(32'hbb6d340d),
	.w4(32'h3a67cfd1),
	.w5(32'h3b008ec1),
	.w6(32'hbb2e4b75),
	.w7(32'hba82d1ec),
	.w8(32'hb8a230fa),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9994723),
	.w1(32'hb993aed2),
	.w2(32'hb96cb2bd),
	.w3(32'hb963e076),
	.w4(32'hb993be82),
	.w5(32'hb94a62d9),
	.w6(32'hb8fddead),
	.w7(32'hb9278b25),
	.w8(32'hb9014638),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66acd3f),
	.w1(32'h36fc3879),
	.w2(32'h37b0dfec),
	.w3(32'hb760fcc2),
	.w4(32'hb6da228b),
	.w5(32'h36ae62ac),
	.w6(32'hb77c48e9),
	.w7(32'hb6c1b299),
	.w8(32'h3626796a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8215ec8),
	.w1(32'h389a455f),
	.w2(32'h38cc5501),
	.w3(32'hb89f0e21),
	.w4(32'hb76575a5),
	.w5(32'hb852a89f),
	.w6(32'hb9205d9c),
	.w7(32'hb8958ec8),
	.w8(32'hb7eacb73),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cafc93),
	.w1(32'h3987b727),
	.w2(32'h39d8b65d),
	.w3(32'h39c0a007),
	.w4(32'h3a05f131),
	.w5(32'h39e979d4),
	.w6(32'h3860cfd4),
	.w7(32'h39d4d0fd),
	.w8(32'h3a1cea1b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959023e),
	.w1(32'h3aa9e377),
	.w2(32'h39ec5162),
	.w3(32'h3a4017b3),
	.w4(32'hb90d2dd6),
	.w5(32'h3aa91a43),
	.w6(32'hb85acc62),
	.w7(32'hba8152fd),
	.w8(32'h3a201451),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69ffa),
	.w1(32'hbb45fbf9),
	.w2(32'h3b6e981e),
	.w3(32'hbb8d41da),
	.w4(32'hbb4cf10a),
	.w5(32'h3b860ba0),
	.w6(32'h3a5c55a7),
	.w7(32'hbb047852),
	.w8(32'h3b8eb9d7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc52abf),
	.w1(32'hbbf33ff1),
	.w2(32'hbb1eaaf0),
	.w3(32'hbb61e47a),
	.w4(32'hbbeb28da),
	.w5(32'hbb15c56a),
	.w6(32'h3ad68c05),
	.w7(32'hba9c6551),
	.w8(32'h3a54d2d9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36d84b),
	.w1(32'hba9144bb),
	.w2(32'hb9e3f85b),
	.w3(32'hb9e939a0),
	.w4(32'hb8a9ec83),
	.w5(32'hb9c3a64f),
	.w6(32'hbaae1212),
	.w7(32'hbad5a5e4),
	.w8(32'hbacc3352),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7c95),
	.w1(32'h3b2dd466),
	.w2(32'h3ab7d575),
	.w3(32'h3a536d3c),
	.w4(32'h3b2132f9),
	.w5(32'h3acf4544),
	.w6(32'h3a6154d3),
	.w7(32'h3acfcb35),
	.w8(32'h3adc2d4b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba651f6),
	.w1(32'hbbd43e6c),
	.w2(32'h3a75cc07),
	.w3(32'hbb7a919b),
	.w4(32'hbba6ccd6),
	.w5(32'h3a6ee761),
	.w6(32'hba257fad),
	.w7(32'hba13440f),
	.w8(32'h3ac02fc4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043411),
	.w1(32'hbb5af2c1),
	.w2(32'hbac1cc55),
	.w3(32'hbaf30f4d),
	.w4(32'hbb21ea19),
	.w5(32'hbac6b717),
	.w6(32'hba59ec21),
	.w7(32'hbac22fdc),
	.w8(32'hba882b74),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba211884),
	.w1(32'hb9d1c7ba),
	.w2(32'hb93c3989),
	.w3(32'hba9babe3),
	.w4(32'hba569a4d),
	.w5(32'hba4d34c1),
	.w6(32'hba9e028d),
	.w7(32'hba8eafd4),
	.w8(32'hba3e6f2e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b0a46),
	.w1(32'hbb81e218),
	.w2(32'h3a709775),
	.w3(32'hba7a0117),
	.w4(32'hbb5f213f),
	.w5(32'h39dcad26),
	.w6(32'h3a0a4fbd),
	.w7(32'hba8ee2bf),
	.w8(32'h39e231c1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944cab2),
	.w1(32'h392b88d6),
	.w2(32'hb83ec293),
	.w3(32'h39d491af),
	.w4(32'h3988a5c5),
	.w5(32'h367a10b2),
	.w6(32'h394501de),
	.w7(32'h387d12f2),
	.w8(32'hb9178c73),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9cc82),
	.w1(32'hbc564351),
	.w2(32'hbc9926b2),
	.w3(32'hbbd9ee05),
	.w4(32'hbc3efd21),
	.w5(32'hbc834183),
	.w6(32'hbb5e7e62),
	.w7(32'h3c08e33c),
	.w8(32'hbb85b796),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c54014),
	.w1(32'hb9d574cd),
	.w2(32'h3a532f1c),
	.w3(32'hba020bc8),
	.w4(32'hb9d6a9e1),
	.w5(32'h3a4baad2),
	.w6(32'h386bb598),
	.w7(32'h3849fc13),
	.w8(32'h3a19f983),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39913de6),
	.w1(32'h3a4c529a),
	.w2(32'h39d344ce),
	.w3(32'h39475e0d),
	.w4(32'h3a24ab01),
	.w5(32'h3987360f),
	.w6(32'h3885e390),
	.w7(32'h39f2f8cb),
	.w8(32'h396b12f6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad63265),
	.w1(32'h3a9427e5),
	.w2(32'hb9526c14),
	.w3(32'h3a006e5a),
	.w4(32'h3a0bcf73),
	.w5(32'hba80d7a9),
	.w6(32'hb9e50a7f),
	.w7(32'hba601a50),
	.w8(32'hbaa98f63),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b667ae),
	.w1(32'hb8a8bf7f),
	.w2(32'h39a1099d),
	.w3(32'hb9035a7a),
	.w4(32'hb9304755),
	.w5(32'h39850bd4),
	.w6(32'h38686a1a),
	.w7(32'hba1d23ef),
	.w8(32'h391520f1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3753f111),
	.w1(32'hb8c4aa8f),
	.w2(32'hb808a69f),
	.w3(32'hb819d17a),
	.w4(32'hb6c030fe),
	.w5(32'hb810bf23),
	.w6(32'hb80c9af7),
	.w7(32'hb8aa1c4e),
	.w8(32'hb8587136),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b71c49),
	.w1(32'hb7b0c473),
	.w2(32'h37ee7eda),
	.w3(32'hb78df1bd),
	.w4(32'hb8093c17),
	.w5(32'h36572006),
	.w6(32'hb658b4e3),
	.w7(32'hb66774dc),
	.w8(32'h37bc9adb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c6b7f),
	.w1(32'hbac898c7),
	.w2(32'hbb0baf8c),
	.w3(32'hba4b59c9),
	.w4(32'hbad99eb2),
	.w5(32'hbb30c732),
	.w6(32'hba5a5579),
	.w7(32'hba7b7b87),
	.w8(32'hbac60b78),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cf8bc),
	.w1(32'hbb1f84f8),
	.w2(32'hba99cd00),
	.w3(32'hbac92c75),
	.w4(32'hbafb5e15),
	.w5(32'hba91f41c),
	.w6(32'hba7af17e),
	.w7(32'hbab4cbdf),
	.w8(32'hba5febe5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38554827),
	.w1(32'h379a103f),
	.w2(32'h377140a4),
	.w3(32'h389d2e94),
	.w4(32'h388092f0),
	.w5(32'h38641019),
	.w6(32'h37823f8d),
	.w7(32'h38ba1722),
	.w8(32'h38835c7e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1def4),
	.w1(32'h3a4d474f),
	.w2(32'h38a145a3),
	.w3(32'h3a99e05c),
	.w4(32'h3adbaa56),
	.w5(32'h39e62616),
	.w6(32'h3a939f33),
	.w7(32'h3ab60a31),
	.w8(32'h3a072377),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d7de8),
	.w1(32'hb9560b5a),
	.w2(32'hb9817dc5),
	.w3(32'hb8d6b173),
	.w4(32'hb9855354),
	.w5(32'hb9b9f0bb),
	.w6(32'hb8e9e05b),
	.w7(32'hb964e998),
	.w8(32'hb98c0bfc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fcd3a),
	.w1(32'hb8125595),
	.w2(32'hb7f7f179),
	.w3(32'hb8e0001d),
	.w4(32'hb8a614b4),
	.w5(32'hb86dd0e4),
	.w6(32'hb8209f78),
	.w7(32'hb884e60f),
	.w8(32'hb79081eb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d25d8),
	.w1(32'hbb1292a5),
	.w2(32'hba99431b),
	.w3(32'h3a31e6b0),
	.w4(32'hb92dbeb1),
	.w5(32'hb6b5a3df),
	.w6(32'h3a5beb92),
	.w7(32'hb893f842),
	.w8(32'hb9408884),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b8a08),
	.w1(32'h37fbf8bb),
	.w2(32'hb989e5a5),
	.w3(32'h3a67c316),
	.w4(32'h3a0120bc),
	.w5(32'h393de9f6),
	.w6(32'h3a92bcc8),
	.w7(32'h3a06872c),
	.w8(32'h3987a82c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6db45f9),
	.w1(32'h37a133eb),
	.w2(32'h384b5145),
	.w3(32'h37feeab5),
	.w4(32'h3825cea9),
	.w5(32'h37a64b1f),
	.w6(32'hb89d333c),
	.w7(32'hb81d9103),
	.w8(32'h37d6008e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba651e3e),
	.w1(32'hbada59c8),
	.w2(32'hba1f8bd6),
	.w3(32'hba7fbc73),
	.w4(32'hbacbb350),
	.w5(32'hba6c60fb),
	.w6(32'hb98a4bb2),
	.w7(32'hba4aee61),
	.w8(32'hba656f8f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891103a),
	.w1(32'h398dd176),
	.w2(32'h3b4b68d1),
	.w3(32'hb9c90a22),
	.w4(32'hb9e8f4e2),
	.w5(32'h3b2a1917),
	.w6(32'h3a8f6cf9),
	.w7(32'h3a3b9c2b),
	.w8(32'h3b381e04),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3dffb),
	.w1(32'h3883cb1d),
	.w2(32'h38a0d8ed),
	.w3(32'h354e9f4b),
	.w4(32'h38f1a783),
	.w5(32'h3942dee9),
	.w6(32'h3924a828),
	.w7(32'h39a4bc83),
	.w8(32'h39df64de),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3746fb3b),
	.w1(32'hb75f0727),
	.w2(32'h37bbc9f1),
	.w3(32'hb6c06942),
	.w4(32'hb41492f8),
	.w5(32'h37e85818),
	.w6(32'hb715a97e),
	.w7(32'h36a0f11c),
	.w8(32'hb6953d3f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0925b9),
	.w1(32'hbb21e39a),
	.w2(32'h3a895a94),
	.w3(32'hbb3a7cf0),
	.w4(32'hbb365353),
	.w5(32'h3a5b70a8),
	.w6(32'hb661f2b7),
	.w7(32'hb9dfd254),
	.w8(32'h3b155e19),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c687f5),
	.w1(32'hba2a158a),
	.w2(32'h38425212),
	.w3(32'h36dfd418),
	.w4(32'hb83a826a),
	.w5(32'h39b72758),
	.w6(32'h3a12841b),
	.w7(32'h3944709b),
	.w8(32'h3a1911bc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba902311),
	.w1(32'hba11ea17),
	.w2(32'h3814973f),
	.w3(32'hba0a011d),
	.w4(32'hb9e19de9),
	.w5(32'h39977e78),
	.w6(32'hb9233ae0),
	.w7(32'hba22f93f),
	.w8(32'hb7a686ec),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b503a17),
	.w1(32'h3b95b716),
	.w2(32'h3a5ad942),
	.w3(32'h3b4a4e62),
	.w4(32'h3b85120e),
	.w5(32'h3a83d9ad),
	.w6(32'h3b3f818d),
	.w7(32'h3b6aaefe),
	.w8(32'h3aab1690),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ba130),
	.w1(32'hbaedd3df),
	.w2(32'h3aa97dec),
	.w3(32'hbbe8cc94),
	.w4(32'hbbf6699d),
	.w5(32'hb94030d2),
	.w6(32'hba950337),
	.w7(32'hbb50543f),
	.w8(32'h3b946c31),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33f341),
	.w1(32'hbaf667a9),
	.w2(32'h3b09debb),
	.w3(32'hbb953126),
	.w4(32'hbb8466c8),
	.w5(32'h3a4d08b1),
	.w6(32'hba94399c),
	.w7(32'hbad51718),
	.w8(32'h3acf6cbe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bf64c),
	.w1(32'hba253f50),
	.w2(32'hb9c4faed),
	.w3(32'h3987234a),
	.w4(32'h38f2dccb),
	.w5(32'hb73eeb10),
	.w6(32'h39b34952),
	.w7(32'h38f6ec4e),
	.w8(32'h3783cf81),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0788c),
	.w1(32'hb6f42e6c),
	.w2(32'h372d9cd6),
	.w3(32'hb819ed50),
	.w4(32'hb7d14a45),
	.w5(32'hb6d668e2),
	.w6(32'hb6cc802c),
	.w7(32'h3623b93a),
	.w8(32'h377bdefe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c938),
	.w1(32'hbaf13ded),
	.w2(32'h3a97b6ed),
	.w3(32'hba34f37b),
	.w4(32'hba88328b),
	.w5(32'h3af66ede),
	.w6(32'h398311ae),
	.w7(32'h3a131604),
	.w8(32'h3b2ede4e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986757d),
	.w1(32'h39c2394d),
	.w2(32'hb9a36cb5),
	.w3(32'hb9d3680d),
	.w4(32'hb8485ac4),
	.w5(32'hb98447e0),
	.w6(32'hba1a6f79),
	.w7(32'hba7d3df9),
	.w8(32'hba50c38c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a02f6),
	.w1(32'h3ac8bda0),
	.w2(32'h3a935046),
	.w3(32'hba729898),
	.w4(32'hba96a02b),
	.w5(32'hb9c80fbf),
	.w6(32'h393048e8),
	.w7(32'hb9b5f9e8),
	.w8(32'h3a59497a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dc715),
	.w1(32'hb943fc0a),
	.w2(32'h3a4d7a3a),
	.w3(32'hb74dbc26),
	.w4(32'hb919f9a3),
	.w5(32'h3aa3fdca),
	.w6(32'h39c6385e),
	.w7(32'h3a15b243),
	.w8(32'h3aa07ac5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b454df),
	.w1(32'h3906eb26),
	.w2(32'h38fc341a),
	.w3(32'h386dd510),
	.w4(32'h3831c050),
	.w5(32'h38cc48ee),
	.w6(32'hb72ab7c9),
	.w7(32'h38659761),
	.w8(32'h39089c21),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35afeabf),
	.w1(32'h38bb8752),
	.w2(32'h3929e378),
	.w3(32'h37af6699),
	.w4(32'hb8398705),
	.w5(32'h385318e0),
	.w6(32'hb7ae8406),
	.w7(32'hb90af1ee),
	.w8(32'hb91e89d5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387e910e),
	.w1(32'h380d953f),
	.w2(32'h3838bf01),
	.w3(32'h385ea1fb),
	.w4(32'h386e4e54),
	.w5(32'h3848fefd),
	.w6(32'h37cca57e),
	.w7(32'h38884690),
	.w8(32'h38ab93cf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99577be),
	.w1(32'hba660122),
	.w2(32'h3a4f2d0c),
	.w3(32'hba3e811a),
	.w4(32'hbac62e66),
	.w5(32'h389d598e),
	.w6(32'h3987c8bd),
	.w7(32'hb925440c),
	.w8(32'h3a52cf71),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08cee1),
	.w1(32'hb93e12a1),
	.w2(32'hba2f973f),
	.w3(32'hbab21150),
	.w4(32'hbb0d8ab5),
	.w5(32'hbae3a799),
	.w6(32'hba91be75),
	.w7(32'hbb289e39),
	.w8(32'hbb09c341),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2b400),
	.w1(32'hba409cab),
	.w2(32'hba4f5adb),
	.w3(32'hb992d249),
	.w4(32'hbabd3514),
	.w5(32'hbae37ad2),
	.w6(32'hba852866),
	.w7(32'hbae79f46),
	.w8(32'hbb2e243a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50d939),
	.w1(32'hba7356ed),
	.w2(32'h38621da3),
	.w3(32'hbaeff4ef),
	.w4(32'hbb12813a),
	.w5(32'hba9b1d8a),
	.w6(32'hb984664a),
	.w7(32'hba263342),
	.w8(32'h38c033ef),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ac07b),
	.w1(32'h3aa652aa),
	.w2(32'h3adbc99d),
	.w3(32'h3aa3f718),
	.w4(32'h39d5b5ab),
	.w5(32'h39db2821),
	.w6(32'h3a616b64),
	.w7(32'h3a820d06),
	.w8(32'h3a492fc9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba580c17),
	.w1(32'hba22a21b),
	.w2(32'hb8dc074c),
	.w3(32'hba44ea99),
	.w4(32'hba29b99d),
	.w5(32'hb90087a3),
	.w6(32'hba0ea606),
	.w7(32'hba38c685),
	.w8(32'hb9f67900),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1c543),
	.w1(32'h39b3587f),
	.w2(32'h39d80144),
	.w3(32'h39d91e13),
	.w4(32'h39d2378d),
	.w5(32'h39c6dadc),
	.w6(32'h39b05ebd),
	.w7(32'h398ab63d),
	.w8(32'h39a02881),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0766d7),
	.w1(32'hbb9696ea),
	.w2(32'hbb6332a1),
	.w3(32'hbb23ce3d),
	.w4(32'hbbb2c330),
	.w5(32'hbbad3446),
	.w6(32'hba97b138),
	.w7(32'hbaebe8bf),
	.w8(32'hbb3f1d99),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a6247),
	.w1(32'h390820cd),
	.w2(32'h37f47111),
	.w3(32'h38c54e20),
	.w4(32'h38a93249),
	.w5(32'hb80e5b7f),
	.w6(32'h38a0ed37),
	.w7(32'h386d1889),
	.w8(32'hb7764140),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e51d8),
	.w1(32'hbb49a4d5),
	.w2(32'hba66e8f4),
	.w3(32'hbacec8f2),
	.w4(32'hbb299410),
	.w5(32'hba4340c7),
	.w6(32'h398f8b33),
	.w7(32'hba5b32ea),
	.w8(32'h394f8be7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395059c6),
	.w1(32'h39a0b32b),
	.w2(32'h39aec485),
	.w3(32'h3992d121),
	.w4(32'h39ae53b4),
	.w5(32'h39a1144d),
	.w6(32'h393cdafc),
	.w7(32'h39ab579a),
	.w8(32'h399aa2ce),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8e19c),
	.w1(32'h3a8d1593),
	.w2(32'h39e98edb),
	.w3(32'h3b0e8103),
	.w4(32'h3ad44646),
	.w5(32'h396ff566),
	.w6(32'h397e67b5),
	.w7(32'h3a0468b2),
	.w8(32'hba6f97c3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888eadd),
	.w1(32'hb80ee48b),
	.w2(32'hb7b2f807),
	.w3(32'hb7d80410),
	.w4(32'hb7f4fcd0),
	.w5(32'h36c30cc6),
	.w6(32'hb74fbdfa),
	.w7(32'h37967180),
	.w8(32'hb6d91d10),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dc637),
	.w1(32'hba1913f8),
	.w2(32'h3a80ac59),
	.w3(32'hbaab1db6),
	.w4(32'h3a1ab27f),
	.w5(32'h3af87249),
	.w6(32'hb933dee5),
	.w7(32'h39d582b1),
	.w8(32'h3aca0c6d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce3fe8),
	.w1(32'hb7c323b9),
	.w2(32'h38006e8b),
	.w3(32'h37bf2928),
	.w4(32'h37bc1472),
	.w5(32'h37fb3d2c),
	.w6(32'hb60c12f9),
	.w7(32'h381451ee),
	.w8(32'h387228ed),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bdedf),
	.w1(32'hbb2de786),
	.w2(32'h3a3f2175),
	.w3(32'hbb33c005),
	.w4(32'hbb44b58e),
	.w5(32'h39b34816),
	.w6(32'hb953648a),
	.w7(32'hba97fcb8),
	.w8(32'h3a2c7e30),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a115ea7),
	.w1(32'h3a2aec28),
	.w2(32'h39c59235),
	.w3(32'h39033728),
	.w4(32'h389e9dd1),
	.w5(32'hb9861734),
	.w6(32'h391e34ea),
	.w7(32'h393012e9),
	.w8(32'h3901c948),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb715ee9a),
	.w1(32'hb9903581),
	.w2(32'hb8f98e96),
	.w3(32'hb90ee6dc),
	.w4(32'hb98634d8),
	.w5(32'hb8d18004),
	.w6(32'hb9b05813),
	.w7(32'hb97aeaae),
	.w8(32'hb93ccd98),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f50367),
	.w1(32'h3782dbb4),
	.w2(32'h3806fc1c),
	.w3(32'h36a86253),
	.w4(32'h37171601),
	.w5(32'h37d16137),
	.w6(32'h36d3cf60),
	.w7(32'h36465656),
	.w8(32'h36bebe36),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d4afcf),
	.w1(32'h389ae29d),
	.w2(32'h39be0e18),
	.w3(32'h3a25c61e),
	.w4(32'h3a0cbafe),
	.w5(32'h3a4a6156),
	.w6(32'h3a82b90e),
	.w7(32'h3a7bed5a),
	.w8(32'h3ab24a9a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf736),
	.w1(32'hbb26eb81),
	.w2(32'h3a59a2b4),
	.w3(32'hbb06cc3b),
	.w4(32'hbb430761),
	.w5(32'h39b60cb0),
	.w6(32'h3926669e),
	.w7(32'hba15daa6),
	.w8(32'h3a513a83),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38562b9e),
	.w1(32'hb97f1e3a),
	.w2(32'h35d8dfe8),
	.w3(32'h3a167832),
	.w4(32'h398c3283),
	.w5(32'h396e0539),
	.w6(32'h39de5ee3),
	.w7(32'h393d3c2c),
	.w8(32'h399195c7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28ee6b),
	.w1(32'hbb992c7e),
	.w2(32'h38c216f4),
	.w3(32'hbab74bbb),
	.w4(32'hbb57b513),
	.w5(32'h39bff9f2),
	.w6(32'h3a9df9fe),
	.w7(32'hba25a000),
	.w8(32'h393a583b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5250c1),
	.w1(32'hbb5ec828),
	.w2(32'h3992008d),
	.w3(32'hbb2c601e),
	.w4(32'hbba5635b),
	.w5(32'hbacfa36c),
	.w6(32'hbadc6aa7),
	.w7(32'hbb47d8e2),
	.w8(32'hba8ab68b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a3ead),
	.w1(32'h3837f727),
	.w2(32'h3639e02a),
	.w3(32'hb7abdc08),
	.w4(32'h383b1919),
	.w5(32'h388b3f5d),
	.w6(32'hb7a30c9e),
	.w7(32'hb835821a),
	.w8(32'h34b92b98),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb735e9a0),
	.w1(32'h37621875),
	.w2(32'h37c09e16),
	.w3(32'hb77b2462),
	.w4(32'h35af90f1),
	.w5(32'h376ff6f0),
	.w6(32'hb76e96de),
	.w7(32'hb69f57d6),
	.w8(32'h37079f88),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7db0456),
	.w1(32'h3826c61b),
	.w2(32'h38ff9c9a),
	.w3(32'hb7f6c88a),
	.w4(32'hb78ef8c0),
	.w5(32'h37b279c3),
	.w6(32'hb8847cf4),
	.w7(32'h37588851),
	.w8(32'h388c4425),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9465d0),
	.w1(32'hbaf878fc),
	.w2(32'hba8fd70a),
	.w3(32'hbaa44264),
	.w4(32'hbafb28a2),
	.w5(32'hba8631e9),
	.w6(32'hbae65672),
	.w7(32'hbaeae2bd),
	.w8(32'hbaa3f8c0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082424),
	.w1(32'hb985e446),
	.w2(32'hb9fc84d9),
	.w3(32'hb9ff86ff),
	.w4(32'hb9df0292),
	.w5(32'hb9dc76c6),
	.w6(32'hb98109d1),
	.w7(32'hb91ab665),
	.w8(32'hb8bb1f2f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bc205),
	.w1(32'hba4d9ccf),
	.w2(32'hba8b2039),
	.w3(32'hb9bd3b76),
	.w4(32'hba570588),
	.w5(32'hbae1d04e),
	.w6(32'hb9ac3e66),
	.w7(32'hba7b5bbc),
	.w8(32'hbabc6abc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92835e9),
	.w1(32'hba29240e),
	.w2(32'hb9c9db64),
	.w3(32'hb7fdcf29),
	.w4(32'hb9e7c7ab),
	.w5(32'hb94692fd),
	.w6(32'h3962e52c),
	.w7(32'hb9707452),
	.w8(32'h3909c2e9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55bb40),
	.w1(32'hba9b444a),
	.w2(32'hb83bbaf3),
	.w3(32'hba6ff5c9),
	.w4(32'hbacbcff4),
	.w5(32'hb9b3638a),
	.w6(32'h394743a3),
	.w7(32'hba0c4887),
	.w8(32'h390b1d94),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39361e7f),
	.w1(32'h3906f112),
	.w2(32'h3aaa1c37),
	.w3(32'h3a0675c2),
	.w4(32'h3a148371),
	.w5(32'h3ae9bbb0),
	.w6(32'h3a167b01),
	.w7(32'h3a39192e),
	.w8(32'h3b08d336),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984eb2b),
	.w1(32'hbab42e8d),
	.w2(32'h38b36b4b),
	.w3(32'hbab74212),
	.w4(32'hbb04ceb4),
	.w5(32'hbaaa2c25),
	.w6(32'hba30d945),
	.w7(32'hbad68c68),
	.w8(32'hba9a5ef2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc7052),
	.w1(32'hbba7d161),
	.w2(32'h3a3ddb15),
	.w3(32'hbba84ec4),
	.w4(32'hbb8effed),
	.w5(32'h3a8f4b94),
	.w6(32'hba92616b),
	.w7(32'hbae4ffdb),
	.w8(32'h3ac9ac72),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c007bd),
	.w1(32'hb665edef),
	.w2(32'h361fe93f),
	.w3(32'h36e32cd1),
	.w4(32'h36b9c855),
	.w5(32'hb6d33355),
	.w6(32'hb6aa435a),
	.w7(32'hb647ab75),
	.w8(32'hb77327cc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e3ff3),
	.w1(32'h37df5790),
	.w2(32'h378368cd),
	.w3(32'hb814acc3),
	.w4(32'hb7b0534f),
	.w5(32'hb821b14e),
	.w6(32'hb8620a41),
	.w7(32'hb8053087),
	.w8(32'hb8218d62),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376ddb52),
	.w1(32'h38009f10),
	.w2(32'h3812d9cc),
	.w3(32'hb75e19d6),
	.w4(32'h370a2a8a),
	.w5(32'h3713dca2),
	.w6(32'hb7c2a711),
	.w7(32'hb72a688b),
	.w8(32'h353ec582),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39082c8e),
	.w1(32'h38844748),
	.w2(32'hb89aeb2b),
	.w3(32'hb821a019),
	.w4(32'hb96fe954),
	.w5(32'hb993f3f9),
	.w6(32'hb8f1be89),
	.w7(32'hb9b5f6d9),
	.w8(32'hb9d5200c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393608cd),
	.w1(32'hb91e15a9),
	.w2(32'h36287d7d),
	.w3(32'h3836decd),
	.w4(32'h390d8c8b),
	.w5(32'hb90366aa),
	.w6(32'h3a3944a1),
	.w7(32'h3a235dff),
	.w8(32'h3a29008a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1199d1),
	.w1(32'hb830d113),
	.w2(32'h399a3ef8),
	.w3(32'h39a0a17d),
	.w4(32'h39e50d6e),
	.w5(32'h398ffb0e),
	.w6(32'h392c74e5),
	.w7(32'h39c9e120),
	.w8(32'h39210bab),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa99c95),
	.w1(32'hba5a0bd2),
	.w2(32'h3a883cef),
	.w3(32'hb9cd7cdc),
	.w4(32'hba9100cc),
	.w5(32'h3a46f4d0),
	.w6(32'h3a0caa7d),
	.w7(32'h3a787b59),
	.w8(32'h3a98c89a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2e351),
	.w1(32'h3838740a),
	.w2(32'hb99432b2),
	.w3(32'h39d4badb),
	.w4(32'h3895bfcd),
	.w5(32'hb9a1c919),
	.w6(32'h389c1b05),
	.w7(32'hb9099831),
	.w8(32'hb9b08766),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee90db),
	.w1(32'hbb28cbb8),
	.w2(32'h39de4def),
	.w3(32'hbaadd5b4),
	.w4(32'hbb28f8bd),
	.w5(32'h389228df),
	.w6(32'h393a2d76),
	.w7(32'h39f3b904),
	.w8(32'h3a799ffe),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29c03a),
	.w1(32'hbb85067f),
	.w2(32'hba9be75f),
	.w3(32'hbb41ee89),
	.w4(32'hbb790283),
	.w5(32'hbac07c83),
	.w6(32'hba9cb06f),
	.w7(32'hbb051477),
	.w8(32'hba317ea2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16739d),
	.w1(32'hbacd898d),
	.w2(32'hba6834dd),
	.w3(32'h39210c00),
	.w4(32'hba42ae2e),
	.w5(32'hba07c9c7),
	.w6(32'h3a030bfd),
	.w7(32'h39370f3c),
	.w8(32'h381c5033),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2536e6),
	.w1(32'h39253a04),
	.w2(32'hbab60e2f),
	.w3(32'h39e474eb),
	.w4(32'h3821cf3e),
	.w5(32'hba993b08),
	.w6(32'hb91a6f95),
	.w7(32'hba2e6ef0),
	.w8(32'hba987fa1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad07e01),
	.w1(32'hba954000),
	.w2(32'h3a242d78),
	.w3(32'h39fe546d),
	.w4(32'h39dc8ca7),
	.w5(32'h3a9e0427),
	.w6(32'h399ca146),
	.w7(32'h380571d8),
	.w8(32'h3a602011),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23b52d),
	.w1(32'h39c5011b),
	.w2(32'hb9184cfa),
	.w3(32'h3b17770c),
	.w4(32'h3b01b1fb),
	.w5(32'h3a44877c),
	.w6(32'h3a855c66),
	.w7(32'h3a21e7e3),
	.w8(32'h35ee2070),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb53b0),
	.w1(32'hba617c88),
	.w2(32'hba7c6a71),
	.w3(32'h3ac4c4a5),
	.w4(32'h3a849b98),
	.w5(32'h39872a45),
	.w6(32'h3aced8d3),
	.w7(32'h3a1f5c77),
	.w8(32'h35ee9e68),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c54415),
	.w1(32'h3875abcf),
	.w2(32'hbaa294f2),
	.w3(32'h3aaf4699),
	.w4(32'h3994574d),
	.w5(32'hbac02220),
	.w6(32'h39d5c9a6),
	.w7(32'hb9f97612),
	.w8(32'hbaf4f77a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c16095),
	.w1(32'h38e2b543),
	.w2(32'h3958f3ff),
	.w3(32'hb8a37a0b),
	.w4(32'hb8104c55),
	.w5(32'h38e517e0),
	.w6(32'hb8ae5b9e),
	.w7(32'hb91e1f9c),
	.w8(32'h38a7b802),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73eeca2),
	.w1(32'hb90518af),
	.w2(32'h38dfc2e4),
	.w3(32'hb96464d5),
	.w4(32'hb98ed0c0),
	.w5(32'hb870add8),
	.w6(32'hb8eb53c7),
	.w7(32'hb88bd341),
	.w8(32'hb75b79e2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63ad6f),
	.w1(32'hbaa67e07),
	.w2(32'hbaa16f24),
	.w3(32'hba7b0aec),
	.w4(32'hba721cf6),
	.w5(32'hba8848ae),
	.w6(32'hba88a2e1),
	.w7(32'hba783ddc),
	.w8(32'hbaae8d5b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ff8305),
	.w1(32'hb9a67fd0),
	.w2(32'hba9f7288),
	.w3(32'h3a4664f3),
	.w4(32'h3a17d1a4),
	.w5(32'hba208138),
	.w6(32'h38f2ebb9),
	.w7(32'hb80428b3),
	.w8(32'hba350271),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae4be1),
	.w1(32'hb8efcac2),
	.w2(32'hb9971091),
	.w3(32'h3987ea5b),
	.w4(32'h39392719),
	.w5(32'hb8e451cf),
	.w6(32'h39c97c5c),
	.w7(32'h39b15f7e),
	.w8(32'h385518c7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36de784c),
	.w1(32'h36efbf47),
	.w2(32'h371ec789),
	.w3(32'hb6c69dee),
	.w4(32'hb6ab09ad),
	.w5(32'hb60e344e),
	.w6(32'hb749eb4c),
	.w7(32'hb77ec6a6),
	.w8(32'hb6f3262b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36395bc0),
	.w1(32'hb7c6a0af),
	.w2(32'hb7a4efb5),
	.w3(32'hb7ff14a7),
	.w4(32'hb7ff9056),
	.w5(32'hb7e4652e),
	.w6(32'hb71360f5),
	.w7(32'hb7903812),
	.w8(32'hb75cd891),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911d103),
	.w1(32'hb9cb74ee),
	.w2(32'hb96b5751),
	.w3(32'hba024944),
	.w4(32'hba73e358),
	.w5(32'hba8ace5a),
	.w6(32'hbac4f9c4),
	.w7(32'hba948244),
	.w8(32'hba6e737c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2818db),
	.w1(32'hbb12b73b),
	.w2(32'hbaa6a930),
	.w3(32'h3901d8ab),
	.w4(32'h3a7885fa),
	.w5(32'h3ab27188),
	.w6(32'hb923e7fd),
	.w7(32'hba4ee93d),
	.w8(32'hba183cec),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9853ddf),
	.w1(32'h385b3628),
	.w2(32'hb8bc24fe),
	.w3(32'hb93a6fab),
	.w4(32'h390ccc8c),
	.w5(32'h38c6ec07),
	.w6(32'hb9690f50),
	.w7(32'hb97f349a),
	.w8(32'hb9753bed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55d9b9),
	.w1(32'h3a0eb8f3),
	.w2(32'hbad1ee34),
	.w3(32'hb8122e39),
	.w4(32'hb9ec86eb),
	.w5(32'hbb1ae19c),
	.w6(32'hba0f4b31),
	.w7(32'hba953489),
	.w8(32'hbb1305ff),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f5995),
	.w1(32'h3af07f95),
	.w2(32'h3a26e396),
	.w3(32'h3af0b031),
	.w4(32'h3afb174c),
	.w5(32'h39e35016),
	.w6(32'h3ab7edbd),
	.w7(32'h3aaefb6e),
	.w8(32'h392290f9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913270b),
	.w1(32'h3a958ff2),
	.w2(32'h3aaa6735),
	.w3(32'hb8467de9),
	.w4(32'h3881e5cd),
	.w5(32'h3a174191),
	.w6(32'hb848d05f),
	.w7(32'hb90bbcdd),
	.w8(32'h394eebff),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63241f),
	.w1(32'h38c426bf),
	.w2(32'h38ee44f1),
	.w3(32'hb94861d9),
	.w4(32'hb8949189),
	.w5(32'hb766f6d5),
	.w6(32'h3885ffce),
	.w7(32'hba120923),
	.w8(32'h37e5548a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9895766),
	.w1(32'hb9c916d5),
	.w2(32'hba51ab43),
	.w3(32'hb9e265bb),
	.w4(32'hb9a944b3),
	.w5(32'hba4d6249),
	.w6(32'hb9885c3e),
	.w7(32'hb98b1d4d),
	.w8(32'hb9efd1db),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule