module layer_10_featuremap_10(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f2cc),
	.w1(32'h3c560439),
	.w2(32'hbb777b5a),
	.w3(32'h3b9e1217),
	.w4(32'h3b719ce6),
	.w5(32'hbc00826d),
	.w6(32'hbbf5cd1e),
	.w7(32'hbaf890c5),
	.w8(32'hba05dea7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd62281),
	.w1(32'h3b8c4962),
	.w2(32'hbb0ad6a0),
	.w3(32'h3aea8b99),
	.w4(32'h3bf18f4e),
	.w5(32'hbb169622),
	.w6(32'h3aa845eb),
	.w7(32'hbaa6b1ed),
	.w8(32'hba98d7a6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b608708),
	.w1(32'h38f50b76),
	.w2(32'hbc2ad64b),
	.w3(32'h3b874491),
	.w4(32'h3a827641),
	.w5(32'hbc4acd78),
	.w6(32'h3bf990f7),
	.w7(32'h3c4a0dba),
	.w8(32'hbbf5b9d6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb2f53),
	.w1(32'h3a18c50e),
	.w2(32'hbb2673b0),
	.w3(32'hbc33d7c1),
	.w4(32'hbc03f1a4),
	.w5(32'hbb18564a),
	.w6(32'hbbf3f958),
	.w7(32'hbc24c830),
	.w8(32'hbc036424),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab42a3),
	.w1(32'h3b6b2dea),
	.w2(32'hbbbae016),
	.w3(32'hbb2a5296),
	.w4(32'hbb8355fc),
	.w5(32'hbc18348e),
	.w6(32'hbbd5e45f),
	.w7(32'hbb73ac90),
	.w8(32'hbc1e3b0d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6190ca),
	.w1(32'hbb2d5226),
	.w2(32'hbbe0e888),
	.w3(32'hbbd9a541),
	.w4(32'hbb7b3352),
	.w5(32'h3c8aca84),
	.w6(32'hbc029796),
	.w7(32'h3a39ded4),
	.w8(32'h3d317b42),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd595c29),
	.w1(32'hbd3e6ccc),
	.w2(32'h3c64f131),
	.w3(32'hbb7a9185),
	.w4(32'hbcdbd01f),
	.w5(32'h3bf138d6),
	.w6(32'h3d85db42),
	.w7(32'h3ce2d3ff),
	.w8(32'h3b0b30aa),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc58c2a),
	.w1(32'h3c6f8ede),
	.w2(32'h3c4e4ae2),
	.w3(32'h3c6f992d),
	.w4(32'h3c014b04),
	.w5(32'hbb9bd21b),
	.w6(32'hb9a7514f),
	.w7(32'hba30e89c),
	.w8(32'h3bcbca16),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c913f09),
	.w1(32'h3c460835),
	.w2(32'h3b910c78),
	.w3(32'h3af9c09f),
	.w4(32'h3a8737c6),
	.w5(32'h3bd76431),
	.w6(32'hbbea2129),
	.w7(32'hbadf9dc7),
	.w8(32'h3b4ce784),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cd6e7),
	.w1(32'hbb5affb6),
	.w2(32'h3c50c9ab),
	.w3(32'h3b97abe6),
	.w4(32'h390b592b),
	.w5(32'h3a994337),
	.w6(32'h3c558f7e),
	.w7(32'h3c19923e),
	.w8(32'hbca0ab98),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d31aad3),
	.w1(32'h3cd9a9ac),
	.w2(32'hbb64c011),
	.w3(32'h3c50a050),
	.w4(32'h3c528788),
	.w5(32'hbc12eadc),
	.w6(32'hbd1188e5),
	.w7(32'hbca90b26),
	.w8(32'hbb15761d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace7ca8),
	.w1(32'hbc0115f2),
	.w2(32'hbb0ba175),
	.w3(32'hbbbd0c49),
	.w4(32'hba8ef7de),
	.w5(32'h3b87fb94),
	.w6(32'hbbc1d540),
	.w7(32'hbc00fe4e),
	.w8(32'h3c72b36c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c288c),
	.w1(32'hbc06f8b9),
	.w2(32'hbbac7fec),
	.w3(32'hbb02c66c),
	.w4(32'hbb836588),
	.w5(32'hbc07c140),
	.w6(32'h3cbe9af2),
	.w7(32'h3c7e4498),
	.w8(32'hbbcbcfd5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ba21),
	.w1(32'h3a86cfed),
	.w2(32'hbbe52990),
	.w3(32'h3b09df65),
	.w4(32'hba3a1c7c),
	.w5(32'h3b08ed52),
	.w6(32'hbb4641b8),
	.w7(32'hbad7b2fa),
	.w8(32'hbc04318b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7b9ab),
	.w1(32'hbb43eb85),
	.w2(32'h3a960b1a),
	.w3(32'hba5c80b7),
	.w4(32'h3aeac41a),
	.w5(32'hbaaa5d0a),
	.w6(32'hbbdd2634),
	.w7(32'hbb99f383),
	.w8(32'h3a003c7a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c328204),
	.w1(32'h3bed1d26),
	.w2(32'h3c0203e5),
	.w3(32'h3bd8413e),
	.w4(32'h3bab8c7d),
	.w5(32'h3bbe43da),
	.w6(32'h3b05a184),
	.w7(32'h3bce4bf2),
	.w8(32'hbb9c3aef),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd92ac5),
	.w1(32'h3c5799dc),
	.w2(32'h3b93e405),
	.w3(32'h3c492afe),
	.w4(32'h3be1f57f),
	.w5(32'h3a75a68a),
	.w6(32'hbc7b0c5c),
	.w7(32'hbc2dc43f),
	.w8(32'h3c1d9165),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972e4ab),
	.w1(32'hbaaefb87),
	.w2(32'h3b880496),
	.w3(32'h3a513434),
	.w4(32'hba9d5400),
	.w5(32'h3b2187f9),
	.w6(32'h3bb6cab7),
	.w7(32'h3b077d2f),
	.w8(32'hbae6ef2d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812697),
	.w1(32'hbbb4025d),
	.w2(32'h3a62a5c4),
	.w3(32'hbaaf5c99),
	.w4(32'hb9907c90),
	.w5(32'hbb6f5c44),
	.w6(32'h39a26800),
	.w7(32'hbb282481),
	.w8(32'hb94fce86),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf439bf),
	.w1(32'h3763847a),
	.w2(32'hb9f1cf40),
	.w3(32'hbbe02594),
	.w4(32'hbba89871),
	.w5(32'hbb4e3fe4),
	.w6(32'hbc3caa2d),
	.w7(32'hbbfb5cd1),
	.w8(32'hbb290d5c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac41cf8),
	.w1(32'hb9ec7723),
	.w2(32'hbbcd459b),
	.w3(32'hbb4eafb0),
	.w4(32'hbb062849),
	.w5(32'hbb4011c6),
	.w6(32'hbb0def03),
	.w7(32'hba95f2c9),
	.w8(32'h3a8eb021),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ce43),
	.w1(32'h3b8572a7),
	.w2(32'h3b99d0e3),
	.w3(32'hbb197cb4),
	.w4(32'h3b9e5efd),
	.w5(32'h3c109c50),
	.w6(32'h3b15e324),
	.w7(32'hbb5a2cae),
	.w8(32'hbb9540ca),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e74ed),
	.w1(32'h3c7523c9),
	.w2(32'h3bff9bb2),
	.w3(32'h3bc4a223),
	.w4(32'h3c1bf6d1),
	.w5(32'hbbfc279b),
	.w6(32'hbbf61ec5),
	.w7(32'hbb84e486),
	.w8(32'hbcc7249b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3c083f),
	.w1(32'h3d00265d),
	.w2(32'h3b3196a3),
	.w3(32'h3bc081a4),
	.w4(32'h3c8d08f3),
	.w5(32'hbad73a06),
	.w6(32'hbd292158),
	.w7(32'hbc9aa51b),
	.w8(32'hbb33fff5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27db81),
	.w1(32'hbb9bcb62),
	.w2(32'hbb95ff81),
	.w3(32'hbaf48903),
	.w4(32'hbb43377c),
	.w5(32'h395086e6),
	.w6(32'hb9e462b7),
	.w7(32'h3af4c964),
	.w8(32'hbb0c956f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3357f),
	.w1(32'hba87faca),
	.w2(32'h3856c5ef),
	.w3(32'h39c288b7),
	.w4(32'hbb948b2d),
	.w5(32'hbbc6c8e0),
	.w6(32'hbb094564),
	.w7(32'hbbd7329a),
	.w8(32'hbc14b90f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83dd7b),
	.w1(32'hbb3286c9),
	.w2(32'hb53d1008),
	.w3(32'hbbf3fcbc),
	.w4(32'hbbc07ea6),
	.w5(32'h33ca1ca3),
	.w6(32'hbbd11b4e),
	.w7(32'hbb3007eb),
	.w8(32'h351c65a1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38275cc8),
	.w1(32'hb92a045f),
	.w2(32'hb8baabdd),
	.w3(32'h390a9141),
	.w4(32'hb8f2c658),
	.w5(32'hb76e159d),
	.w6(32'h3905e4c5),
	.w7(32'hb8cdceb1),
	.w8(32'hb7f78c67),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a354b2),
	.w1(32'hb55ca960),
	.w2(32'hb72b6647),
	.w3(32'h376693e5),
	.w4(32'h36a4b322),
	.w5(32'h346c1071),
	.w6(32'hb67181ba),
	.w7(32'h3737db6b),
	.w8(32'h378c744f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b87cf),
	.w1(32'hb93c4fae),
	.w2(32'hb8b8fd01),
	.w3(32'h39047a00),
	.w4(32'hb94c1df1),
	.w5(32'hb917b528),
	.w6(32'h3915b3ef),
	.w7(32'hb9286374),
	.w8(32'hb8e0f6a7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3502b2bc),
	.w1(32'h3583307a),
	.w2(32'hb5adbc07),
	.w3(32'h3683825f),
	.w4(32'h36994444),
	.w5(32'h3621da40),
	.w6(32'h35f766a1),
	.w7(32'h36660aa6),
	.w8(32'hb5f3a167),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e0954d),
	.w1(32'hb520d613),
	.w2(32'hb65de828),
	.w3(32'hb61ce508),
	.w4(32'hb63de854),
	.w5(32'hb699083b),
	.w6(32'hb7030ccb),
	.w7(32'hb6259673),
	.w8(32'h36d2a92e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a19fd5),
	.w1(32'h36a45c4b),
	.w2(32'hb7ab562d),
	.w3(32'h38889111),
	.w4(32'h36af05c0),
	.w5(32'hb783e12d),
	.w6(32'h37cabc56),
	.w7(32'hb80792df),
	.w8(32'hb7cc1a59),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3781771f),
	.w1(32'hb7627833),
	.w2(32'hb7f07a5c),
	.w3(32'h37b6c7ee),
	.w4(32'hb8097446),
	.w5(32'hb85160b6),
	.w6(32'h37d93350),
	.w7(32'hb7bda138),
	.w8(32'hb835b00b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f5a105),
	.w1(32'hb611e768),
	.w2(32'hb73803be),
	.w3(32'h373a8db5),
	.w4(32'h37b211e6),
	.w5(32'hb5f1fab5),
	.w6(32'h370b368f),
	.w7(32'h36db4b65),
	.w8(32'hb6ca0d00),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38935710),
	.w1(32'h38396dd5),
	.w2(32'h377bbce9),
	.w3(32'h3804d676),
	.w4(32'h38260d79),
	.w5(32'hb70b02bb),
	.w6(32'hb8231041),
	.w7(32'hb7a6b7f6),
	.w8(32'hb7d4eeae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913af8d),
	.w1(32'h396607be),
	.w2(32'h393192fc),
	.w3(32'hb8ed962a),
	.w4(32'h3897fd28),
	.w5(32'h3842f128),
	.w6(32'hb92ea72d),
	.w7(32'hb82d716f),
	.w8(32'hb904f48b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb668e052),
	.w1(32'hb982c89d),
	.w2(32'hb91d6418),
	.w3(32'h39150f2d),
	.w4(32'hb98346e1),
	.w5(32'hb9805720),
	.w6(32'h39593d33),
	.w7(32'hb93ee477),
	.w8(32'hb981cb99),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938a4e7),
	.w1(32'hb9828085),
	.w2(32'hb97ac8e8),
	.w3(32'h39954110),
	.w4(32'hb96afcc3),
	.w5(32'hb98b6fa5),
	.w6(32'h394ec0ce),
	.w7(32'hb975c730),
	.w8(32'hb9a3306a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371c6f53),
	.w1(32'hb880d77c),
	.w2(32'hb7a9a1cc),
	.w3(32'h37dfc71a),
	.w4(32'hb8614043),
	.w5(32'hb7afa42a),
	.w6(32'h3794099d),
	.w7(32'hb82be7da),
	.w8(32'hb8027cf0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8015fc1),
	.w1(32'hb743bd6e),
	.w2(32'hb703b6df),
	.w3(32'hb8033b63),
	.w4(32'hb713b145),
	.w5(32'h360ff926),
	.w6(32'hb7369ceb),
	.w7(32'h36ed68f8),
	.w8(32'h36d15fd5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb752e32d),
	.w1(32'hb68ac301),
	.w2(32'hb73fb9db),
	.w3(32'hb656686a),
	.w4(32'h371535a2),
	.w5(32'hb6f7948d),
	.w6(32'h3612ac6e),
	.w7(32'h35d64074),
	.w8(32'hb71f4980),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8234e94),
	.w1(32'hb7c26aec),
	.w2(32'hb8222680),
	.w3(32'hb8542365),
	.w4(32'hb6f79ddd),
	.w5(32'hb72f4d32),
	.w6(32'hb862dc8c),
	.w7(32'hb83a5e53),
	.w8(32'hb7029e1c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391af80d),
	.w1(32'hb8439b81),
	.w2(32'h35d682cd),
	.w3(32'h38912a2a),
	.w4(32'hb7a7ff5e),
	.w5(32'hb80813a6),
	.w6(32'hb8210982),
	.w7(32'hb903c735),
	.w8(32'h372b37ec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b47fb),
	.w1(32'hb873e9f7),
	.w2(32'hb80944b4),
	.w3(32'h38dc6405),
	.w4(32'hb8dc561f),
	.w5(32'hb8780003),
	.w6(32'h38a0c2b7),
	.w7(32'hb8fc6242),
	.w8(32'hb89d0256),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39403734),
	.w1(32'hb84654d1),
	.w2(32'hb8714e0d),
	.w3(32'h3902e51d),
	.w4(32'hb8f8a1cf),
	.w5(32'hb8b67276),
	.w6(32'h382279a7),
	.w7(32'hb91401e1),
	.w8(32'hb900e615),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807755d),
	.w1(32'hb721545e),
	.w2(32'h37f9fbd2),
	.w3(32'hb61cd63d),
	.w4(32'hb8a6b287),
	.w5(32'hb68710d5),
	.w6(32'hb7f57f7a),
	.w7(32'hb8e6dcf9),
	.w8(32'hb8527485),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39406a57),
	.w1(32'h39400eef),
	.w2(32'h39a18634),
	.w3(32'hb7e36231),
	.w4(32'h3924bbf0),
	.w5(32'h3922a2ba),
	.w6(32'hb9649cbd),
	.w7(32'hb8f303a3),
	.w8(32'h3915924b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76cb93a),
	.w1(32'hb6cea13e),
	.w2(32'h36a7669c),
	.w3(32'hb75e89b3),
	.w4(32'hb6583db8),
	.w5(32'hb6a57430),
	.w6(32'h359c186b),
	.w7(32'h3703bad1),
	.w8(32'h369efde2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7439875),
	.w1(32'hb70e21b6),
	.w2(32'hb793e468),
	.w3(32'hb84f6449),
	.w4(32'hb8313c16),
	.w5(32'hb7f09cd7),
	.w6(32'hb6a77640),
	.w7(32'hb6dae3c5),
	.w8(32'hb76ed12f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7958fe5),
	.w1(32'hb7774376),
	.w2(32'hb76e541d),
	.w3(32'hb6a796d1),
	.w4(32'hb4f3060d),
	.w5(32'hb7abccc9),
	.w6(32'hb7de2268),
	.w7(32'hb7686a99),
	.w8(32'hb6e6ae01),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3c4dc),
	.w1(32'h36c05998),
	.w2(32'hb7690347),
	.w3(32'h38e404bd),
	.w4(32'hb632353f),
	.w5(32'hb7e6c9d7),
	.w6(32'h382038ea),
	.w7(32'hb85788f5),
	.w8(32'hb80bb63b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e38275),
	.w1(32'h372ad559),
	.w2(32'h3736e3ac),
	.w3(32'h378ac07a),
	.w4(32'h36362bce),
	.w5(32'h3560d12a),
	.w6(32'hb7357c82),
	.w7(32'hb7739c0e),
	.w8(32'hb717ea5f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39369850),
	.w1(32'h38e31ceb),
	.w2(32'h391aa139),
	.w3(32'h38a5bee9),
	.w4(32'h3907e205),
	.w5(32'h38a263e9),
	.w6(32'hb89f8110),
	.w7(32'hb8d67836),
	.w8(32'h379bdcbb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c66a10),
	.w1(32'h37483e27),
	.w2(32'h37c75820),
	.w3(32'h3817db27),
	.w4(32'h37c61a31),
	.w5(32'h37f55906),
	.w6(32'h35b724e6),
	.w7(32'hb7161376),
	.w8(32'h37d070e1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36387742),
	.w1(32'hb62d4a61),
	.w2(32'hb6afe78d),
	.w3(32'hb71a1bf6),
	.w4(32'hb7461ebe),
	.w5(32'hb7063154),
	.w6(32'hb60faaf6),
	.w7(32'hb56ccd9d),
	.w8(32'h36372913),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f588e1),
	.w1(32'h3738aae2),
	.w2(32'hb59e7a8e),
	.w3(32'hb75604f0),
	.w4(32'hb6548d88),
	.w5(32'h3687120d),
	.w6(32'hb63ca591),
	.w7(32'hb60e204d),
	.w8(32'h35c9bb96),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371a2875),
	.w1(32'hb7159435),
	.w2(32'hb62d18e3),
	.w3(32'h379a6d22),
	.w4(32'h36897193),
	.w5(32'hb6b4384f),
	.w6(32'h379a275a),
	.w7(32'h36c56e83),
	.w8(32'h36a28b8f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79be652),
	.w1(32'h36cd6ed3),
	.w2(32'hb6fddf85),
	.w3(32'hb786174c),
	.w4(32'h359ea28a),
	.w5(32'hb6e9be46),
	.w6(32'hb665033b),
	.w7(32'hb6450f66),
	.w8(32'hb7315e75),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a821e),
	.w1(32'hb6a29551),
	.w2(32'hb79579eb),
	.w3(32'hb5d3fbfb),
	.w4(32'h37397db7),
	.w5(32'hb77141d1),
	.w6(32'hb6e84a5b),
	.w7(32'hb76e78cd),
	.w8(32'hb73faf29),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8d0fa),
	.w1(32'h386fe0f5),
	.w2(32'h38a223b8),
	.w3(32'h385f0d4d),
	.w4(32'h3890318e),
	.w5(32'h37cb485b),
	.w6(32'hb7ba7654),
	.w7(32'h37f8a313),
	.w8(32'h388fc8aa),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6870ec5),
	.w1(32'hb7c91356),
	.w2(32'h37969ca7),
	.w3(32'hb7a78abf),
	.w4(32'hb8812efd),
	.w5(32'h379cfdfe),
	.w6(32'hb82c6a86),
	.w7(32'hb8275989),
	.w8(32'h38cd8209),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69b208f),
	.w1(32'h372156a6),
	.w2(32'h35d41cba),
	.w3(32'hb6cafb64),
	.w4(32'hb4fccfb9),
	.w5(32'h364a9af4),
	.w6(32'h359b8d35),
	.w7(32'h369e466d),
	.w8(32'h36430b04),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3385b6b0),
	.w1(32'hb5fd1b78),
	.w2(32'hb4d3f915),
	.w3(32'h367820f6),
	.w4(32'hb5bc22b1),
	.w5(32'h36a6e6e7),
	.w6(32'hb52dbeee),
	.w7(32'hb69badb4),
	.w8(32'h351fc4ad),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c79408),
	.w1(32'hb67a9dcc),
	.w2(32'hb68864a3),
	.w3(32'hb681b382),
	.w4(32'h35378dfd),
	.w5(32'h356d785c),
	.w6(32'h340f4219),
	.w7(32'hb202e45c),
	.w8(32'hb60a3ee0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60d1981),
	.w1(32'hb6621817),
	.w2(32'h370541d2),
	.w3(32'hb49ff4ab),
	.w4(32'hb5bb7950),
	.w5(32'h370bc860),
	.w6(32'hb49b44aa),
	.w7(32'hb4fbf77f),
	.w8(32'h3715c591),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39275b78),
	.w1(32'h38bd16d5),
	.w2(32'h36cda37c),
	.w3(32'h391de215),
	.w4(32'h3830fa91),
	.w5(32'h3741bb86),
	.w6(32'h37ee3c6f),
	.w7(32'hb89ad78e),
	.w8(32'hb889b5f9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992182d),
	.w1(32'h37a064e6),
	.w2(32'hb87d7563),
	.w3(32'h395e1d0f),
	.w4(32'h369dbd57),
	.w5(32'hb8334132),
	.w6(32'h381bafa2),
	.w7(32'hb901ab20),
	.w8(32'hb8e24338),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930abb4),
	.w1(32'h38c7ef0d),
	.w2(32'h384b0c15),
	.w3(32'h394b41fa),
	.w4(32'h38752b10),
	.w5(32'h382e1af4),
	.w6(32'h3751eb07),
	.w7(32'hb7562a36),
	.w8(32'h3856823d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397336cd),
	.w1(32'hb92aab70),
	.w2(32'hb8c6425d),
	.w3(32'h397733e9),
	.w4(32'hb974f865),
	.w5(32'hb9662222),
	.w6(32'h3981762c),
	.w7(32'hb93f4770),
	.w8(32'hb95b9b82),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61f94ec),
	.w1(32'h36ba1bcd),
	.w2(32'hb688726d),
	.w3(32'hb6887801),
	.w4(32'h37194fcd),
	.w5(32'hb6838a75),
	.w6(32'h352e6f1d),
	.w7(32'h370e9f41),
	.w8(32'hb65aece9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6202d15),
	.w1(32'hb708e57f),
	.w2(32'hb6a886bf),
	.w3(32'hb5a0cbd1),
	.w4(32'hb7334ad9),
	.w5(32'hb70cea02),
	.w6(32'h35bf450a),
	.w7(32'hb6c2570a),
	.w8(32'hb68a0d34),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb009674a),
	.w1(32'h34cb026e),
	.w2(32'h36733e74),
	.w3(32'hb5edc0e6),
	.w4(32'hb5b31773),
	.w5(32'h3726053b),
	.w6(32'h368613f3),
	.w7(32'h346c9c1c),
	.w8(32'h363e634c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829f105),
	.w1(32'h37dcde31),
	.w2(32'h37d76013),
	.w3(32'h38197fdd),
	.w4(32'h38230b95),
	.w5(32'h3818cfcf),
	.w6(32'hb720e4ec),
	.w7(32'h35e8e0d0),
	.w8(32'h380feb4a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3333c568),
	.w1(32'hb4ad26ab),
	.w2(32'hb720f0cc),
	.w3(32'hb4992a2e),
	.w4(32'hb6a9efbc),
	.w5(32'hb71bc4f9),
	.w6(32'h3698fa6c),
	.w7(32'h365e8993),
	.w8(32'h35fca586),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390970b3),
	.w1(32'h38f7671d),
	.w2(32'h38ca6ae2),
	.w3(32'h38377967),
	.w4(32'h38d24c35),
	.w5(32'h38150323),
	.w6(32'hb7824d82),
	.w7(32'hb6ae274e),
	.w8(32'hb7d95a38),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ff56e),
	.w1(32'h391ba712),
	.w2(32'h395bbb6d),
	.w3(32'h37a70027),
	.w4(32'h38fc0290),
	.w5(32'h39092e2b),
	.w6(32'hb7a585cc),
	.w7(32'h379863d0),
	.w8(32'hb79bce9a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927e797),
	.w1(32'hb7db6c67),
	.w2(32'h37b17710),
	.w3(32'h390a8335),
	.w4(32'hb823af2d),
	.w5(32'hb7bd8749),
	.w6(32'h385706be),
	.w7(32'hb8b37978),
	.w8(32'hb868b803),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7b457),
	.w1(32'h37b50090),
	.w2(32'hb67a373c),
	.w3(32'h38eba2d8),
	.w4(32'h36bb56ad),
	.w5(32'hb707f510),
	.w6(32'h3848db60),
	.w7(32'hb7baa06c),
	.w8(32'hb72324d8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894d108),
	.w1(32'h35b99eb6),
	.w2(32'hb7c0ae78),
	.w3(32'h38d1c9dd),
	.w4(32'h37e8504a),
	.w5(32'hb7772120),
	.w6(32'h3852804b),
	.w7(32'hb7c9892f),
	.w8(32'hb8443bd7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f8a5d8),
	.w1(32'hb7b605cc),
	.w2(32'hb7802897),
	.w3(32'h37f7e13c),
	.w4(32'hb807b832),
	.w5(32'hb7798c51),
	.w6(32'h37c8278a),
	.w7(32'hb808693a),
	.w8(32'hb742fca8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6bd60),
	.w1(32'h38ab4024),
	.w2(32'h38b9ddee),
	.w3(32'h389c9228),
	.w4(32'h389b11cd),
	.w5(32'h386e6af9),
	.w6(32'hb7998c4e),
	.w7(32'hb7fd0d0a),
	.w8(32'h380a7dc3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5dd91d0),
	.w1(32'hb6174847),
	.w2(32'h365e5723),
	.w3(32'hb6395967),
	.w4(32'hb6a0e7d6),
	.w5(32'h36b3edb1),
	.w6(32'h34b02d8b),
	.w7(32'hb6592174),
	.w8(32'h372edaac),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb650f425),
	.w1(32'hb69db24d),
	.w2(32'h3698d970),
	.w3(32'hb727ce8d),
	.w4(32'hb72ef742),
	.w5(32'hb721d62e),
	.w6(32'h36426fd0),
	.w7(32'h339252da),
	.w8(32'hb586f245),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4e8a9da),
	.w1(32'h371181a3),
	.w2(32'hb5dafb6c),
	.w3(32'hb5f53a76),
	.w4(32'hb6f5f8c2),
	.w5(32'h35bbf0e2),
	.w6(32'hb6d23eec),
	.w7(32'h31c6030b),
	.w8(32'hb658073a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ef9207),
	.w1(32'hb799f3ad),
	.w2(32'hb7699606),
	.w3(32'h371ef66b),
	.w4(32'hb78affd6),
	.w5(32'hb75616d9),
	.w6(32'h36caf9c4),
	.w7(32'hb774dc52),
	.w8(32'hb77f4545),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a37ab4),
	.w1(32'hb890c87e),
	.w2(32'hb7243f4f),
	.w3(32'h37843055),
	.w4(32'hb87d7623),
	.w5(32'hb848f4fe),
	.w6(32'h3823d708),
	.w7(32'hb85b02d8),
	.w8(32'hb8aa9940),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb660380d),
	.w1(32'h36f796dc),
	.w2(32'h3691fa58),
	.w3(32'hb68a1d99),
	.w4(32'h361dbd55),
	.w5(32'hb6d61a55),
	.w6(32'hb7101dee),
	.w7(32'hb6eec704),
	.w8(32'hb704d22f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381c3a50),
	.w1(32'hb786a9a6),
	.w2(32'h3794099e),
	.w3(32'h37b77755),
	.w4(32'hb8011bd3),
	.w5(32'h3754feef),
	.w6(32'hb6f4c848),
	.w7(32'hb87acc14),
	.w8(32'hb598528d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943df7f),
	.w1(32'h38f8d77f),
	.w2(32'h391eb06c),
	.w3(32'h38cf4c25),
	.w4(32'h389b9342),
	.w5(32'h38a83e4a),
	.w6(32'hb752ea01),
	.w7(32'hb8a5a2fb),
	.w8(32'h38aa472c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381957e8),
	.w1(32'hb8bb5083),
	.w2(32'hb7e33fc7),
	.w3(32'h3887c90e),
	.w4(32'hb8967a24),
	.w5(32'hb80ff38f),
	.w6(32'h374e3fd6),
	.w7(32'hb8ebdbd1),
	.w8(32'hb8b3caef),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f264f8),
	.w1(32'h39312d40),
	.w2(32'h38aeff59),
	.w3(32'h3912f83f),
	.w4(32'h38e7786c),
	.w5(32'h34a76a62),
	.w6(32'hb821a5a6),
	.w7(32'hb7a6179f),
	.w8(32'hb7c4435c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e39e3),
	.w1(32'hb89d9bd4),
	.w2(32'hb8df0b2b),
	.w3(32'h38d7d287),
	.w4(32'hb80a0b7b),
	.w5(32'hb8c94c51),
	.w6(32'h3893b49e),
	.w7(32'hb83a6b44),
	.w8(32'hb8b8b042),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39373337),
	.w1(32'h381237df),
	.w2(32'h36948434),
	.w3(32'h391ff535),
	.w4(32'hb71f738d),
	.w5(32'hb7315673),
	.w6(32'h38684f52),
	.w7(32'hb8a118fe),
	.w8(32'hb7981d15),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899d4f3),
	.w1(32'hb7812780),
	.w2(32'hb83c12c4),
	.w3(32'h38bc4f43),
	.w4(32'hb768d3e1),
	.w5(32'hb8ad595b),
	.w6(32'h38932b16),
	.w7(32'hb8774290),
	.w8(32'hb8955ee8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aaa2c6),
	.w1(32'hb8cc7d30),
	.w2(32'hb848e4b1),
	.w3(32'h39015442),
	.w4(32'hb8decc30),
	.w5(32'hb88b1fd8),
	.w6(32'h38907927),
	.w7(32'hb91277ba),
	.w8(32'hb909d3a8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bb86bc),
	.w1(32'hb6da75a4),
	.w2(32'h368d1c9a),
	.w3(32'hb84de8dc),
	.w4(32'hb7e03768),
	.w5(32'hb6e4a0fb),
	.w6(32'hb6b158c2),
	.w7(32'hb69536a6),
	.w8(32'hb5f929f3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dfe63b),
	.w1(32'h38512db4),
	.w2(32'h38882d3f),
	.w3(32'h371c9468),
	.w4(32'hb636c032),
	.w5(32'hb7cf9cf9),
	.w6(32'hb8a15817),
	.w7(32'hb917cd96),
	.w8(32'hb6924821),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d97c7),
	.w1(32'h38e117f3),
	.w2(32'hb7aa3eeb),
	.w3(32'h391d123e),
	.w4(32'h38a57cf1),
	.w5(32'hb8f1a717),
	.w6(32'h375f2a2c),
	.w7(32'hb8913ad4),
	.w8(32'hb8dd2bcf),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39717498),
	.w1(32'h39790f90),
	.w2(32'h39873778),
	.w3(32'hb88367ba),
	.w4(32'h393e5ed4),
	.w5(32'h3946415b),
	.w6(32'hb85074eb),
	.w7(32'hb88b43ef),
	.w8(32'hb411ec5e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eff222),
	.w1(32'hb9acde81),
	.w2(32'hb9a5dba6),
	.w3(32'hb8be0994),
	.w4(32'hb99d1eb8),
	.w5(32'hb9ba13dd),
	.w6(32'hb84d1c87),
	.w7(32'hb9942d1c),
	.w8(32'hb9c4dfe9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39238946),
	.w1(32'hb9561c27),
	.w2(32'hb8cf7a78),
	.w3(32'h38d6d828),
	.w4(32'hb995b9e3),
	.w5(32'hb94bb5f0),
	.w6(32'h3912f634),
	.w7(32'hb91efb0f),
	.w8(32'hb91757ea),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a8865),
	.w1(32'h39503543),
	.w2(32'h38e2dc00),
	.w3(32'h3860ce0c),
	.w4(32'h3931503e),
	.w5(32'h38d63136),
	.w6(32'hb8fce084),
	.w7(32'hb7a3ece6),
	.w8(32'h37eed7cc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8389b60),
	.w1(32'hb8933c4c),
	.w2(32'hb85d252a),
	.w3(32'hb4553799),
	.w4(32'hb8838825),
	.w5(32'hb89c8cc2),
	.w6(32'h35991b48),
	.w7(32'h3720ad14),
	.w8(32'hb8569ae1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994b641),
	.w1(32'h3983415a),
	.w2(32'h39d35e30),
	.w3(32'hb8864930),
	.w4(32'h3960aac5),
	.w5(32'h392d3619),
	.w6(32'h36da70c2),
	.w7(32'h38afd982),
	.w8(32'hb8f3b4b4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803e7ad),
	.w1(32'hb7977dbd),
	.w2(32'hb80f7d38),
	.w3(32'h37d75e3d),
	.w4(32'h379dfd36),
	.w5(32'hb806c47a),
	.w6(32'h37837510),
	.w7(32'h3774ed6e),
	.w8(32'hb8910b32),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37146ff0),
	.w1(32'hb6d3ac2b),
	.w2(32'hb7184f17),
	.w3(32'h3731afd6),
	.w4(32'hb708fe60),
	.w5(32'hb716c7dd),
	.w6(32'h36aedbca),
	.w7(32'hb70a2481),
	.w8(32'hb7093bd1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8e223),
	.w1(32'h380781ab),
	.w2(32'hb745a7fb),
	.w3(32'h380bc073),
	.w4(32'h36b775a0),
	.w5(32'hb79d9e0a),
	.w6(32'h37a5a6c8),
	.w7(32'hb630673c),
	.w8(32'hb810e250),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a46aed),
	.w1(32'hb8595d9d),
	.w2(32'hb887365d),
	.w3(32'h38d74623),
	.w4(32'hb85d0497),
	.w5(32'hb87b6eee),
	.w6(32'h377c313e),
	.w7(32'hb8de2735),
	.w8(32'hb86123c6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39008508),
	.w1(32'hb8943cfa),
	.w2(32'hb838d0ca),
	.w3(32'h388f32ad),
	.w4(32'hb9019272),
	.w5(32'hb8cdf93b),
	.w6(32'h38f95d73),
	.w7(32'hb89af77a),
	.w8(32'hb89ab12a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3856d784),
	.w1(32'hb823aae9),
	.w2(32'hb6c6019c),
	.w3(32'h381b5553),
	.w4(32'hb8a02477),
	.w5(32'h3696b327),
	.w6(32'hb776e450),
	.w7(32'hb88076c3),
	.w8(32'hb7f44c73),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388310ba),
	.w1(32'h3718ec7d),
	.w2(32'h35ea8b02),
	.w3(32'h360537bc),
	.w4(32'hb81ec387),
	.w5(32'hb5deb77a),
	.w6(32'hb724e3e4),
	.w7(32'hb860cabc),
	.w8(32'hb7e19bd6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797fb03),
	.w1(32'h3759032a),
	.w2(32'h38c48773),
	.w3(32'hb79b2afd),
	.w4(32'h371b3e0d),
	.w5(32'h38ed956d),
	.w6(32'hb826348c),
	.w7(32'hb80620d0),
	.w8(32'h3810f80c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2291a),
	.w1(32'h3876b90c),
	.w2(32'h37fa5ac6),
	.w3(32'h37a4f2e3),
	.w4(32'hb6a03ec3),
	.w5(32'h380744f5),
	.w6(32'hb7b6ca3b),
	.w7(32'hb837c541),
	.w8(32'h373a54df),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837611f),
	.w1(32'hb81c8269),
	.w2(32'hb7cf69ac),
	.w3(32'h37db1441),
	.w4(32'hb878ce2f),
	.w5(32'hb84c854e),
	.w6(32'h37b487b1),
	.w7(32'hb87a289d),
	.w8(32'hb8166bf5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb612ce9f),
	.w1(32'h368ace6d),
	.w2(32'h369977e0),
	.w3(32'hb630e99d),
	.w4(32'h362ec94c),
	.w5(32'h368e2ad9),
	.w6(32'hb3c3a391),
	.w7(32'h33afbccc),
	.w8(32'hb5679cec),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d5745a),
	.w1(32'hb5c96d45),
	.w2(32'h3645cad9),
	.w3(32'h34c506e4),
	.w4(32'h31280418),
	.w5(32'h3656558c),
	.w6(32'h36937651),
	.w7(32'h36c82e8b),
	.w8(32'h360c9820),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4af3f91),
	.w1(32'h35873d71),
	.w2(32'h350d6d28),
	.w3(32'h35bb92c4),
	.w4(32'h36079962),
	.w5(32'h36d31d38),
	.w6(32'hb6959830),
	.w7(32'hb6a38962),
	.w8(32'hb6f16c9d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368351f6),
	.w1(32'h36a4490c),
	.w2(32'hb66ccc20),
	.w3(32'h36e2196f),
	.w4(32'h36bc035a),
	.w5(32'h3536a55e),
	.w6(32'hb68d50d6),
	.w7(32'hb68e4090),
	.w8(32'h367b8333),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4c512),
	.w1(32'hb85f58cd),
	.w2(32'hb7dc7dc0),
	.w3(32'h38803932),
	.w4(32'hb87563e8),
	.w5(32'hb868562b),
	.w6(32'h37db7c3d),
	.w7(32'hb8970475),
	.w8(32'hb891db6a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4de81e9),
	.w1(32'h37289ac5),
	.w2(32'h374542f8),
	.w3(32'hb6f2d82b),
	.w4(32'h36903073),
	.w5(32'h3731e7f9),
	.w6(32'hb5049243),
	.w7(32'h378c13dc),
	.w8(32'h37174b77),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f4f1ad),
	.w1(32'h384a920d),
	.w2(32'h388018f0),
	.w3(32'h370f87e8),
	.w4(32'h3813eee0),
	.w5(32'h3826e111),
	.w6(32'hb8811efd),
	.w7(32'hb7b2d8ba),
	.w8(32'h37e2218f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e25b6e),
	.w1(32'hb8fb9c6c),
	.w2(32'hb87c3574),
	.w3(32'h38f44a81),
	.w4(32'hb90ab86e),
	.w5(32'hb8a25215),
	.w6(32'h38d0799c),
	.w7(32'hb90c6d23),
	.w8(32'hb8ed2541),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360a738d),
	.w1(32'hb681d33c),
	.w2(32'hb6f2e364),
	.w3(32'h371fe0a1),
	.w4(32'hb72e7f4f),
	.w5(32'hb70f4940),
	.w6(32'h361f9dec),
	.w7(32'hb705d872),
	.w8(32'hb70c5942),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ce1205),
	.w1(32'hb68da85b),
	.w2(32'h35b90980),
	.w3(32'hb6daaee4),
	.w4(32'hb6f84921),
	.w5(32'hb3e07a82),
	.w6(32'hb6e6a118),
	.w7(32'hb68e99bf),
	.w8(32'hb69170e8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e65963),
	.w1(32'hb62e2d04),
	.w2(32'hb695865e),
	.w3(32'hb62b5a8f),
	.w4(32'hb59bad9a),
	.w5(32'hb77ecae9),
	.w6(32'hb73c4399),
	.w7(32'h340c94d2),
	.w8(32'hb7265f29),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c7d9bc),
	.w1(32'hb7447933),
	.w2(32'hb6f14dde),
	.w3(32'hb7ec4c3a),
	.w4(32'hb7792eb6),
	.w5(32'hb6025bdb),
	.w6(32'hb7abf6e5),
	.w7(32'hb6aa8e6b),
	.w8(32'h33848604),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398116c5),
	.w1(32'h393f10be),
	.w2(32'h37860e0e),
	.w3(32'h392299dd),
	.w4(32'h39079dc3),
	.w5(32'hb700b938),
	.w6(32'hb7975278),
	.w7(32'h3893bf0f),
	.w8(32'h3680a08f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f46428),
	.w1(32'hb66ec914),
	.w2(32'h369b92fd),
	.w3(32'h38f59cb8),
	.w4(32'h380a3d18),
	.w5(32'h38260a80),
	.w6(32'h384b30a8),
	.w7(32'hb85e0e3b),
	.w8(32'h381e59e5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376925e1),
	.w1(32'h3717cdb6),
	.w2(32'h37efcedb),
	.w3(32'h359ca414),
	.w4(32'h3788b2db),
	.w5(32'h380ce761),
	.w6(32'h362eac74),
	.w7(32'h356bef74),
	.w8(32'h37eb05a3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377bd085),
	.w1(32'h36b79e57),
	.w2(32'h32a28941),
	.w3(32'h374ea61c),
	.w4(32'h351a015e),
	.w5(32'hb6da89e2),
	.w6(32'h37ca7809),
	.w7(32'h378f1380),
	.w8(32'hb783f2f6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380df118),
	.w1(32'hb782bbba),
	.w2(32'h34858178),
	.w3(32'h37fdec18),
	.w4(32'hb8060825),
	.w5(32'hb72305ec),
	.w6(32'h36ab0d7d),
	.w7(32'hb841f787),
	.w8(32'hb7d5bea5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38763a95),
	.w1(32'hb5f33319),
	.w2(32'h36a6955f),
	.w3(32'h381a0078),
	.w4(32'hb8054b06),
	.w5(32'h368da2b1),
	.w6(32'h37a27be0),
	.w7(32'hb81e3bf6),
	.w8(32'h3680e3ca),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7e7cc),
	.w1(32'hb7c09d56),
	.w2(32'h3664cf1e),
	.w3(32'h38f56087),
	.w4(32'hb874ad4f),
	.w5(32'hb7c891c3),
	.w6(32'h38d375d7),
	.w7(32'hb88a223e),
	.w8(32'hb7fda7a0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b1a58),
	.w1(32'h3927356d),
	.w2(32'h39593e3a),
	.w3(32'h390ac429),
	.w4(32'h3950db2f),
	.w5(32'h375babc7),
	.w6(32'hb78c8609),
	.w7(32'hb8bb4cc0),
	.w8(32'h376e2d40),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372f964f),
	.w1(32'hb8b2bc0c),
	.w2(32'hb7f0f4f2),
	.w3(32'h37874f43),
	.w4(32'hb8af56e1),
	.w5(32'hb81b874a),
	.w6(32'h36baaf1e),
	.w7(32'hb8d99ba9),
	.w8(32'hb8956286),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38942f51),
	.w1(32'h384911cd),
	.w2(32'h385140be),
	.w3(32'h3839cbc4),
	.w4(32'h3776b0b6),
	.w5(32'h36c6c8eb),
	.w6(32'hb612df09),
	.w7(32'hb7370d12),
	.w8(32'h3800ee49),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38917a09),
	.w1(32'h38b6651a),
	.w2(32'h39084de4),
	.w3(32'h36f20e7f),
	.w4(32'h38800d06),
	.w5(32'h3708c5e8),
	.w6(32'hb88a60d6),
	.w7(32'hb9155f65),
	.w8(32'h38a6fa33),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381d5f97),
	.w1(32'h35753e4a),
	.w2(32'h38344d78),
	.w3(32'h37c35c93),
	.w4(32'hb7fab61e),
	.w5(32'h3711ba3b),
	.w6(32'hb65fd136),
	.w7(32'hb833c157),
	.w8(32'hb73e3992),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f7b1a),
	.w1(32'h3704378d),
	.w2(32'h3718ec01),
	.w3(32'h381f9662),
	.w4(32'h37cfc3f3),
	.w5(32'hb68ed5cb),
	.w6(32'h37356c14),
	.w7(32'hb8119d95),
	.w8(32'hb7c4cf8d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ac7c9),
	.w1(32'hb71a0fe5),
	.w2(32'hb6f09311),
	.w3(32'h37f2eaf8),
	.w4(32'hb771e65a),
	.w5(32'hb727fecd),
	.w6(32'h377a27ba),
	.w7(32'hb7c97dc0),
	.w8(32'hb7b16c25),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d65f61),
	.w1(32'hb98fff3e),
	.w2(32'hb92fe9a8),
	.w3(32'h3913ed86),
	.w4(32'hb989a860),
	.w5(32'hb95d7782),
	.w6(32'h388c3b44),
	.w7(32'hb9a509b2),
	.w8(32'hb96851e4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e0194a),
	.w1(32'hb7664b71),
	.w2(32'h372fdced),
	.w3(32'h380b79b4),
	.w4(32'hb7173f9d),
	.w5(32'h372f9dee),
	.w6(32'h37582e74),
	.w7(32'hb7b6d618),
	.w8(32'hb74e4b33),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33135aa5),
	.w1(32'h36568d86),
	.w2(32'hb6b708e3),
	.w3(32'h33d47ac9),
	.w4(32'h36a09ea5),
	.w5(32'hb6bb7c9a),
	.w6(32'hb615a903),
	.w7(32'h322ce725),
	.w8(32'hb6bbc5cf),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a4426f),
	.w1(32'hb6bca141),
	.w2(32'hb4218504),
	.w3(32'hb5c385bd),
	.w4(32'hb68f5116),
	.w5(32'hb617a89c),
	.w6(32'hb67dcc09),
	.w7(32'hb6bffb45),
	.w8(32'hb6cfe1ad),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc88b1),
	.w1(32'hb6ce99e9),
	.w2(32'h35f54084),
	.w3(32'h376ad7f4),
	.w4(32'h37326b9f),
	.w5(32'h377b6ca6),
	.w6(32'hb708bfc4),
	.w7(32'h376c5d77),
	.w8(32'hb7208d78),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a308d),
	.w1(32'hb87e6111),
	.w2(32'h375cb296),
	.w3(32'h3850e09d),
	.w4(32'hb8a33474),
	.w5(32'hb765b94b),
	.w6(32'h37982a07),
	.w7(32'hb8cd9d49),
	.w8(32'hb8ec9d53),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397668ef),
	.w1(32'h3885be2f),
	.w2(32'h37699ab5),
	.w3(32'h394cef10),
	.w4(32'h380ab09c),
	.w5(32'h3598f3c1),
	.w6(32'h3884a0ef),
	.w7(32'hb879400e),
	.w8(32'hb82fe3cc),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d745df),
	.w1(32'hb3d3f909),
	.w2(32'h36382710),
	.w3(32'hb63ef59f),
	.w4(32'hb55a3622),
	.w5(32'hb5bc006a),
	.w6(32'h3555ba12),
	.w7(32'h362032ef),
	.w8(32'hb64bf101),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f47f4),
	.w1(32'hb7851c4a),
	.w2(32'hb80ec7a7),
	.w3(32'h38fd08c6),
	.w4(32'hb8078a76),
	.w5(32'hb83e125e),
	.w6(32'h37ce754d),
	.w7(32'hb8b649af),
	.w8(32'hb89fc287),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389bec3f),
	.w1(32'hb8a74747),
	.w2(32'hb88104d4),
	.w3(32'h386d5650),
	.w4(32'hb87f1f50),
	.w5(32'hb88de87f),
	.w6(32'h37aff819),
	.w7(32'hb8b9e15e),
	.w8(32'hb8a8d1e2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1c491),
	.w1(32'h394ff874),
	.w2(32'h391d8e46),
	.w3(32'h38d5485d),
	.w4(32'h390443f7),
	.w5(32'h389669cf),
	.w6(32'hb8b5ad3f),
	.w7(32'h37ac2b8b),
	.w8(32'h38307ddf),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925d49e),
	.w1(32'hb8e8c660),
	.w2(32'hb7d87548),
	.w3(32'h39377177),
	.w4(32'hb8f4e03a),
	.w5(32'hb8236e5b),
	.w6(32'h390bcdfa),
	.w7(32'hb909faf5),
	.w8(32'hb87a0f5d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8065014),
	.w1(32'hb8629cc9),
	.w2(32'hb8457d0f),
	.w3(32'h37053f6d),
	.w4(32'hb8754d12),
	.w5(32'hb844401c),
	.w6(32'h3317055c),
	.w7(32'hb7d4cf21),
	.w8(32'hb84a3668),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813441a),
	.w1(32'hb7ccba58),
	.w2(32'hbb0fd47a),
	.w3(32'hb891b5cb),
	.w4(32'hb79d68c3),
	.w5(32'h3b41aadf),
	.w6(32'hb88c5fab),
	.w7(32'hb7d87323),
	.w8(32'h3aab3a09),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1da083),
	.w1(32'hbb3a6387),
	.w2(32'h3b03e095),
	.w3(32'h3ba4eacc),
	.w4(32'h397db229),
	.w5(32'hbc3a9267),
	.w6(32'h3b9d2ac9),
	.w7(32'hbb38a0de),
	.w8(32'hbc3b77c5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83ed68),
	.w1(32'hbbc9cd96),
	.w2(32'hbb998eab),
	.w3(32'hbc6fcb26),
	.w4(32'hbbdc5d7d),
	.w5(32'h3b287f92),
	.w6(32'hbc14c97b),
	.w7(32'h3bbcebae),
	.w8(32'h3924cea8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65cf06),
	.w1(32'h38cc3f77),
	.w2(32'h3d8490a3),
	.w3(32'h3c11395c),
	.w4(32'h3b12ca06),
	.w5(32'h3ce38299),
	.w6(32'h39aeffcf),
	.w7(32'h3ae2aeff),
	.w8(32'hbd02e577),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd34a1b),
	.w1(32'h3d5d0801),
	.w2(32'hba6e9dd3),
	.w3(32'h3b719c01),
	.w4(32'hbc9c3e16),
	.w5(32'hbc2f3af6),
	.w6(32'hbdcad21a),
	.w7(32'hbdab57b8),
	.w8(32'h3a455f08),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf1968),
	.w1(32'h3c50b92e),
	.w2(32'hbaff9727),
	.w3(32'hb9113294),
	.w4(32'h3b1382a4),
	.w5(32'h3b85d95a),
	.w6(32'h3c0aa85c),
	.w7(32'h3b99fa26),
	.w8(32'h3c043d86),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68e621),
	.w1(32'hbb667749),
	.w2(32'h3d812e00),
	.w3(32'h3c400f85),
	.w4(32'h3c5ceae7),
	.w5(32'h3cd3c919),
	.w6(32'h3c43036b),
	.w7(32'h3b9996fd),
	.w8(32'hbd222e5f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ddcb587),
	.w1(32'h3d53689f),
	.w2(32'h3c1e82f0),
	.w3(32'hbb9a1bce),
	.w4(32'hbcbcd4e1),
	.w5(32'hbbc87199),
	.w6(32'hbdf63991),
	.w7(32'hbdb2a820),
	.w8(32'hbbe8cf04),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f9f47),
	.w1(32'hbbff2ae3),
	.w2(32'hbd05b9e4),
	.w3(32'hbbda0bdb),
	.w4(32'hbbf8916c),
	.w5(32'hbbe9baac),
	.w6(32'hbc393b03),
	.w7(32'hbc110ffe),
	.w8(32'h3ca01f30),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5dd440),
	.w1(32'hbcdb36e2),
	.w2(32'h3b990396),
	.w3(32'h3a974d6c),
	.w4(32'h3c6bff7f),
	.w5(32'hbaebfa73),
	.w6(32'h3d69fb25),
	.w7(32'h3d4607bb),
	.w8(32'h3ae38f91),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf971d9),
	.w1(32'hba1e3242),
	.w2(32'h3d3cf852),
	.w3(32'h3c5a0e70),
	.w4(32'h3b95fa74),
	.w5(32'h3c83aba2),
	.w6(32'h3c1d7600),
	.w7(32'hba2b020d),
	.w8(32'hbd120492),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db9dfc4),
	.w1(32'h3d39b42e),
	.w2(32'hbb81301d),
	.w3(32'hbb48dfc2),
	.w4(32'hbc4e3f0a),
	.w5(32'hbb89e618),
	.w6(32'hbdbc4459),
	.w7(32'hbd7a33e4),
	.w8(32'h3b8ecb88),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db73b),
	.w1(32'hbafdd3c3),
	.w2(32'hbbbc5897),
	.w3(32'hbbbea90c),
	.w4(32'hbbf2605e),
	.w5(32'hbc0b4e79),
	.w6(32'h3bdf89b2),
	.w7(32'hba2559e2),
	.w8(32'hbbd5a085),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5d6a7),
	.w1(32'h3c2b6f24),
	.w2(32'h3bdf0df1),
	.w3(32'hbc16cccf),
	.w4(32'h3b8b3530),
	.w5(32'h3bcdf914),
	.w6(32'hbc116089),
	.w7(32'hbbe4009f),
	.w8(32'hba718221),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b300314),
	.w1(32'h3b33aaed),
	.w2(32'hbb7ad5c4),
	.w3(32'hbb83a0cf),
	.w4(32'hbb868bdb),
	.w5(32'hba9e6667),
	.w6(32'hbc24d791),
	.w7(32'hbc1da3fb),
	.w8(32'hbb429130),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb63f99),
	.w1(32'hbbf43acf),
	.w2(32'h3ae25f87),
	.w3(32'h39830800),
	.w4(32'h3b8c1be3),
	.w5(32'hb9f101b3),
	.w6(32'h3a526e30),
	.w7(32'h3bb11aa4),
	.w8(32'h3bae7b6f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803057c),
	.w1(32'h3bec1ea5),
	.w2(32'hbd775366),
	.w3(32'h3bf736cf),
	.w4(32'h39a52309),
	.w5(32'hbc9c3895),
	.w6(32'h3baff5a3),
	.w7(32'h3ad80568),
	.w8(32'h3d205eea),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdbdbfb7),
	.w1(32'hbd3a6c8a),
	.w2(32'h3b9cbdad),
	.w3(32'h3c09d917),
	.w4(32'h3ca6145c),
	.w5(32'h3bac42bd),
	.w6(32'h3de2f3c7),
	.w7(32'h3d9f2c21),
	.w8(32'h3ac4c0de),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83aba1),
	.w1(32'h3b50d482),
	.w2(32'hbb105366),
	.w3(32'h3ba55c1c),
	.w4(32'h3b87f587),
	.w5(32'h3ba5548e),
	.w6(32'h3bb8d798),
	.w7(32'h3afa5bc2),
	.w8(32'h3b04fc0f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55099b),
	.w1(32'hb816c30d),
	.w2(32'hbb73d253),
	.w3(32'h3a3554eb),
	.w4(32'hbb506285),
	.w5(32'hbb1f7c46),
	.w6(32'h3b9bf68d),
	.w7(32'hba780a3d),
	.w8(32'h3b023481),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3137c6),
	.w1(32'hba4118e5),
	.w2(32'hbbed2a01),
	.w3(32'h3c7f5a3b),
	.w4(32'h3c418a28),
	.w5(32'hbb8cd299),
	.w6(32'h3c3d35b2),
	.w7(32'h3c0998e9),
	.w8(32'hbae39d0f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf93b4c),
	.w1(32'hbbf0ec5c),
	.w2(32'hbd8fd6d8),
	.w3(32'hbb6ce93d),
	.w4(32'h3baee6bb),
	.w5(32'hbcdf0b37),
	.w6(32'hbad71257),
	.w7(32'hbba08409),
	.w8(32'h3d24cf71),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdddae7c),
	.w1(32'hbd5fabe2),
	.w2(32'hbbb4f19d),
	.w3(32'h3be99e1e),
	.w4(32'h3cdd239b),
	.w5(32'h3ab6c372),
	.w6(32'h3dfb2023),
	.w7(32'h3dcd3f6a),
	.w8(32'hbb72acb8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfac0f),
	.w1(32'hb94d72db),
	.w2(32'hbb1291f7),
	.w3(32'hbca64310),
	.w4(32'hbc1f5c0d),
	.w5(32'hbbe68ca3),
	.w6(32'hbc72c67d),
	.w7(32'hbc1214d7),
	.w8(32'hbb8806ec),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6fed3),
	.w1(32'h3b17c181),
	.w2(32'hbbc90e06),
	.w3(32'hba68f843),
	.w4(32'h39f5d9a2),
	.w5(32'h3b2c1b33),
	.w6(32'h3b71c801),
	.w7(32'h3b888e7c),
	.w8(32'h3bf0d602),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb48a6f),
	.w1(32'h3b34e183),
	.w2(32'hbbef4e86),
	.w3(32'h3b753a66),
	.w4(32'h3bb8f3ea),
	.w5(32'hbc2b1fa1),
	.w6(32'h3bcf0fdc),
	.w7(32'h3bc4f550),
	.w8(32'hbbca2e18),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0c7d),
	.w1(32'hbb74b01a),
	.w2(32'hbc00f3a3),
	.w3(32'hbad0e88a),
	.w4(32'hbc17e508),
	.w5(32'hbbfcb465),
	.w6(32'h3b2702d4),
	.w7(32'hbb03babf),
	.w8(32'hbad2a4a8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae32370),
	.w1(32'h3a7eace0),
	.w2(32'hbbabbde4),
	.w3(32'hbc4dfb62),
	.w4(32'hba44d6c6),
	.w5(32'hbbb09e13),
	.w6(32'h3b4648cd),
	.w7(32'h3b9640f7),
	.w8(32'hbbea9c14),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad8526),
	.w1(32'hbb6b97b1),
	.w2(32'hbc1db39f),
	.w3(32'hbbfdff45),
	.w4(32'hbc10985a),
	.w5(32'hbc0c8beb),
	.w6(32'hbba4ea03),
	.w7(32'hbb68bd22),
	.w8(32'hbc232c6e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd134af),
	.w1(32'hbb872649),
	.w2(32'h3be19921),
	.w3(32'hbbe26524),
	.w4(32'hbc843c58),
	.w5(32'h3ab56579),
	.w6(32'hbbde7174),
	.w7(32'hbc9dce23),
	.w8(32'hbb429661),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3ddb),
	.w1(32'h3bed32a6),
	.w2(32'h3c833c97),
	.w3(32'h3c27a070),
	.w4(32'h3c805cc8),
	.w5(32'hbab334f2),
	.w6(32'h3c407953),
	.w7(32'h3c7f0671),
	.w8(32'hbc1d9e5b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83832f),
	.w1(32'h3ba75b60),
	.w2(32'hbb089ba1),
	.w3(32'hbc378420),
	.w4(32'hbb9bb523),
	.w5(32'hbb6159d7),
	.w6(32'hbc93e155),
	.w7(32'hbb2c51cc),
	.w8(32'h3becdeaf),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1fbf1),
	.w1(32'hbbf485e2),
	.w2(32'h3c4b9d99),
	.w3(32'h3a42e981),
	.w4(32'hbc2568f2),
	.w5(32'hbbc38c85),
	.w6(32'h3b936c32),
	.w7(32'hbaee5f07),
	.w8(32'h3ab595a9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4796c),
	.w1(32'h3c5b36db),
	.w2(32'h3bb4c172),
	.w3(32'hbc673328),
	.w4(32'hbb331644),
	.w5(32'hbb882f4c),
	.w6(32'hbbe33c51),
	.w7(32'h3ae8763b),
	.w8(32'h3b16207f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ae469),
	.w1(32'h3be29468),
	.w2(32'hbc65ee5a),
	.w3(32'hbad740e6),
	.w4(32'h3b215752),
	.w5(32'hbb34109f),
	.w6(32'hba460cb9),
	.w7(32'h3a84a61b),
	.w8(32'h3b2800da),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258f45),
	.w1(32'hbbcc8d48),
	.w2(32'hb9a04591),
	.w3(32'h3afe807c),
	.w4(32'hbb8d2ade),
	.w5(32'hbb329e35),
	.w6(32'h3b782c5b),
	.w7(32'hbbbb03ba),
	.w8(32'hba5f9cf8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fae2ca),
	.w1(32'h3bd4ad3e),
	.w2(32'hbb3a1c0d),
	.w3(32'h3bce9940),
	.w4(32'h3c08dba2),
	.w5(32'h3a8099b4),
	.w6(32'h3b8a4934),
	.w7(32'h3b473ad8),
	.w8(32'h3b7729dc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5e409),
	.w1(32'h3b934214),
	.w2(32'hbb25c453),
	.w3(32'h3c239f1f),
	.w4(32'h3b2da669),
	.w5(32'h3c0a1c55),
	.w6(32'h3c4cd4fd),
	.w7(32'h3ba1f11c),
	.w8(32'hbb2372dd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f91d5),
	.w1(32'hbb6ab7a1),
	.w2(32'h3c11f263),
	.w3(32'h3b3979e2),
	.w4(32'h3b6ffd62),
	.w5(32'h3c1b519f),
	.w6(32'hbb978149),
	.w7(32'hbb9bf570),
	.w8(32'h3bbf66fe),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1516b4),
	.w1(32'h3b9046d6),
	.w2(32'h3c2ea507),
	.w3(32'h3bf9b50e),
	.w4(32'h3bbd172e),
	.w5(32'h3c3068fb),
	.w6(32'h3bbb99f8),
	.w7(32'h3bd3ed53),
	.w8(32'h3baab946),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a2021),
	.w1(32'h3c387532),
	.w2(32'h3b6640c3),
	.w3(32'h3adce77f),
	.w4(32'hbb8abca6),
	.w5(32'h39e0d71c),
	.w6(32'hbbe9bd73),
	.w7(32'hbc4498fa),
	.w8(32'h3b0c085e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff70d2),
	.w1(32'h3ad48a96),
	.w2(32'h3b6a33bc),
	.w3(32'h3bb566d4),
	.w4(32'h3aab8754),
	.w5(32'h3bfa2eaa),
	.w6(32'h3bcd2852),
	.w7(32'h3b933c54),
	.w8(32'h3a4883de),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab791d8),
	.w1(32'hbb208205),
	.w2(32'h3b637508),
	.w3(32'h3b03c230),
	.w4(32'h3aec3888),
	.w5(32'h3b9a3287),
	.w6(32'h3ae3ec95),
	.w7(32'hbb4ef4b7),
	.w8(32'h3b6447d8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba992397),
	.w1(32'h3aadf8a3),
	.w2(32'h3bfc48c9),
	.w3(32'hba369b28),
	.w4(32'h3b8ecab8),
	.w5(32'hba7d96b9),
	.w6(32'hbb1b336d),
	.w7(32'h3b559e97),
	.w8(32'hbbe6207e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beddc8d),
	.w1(32'h3c1cddff),
	.w2(32'hbc0bebcc),
	.w3(32'hbb1ec047),
	.w4(32'hbb1a9ca4),
	.w5(32'hbc2aacd6),
	.w6(32'hbc001fb1),
	.w7(32'hbc91ced8),
	.w8(32'hbc1282c4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc52e8),
	.w1(32'hbbb448c1),
	.w2(32'hb9c48482),
	.w3(32'hbc00feae),
	.w4(32'hbc2ae946),
	.w5(32'h3a7db12d),
	.w6(32'hbba2ac95),
	.w7(32'hbb5cffd9),
	.w8(32'h3b3e6d3f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba743c4a),
	.w1(32'hbb689f4c),
	.w2(32'h3b825fcc),
	.w3(32'h3b935d06),
	.w4(32'hb9cabe1a),
	.w5(32'hbb4802fa),
	.w6(32'h3c0c1e19),
	.w7(32'hbbbe3d16),
	.w8(32'hbaafc20c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be89f77),
	.w1(32'hb9223096),
	.w2(32'hbd662f34),
	.w3(32'h3b89a05f),
	.w4(32'h3c0b1f44),
	.w5(32'hbcd4027c),
	.w6(32'hb828d0f1),
	.w7(32'h3ba17cf8),
	.w8(32'h3cbbcb61),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda8fcdb),
	.w1(32'hbd5e9d9a),
	.w2(32'h3c06e54b),
	.w3(32'h3abb545c),
	.w4(32'h3bd065c9),
	.w5(32'h3c102493),
	.w6(32'h3dad28c0),
	.w7(32'h3d7497db),
	.w8(32'h3c05f77f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad826d3),
	.w1(32'hba516b51),
	.w2(32'hbb0a569d),
	.w3(32'hbb8d1fdc),
	.w4(32'hbbf8ab16),
	.w5(32'hb930f86f),
	.w6(32'hbb4b1270),
	.w7(32'hbb7f77ff),
	.w8(32'h3b7c0eaf),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866354d),
	.w1(32'h3b9fb7d2),
	.w2(32'hbc45d43c),
	.w3(32'h3baa6c2c),
	.w4(32'h391fc8f5),
	.w5(32'h3b00ceba),
	.w6(32'h3a228b76),
	.w7(32'hbbc17454),
	.w8(32'h39c0cdbe),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f1df4),
	.w1(32'h3b5c3bbd),
	.w2(32'h3b9daa6d),
	.w3(32'h3c1bde4c),
	.w4(32'h3b8ec4eb),
	.w5(32'hbb01a77f),
	.w6(32'h3be568ab),
	.w7(32'h3abcae8d),
	.w8(32'hbb7e9e33),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf772d),
	.w1(32'h3ab5f06b),
	.w2(32'hbb21eea5),
	.w3(32'h3bb27bbd),
	.w4(32'h3ba0166a),
	.w5(32'h3afd60f2),
	.w6(32'h3b65117a),
	.w7(32'h3c1a323b),
	.w8(32'h3a9b2684),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc380361),
	.w1(32'hbb91dace),
	.w2(32'hbba536b0),
	.w3(32'hbc046810),
	.w4(32'hbadc7bda),
	.w5(32'hbb886df9),
	.w6(32'hbc143ed5),
	.w7(32'hbbb5626d),
	.w8(32'hbb97dbe1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee4683),
	.w1(32'h3ab7790d),
	.w2(32'h3cfa91b8),
	.w3(32'hbb602453),
	.w4(32'h3b6b554a),
	.w5(32'h3ca96f90),
	.w6(32'h3ab5e342),
	.w7(32'h3b287aed),
	.w8(32'hbc0b0e5e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d51f873),
	.w1(32'h3c818e28),
	.w2(32'h3afe2180),
	.w3(32'h3b39c6c6),
	.w4(32'hbc9a2bbf),
	.w5(32'hbac2b66c),
	.w6(32'hbd5297c7),
	.w7(32'hbd3e7893),
	.w8(32'hbb8e97c7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade3e3d),
	.w1(32'hbaa651e9),
	.w2(32'hbb17d524),
	.w3(32'h3be31647),
	.w4(32'h393704f4),
	.w5(32'h3b8167cb),
	.w6(32'h3c04c114),
	.w7(32'h3a33391c),
	.w8(32'h3c61c0a4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e4af),
	.w1(32'hbb0cd4f2),
	.w2(32'hbb3fde2c),
	.w3(32'h39afdadd),
	.w4(32'h3bb16f8a),
	.w5(32'h3a755b97),
	.w6(32'h3c5b1ad1),
	.w7(32'h3bc790e3),
	.w8(32'h3a4adbc7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc065bf9),
	.w1(32'hb9d74c08),
	.w2(32'hbacd8c61),
	.w3(32'h3af267ba),
	.w4(32'hbbe3c452),
	.w5(32'h3b81b8c2),
	.w6(32'h3ab02695),
	.w7(32'hba4f1ff7),
	.w8(32'hbb030475),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8874a5),
	.w1(32'hbc0dde93),
	.w2(32'h3b88840d),
	.w3(32'hbb48e8c7),
	.w4(32'hbb20142e),
	.w5(32'h3a9d9fc7),
	.w6(32'hb9847163),
	.w7(32'h3c046038),
	.w8(32'hb9a1b056),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b707ac6),
	.w1(32'hbb8bf17c),
	.w2(32'h3b63ac33),
	.w3(32'h3bbb810e),
	.w4(32'hbadda769),
	.w5(32'h3b93e7aa),
	.w6(32'h3c18a05c),
	.w7(32'h3b9db79b),
	.w8(32'h3b2e3bf5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b764),
	.w1(32'hbc018c00),
	.w2(32'hbb50d382),
	.w3(32'hba6f4ff9),
	.w4(32'h399ae96e),
	.w5(32'hbabedd3d),
	.w6(32'h3bbdddd3),
	.w7(32'h3bc3a8b9),
	.w8(32'hbb137cfd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aab23),
	.w1(32'hbb44a8cc),
	.w2(32'hbbbe1fbe),
	.w3(32'h3ac7c8f2),
	.w4(32'hbbbd464b),
	.w5(32'hbc46fda5),
	.w6(32'hbb2e5145),
	.w7(32'h3ba1756e),
	.w8(32'hbb9c6fff),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2cdd),
	.w1(32'hba8b3c3d),
	.w2(32'h3c0d9c3b),
	.w3(32'hbc61d399),
	.w4(32'hbc57653c),
	.w5(32'h3c97091a),
	.w6(32'hbb037671),
	.w7(32'hbb69f5c3),
	.w8(32'h3c1c410d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c924d66),
	.w1(32'h3c9d5dac),
	.w2(32'h3bdcfbef),
	.w3(32'h3cb8188e),
	.w4(32'h3ca0b713),
	.w5(32'hbb3ef8c5),
	.w6(32'h3c20a4fb),
	.w7(32'h3bd64fa8),
	.w8(32'h3b5962ea),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50a4f9),
	.w1(32'h3c449950),
	.w2(32'h3a2cf685),
	.w3(32'h3b178cfa),
	.w4(32'h3bda1996),
	.w5(32'h3b87abaf),
	.w6(32'h3b8ac539),
	.w7(32'h3bb848b2),
	.w8(32'h3aeb5125),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c9775),
	.w1(32'hbb2eeeda),
	.w2(32'hbb6d9d71),
	.w3(32'hbb8cb0a5),
	.w4(32'hbb697bb9),
	.w5(32'hbaedeadf),
	.w6(32'hbc19f050),
	.w7(32'hbbba20ac),
	.w8(32'h3b85e041),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8eb981),
	.w1(32'hbc3740b8),
	.w2(32'h3b9f67a1),
	.w3(32'hbad86a71),
	.w4(32'hbbfc29a7),
	.w5(32'h3bd0b96f),
	.w6(32'h3c3c4959),
	.w7(32'hbaead801),
	.w8(32'hbafcaeb5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ed79),
	.w1(32'hba8e29ff),
	.w2(32'hbbca2313),
	.w3(32'h3bbe338d),
	.w4(32'h3bb11024),
	.w5(32'h3bd510a7),
	.w6(32'hba94aa76),
	.w7(32'h39131d2b),
	.w8(32'h3c2571df),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3095e8),
	.w1(32'h3bc0596d),
	.w2(32'hb9a6af05),
	.w3(32'h3c3637c7),
	.w4(32'h3b0bc11f),
	.w5(32'hba3a4c22),
	.w6(32'h3c02503b),
	.w7(32'h3b6905a5),
	.w8(32'h3bb4455d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab105f),
	.w1(32'hbb13fdd5),
	.w2(32'hbb39c4b7),
	.w3(32'hbb6fa620),
	.w4(32'hbb871ca3),
	.w5(32'hbbc67fec),
	.w6(32'h3b9dbec6),
	.w7(32'h378e522c),
	.w8(32'hbb978617),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87c419),
	.w1(32'h3ba72e23),
	.w2(32'hbbb13d4c),
	.w3(32'h3c276beb),
	.w4(32'h3c2b7b49),
	.w5(32'hbc1363ed),
	.w6(32'h3baf5497),
	.w7(32'h3bf50381),
	.w8(32'hbc3467b5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2affe9),
	.w1(32'hbc109e35),
	.w2(32'h3b563f68),
	.w3(32'hbc030cad),
	.w4(32'hbb34171d),
	.w5(32'h3ba9848b),
	.w6(32'h3aae1807),
	.w7(32'h3bb54bd9),
	.w8(32'h3c2fb0f6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a1592),
	.w1(32'h3bb7f6b9),
	.w2(32'hbbaeab54),
	.w3(32'h3c54a118),
	.w4(32'hbbda5922),
	.w5(32'hbb052f71),
	.w6(32'h3c9d8a18),
	.w7(32'hbbaf97e2),
	.w8(32'hbb3a8eff),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe614eb),
	.w1(32'hba5e48d9),
	.w2(32'h3ab788ec),
	.w3(32'h3ada3151),
	.w4(32'h3a87c6ed),
	.w5(32'hbbc7a3f3),
	.w6(32'h3b05e496),
	.w7(32'hbb4fd923),
	.w8(32'hbb54f90a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eeb8c9),
	.w1(32'hbc078e0a),
	.w2(32'hbc049cc6),
	.w3(32'hb928ba1a),
	.w4(32'hbb8c8881),
	.w5(32'hbb854302),
	.w6(32'h3aad10fc),
	.w7(32'hba2adb6c),
	.w8(32'hbb5170a9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e3143),
	.w1(32'hbbbfe573),
	.w2(32'hb875bd93),
	.w3(32'hbbe3ae5b),
	.w4(32'hbad2d2b9),
	.w5(32'h3b006668),
	.w6(32'h3c3b71ae),
	.w7(32'h3b305eb6),
	.w8(32'h3bc47620),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97b7fc),
	.w1(32'h3baabd1e),
	.w2(32'hbb565184),
	.w3(32'h3be34b58),
	.w4(32'h3c1ec928),
	.w5(32'hbb553fc8),
	.w6(32'h3cad27f5),
	.w7(32'h3c1a0509),
	.w8(32'h3a5ad6e3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc169c63),
	.w1(32'hbb19bd0e),
	.w2(32'hbb83be08),
	.w3(32'h3a822460),
	.w4(32'h3bab078d),
	.w5(32'hbc148938),
	.w6(32'h3c67904b),
	.w7(32'h3c661123),
	.w8(32'hbc39e426),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba976d0),
	.w1(32'hbb917a74),
	.w2(32'hbb91f90c),
	.w3(32'hbbf09a6c),
	.w4(32'hbb6aafc8),
	.w5(32'hbbe8160b),
	.w6(32'hbc214f70),
	.w7(32'hbb17f9d0),
	.w8(32'hbc34a7b9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2798f8),
	.w1(32'hbb956756),
	.w2(32'hbc4958b3),
	.w3(32'hbbaf0852),
	.w4(32'h3a73bf98),
	.w5(32'hbbe18513),
	.w6(32'hbb6e76f2),
	.w7(32'h3bea8a62),
	.w8(32'hbb8d4599),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49bac9),
	.w1(32'hbbcf3667),
	.w2(32'hbb3198bf),
	.w3(32'hbc2be86e),
	.w4(32'hbc1f83a5),
	.w5(32'hba3c209f),
	.w6(32'h3be05dae),
	.w7(32'h3b89fd98),
	.w8(32'h3c0e6e33),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4df5e6),
	.w1(32'hbad4af7c),
	.w2(32'hbc3fc291),
	.w3(32'hbb4ab2fd),
	.w4(32'hbb3a055c),
	.w5(32'hbb878373),
	.w6(32'h3b6997c7),
	.w7(32'h3aef3671),
	.w8(32'hbbadb2f1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf450e9),
	.w1(32'hbae5ce4d),
	.w2(32'h3ae91740),
	.w3(32'hbbdfe20c),
	.w4(32'hbb82f56c),
	.w5(32'hbbdf5c71),
	.w6(32'hbb53e1ca),
	.w7(32'hbb77064a),
	.w8(32'hb9b5a8fa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a30f3),
	.w1(32'hbb71a8bf),
	.w2(32'h3ae6840d),
	.w3(32'h3b339b7d),
	.w4(32'hbabef737),
	.w5(32'hbba56cd7),
	.w6(32'hbb2ce3c0),
	.w7(32'hb9cea5f4),
	.w8(32'hbbd2a482),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9463a3),
	.w1(32'h3c15555e),
	.w2(32'hbb488c2b),
	.w3(32'h3b933601),
	.w4(32'h3b0d0882),
	.w5(32'hbaa097df),
	.w6(32'h3b9d0025),
	.w7(32'hbb308fa4),
	.w8(32'hbab475c9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ff5fd8),
	.w1(32'hbb2bbd8e),
	.w2(32'hb9bc8144),
	.w3(32'hbb821dd1),
	.w4(32'hba28bbfd),
	.w5(32'hb81e9777),
	.w6(32'hbb6c756e),
	.w7(32'hbc6b2511),
	.w8(32'h39f1a648),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f98f6),
	.w1(32'h3b70ecd1),
	.w2(32'hbac65a03),
	.w3(32'h393430e3),
	.w4(32'h3b2d13b1),
	.w5(32'hbbcbc21e),
	.w6(32'h3a9cf21f),
	.w7(32'h3bdb97cc),
	.w8(32'h3b4647fb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2b3e4),
	.w1(32'hbb86e02b),
	.w2(32'hbb8daf24),
	.w3(32'hbc1832c5),
	.w4(32'hbb979850),
	.w5(32'hbba264a9),
	.w6(32'hbbab122b),
	.w7(32'h3b78e0e9),
	.w8(32'h3b839971),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4825),
	.w1(32'hbbd7322c),
	.w2(32'h3bfee70c),
	.w3(32'hbc2c4642),
	.w4(32'hbc563a05),
	.w5(32'hbabee816),
	.w6(32'h3b013a25),
	.w7(32'hbb05766b),
	.w8(32'h3b53fa4a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d09ac),
	.w1(32'h3c1b1bbe),
	.w2(32'hbbc717ac),
	.w3(32'h3bb086c5),
	.w4(32'h3a25ce34),
	.w5(32'hbca056bb),
	.w6(32'hbaf704b7),
	.w7(32'hbb11f875),
	.w8(32'hbbf97890),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc790c16),
	.w1(32'hbbbd00fa),
	.w2(32'hbb7c8faf),
	.w3(32'hbcf2db9d),
	.w4(32'hbc7be1ff),
	.w5(32'hbbad10fb),
	.w6(32'hbc10de75),
	.w7(32'hbb5684a9),
	.w8(32'hb81b1d89),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f57f3),
	.w1(32'h3ace4c3c),
	.w2(32'hbb9a2cdf),
	.w3(32'h3bbd2da0),
	.w4(32'hbb236e3f),
	.w5(32'hbb8fe423),
	.w6(32'h3bae282e),
	.w7(32'h3ba878a0),
	.w8(32'h3a7f4f1b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f719d),
	.w1(32'hbb79981c),
	.w2(32'h3bd8185d),
	.w3(32'hba861c06),
	.w4(32'h3a96a2b9),
	.w5(32'h39f57c66),
	.w6(32'hbb607315),
	.w7(32'hbbc94901),
	.w8(32'h3b83f41b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80724c),
	.w1(32'h3b4bd776),
	.w2(32'h3c993738),
	.w3(32'h39f085d9),
	.w4(32'h3b3ec80e),
	.w5(32'h3c05a9ef),
	.w6(32'h3af96b32),
	.w7(32'h3b37ebee),
	.w8(32'hbbb6f441),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4fdc4),
	.w1(32'h3c9ddf73),
	.w2(32'h3d16587e),
	.w3(32'h3bf8e2f8),
	.w4(32'h3a5c4658),
	.w5(32'h3ca42405),
	.w6(32'hbc89a08f),
	.w7(32'hbc788ebd),
	.w8(32'hbc08b0de),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5452d4),
	.w1(32'h3ce7875d),
	.w2(32'h3af2547a),
	.w3(32'h3c0d5737),
	.w4(32'hbb038878),
	.w5(32'hba8e0345),
	.w6(32'hbd1ee6c3),
	.w7(32'hbcfc25e8),
	.w8(32'hbc1fcda9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd265a),
	.w1(32'h3a557931),
	.w2(32'h3b65f3d7),
	.w3(32'hba884d0b),
	.w4(32'h3c06a9c3),
	.w5(32'hbc0c9760),
	.w6(32'h3b7127df),
	.w7(32'h3c405d57),
	.w8(32'hbb93a99b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cf908),
	.w1(32'hb9464962),
	.w2(32'hbbf4dfa9),
	.w3(32'hbc3f305d),
	.w4(32'h3ad825a0),
	.w5(32'hbad20068),
	.w6(32'hbc10a0c9),
	.w7(32'hba9d8f67),
	.w8(32'h3b2b5c1c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00bc8),
	.w1(32'h3bae02e1),
	.w2(32'h3ba785d3),
	.w3(32'h3aceb466),
	.w4(32'h3c11df6a),
	.w5(32'h3b9a9935),
	.w6(32'h3aa47d4f),
	.w7(32'h3b9f9227),
	.w8(32'h3b8283c0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba734218),
	.w1(32'h3c15281d),
	.w2(32'h3bc3dedc),
	.w3(32'h3bf03399),
	.w4(32'hbae50c46),
	.w5(32'h3bd0b18d),
	.w6(32'h3c4f9586),
	.w7(32'h3acdd017),
	.w8(32'h3bf3c7a0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5838a),
	.w1(32'h3a6896fd),
	.w2(32'hbc279048),
	.w3(32'h3b85f7f5),
	.w4(32'h3a20b4ed),
	.w5(32'hbbdcf2de),
	.w6(32'h3b451f33),
	.w7(32'h3bece84b),
	.w8(32'h3b347624),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule