module layer_8_featuremap_48(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb4af),
	.w1(32'hbb2906f2),
	.w2(32'hbad6ed97),
	.w3(32'hba43960c),
	.w4(32'hbbcb1d6a),
	.w5(32'hbbaf6d3a),
	.w6(32'hbb6130a4),
	.w7(32'hbb3f86fb),
	.w8(32'hbafc34df),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999d2b),
	.w1(32'h3a981bdd),
	.w2(32'h3b77b10f),
	.w3(32'hbb0183b8),
	.w4(32'hba7e7b52),
	.w5(32'hba6f296c),
	.w6(32'h3a11560e),
	.w7(32'h39b46e37),
	.w8(32'hbae2b597),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c824),
	.w1(32'h387e7f2f),
	.w2(32'h3ae6df4f),
	.w3(32'hbab36fcf),
	.w4(32'h3a124b3b),
	.w5(32'hb96dec12),
	.w6(32'h3ab86ae6),
	.w7(32'h3a770043),
	.w8(32'h3c7550cf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02bdbd),
	.w1(32'h3c61844c),
	.w2(32'h3d0e123d),
	.w3(32'hbafe243a),
	.w4(32'h3bc2628a),
	.w5(32'h3c794afb),
	.w6(32'h3c0f9373),
	.w7(32'h3bc5ccb1),
	.w8(32'hbb641e0a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17a475),
	.w1(32'h3b0dfe17),
	.w2(32'h3b01dc8a),
	.w3(32'hbbac0858),
	.w4(32'h39c7b860),
	.w5(32'hba19caf7),
	.w6(32'h39c122dd),
	.w7(32'hbaa14f7f),
	.w8(32'hbcc38d6e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd22347a),
	.w1(32'h3bfdd965),
	.w2(32'h3d2cfe79),
	.w3(32'hbc8162ec),
	.w4(32'h3a27e6e3),
	.w5(32'h3c836d89),
	.w6(32'hba8f1226),
	.w7(32'h3c604682),
	.w8(32'hbaf37ee3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf9df3),
	.w1(32'hba374b2c),
	.w2(32'h3b253a3e),
	.w3(32'hbad6df63),
	.w4(32'hba893726),
	.w5(32'hbb2a55b7),
	.w6(32'h3a6b8d64),
	.w7(32'hb688b566),
	.w8(32'hbb7f1367),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33be36),
	.w1(32'h3aa213c8),
	.w2(32'h3a2274c0),
	.w3(32'hbbad5abf),
	.w4(32'hbac279b5),
	.w5(32'hbb3b4fbf),
	.w6(32'hbaa259ec),
	.w7(32'hbb35f82e),
	.w8(32'hbb8fe11c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ecaeb),
	.w1(32'hbab5d534),
	.w2(32'hba538026),
	.w3(32'hbb7f0eb0),
	.w4(32'hbb2249cb),
	.w5(32'hbbcc1910),
	.w6(32'hb8dcb6d9),
	.w7(32'hbb5ad934),
	.w8(32'hb909091d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaeb1e6),
	.w1(32'hbbc0c29d),
	.w2(32'hbbcd7c7b),
	.w3(32'hbc10074f),
	.w4(32'hbaa7cdd3),
	.w5(32'h3b954c3d),
	.w6(32'h3bf011c5),
	.w7(32'hbb94a0dc),
	.w8(32'hbb29b939),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f4cee),
	.w1(32'hbae679cf),
	.w2(32'hbabcad53),
	.w3(32'hbaf31302),
	.w4(32'hb937906d),
	.w5(32'hbb727f2c),
	.w6(32'h3a81e742),
	.w7(32'hbaf9f9f0),
	.w8(32'hbb86be4b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a695d),
	.w1(32'h3a0e35e6),
	.w2(32'h3b9fa265),
	.w3(32'hbb58d138),
	.w4(32'hba6d8d07),
	.w5(32'hbabf097c),
	.w6(32'h38c1475b),
	.w7(32'h3a0ed962),
	.w8(32'hbb52c5d9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd04ae),
	.w1(32'hba98c94c),
	.w2(32'h36710730),
	.w3(32'hbb17f79a),
	.w4(32'hbab3078e),
	.w5(32'hbb847fe4),
	.w6(32'h3a74ceb6),
	.w7(32'hbad38a87),
	.w8(32'hbcd50767),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e1e86),
	.w1(32'h3c06b369),
	.w2(32'h3d3e83b1),
	.w3(32'hbc883aed),
	.w4(32'hba32ef34),
	.w5(32'h3c871a15),
	.w6(32'hbb0119ac),
	.w7(32'h3c699580),
	.w8(32'hbc88f715),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03dd70),
	.w1(32'h3ba1b4f3),
	.w2(32'h3cedb8e8),
	.w3(32'hbc71aa51),
	.w4(32'h3aa7539d),
	.w5(32'h3c3e059a),
	.w6(32'h3ac3bb46),
	.w7(32'h3c161e5b),
	.w8(32'hbaf2e41e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925141),
	.w1(32'hba3ff548),
	.w2(32'h397dd00a),
	.w3(32'h3b1539bd),
	.w4(32'hbb9a8d90),
	.w5(32'hbbcecade),
	.w6(32'hbbc7436d),
	.w7(32'hbb425a9e),
	.w8(32'h3c68c733),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cec3854),
	.w1(32'hbc11bb8c),
	.w2(32'hbc2da83b),
	.w3(32'hbb36b4d9),
	.w4(32'h3bf01d24),
	.w5(32'h3cb0dba6),
	.w6(32'hbb82e604),
	.w7(32'hbb58c88d),
	.w8(32'hbb1a5532),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd56dd5),
	.w1(32'hbaf6c1db),
	.w2(32'hb982ebf4),
	.w3(32'hba5e48b1),
	.w4(32'hbaa940b4),
	.w5(32'hbb82e684),
	.w6(32'h3b5e6271),
	.w7(32'hba412593),
	.w8(32'hbbbda882),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc503567),
	.w1(32'h3b1b724a),
	.w2(32'hbbd7f2b9),
	.w3(32'hbb7e023d),
	.w4(32'hbb3fc077),
	.w5(32'hbc44b37c),
	.w6(32'hbb35d72c),
	.w7(32'hbc5915c5),
	.w8(32'hbbad6b84),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00b38c),
	.w1(32'h3b77d752),
	.w2(32'hbcd1ffdb),
	.w3(32'h3c1e09b4),
	.w4(32'hbc3afdde),
	.w5(32'hbc5e6fab),
	.w6(32'hbb7dba24),
	.w7(32'hbc610a3b),
	.w8(32'hbba23331),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13261e),
	.w1(32'hbb7ae356),
	.w2(32'hbc251a83),
	.w3(32'hbb319c27),
	.w4(32'hbb4c9e37),
	.w5(32'hbb70cd87),
	.w6(32'hbb8ddc52),
	.w7(32'hbb9da94f),
	.w8(32'hbb61f2ff),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc047f37),
	.w1(32'h3b2a82ac),
	.w2(32'h3bde0a68),
	.w3(32'hbb5b2462),
	.w4(32'h3b0d6cd7),
	.w5(32'h3b84c108),
	.w6(32'h3c0d0989),
	.w7(32'h3bdc0eea),
	.w8(32'h3cdfa9bb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4ccca7),
	.w1(32'hbc142d08),
	.w2(32'hbd330423),
	.w3(32'h3ca1d220),
	.w4(32'hbc44af94),
	.w5(32'hbcdcdba6),
	.w6(32'hbc5f2b67),
	.w7(32'hbcc9efb3),
	.w8(32'hbb83b6ae),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5efc66),
	.w1(32'h3ad5330e),
	.w2(32'hbc46a481),
	.w3(32'hbb05800d),
	.w4(32'hbbedb435),
	.w5(32'hbc7db631),
	.w6(32'hbb2cc15b),
	.w7(32'hbc6de31b),
	.w8(32'hbbb857a0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a9716),
	.w1(32'hba2ba4b0),
	.w2(32'hbc54fa79),
	.w3(32'hbbf69920),
	.w4(32'hba92a53c),
	.w5(32'h3a8659bf),
	.w6(32'hbc03873c),
	.w7(32'hba501dd7),
	.w8(32'h3cb8790a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d44a15d),
	.w1(32'hbc005a1d),
	.w2(32'hbd207b6e),
	.w3(32'h3cb0dea1),
	.w4(32'hbc180721),
	.w5(32'hbcb91309),
	.w6(32'hbc11132b),
	.w7(32'hbca5392e),
	.w8(32'h3cacdd10),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2b164b),
	.w1(32'hbbc585cd),
	.w2(32'hbd069c0d),
	.w3(32'h3c9d21f2),
	.w4(32'hbbe876e0),
	.w5(32'hbc983832),
	.w6(32'hbbe1e9c9),
	.w7(32'hbc8aec76),
	.w8(32'h3b90adbc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28c179),
	.w1(32'h3a244644),
	.w2(32'hbc2c00ae),
	.w3(32'hbb32a1fc),
	.w4(32'h3a86b489),
	.w5(32'hbaf7080b),
	.w6(32'hbb1409fa),
	.w7(32'hbbbf6f63),
	.w8(32'hbc0e79bc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba709681),
	.w1(32'hbae80bcb),
	.w2(32'hbce52085),
	.w3(32'hbb45c6ff),
	.w4(32'hbcf4d95b),
	.w5(32'hbcc3e29f),
	.w6(32'hbd146d21),
	.w7(32'hbd16146e),
	.w8(32'hbaf116ad),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaf67e),
	.w1(32'h39ab256f),
	.w2(32'h3b55e8f3),
	.w3(32'hbab96211),
	.w4(32'h3a66c065),
	.w5(32'h3a11a0fd),
	.w6(32'h3a9b2b05),
	.w7(32'h3abe318c),
	.w8(32'hbc5bf35b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074eed),
	.w1(32'hbc3e4525),
	.w2(32'h3c9ecd85),
	.w3(32'h3d016f29),
	.w4(32'h3b2489f5),
	.w5(32'hbc20e87c),
	.w6(32'h3b961e71),
	.w7(32'h3cc04ec6),
	.w8(32'hbbc673b7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41f680),
	.w1(32'hbc0ed499),
	.w2(32'hbc8c0956),
	.w3(32'hbc02d7ea),
	.w4(32'hbaaadb4d),
	.w5(32'hb8135bf0),
	.w6(32'hbbadd081),
	.w7(32'h39bfd662),
	.w8(32'hbbf4ea79),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf82d10),
	.w1(32'hbb4b72ab),
	.w2(32'h3d095a48),
	.w3(32'hbc059204),
	.w4(32'hbc872e0a),
	.w5(32'hbc24f3f0),
	.w6(32'hbc18bb95),
	.w7(32'hb8bd7faa),
	.w8(32'h3ae4e9d8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44cec1),
	.w1(32'hbb9e09c5),
	.w2(32'hba215e75),
	.w3(32'h3b4ced7f),
	.w4(32'h3b2d5f2f),
	.w5(32'h3aafe085),
	.w6(32'h3b50ee40),
	.w7(32'h3b82a5b0),
	.w8(32'hbcb6dda9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd13d9b0),
	.w1(32'h3c015268),
	.w2(32'h3d29a594),
	.w3(32'hbc59f7cd),
	.w4(32'h395553d3),
	.w5(32'h3c771ba0),
	.w6(32'hba89130e),
	.w7(32'h3c55d9a7),
	.w8(32'hba0d761f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06703),
	.w1(32'h3a30bc22),
	.w2(32'hbbad370c),
	.w3(32'hbb459a53),
	.w4(32'hbbde17b0),
	.w5(32'hbc4a3561),
	.w6(32'hbb878417),
	.w7(32'hbc2ae1b5),
	.w8(32'hbb8cd003),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db20a),
	.w1(32'hbbf81722),
	.w2(32'hbc5ff3bc),
	.w3(32'hbc251922),
	.w4(32'hbbca4a20),
	.w5(32'hbb13c707),
	.w6(32'hbc06efd0),
	.w7(32'hba6415a8),
	.w8(32'hbb6c34ab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda6d94),
	.w1(32'h3ac348de),
	.w2(32'h3b747404),
	.w3(32'hbad91c96),
	.w4(32'h3b2a6f5e),
	.w5(32'h3afcca13),
	.w6(32'h3b42f9b2),
	.w7(32'h3b228e8f),
	.w8(32'hbd020ce1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8508c1),
	.w1(32'h3bd7bbf2),
	.w2(32'h3d5712c5),
	.w3(32'hbcff07d6),
	.w4(32'h3a699180),
	.w5(32'h3caa3802),
	.w6(32'h39c8e6a9),
	.w7(32'h3c6f20d9),
	.w8(32'h3b219b96),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c54d1),
	.w1(32'hbab54495),
	.w2(32'hbc2a4893),
	.w3(32'h3aca32f2),
	.w4(32'h3b17423f),
	.w5(32'hb8f21900),
	.w6(32'h394f0c60),
	.w7(32'hbaf8a5f5),
	.w8(32'h3c2c1845),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fc633),
	.w1(32'hbb5e83b1),
	.w2(32'hbc87998a),
	.w3(32'h3c0cd92c),
	.w4(32'hbb7009aa),
	.w5(32'hbc1826c8),
	.w6(32'hbb6a7f1d),
	.w7(32'hbc08ff32),
	.w8(32'hb94bab5d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82cadb9),
	.w1(32'h38c7d0b7),
	.w2(32'h37351321),
	.w3(32'hb89d3401),
	.w4(32'h38ab08bd),
	.w5(32'h381b5a84),
	.w6(32'hb932b3cd),
	.w7(32'hb76525dd),
	.w8(32'hb693fd8c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98acc69),
	.w1(32'hb97cde5c),
	.w2(32'hb9b60902),
	.w3(32'hb9ace9d3),
	.w4(32'hb9b7da7a),
	.w5(32'hb9c1b97e),
	.w6(32'hb96d2d1f),
	.w7(32'hb962839e),
	.w8(32'hb9b738d9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cb9cc),
	.w1(32'hba0f3cd5),
	.w2(32'hba5ea828),
	.w3(32'hba7336ce),
	.w4(32'hba5a395c),
	.w5(32'hba90328a),
	.w6(32'hba8cd529),
	.w7(32'hba82d0f7),
	.w8(32'hba966dbe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5b10e),
	.w1(32'h3a1203e0),
	.w2(32'h3a63ed2d),
	.w3(32'h3b164775),
	.w4(32'h3a7ec22f),
	.w5(32'h3a7e3af8),
	.w6(32'h3b212dc2),
	.w7(32'h3ac9a3d4),
	.w8(32'h3a88caa2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399133c4),
	.w1(32'h3a2d7d9b),
	.w2(32'h3a4cb63d),
	.w3(32'h3a3121fd),
	.w4(32'h3a75fbf1),
	.w5(32'h3a825f5d),
	.w6(32'h3a3b6076),
	.w7(32'h3a710a6e),
	.w8(32'h3a88d9c3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb35609f5),
	.w1(32'hb78eb2e8),
	.w2(32'h3713986d),
	.w3(32'hb7b4f60d),
	.w4(32'hb7b3edd2),
	.w5(32'h374d37ba),
	.w6(32'h373d9ea9),
	.w7(32'h37c1d3a7),
	.w8(32'h358a154d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90162aa),
	.w1(32'hbabb7e06),
	.w2(32'hbae6aefc),
	.w3(32'hba71c014),
	.w4(32'hbafef213),
	.w5(32'hbb4ce99b),
	.w6(32'hba04d802),
	.w7(32'hbaa5f196),
	.w8(32'hbb18ffe2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddfa3b),
	.w1(32'h393563dc),
	.w2(32'h396b33f5),
	.w3(32'h38994d3f),
	.w4(32'h3920a904),
	.w5(32'h39766095),
	.w6(32'h390dc830),
	.w7(32'h392cb824),
	.w8(32'h397054c1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bcbf3),
	.w1(32'h3acb9522),
	.w2(32'h3a91c487),
	.w3(32'h3b2854f7),
	.w4(32'h3adf395f),
	.w5(32'h3a4f25ac),
	.w6(32'h3ad4ca08),
	.w7(32'h3a8b425a),
	.w8(32'h39c3e7c4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee932a),
	.w1(32'h3a1da69f),
	.w2(32'h3a9d575c),
	.w3(32'h3a0aadcd),
	.w4(32'h3a4301e3),
	.w5(32'h3a83cb06),
	.w6(32'h3991a9ba),
	.w7(32'h3a1a7a92),
	.w8(32'h3a830acd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba818438),
	.w1(32'hba891efe),
	.w2(32'hba6b9a10),
	.w3(32'hb9a2a91d),
	.w4(32'hba5d11e0),
	.w5(32'hba28e579),
	.w6(32'h39a5e12a),
	.w7(32'hb9cc796a),
	.w8(32'hb9c37182),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7173de),
	.w1(32'hba8c0bac),
	.w2(32'hbb15d31f),
	.w3(32'hbb0e7fd1),
	.w4(32'hbac81e52),
	.w5(32'hbb231d7a),
	.w6(32'hbb05c44b),
	.w7(32'hbb2b501d),
	.w8(32'hbb2ddeae),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892c84a),
	.w1(32'h38ded179),
	.w2(32'hba42b019),
	.w3(32'hb806aaa8),
	.w4(32'h39177321),
	.w5(32'hba7d280d),
	.w6(32'hba09f79f),
	.w7(32'hb863efe0),
	.w8(32'hb9d83206),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861222b),
	.w1(32'hb8114869),
	.w2(32'h37e071e1),
	.w3(32'h387db68c),
	.w4(32'hb7c0bf47),
	.w5(32'h37e7aca9),
	.w6(32'hb7c4b3f0),
	.w7(32'h36b6cbfb),
	.w8(32'hb48a0879),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd5522),
	.w1(32'h3a984e6f),
	.w2(32'hb8b9e126),
	.w3(32'hb95da67b),
	.w4(32'hb95bc2bd),
	.w5(32'hba493c03),
	.w6(32'hba3b77ff),
	.w7(32'h3a1edf96),
	.w8(32'hba998735),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9475dd0),
	.w1(32'h38d804d4),
	.w2(32'h38f235d3),
	.w3(32'hb9bec241),
	.w4(32'hb7509aa0),
	.w5(32'h390b6af9),
	.w6(32'hb9969eaa),
	.w7(32'hb97907c4),
	.w8(32'h37d8a940),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9516b60),
	.w1(32'hb851b416),
	.w2(32'hba6a1b0e),
	.w3(32'hba8ef31d),
	.w4(32'hb9a413d0),
	.w5(32'hba449788),
	.w6(32'hbaebf9c7),
	.w7(32'hbaadd096),
	.w8(32'hba368401),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a4858f),
	.w1(32'hb885eeac),
	.w2(32'hb9372149),
	.w3(32'hb90945a7),
	.w4(32'hb8da4844),
	.w5(32'hb9434335),
	.w6(32'hb9217e72),
	.w7(32'hb914efdb),
	.w8(32'hb950f986),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d4d303),
	.w1(32'hb98715b7),
	.w2(32'hb9f557e3),
	.w3(32'hb96b307b),
	.w4(32'hb9b764eb),
	.w5(32'hba1da5f0),
	.w6(32'hba11e6c9),
	.w7(32'hba3dc3f6),
	.w8(32'hba2f1f9e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2003df),
	.w1(32'hba4837ff),
	.w2(32'hbaee47ce),
	.w3(32'hbad44979),
	.w4(32'hbab1b104),
	.w5(32'hbb018a72),
	.w6(32'hbb072b53),
	.w7(32'hbb0fd1d0),
	.w8(32'hbb1c6ea5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c25f4c),
	.w1(32'h3910f0ad),
	.w2(32'h394806a8),
	.w3(32'h3907a054),
	.w4(32'h390a737a),
	.w5(32'h38cb61c2),
	.w6(32'h389db475),
	.w7(32'h391cf120),
	.w8(32'h37b1b142),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918d52e),
	.w1(32'h397509ba),
	.w2(32'h395b9ca1),
	.w3(32'h385dc006),
	.w4(32'h3947d9a3),
	.w5(32'h3944b524),
	.w6(32'hb72991c8),
	.w7(32'h39086e4d),
	.w8(32'h3906bf84),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d80897),
	.w1(32'h37f40a11),
	.w2(32'hb91a669b),
	.w3(32'h38287b4c),
	.w4(32'h395c1484),
	.w5(32'h38a6c459),
	.w6(32'h394a7693),
	.w7(32'h39a7988d),
	.w8(32'h3988326f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a350f),
	.w1(32'h388a680a),
	.w2(32'h387a0211),
	.w3(32'h38234637),
	.w4(32'h37a1726f),
	.w5(32'h37f81235),
	.w6(32'h3748608f),
	.w7(32'h36e82c38),
	.w8(32'h372faa61),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3796c2a3),
	.w1(32'h37ce0f39),
	.w2(32'hba0976e3),
	.w3(32'hb997842c),
	.w4(32'hb9c1fa99),
	.w5(32'hba3950bf),
	.w6(32'hba47a120),
	.w7(32'hba5a109f),
	.w8(32'hba70939b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6399c5),
	.w1(32'hba3d125a),
	.w2(32'hba9c904c),
	.w3(32'hbaf7f282),
	.w4(32'hba8e4e65),
	.w5(32'hba5a0704),
	.w6(32'hbaf8fa40),
	.w7(32'hbad5c9e1),
	.w8(32'hba6b4a44),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a937b9b),
	.w1(32'hb9a50ab9),
	.w2(32'hba190180),
	.w3(32'h3a017cda),
	.w4(32'hba06e40e),
	.w5(32'hba923965),
	.w6(32'hba7ae435),
	.w7(32'hbad69026),
	.w8(32'hbb10cc32),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e411e1),
	.w1(32'h3a2b8013),
	.w2(32'hb859e909),
	.w3(32'hb9d26b07),
	.w4(32'h399367a4),
	.w5(32'hb99be817),
	.w6(32'hb9cf38ca),
	.w7(32'hb9348518),
	.w8(32'hb8f97405),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc3e9e),
	.w1(32'hba164b67),
	.w2(32'hba88c87e),
	.w3(32'hbaab01a5),
	.w4(32'hbab612b1),
	.w5(32'hbac2580a),
	.w6(32'hbaf59754),
	.w7(32'hbaf80d38),
	.w8(32'hbaf5a864),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38314b16),
	.w1(32'h3966c748),
	.w2(32'h3a0f4672),
	.w3(32'hb7a2d507),
	.w4(32'h39bc4243),
	.w5(32'h3a263596),
	.w6(32'h38323bfb),
	.w7(32'h398de231),
	.w8(32'h3a1cb91d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391aa131),
	.w1(32'h394c727a),
	.w2(32'h39c9e7b4),
	.w3(32'hb9168300),
	.w4(32'hb9b93a11),
	.w5(32'hb7d61d9c),
	.w6(32'hba5b83a5),
	.w7(32'hba3a936f),
	.w8(32'hb930613a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c20ddf),
	.w1(32'h39b9e814),
	.w2(32'h39a8aa78),
	.w3(32'hb7baeaea),
	.w4(32'hb93e784d),
	.w5(32'hb90425e0),
	.w6(32'hba0b1383),
	.w7(32'hba1e0ec4),
	.w8(32'hba0d2ba8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ce00f),
	.w1(32'hbb122281),
	.w2(32'hbb8ee1d2),
	.w3(32'hbb87269c),
	.w4(32'hbb7aeb74),
	.w5(32'hbba24fe6),
	.w6(32'hbb685bf3),
	.w7(32'hbb76ca2c),
	.w8(32'hbba52ac3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f574c),
	.w1(32'hb674b9e9),
	.w2(32'h34f15a67),
	.w3(32'hb5d2f385),
	.w4(32'h35799526),
	.w5(32'h36b94452),
	.w6(32'h368dd8ef),
	.w7(32'h369b92b9),
	.w8(32'h35a2e0a7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1789b),
	.w1(32'hb956386e),
	.w2(32'hbab4075a),
	.w3(32'hbabebb40),
	.w4(32'hba396659),
	.w5(32'hba88bebc),
	.w6(32'hbb1177a1),
	.w7(32'hbaed972c),
	.w8(32'hbad1ba37),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c9c9f1),
	.w1(32'hb8bce4a1),
	.w2(32'hb963c513),
	.w3(32'hb7c0c62e),
	.w4(32'hb9375cc3),
	.w5(32'hb999c657),
	.w6(32'hb792f783),
	.w7(32'hb96f16b7),
	.w8(32'hb9bbd74d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981225f),
	.w1(32'hb92907ac),
	.w2(32'hb92bf45a),
	.w3(32'hb97f8961),
	.w4(32'hb9a8d6ee),
	.w5(32'hb95edcb2),
	.w6(32'hb9d4e99f),
	.w7(32'hb9b52ca0),
	.w8(32'hb91d99e6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d45a85),
	.w1(32'h39fb7490),
	.w2(32'hb99c1d4b),
	.w3(32'hb9a89430),
	.w4(32'hb9a4cd6f),
	.w5(32'hb9580ff2),
	.w6(32'hb9db2c27),
	.w7(32'hba8cbe17),
	.w8(32'hba0a233b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c1e9),
	.w1(32'hbada285e),
	.w2(32'hba9c12d0),
	.w3(32'hbad8d44f),
	.w4(32'hba93ae16),
	.w5(32'hba3b079d),
	.w6(32'hbaba7fc4),
	.w7(32'hba110ce6),
	.w8(32'hba069dc7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fb057b),
	.w1(32'h36a53585),
	.w2(32'h37cda6ca),
	.w3(32'hb75ad69c),
	.w4(32'h37a745bf),
	.w5(32'h3795b7c4),
	.w6(32'hb8446031),
	.w7(32'hb7378f00),
	.w8(32'h380ed451),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958e823),
	.w1(32'h38c1674c),
	.w2(32'hb9a014ce),
	.w3(32'hb9e7cc25),
	.w4(32'hb9f5c877),
	.w5(32'hba3504c8),
	.w6(32'hb998b9ce),
	.w7(32'hb9b48f76),
	.w8(32'hba222919),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a43f7),
	.w1(32'hba3d4b1c),
	.w2(32'hba3ff489),
	.w3(32'h39f773ee),
	.w4(32'hba7a36c2),
	.w5(32'hb93753b4),
	.w6(32'h3a8f69ed),
	.w7(32'h39f56a28),
	.w8(32'h39444fd1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f22c9),
	.w1(32'h3a2e188d),
	.w2(32'h39935e7c),
	.w3(32'hba157565),
	.w4(32'h39b65948),
	.w5(32'h38d8cede),
	.w6(32'hba346474),
	.w7(32'h388f316d),
	.w8(32'hb825841f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b989bf),
	.w1(32'h3a096512),
	.w2(32'hbaa42b69),
	.w3(32'hbb10872a),
	.w4(32'hb9ef1faa),
	.w5(32'hbaa7f40a),
	.w6(32'hbb313422),
	.w7(32'hbb4dcfc6),
	.w8(32'hbb3cd439),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d396ae),
	.w1(32'h393c8b8d),
	.w2(32'hb9c59ec4),
	.w3(32'hb9bfb81c),
	.w4(32'hb9e17353),
	.w5(32'hb9804bc5),
	.w6(32'hba5c1594),
	.w7(32'hba94e386),
	.w8(32'hba8bd03f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a756c5),
	.w1(32'h38c5efb5),
	.w2(32'h3911188e),
	.w3(32'h3933eecb),
	.w4(32'h3902cfd4),
	.w5(32'h39594d9b),
	.w6(32'h39750203),
	.w7(32'h3947be23),
	.w8(32'h398ca0ab),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375e13bc),
	.w1(32'h33f5ed30),
	.w2(32'h36c73b33),
	.w3(32'h37404482),
	.w4(32'h362fc63b),
	.w5(32'h369c6ddb),
	.w6(32'h37549f58),
	.w7(32'h3587f300),
	.w8(32'hb7117021),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e310dd),
	.w1(32'h39636c10),
	.w2(32'h3a0e9c91),
	.w3(32'h39f3ac55),
	.w4(32'h3956f379),
	.w5(32'h3a0de189),
	.w6(32'h38f3a710),
	.w7(32'h39557abe),
	.w8(32'h39ca6095),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fc5da3),
	.w1(32'h3838fa6f),
	.w2(32'hb918571f),
	.w3(32'h389b929b),
	.w4(32'h380fa31a),
	.w5(32'hb93eb15c),
	.w6(32'h378b6ed3),
	.w7(32'h381e1144),
	.w8(32'h3881e12c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39436888),
	.w1(32'h395eabaf),
	.w2(32'h39230599),
	.w3(32'h39920ed3),
	.w4(32'h39620cc3),
	.w5(32'h393e8d42),
	.w6(32'h399f20f7),
	.w7(32'h3998fd91),
	.w8(32'h3986b6af),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21bbde),
	.w1(32'h3a21344d),
	.w2(32'h3ab80989),
	.w3(32'hba9555e7),
	.w4(32'h3a178866),
	.w5(32'h3a8140b6),
	.w6(32'hba5bcf75),
	.w7(32'h39434468),
	.w8(32'h3acc4e79),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c8762),
	.w1(32'h39c3e04a),
	.w2(32'h398f5a93),
	.w3(32'h38e71854),
	.w4(32'h3a69d914),
	.w5(32'h3a7303ce),
	.w6(32'h39674dd1),
	.w7(32'h3a44d0a7),
	.w8(32'h3a8f6b04),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38212e),
	.w1(32'h3b0bdcbd),
	.w2(32'h3af237f8),
	.w3(32'h3b2d4dcb),
	.w4(32'h3aaac5c7),
	.w5(32'h3abc5fc8),
	.w6(32'h3a9034b5),
	.w7(32'h39d0d9fd),
	.w8(32'h39a97ace),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b847bf2),
	.w1(32'h3b1840d3),
	.w2(32'h3b6b7ec6),
	.w3(32'h3b918b01),
	.w4(32'h3b1cb716),
	.w5(32'h3b18b720),
	.w6(32'h3b36ec8f),
	.w7(32'h3b172df3),
	.w8(32'h3ae37ae5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fa649),
	.w1(32'hba3dd5d6),
	.w2(32'hb8cb6af7),
	.w3(32'hba39cf65),
	.w4(32'hb95369f5),
	.w5(32'h39fb2963),
	.w6(32'hb7dbe770),
	.w7(32'h39d6eb8a),
	.w8(32'h3a675f0c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46366e),
	.w1(32'hba2659eb),
	.w2(32'hba531e6f),
	.w3(32'hba8208c0),
	.w4(32'hba400063),
	.w5(32'hba71b6df),
	.w6(32'hba65560d),
	.w7(32'hba10dc75),
	.w8(32'hba544ec1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7206f2d),
	.w1(32'hb7330e56),
	.w2(32'hb7488546),
	.w3(32'h370258aa),
	.w4(32'hb4e89966),
	.w5(32'hb626c68a),
	.w6(32'h36855f7a),
	.w7(32'hb7916dac),
	.w8(32'hb68d9d3d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875803b),
	.w1(32'hb7841c1d),
	.w2(32'hb7d3df00),
	.w3(32'h38475652),
	.w4(32'hb7c60939),
	.w5(32'hb814a54a),
	.w6(32'h3877a137),
	.w7(32'hb7d1a995),
	.w8(32'hb765ee80),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e1316a),
	.w1(32'h372547e2),
	.w2(32'h36c06355),
	.w3(32'h376f1e7d),
	.w4(32'h365d42b8),
	.w5(32'h35f516ff),
	.w6(32'h37c10ae2),
	.w7(32'h35e3cc7b),
	.w8(32'h3760816c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89ad410),
	.w1(32'h392f2644),
	.w2(32'hb8a0243d),
	.w3(32'hb9aa1bb4),
	.w4(32'h38bc727e),
	.w5(32'h386a964a),
	.w6(32'hb8e982ad),
	.w7(32'hb8142214),
	.w8(32'h39611337),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f24fe2),
	.w1(32'hb92dc2c2),
	.w2(32'hb9af3999),
	.w3(32'h3a23c923),
	.w4(32'h39a7ab19),
	.w5(32'hb8ced9da),
	.w6(32'h3a6f118a),
	.w7(32'h3a347de9),
	.w8(32'h3a36c911),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cafee8),
	.w1(32'h3b09808a),
	.w2(32'hba026bb1),
	.w3(32'hbac75f9a),
	.w4(32'hb99a0e14),
	.w5(32'hbabd2fff),
	.w6(32'hbb22231a),
	.w7(32'hb9943796),
	.w8(32'hb9c22b6f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02667c),
	.w1(32'hb9f432dc),
	.w2(32'hb9fb3980),
	.w3(32'hba737500),
	.w4(32'hba5d5cd8),
	.w5(32'hba2fa08b),
	.w6(32'hba8750ff),
	.w7(32'hba96f7cf),
	.w8(32'hba926395),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b9b917),
	.w1(32'h38a905b0),
	.w2(32'h38f3f3b9),
	.w3(32'hb8c9a2c7),
	.w4(32'hb778d89c),
	.w5(32'h38733d8c),
	.w6(32'h38a309be),
	.w7(32'h383d8973),
	.w8(32'h39df5a37),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cba90),
	.w1(32'hba9d4c97),
	.w2(32'hbb48a09c),
	.w3(32'hbb3e312d),
	.w4(32'hbb39da87),
	.w5(32'hbb871583),
	.w6(32'hbb9398e9),
	.w7(32'hbba660b5),
	.w8(32'hbbd3a5ae),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374a82),
	.w1(32'h3b502e93),
	.w2(32'h38a02ef3),
	.w3(32'h3b09ca16),
	.w4(32'h3b88deeb),
	.w5(32'h3b7a0433),
	.w6(32'h3a484b3e),
	.w7(32'h3b50b09b),
	.w8(32'h3a60db37),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9143006),
	.w1(32'hba382f6a),
	.w2(32'hba3194f0),
	.w3(32'h39d8f03c),
	.w4(32'hb84c725e),
	.w5(32'h3930efca),
	.w6(32'h3a72929d),
	.w7(32'h3a5522a6),
	.w8(32'h3aaa6106),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802f72),
	.w1(32'h3b28333d),
	.w2(32'h3b15d2ef),
	.w3(32'h3aa6099a),
	.w4(32'h3b3c76fe),
	.w5(32'h3b342749),
	.w6(32'h3af553d2),
	.w7(32'h3ad5b935),
	.w8(32'h3b06e1fa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9391fed),
	.w1(32'h39af911e),
	.w2(32'hba39252d),
	.w3(32'h3a9445bb),
	.w4(32'h38486606),
	.w5(32'hb9b0c25c),
	.w6(32'h3aa038df),
	.w7(32'hb9c7da26),
	.w8(32'hba352833),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2be5e9),
	.w1(32'hbb8e34ed),
	.w2(32'h3b004bd7),
	.w3(32'hbb16b1fb),
	.w4(32'hbbfd2e90),
	.w5(32'hbb62662f),
	.w6(32'h3a0004b9),
	.w7(32'h3b176757),
	.w8(32'hba98f477),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba596409),
	.w1(32'hb9b1176d),
	.w2(32'hbaa1af38),
	.w3(32'hb99c8a5a),
	.w4(32'h3a2ca2c0),
	.w5(32'hba9409cd),
	.w6(32'hbaccea91),
	.w7(32'hbab5d990),
	.w8(32'h394a56b5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bde78),
	.w1(32'h3abc1654),
	.w2(32'hbabbb3fc),
	.w3(32'h39ec64d9),
	.w4(32'h3ad31fa0),
	.w5(32'h398d7813),
	.w6(32'hba0a6f38),
	.w7(32'hbac64fb2),
	.w8(32'h39ceec2d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9697d04),
	.w1(32'h38e30b3b),
	.w2(32'hba428714),
	.w3(32'hb8830ea2),
	.w4(32'h39877717),
	.w5(32'hb7dc46b8),
	.w6(32'h3a0f248a),
	.w7(32'hba3554d8),
	.w8(32'h3a27cc99),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29271c),
	.w1(32'h394fec82),
	.w2(32'h38e01955),
	.w3(32'h3a39e470),
	.w4(32'h3a0aa656),
	.w5(32'h3a1ff90f),
	.w6(32'h3a1ebc0a),
	.w7(32'h39ef3377),
	.w8(32'h3aa4b72e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999f641),
	.w1(32'hb9fedf05),
	.w2(32'hba89c433),
	.w3(32'hba35516a),
	.w4(32'hb952efdc),
	.w5(32'hb91229d7),
	.w6(32'hba8e2e2b),
	.w7(32'hba453b7b),
	.w8(32'hbb41d73b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec4713),
	.w1(32'h3af0023d),
	.w2(32'h3b1575c9),
	.w3(32'hbb558a8b),
	.w4(32'h3a86b818),
	.w5(32'h3a692660),
	.w6(32'hbb0db2b8),
	.w7(32'h3ae9f397),
	.w8(32'h3b1caae2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a8d80),
	.w1(32'h3ac6782f),
	.w2(32'hb9e5397c),
	.w3(32'h3a8e446a),
	.w4(32'h3acc2ce0),
	.w5(32'h39a6c032),
	.w6(32'h3aead6ae),
	.w7(32'h38870d3c),
	.w8(32'hbb098215),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d6943),
	.w1(32'h3bc52906),
	.w2(32'h3b7a5864),
	.w3(32'h39b9ac90),
	.w4(32'h3a836387),
	.w5(32'h3a56e61e),
	.w6(32'h3b83cbcf),
	.w7(32'h3bab6f1b),
	.w8(32'hb7eb605d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0cb67),
	.w1(32'hbb0c7792),
	.w2(32'hbb964f1f),
	.w3(32'h3aff8eea),
	.w4(32'hbaf4b666),
	.w5(32'hbacfe5b1),
	.w6(32'hbb042675),
	.w7(32'hbb3fab44),
	.w8(32'hbb52a343),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933f48),
	.w1(32'h386f2235),
	.w2(32'hbafbd93d),
	.w3(32'hbaab6fb3),
	.w4(32'hba65097d),
	.w5(32'hbb997ca1),
	.w6(32'hba281116),
	.w7(32'hb98c04a2),
	.w8(32'hbb097b10),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47d76b),
	.w1(32'hbb626a03),
	.w2(32'hbaec2be5),
	.w3(32'h3a8ffd50),
	.w4(32'hbac9ac21),
	.w5(32'h3881a525),
	.w6(32'hbbe2b171),
	.w7(32'hbb133374),
	.w8(32'hba650db4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d75999),
	.w1(32'h3a6aedac),
	.w2(32'hb9d58f44),
	.w3(32'h3a8d2b54),
	.w4(32'h3ad13ed5),
	.w5(32'h3a206cb3),
	.w6(32'h392b2275),
	.w7(32'hb9e6e41a),
	.w8(32'hbad4c26a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bc9a0),
	.w1(32'h3a295e5f),
	.w2(32'h39eeebf2),
	.w3(32'hbaceecac),
	.w4(32'hba217e1e),
	.w5(32'hbabbdf6a),
	.w6(32'hbadd65f4),
	.w7(32'hba99fa20),
	.w8(32'hbb25032e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e4733),
	.w1(32'hbb559ee4),
	.w2(32'h3afa6668),
	.w3(32'hbb394726),
	.w4(32'hbb6751b6),
	.w5(32'hbb43fe38),
	.w6(32'hbadf813a),
	.w7(32'h3b4513c6),
	.w8(32'h38c8f02b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a734),
	.w1(32'h3aa977cf),
	.w2(32'h3a8dc2c4),
	.w3(32'h39e5d7a3),
	.w4(32'h3a22362f),
	.w5(32'h3a2bd311),
	.w6(32'h3b2b61f0),
	.w7(32'h3a2772fd),
	.w8(32'h3b43fafd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b8497),
	.w1(32'hba370cee),
	.w2(32'hbab93e69),
	.w3(32'hba375854),
	.w4(32'hb9361a78),
	.w5(32'h38b94116),
	.w6(32'h39b5dfbc),
	.w7(32'hba5dfb12),
	.w8(32'hbba97023),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fcd60),
	.w1(32'hbb84a879),
	.w2(32'hbb0ded8e),
	.w3(32'hbb0564ea),
	.w4(32'hbaad1013),
	.w5(32'h3ab4eed8),
	.w6(32'hbbf1bed5),
	.w7(32'hbb58637e),
	.w8(32'h3a8413aa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule