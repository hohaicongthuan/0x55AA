module layer_10_featuremap_86(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9961ce),
	.w1(32'h3adb7ad0),
	.w2(32'hbb1b1467),
	.w3(32'hbb60058d),
	.w4(32'hb9ebb529),
	.w5(32'hbb94fd5c),
	.w6(32'h38f653f9),
	.w7(32'hbb1ab556),
	.w8(32'hbc45b612),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08fa7),
	.w1(32'hba221d1f),
	.w2(32'hb9490454),
	.w3(32'hbb7bd296),
	.w4(32'hbaa4c094),
	.w5(32'h3b308d41),
	.w6(32'h3bdfce7a),
	.w7(32'h3bdc0879),
	.w8(32'hbb6ec9d3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9f351),
	.w1(32'hbb702211),
	.w2(32'hbacd9eab),
	.w3(32'h3d4e3dbd),
	.w4(32'h3c923c7a),
	.w5(32'h3ad9a57f),
	.w6(32'h3c2178e0),
	.w7(32'hba96d1bb),
	.w8(32'hbbb5d6a3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd1f7),
	.w1(32'hbb97c187),
	.w2(32'hbb1c0cec),
	.w3(32'hbb32b578),
	.w4(32'hbbf56387),
	.w5(32'hbb6c0ec5),
	.w6(32'hbba6fc53),
	.w7(32'h3a35567c),
	.w8(32'hbc06d945),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee2ef6),
	.w1(32'hbc1fc0f4),
	.w2(32'hbc1c8ac1),
	.w3(32'hbb4813e7),
	.w4(32'h3ae83a18),
	.w5(32'h3abcfc48),
	.w6(32'h3910b6cb),
	.w7(32'h3b8cab2f),
	.w8(32'h3b77c5bc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3d1e4),
	.w1(32'h3a86f9cd),
	.w2(32'h3bddfc2b),
	.w3(32'hbb331f3a),
	.w4(32'hbade5849),
	.w5(32'hbb9e39c4),
	.w6(32'h3bc4c533),
	.w7(32'hba0bb725),
	.w8(32'hbc4ffe6a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb705fc3),
	.w1(32'hbbcbe4cf),
	.w2(32'hba56f4b5),
	.w3(32'h3b02ec12),
	.w4(32'h3bfc7181),
	.w5(32'hbbcb1b04),
	.w6(32'h3b3813f4),
	.w7(32'h3bb1e732),
	.w8(32'h3b27df77),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a457b),
	.w1(32'hba687c72),
	.w2(32'h3c2e7fdf),
	.w3(32'h3bdb4188),
	.w4(32'h3c6e3d71),
	.w5(32'h3ab640f2),
	.w6(32'hbb572cc8),
	.w7(32'h3bd5b6a0),
	.w8(32'hbc90a702),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ead3),
	.w1(32'h3b8aac89),
	.w2(32'h3c7e6bf3),
	.w3(32'hbbbe06ce),
	.w4(32'hbb9573b8),
	.w5(32'h3bac09b7),
	.w6(32'h3b2cdb07),
	.w7(32'hbc07c7b3),
	.w8(32'h3995cdc3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12a290),
	.w1(32'hbb445a7f),
	.w2(32'hbbd92b9f),
	.w3(32'hbb91cfe3),
	.w4(32'hbc0562c6),
	.w5(32'hbc109ac8),
	.w6(32'hbbdafbae),
	.w7(32'h3aa6b42c),
	.w8(32'h3b64e9b7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28488),
	.w1(32'h3b11ea76),
	.w2(32'hba3be49e),
	.w3(32'h398fa26e),
	.w4(32'h3bd1b5ad),
	.w5(32'h3a784f79),
	.w6(32'hbaff88ff),
	.w7(32'hb9d42f08),
	.w8(32'h3b1427a5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d1f1b),
	.w1(32'hb9986345),
	.w2(32'hbb5ebb2d),
	.w3(32'hbb85613f),
	.w4(32'h3b250553),
	.w5(32'h3aee5d88),
	.w6(32'h3a8b15dc),
	.w7(32'h3b921a07),
	.w8(32'h3c21545c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13f1d0),
	.w1(32'hbaf85305),
	.w2(32'h3b138b29),
	.w3(32'h3c2d09fb),
	.w4(32'hbb7b7b77),
	.w5(32'h3ab9becf),
	.w6(32'h3a719836),
	.w7(32'hbbfbe695),
	.w8(32'hbbf5299d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054d8d),
	.w1(32'hb98ccc9e),
	.w2(32'h3ba56cae),
	.w3(32'hbb7b7207),
	.w4(32'hb87f44ee),
	.w5(32'hb9a7b086),
	.w6(32'h3b48222e),
	.w7(32'hb9002802),
	.w8(32'hbad960e0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43ee5d),
	.w1(32'hba012f52),
	.w2(32'h3b190886),
	.w3(32'hbb3bd015),
	.w4(32'hbc0532b2),
	.w5(32'hbc1071a6),
	.w6(32'hbc2c1729),
	.w7(32'hbc2ad57a),
	.w8(32'hbbaea1b3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4266),
	.w1(32'hbafa4219),
	.w2(32'hbad2292d),
	.w3(32'hbbab2ba5),
	.w4(32'h3b135702),
	.w5(32'hbc4e6e0e),
	.w6(32'hbc238d2d),
	.w7(32'h3b737776),
	.w8(32'hbc50f1ac),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd8c20),
	.w1(32'hb9a4c44c),
	.w2(32'hbb96acdc),
	.w3(32'hbacd3251),
	.w4(32'h389fb3eb),
	.w5(32'h39e097b4),
	.w6(32'h3a962841),
	.w7(32'h3c1d0c35),
	.w8(32'h3b5bfea2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a918da),
	.w1(32'h3b8bcccb),
	.w2(32'hbc46f487),
	.w3(32'h3aa0368a),
	.w4(32'h3bbc9262),
	.w5(32'hbb83ad2b),
	.w6(32'hbc6b7073),
	.w7(32'h3a933ae7),
	.w8(32'hbbbd1407),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10adc2),
	.w1(32'h3b85946c),
	.w2(32'hbaa669f2),
	.w3(32'h3be0ec2c),
	.w4(32'h3c718410),
	.w5(32'hbc0d4501),
	.w6(32'h3bb62b5e),
	.w7(32'hbc02f002),
	.w8(32'hbb934d5e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15048f),
	.w1(32'h3bd19d91),
	.w2(32'hbc217896),
	.w3(32'hbaa48f12),
	.w4(32'hbac0c7b2),
	.w5(32'h3c4adc73),
	.w6(32'hb9bd9e38),
	.w7(32'hbc09046d),
	.w8(32'hbab84e7f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ceada),
	.w1(32'h3a0b09f4),
	.w2(32'h3b41ee26),
	.w3(32'h3a97a7ab),
	.w4(32'hbb3dd390),
	.w5(32'h3c52577d),
	.w6(32'h3a203eed),
	.w7(32'hbbd23cb7),
	.w8(32'hbb993777),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b7f0a),
	.w1(32'h3b1d8b3e),
	.w2(32'hbbeafc9b),
	.w3(32'hbb2bae1a),
	.w4(32'h3ae775b2),
	.w5(32'hbbbdc056),
	.w6(32'h3ab8f910),
	.w7(32'h3a939593),
	.w8(32'h3b759654),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b179a),
	.w1(32'hbace1157),
	.w2(32'h3b2286ab),
	.w3(32'hbb2c442b),
	.w4(32'hbc1923ac),
	.w5(32'hbbf5a402),
	.w6(32'h3b07d58c),
	.w7(32'hbbd65fa1),
	.w8(32'hbc1aead4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805ac6),
	.w1(32'h3b163a5e),
	.w2(32'hbc8bd03c),
	.w3(32'hbc0f1f4d),
	.w4(32'hbc5b822f),
	.w5(32'h3a16a333),
	.w6(32'hbbcfe5f1),
	.w7(32'h3c3106a8),
	.w8(32'hbc83db1c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f805),
	.w1(32'hbc113e8e),
	.w2(32'h3cc408b0),
	.w3(32'hbc344ec6),
	.w4(32'hbc447497),
	.w5(32'hbbcc37a6),
	.w6(32'h3b97e9c9),
	.w7(32'h3b11b6ee),
	.w8(32'hbc979387),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8e64),
	.w1(32'hbc1318c3),
	.w2(32'h3b6c6795),
	.w3(32'h3c1206c2),
	.w4(32'h3c607dd3),
	.w5(32'hba8ca663),
	.w6(32'h3aad7bd0),
	.w7(32'h3c12f960),
	.w8(32'hbbaef0fa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf3e85),
	.w1(32'h3bf64052),
	.w2(32'h3bdfa926),
	.w3(32'hbb06080f),
	.w4(32'h3bb0963d),
	.w5(32'h3b7bd4a1),
	.w6(32'h3b66aa33),
	.w7(32'hba8a4cc9),
	.w8(32'hbb58ea63),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95576d),
	.w1(32'hbbf7a772),
	.w2(32'h3bc70838),
	.w3(32'h3ae1dd05),
	.w4(32'h3c0e070e),
	.w5(32'h3b8e0353),
	.w6(32'h3b5246f0),
	.w7(32'h3b804056),
	.w8(32'h3a98fc1b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e4e01),
	.w1(32'hba44069a),
	.w2(32'hb9f56c42),
	.w3(32'hbb719851),
	.w4(32'h3a390bf5),
	.w5(32'h3b442d54),
	.w6(32'h38c262c6),
	.w7(32'hbac73ef2),
	.w8(32'h3b6e18c2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31f6fc),
	.w1(32'hbc8f8ce4),
	.w2(32'hbbe3c85d),
	.w3(32'hbc159755),
	.w4(32'h3b1693c2),
	.w5(32'hbc5f1ecc),
	.w6(32'h3c06df5c),
	.w7(32'h3b4f7ce3),
	.w8(32'hbbb152cf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00c36),
	.w1(32'hbbce402a),
	.w2(32'hbbeefa97),
	.w3(32'h3b0aa864),
	.w4(32'hbbdd3fd6),
	.w5(32'hba221f54),
	.w6(32'hb9aa6e55),
	.w7(32'hb96de2fa),
	.w8(32'h3bb57028),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ffe9e),
	.w1(32'hba5eaa13),
	.w2(32'h3b33f592),
	.w3(32'hb8d7d8aa),
	.w4(32'h3b51b139),
	.w5(32'h3b3ddcc9),
	.w6(32'h3b443fc5),
	.w7(32'hbae1de93),
	.w8(32'hbb857fa8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c0a93),
	.w1(32'hbbbcc974),
	.w2(32'hbb706a0d),
	.w3(32'hbb282166),
	.w4(32'hbbb00fed),
	.w5(32'h3b837597),
	.w6(32'hbba28169),
	.w7(32'hba778aae),
	.w8(32'hbbb47d7c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94381),
	.w1(32'hbb12db5a),
	.w2(32'hbb5dbf22),
	.w3(32'hbb3c85bb),
	.w4(32'hbb536b04),
	.w5(32'hbb05c52a),
	.w6(32'hbab22a61),
	.w7(32'hbc2d04e6),
	.w8(32'h3a7486a2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8765d),
	.w1(32'hba03f262),
	.w2(32'hbbb7fa88),
	.w3(32'hbb7d9bd2),
	.w4(32'hba5891b4),
	.w5(32'hbb1923e4),
	.w6(32'h3b5af8fc),
	.w7(32'hbbc6059f),
	.w8(32'hbc2812ae),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1048d3),
	.w1(32'h3bed3972),
	.w2(32'hbb4176f7),
	.w3(32'hbb5f2e31),
	.w4(32'hb9c4b07b),
	.w5(32'h3b0d1288),
	.w6(32'h3ce8d96e),
	.w7(32'h3af91342),
	.w8(32'h3b41f9b4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ea0b5),
	.w1(32'h3ae28510),
	.w2(32'h3c02eec5),
	.w3(32'hbcc8a567),
	.w4(32'hbca74575),
	.w5(32'h3d339d85),
	.w6(32'hbc83eac3),
	.w7(32'hbc7e566f),
	.w8(32'h3ca92781),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60497f),
	.w1(32'h3b01eede),
	.w2(32'h3ba912cf),
	.w3(32'h3bcb61ce),
	.w4(32'hbb0832c2),
	.w5(32'hbb957816),
	.w6(32'h3bd9335e),
	.w7(32'h3b8517db),
	.w8(32'hbbf94287),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b2d6a),
	.w1(32'hbbb16add),
	.w2(32'hba9f20c3),
	.w3(32'hba8a436f),
	.w4(32'hba91f779),
	.w5(32'hbc301a56),
	.w6(32'h3c45384f),
	.w7(32'h3bb86dc4),
	.w8(32'hbc5fdca5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813cf4),
	.w1(32'hba0699a9),
	.w2(32'hbb1032c5),
	.w3(32'hbad60601),
	.w4(32'hba21a63d),
	.w5(32'hbb30619b),
	.w6(32'h3a9c23f8),
	.w7(32'h3b96a050),
	.w8(32'h3bca5b0c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967faac),
	.w1(32'h3b8543d2),
	.w2(32'h3a887e97),
	.w3(32'h3c109c16),
	.w4(32'h3b10c04b),
	.w5(32'hbb85afa5),
	.w6(32'hb8e918df),
	.w7(32'hbb1dbc40),
	.w8(32'h3a694002),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ab74f),
	.w1(32'h39c291d4),
	.w2(32'h3ab62caa),
	.w3(32'h39ca68ef),
	.w4(32'h3c887bc8),
	.w5(32'hbb270adc),
	.w6(32'h39046430),
	.w7(32'hbb24e9ff),
	.w8(32'hbc573c07),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f0d5e),
	.w1(32'h3a27734a),
	.w2(32'hbb247bba),
	.w3(32'hb9e2a9ab),
	.w4(32'hbb88bc2b),
	.w5(32'hbab61f18),
	.w6(32'hbb0e7cd3),
	.w7(32'hbb20980a),
	.w8(32'h39bc4c10),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddcbc5),
	.w1(32'hba127f84),
	.w2(32'hbbc6bdd2),
	.w3(32'h3b2432f7),
	.w4(32'h3bae7261),
	.w5(32'hbc430984),
	.w6(32'hbc00925b),
	.w7(32'h3cdb39c4),
	.w8(32'hbc852f97),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd45fec),
	.w1(32'h3be9745f),
	.w2(32'h3ac812f8),
	.w3(32'hbb44d94a),
	.w4(32'hbba097b9),
	.w5(32'h3c618437),
	.w6(32'hbc1c246e),
	.w7(32'hbc0ba125),
	.w8(32'hbb81ace0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba71f93),
	.w1(32'hba707d96),
	.w2(32'hbbd92b2e),
	.w3(32'hbc1a48f6),
	.w4(32'hbc372243),
	.w5(32'hbbd736ee),
	.w6(32'hbcc0cbff),
	.w7(32'hbc021664),
	.w8(32'hbc56efe3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797760),
	.w1(32'hbbbf183f),
	.w2(32'h3935421e),
	.w3(32'hbb1b14b9),
	.w4(32'h3b95c6b5),
	.w5(32'h3b3fd841),
	.w6(32'hbb095f5d),
	.w7(32'h3b9ce884),
	.w8(32'hbc282be0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227d58),
	.w1(32'h3b6b67b8),
	.w2(32'hbc0e7643),
	.w3(32'h3c285eb2),
	.w4(32'h3c79cfd1),
	.w5(32'h3c03a37d),
	.w6(32'hbbe43c1d),
	.w7(32'hbb63bd1e),
	.w8(32'hbbb6fc8e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba353268),
	.w1(32'hbba11411),
	.w2(32'h3c30ff9d),
	.w3(32'hbb1b26fd),
	.w4(32'hbb9addfa),
	.w5(32'hba44c2dd),
	.w6(32'hb8b3b40e),
	.w7(32'hbb1e05f0),
	.w8(32'hbb5ff8e5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaed212),
	.w1(32'hbb53793b),
	.w2(32'h3aa87d60),
	.w3(32'hbc3971cb),
	.w4(32'hbb5ffb62),
	.w5(32'hbba5e9c9),
	.w6(32'h39a5cec2),
	.w7(32'hb9cc39d1),
	.w8(32'hbab81206),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa51fc),
	.w1(32'hbc12d84e),
	.w2(32'hbaa919bd),
	.w3(32'hbadf3ee4),
	.w4(32'hb9d9a06f),
	.w5(32'hb9a5505e),
	.w6(32'h37d69127),
	.w7(32'h39446e0b),
	.w8(32'hba96e5bf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39e090),
	.w1(32'hbc19e371),
	.w2(32'hbbe1e99b),
	.w3(32'hbc513b9c),
	.w4(32'hbb269ca7),
	.w5(32'hbc1bddd8),
	.w6(32'hbc3b1eb2),
	.w7(32'hbaddde2f),
	.w8(32'hbc53bb1a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab38c6),
	.w1(32'hbb804e13),
	.w2(32'hba03e863),
	.w3(32'h3a8e3abb),
	.w4(32'hbba9d46b),
	.w5(32'h3c2801de),
	.w6(32'h3b734a87),
	.w7(32'hbb5932ef),
	.w8(32'hbb9aeeac),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43000f),
	.w1(32'hbc4712b1),
	.w2(32'hbc88d23d),
	.w3(32'h3bfd7a87),
	.w4(32'h3ba4404f),
	.w5(32'hbac484a0),
	.w6(32'hbbeace4a),
	.w7(32'h3b134992),
	.w8(32'hbc8223f9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a857),
	.w1(32'h3a0af4df),
	.w2(32'hbb91f5cf),
	.w3(32'h3c3e40f5),
	.w4(32'hbb59c530),
	.w5(32'hba53fe90),
	.w6(32'hbb1637dc),
	.w7(32'h3b1e030f),
	.w8(32'hbbcf748d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab05214),
	.w1(32'h3a99607d),
	.w2(32'hbb3854ec),
	.w3(32'h3b0e58ac),
	.w4(32'hbaf000b1),
	.w5(32'hbc832857),
	.w6(32'hbb87d982),
	.w7(32'h3ab90f83),
	.w8(32'h3b904663),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db343b9),
	.w1(32'hb9f6c3ca),
	.w2(32'h3b7f3504),
	.w3(32'h3a078e55),
	.w4(32'hb8f9823a),
	.w5(32'h3bd59a62),
	.w6(32'hbc633485),
	.w7(32'hbc0a0ff4),
	.w8(32'hbb7e8511),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d29e40),
	.w1(32'h3bd2e9b3),
	.w2(32'hbb83eb9c),
	.w3(32'hbc6fae1b),
	.w4(32'hb8ff9c71),
	.w5(32'h3b8a9c4e),
	.w6(32'h3c1f36a7),
	.w7(32'h3acbabe5),
	.w8(32'hbc8dd64a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae94f5),
	.w1(32'h3c2b4dd1),
	.w2(32'h3ae7156c),
	.w3(32'h3b993cfe),
	.w4(32'h39b2113f),
	.w5(32'hbb6145da),
	.w6(32'hbae3d7da),
	.w7(32'hbb9904ff),
	.w8(32'h3b2fd0cd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796304),
	.w1(32'hbafa7273),
	.w2(32'h3b2ced62),
	.w3(32'hb99bea28),
	.w4(32'hbb208897),
	.w5(32'hbb42a235),
	.w6(32'hbb77eb34),
	.w7(32'hbc4368f3),
	.w8(32'hbb8693a4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15fada),
	.w1(32'h39440f18),
	.w2(32'h3bbcf0f8),
	.w3(32'h3b1653e7),
	.w4(32'h3bafafb7),
	.w5(32'hb9391838),
	.w6(32'hbbc9ff7d),
	.w7(32'h3bc6d8d1),
	.w8(32'hba8675cd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd877b3),
	.w1(32'hbbe81a5a),
	.w2(32'hbaac126a),
	.w3(32'h3b2bd5c1),
	.w4(32'hbb01e962),
	.w5(32'hbd865430),
	.w6(32'hbba93d5a),
	.w7(32'h3a81d5a1),
	.w8(32'hbb2f8be4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d83e),
	.w1(32'hbc0dab2e),
	.w2(32'hbb2e386f),
	.w3(32'hbc956908),
	.w4(32'hbb7d09ab),
	.w5(32'h3b7fd7f3),
	.w6(32'hbaff7fc2),
	.w7(32'h3bbc852d),
	.w8(32'hbaf99179),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17c594),
	.w1(32'h3d4d470f),
	.w2(32'hbdb74bd2),
	.w3(32'hbc2cb30d),
	.w4(32'h3c040d6f),
	.w5(32'h3c428821),
	.w6(32'hbbfcd7f4),
	.w7(32'hbbe04ead),
	.w8(32'h3af29cea),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28ccfe),
	.w1(32'hbc1d8881),
	.w2(32'h3af3362e),
	.w3(32'h3af82c8f),
	.w4(32'hbb022abc),
	.w5(32'hbc604695),
	.w6(32'h3ad29739),
	.w7(32'hbc4a7978),
	.w8(32'h3c1edf60),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba866139),
	.w1(32'hbbee89ea),
	.w2(32'h3b83a566),
	.w3(32'h3aba907a),
	.w4(32'h39719fd5),
	.w5(32'h377f7120),
	.w6(32'hbd2e31e1),
	.w7(32'hbc9e4020),
	.w8(32'hbc261a80),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc733367),
	.w1(32'hbbae1b23),
	.w2(32'hbc74d53e),
	.w3(32'hbb95df71),
	.w4(32'h3cee370a),
	.w5(32'hbca3bea7),
	.w6(32'h3b0b3ab2),
	.w7(32'h3cbd22b9),
	.w8(32'hbba77d11),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0c31),
	.w1(32'h3d2227ef),
	.w2(32'hbbd8dff2),
	.w3(32'hbc72f929),
	.w4(32'hbbaaeab9),
	.w5(32'hbb1f20a9),
	.w6(32'hbb611ec5),
	.w7(32'hbc292ce2),
	.w8(32'hbc83c3e5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a6c9c),
	.w1(32'h3c8cc916),
	.w2(32'h3a8df7f6),
	.w3(32'h3aed346f),
	.w4(32'h3ad0ceff),
	.w5(32'hbbdbc100),
	.w6(32'hbbb39077),
	.w7(32'hbc8f2252),
	.w8(32'hbc230bf8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce73e8),
	.w1(32'hbb350614),
	.w2(32'h3c4fb62c),
	.w3(32'hbba082d5),
	.w4(32'hbc1b07fc),
	.w5(32'hbb2fb4cb),
	.w6(32'h39afb113),
	.w7(32'hbb852ba7),
	.w8(32'hbcca6dc1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb57670),
	.w1(32'hbc7961f4),
	.w2(32'h3b339f99),
	.w3(32'h3b7e567e),
	.w4(32'h3c86790b),
	.w5(32'hbb4a9b6e),
	.w6(32'h3bf6ec3c),
	.w7(32'hbc542ed8),
	.w8(32'hba838007),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd5135),
	.w1(32'h3aaf8c2e),
	.w2(32'h3b90fd39),
	.w3(32'hbab2120b),
	.w4(32'h3a2d411a),
	.w5(32'hbc82a8ed),
	.w6(32'hba0f6644),
	.w7(32'hbc043071),
	.w8(32'hbab4cbd7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd791aa4),
	.w1(32'h3a0782d4),
	.w2(32'hbaefdb3d),
	.w3(32'hbb9590ac),
	.w4(32'hbabb5127),
	.w5(32'hbcb12fa5),
	.w6(32'hba8cfafb),
	.w7(32'h3b839566),
	.w8(32'h3aceab53),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ad49),
	.w1(32'h39b83704),
	.w2(32'h3d10ec8e),
	.w3(32'hbb3ebe66),
	.w4(32'h3b41c21b),
	.w5(32'hbac1f78c),
	.w6(32'hbccc8353),
	.w7(32'h3b85adc9),
	.w8(32'hbbb51fa8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919afff),
	.w1(32'hbb35a83e),
	.w2(32'hbaf8f5b7),
	.w3(32'h3c77e25f),
	.w4(32'hbd8e8f6e),
	.w5(32'h3c0e56f8),
	.w6(32'hbb8a0807),
	.w7(32'h3b11fd00),
	.w8(32'hbc172a4e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba5ab9),
	.w1(32'hba92c0d1),
	.w2(32'hbab3dedb),
	.w3(32'h3a868cf8),
	.w4(32'h3c1cff3d),
	.w5(32'hbab5ed97),
	.w6(32'hbd3bf417),
	.w7(32'hbc359bdb),
	.w8(32'hbcd632cc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f38eb),
	.w1(32'h3d200cf1),
	.w2(32'hbb84963e),
	.w3(32'hbb2c3aff),
	.w4(32'h3b858c29),
	.w5(32'h3b8b66b1),
	.w6(32'hbc34c5c2),
	.w7(32'h3ba57547),
	.w8(32'hbb3d497e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202258),
	.w1(32'hbbae7655),
	.w2(32'h3b91ea0f),
	.w3(32'hbd3eb3ba),
	.w4(32'hbbfcfe3e),
	.w5(32'h3c1cc805),
	.w6(32'hbba5cb7f),
	.w7(32'h3d19290d),
	.w8(32'h3c95787f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b2978),
	.w1(32'hbbf610ea),
	.w2(32'hbb1671fb),
	.w3(32'hbc112784),
	.w4(32'h3ade9b7e),
	.w5(32'hbc033ac6),
	.w6(32'hbb1cb73d),
	.w7(32'hbbb9996c),
	.w8(32'hbc4ab0f0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4302c5),
	.w1(32'h3b21c8ed),
	.w2(32'h3bd11a28),
	.w3(32'hbc05a6c5),
	.w4(32'hbc670b62),
	.w5(32'hbbd472fa),
	.w6(32'h3b96d4c3),
	.w7(32'hbcc71374),
	.w8(32'h3a647ebc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e710b5),
	.w1(32'hbc0c7434),
	.w2(32'h3b31cec1),
	.w3(32'h3b9323ef),
	.w4(32'hbc21ec21),
	.w5(32'hb9b70bbe),
	.w6(32'h3c00159f),
	.w7(32'hba2c2cae),
	.w8(32'hba0e7b1b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e2bff),
	.w1(32'h3bf230cc),
	.w2(32'hbb391a0a),
	.w3(32'h3ba7114f),
	.w4(32'h3bd279b2),
	.w5(32'h3b5b96a2),
	.w6(32'hbbea00cc),
	.w7(32'hbb89d34d),
	.w8(32'hbb8be093),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0b8fb),
	.w1(32'h3c9baca1),
	.w2(32'h3bead443),
	.w3(32'h3ce34594),
	.w4(32'hbbccebc9),
	.w5(32'h3b753ca4),
	.w6(32'h3a881f9e),
	.w7(32'hbc06de3e),
	.w8(32'h3b5a0215),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27145),
	.w1(32'hbb3e2b17),
	.w2(32'h3a9d8b08),
	.w3(32'h3bc3ddfd),
	.w4(32'h3b122449),
	.w5(32'h3b46e369),
	.w6(32'hbb58973f),
	.w7(32'hbaada585),
	.w8(32'h3aa051dc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4e625),
	.w1(32'h3b5e840e),
	.w2(32'hbcc4cb11),
	.w3(32'h3b8826a4),
	.w4(32'h3ca8d181),
	.w5(32'hbaf31a0c),
	.w6(32'hbb479c2d),
	.w7(32'hba148073),
	.w8(32'h3b612cd7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb2275),
	.w1(32'h3ac38a2a),
	.w2(32'hbb56395e),
	.w3(32'hbb08e074),
	.w4(32'hba886e58),
	.w5(32'h3b56efac),
	.w6(32'hba3999b4),
	.w7(32'h3cfac6a1),
	.w8(32'hbacb8825),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f07d),
	.w1(32'h3d11d03a),
	.w2(32'h3c16ba82),
	.w3(32'hbbf391e0),
	.w4(32'hbb8fb306),
	.w5(32'h3a9df1e4),
	.w6(32'hba99eb70),
	.w7(32'hbbea924d),
	.w8(32'hb8dea634),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c208),
	.w1(32'hbace60b7),
	.w2(32'h3b4f5fe8),
	.w3(32'hba0badec),
	.w4(32'h39afb5b7),
	.w5(32'h3c7f9748),
	.w6(32'hb9d066f3),
	.w7(32'hbb3d0a31),
	.w8(32'h3ad558bf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52dcbf),
	.w1(32'hba935848),
	.w2(32'h3adbe4f1),
	.w3(32'hbb8dbd94),
	.w4(32'hba0b817e),
	.w5(32'h39a7c68f),
	.w6(32'hbc128da3),
	.w7(32'hbc0d6f4f),
	.w8(32'hbbd6957c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b30ed),
	.w1(32'h3bf95769),
	.w2(32'h3b04aad9),
	.w3(32'h3bc79fe7),
	.w4(32'h3b16caa2),
	.w5(32'hba084f68),
	.w6(32'hbbceb969),
	.w7(32'hbb0de46c),
	.w8(32'hbbc06ab1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb270f8),
	.w1(32'hba9a4926),
	.w2(32'hba3fd20b),
	.w3(32'h3ad6bd56),
	.w4(32'hba4f2636),
	.w5(32'h3a110042),
	.w6(32'h3c929421),
	.w7(32'h392eb2af),
	.w8(32'hbb61df31),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a9cd),
	.w1(32'hb9c3ae9e),
	.w2(32'hbb541c26),
	.w3(32'hbc04fe97),
	.w4(32'hbb5679ab),
	.w5(32'hbca2ba87),
	.w6(32'hbbb7598f),
	.w7(32'hbbb13756),
	.w8(32'hbc22d03d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9af19),
	.w1(32'h3b195e44),
	.w2(32'h3b967ac4),
	.w3(32'hbc1ca49b),
	.w4(32'h3ac995f4),
	.w5(32'hbb408e05),
	.w6(32'hbbadefe5),
	.w7(32'hbb2df56a),
	.w8(32'hbbeba6cc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48631c),
	.w1(32'h3c745e52),
	.w2(32'hbcec325d),
	.w3(32'h36165c8e),
	.w4(32'h3b833c03),
	.w5(32'hbacc8515),
	.w6(32'hbc0cdac0),
	.w7(32'hbbb5d433),
	.w8(32'hbc424887),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca88f5),
	.w1(32'hba3aa4a3),
	.w2(32'hbb4c5724),
	.w3(32'hbbbf54f6),
	.w4(32'hbb6cfb28),
	.w5(32'hbab0d8f0),
	.w6(32'h39cb0442),
	.w7(32'h3b9f735d),
	.w8(32'h3c3e20ae),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66875e),
	.w1(32'hba23a1e2),
	.w2(32'hb984ab01),
	.w3(32'h3bcf5f96),
	.w4(32'h3c038dfd),
	.w5(32'hbc31e10e),
	.w6(32'h3c30abf2),
	.w7(32'h3ba2c749),
	.w8(32'h3b2733ec),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994f6c7),
	.w1(32'h3cebb8b6),
	.w2(32'hba876228),
	.w3(32'h3cf7fdbf),
	.w4(32'hb99ff5f8),
	.w5(32'hbb413416),
	.w6(32'hbb1d1b83),
	.w7(32'h3ae63409),
	.w8(32'h38a1aec7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0c09f),
	.w1(32'hbb9c60b8),
	.w2(32'hbbb433ac),
	.w3(32'h39fe121a),
	.w4(32'h3b99d6e0),
	.w5(32'hbb1a430a),
	.w6(32'hbc04a4e8),
	.w7(32'hbbe510e3),
	.w8(32'h3b2f4f63),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3887d1),
	.w1(32'hbca14d9f),
	.w2(32'hbc1dc088),
	.w3(32'hbb9f8d6d),
	.w4(32'hbc3be088),
	.w5(32'hbc264282),
	.w6(32'hbb8865f6),
	.w7(32'h3b6c2902),
	.w8(32'hbd0b31f5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc238406),
	.w1(32'h3b2402e5),
	.w2(32'h3caf2526),
	.w3(32'hbc0a8ae6),
	.w4(32'hba9dadb9),
	.w5(32'h3cfe1065),
	.w6(32'h3a4aee87),
	.w7(32'hbc890e3c),
	.w8(32'h3c1bcc96),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d04fd),
	.w1(32'h3bc5e875),
	.w2(32'h3b7bb232),
	.w3(32'hbba6d995),
	.w4(32'hbc4caf94),
	.w5(32'h3abddaaa),
	.w6(32'h3a234dd9),
	.w7(32'hbb124424),
	.w8(32'hbb743113),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b6e7),
	.w1(32'hbb467ebf),
	.w2(32'hbc735f16),
	.w3(32'hbb386141),
	.w4(32'hbba6da2b),
	.w5(32'hbaa40e6e),
	.w6(32'hbcac2043),
	.w7(32'hbbaa4efc),
	.w8(32'hbb4bf296),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc458651),
	.w1(32'hba8a63ca),
	.w2(32'h3cd4d4ba),
	.w3(32'h3af8b205),
	.w4(32'hbbfe4fd5),
	.w5(32'h3b539054),
	.w6(32'hbc8182d2),
	.w7(32'hbbabf0d5),
	.w8(32'h3c17c2da),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd57632),
	.w1(32'h3a4c6d1f),
	.w2(32'h3c9643f1),
	.w3(32'h3913879d),
	.w4(32'hba41b3d5),
	.w5(32'h3989b5a8),
	.w6(32'hba0e9b51),
	.w7(32'hbaeda7cc),
	.w8(32'h3b6bc52a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a431981),
	.w1(32'h3d162c41),
	.w2(32'h3bd6ef8b),
	.w3(32'hbc0b4760),
	.w4(32'hbab4ab88),
	.w5(32'h3c2c5d4b),
	.w6(32'hbb19d3e3),
	.w7(32'hbbefc40e),
	.w8(32'h3aca53f4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0467dd),
	.w1(32'h3b1d19e9),
	.w2(32'h39f6f9f0),
	.w3(32'h3a3e55e5),
	.w4(32'h3b3fa664),
	.w5(32'h3b0fcb33),
	.w6(32'hbb8be866),
	.w7(32'hbb80bc37),
	.w8(32'hba4f11b3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeff52a),
	.w1(32'h3af3df0c),
	.w2(32'h3b52f256),
	.w3(32'hbb26c52b),
	.w4(32'hb7ebd73b),
	.w5(32'h39981249),
	.w6(32'h3a6f7e12),
	.w7(32'h38d23308),
	.w8(32'h39870adb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9ccda),
	.w1(32'h3acd3d7b),
	.w2(32'h3b8315e7),
	.w3(32'hbb516c4c),
	.w4(32'hb9a59d46),
	.w5(32'hbb123ad7),
	.w6(32'hba4b00bc),
	.w7(32'hbb1398c6),
	.w8(32'hbb15716e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c282d),
	.w1(32'h3af7fc42),
	.w2(32'hbb539ad3),
	.w3(32'h3bcfb425),
	.w4(32'hb925e816),
	.w5(32'hba3ad235),
	.w6(32'hbb2f5463),
	.w7(32'hbb8bc435),
	.w8(32'hbbad6317),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53223a),
	.w1(32'hbaa876f7),
	.w2(32'hbb1b6408),
	.w3(32'hba6988fa),
	.w4(32'h39efd3c4),
	.w5(32'hbb257e21),
	.w6(32'hbac9ec6f),
	.w7(32'hbb4097c6),
	.w8(32'h3b2248dd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278f36),
	.w1(32'h3bc3ea8c),
	.w2(32'h3af33f95),
	.w3(32'h3b82142c),
	.w4(32'hba52b754),
	.w5(32'h3af34ede),
	.w6(32'h3acd04a6),
	.w7(32'hbb931ff0),
	.w8(32'hbbb7f442),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87240e),
	.w1(32'hbb9b978d),
	.w2(32'hbb47c51c),
	.w3(32'hbae399f6),
	.w4(32'hbab170f7),
	.w5(32'h3b0c28b1),
	.w6(32'h393b2f74),
	.w7(32'h3b9ee8a0),
	.w8(32'hba9393b9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390a83),
	.w1(32'h3af58528),
	.w2(32'hbb503575),
	.w3(32'hbbd10a0f),
	.w4(32'hbb25e43e),
	.w5(32'h3b76a397),
	.w6(32'hbb33e75e),
	.w7(32'hbc1b7e36),
	.w8(32'hbc5d51cf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaa0ef),
	.w1(32'h3b12296c),
	.w2(32'hbb7b5011),
	.w3(32'h3c85a664),
	.w4(32'hbafc5dab),
	.w5(32'hbac63550),
	.w6(32'h39abae64),
	.w7(32'h3b5e32b3),
	.w8(32'hbc04ad90),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbdafc),
	.w1(32'hbb4d4397),
	.w2(32'h3a7d775f),
	.w3(32'h3b18b4c9),
	.w4(32'hbb48fd7a),
	.w5(32'hbbfa92e9),
	.w6(32'hbafc1ddb),
	.w7(32'hbb5a6586),
	.w8(32'hbaa20890),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33c0b3),
	.w1(32'hba86c725),
	.w2(32'hb9658d11),
	.w3(32'hbb528c57),
	.w4(32'h3ad00c45),
	.w5(32'hbbb40cef),
	.w6(32'h3a976f00),
	.w7(32'h3aafa981),
	.w8(32'h3b09078f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbd0ba),
	.w1(32'h3b15abb2),
	.w2(32'hba90de8b),
	.w3(32'h3b4826ed),
	.w4(32'h3a06d9f7),
	.w5(32'h3abd40b9),
	.w6(32'h3b9415d4),
	.w7(32'hbb38c784),
	.w8(32'h3b27ef45),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a073088),
	.w1(32'h3b8faa4e),
	.w2(32'hba62361a),
	.w3(32'h3bff5496),
	.w4(32'h3b0616cf),
	.w5(32'hb990017d),
	.w6(32'hbb1d4b9a),
	.w7(32'h3ba05443),
	.w8(32'hba425636),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb9018),
	.w1(32'hbb2939a3),
	.w2(32'hbc41d188),
	.w3(32'h3bdab9d5),
	.w4(32'h3af3a991),
	.w5(32'h399e87b9),
	.w6(32'hbb6f98db),
	.w7(32'h3a038dc4),
	.w8(32'h3b058ec0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc90607),
	.w1(32'hbb8a0a43),
	.w2(32'hb8c8d63a),
	.w3(32'hbb6bafbe),
	.w4(32'hbaec0149),
	.w5(32'hbb04fb2f),
	.w6(32'hbb36e7d8),
	.w7(32'hbb3c66bd),
	.w8(32'hbc0c23db),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce0469),
	.w1(32'h3a8d4232),
	.w2(32'hba580280),
	.w3(32'h3a71feaf),
	.w4(32'h3a52a699),
	.w5(32'hba92a81f),
	.w6(32'h3bcbb5d8),
	.w7(32'h3c930e1f),
	.w8(32'hbb25a662),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f199fd),
	.w1(32'h3b464184),
	.w2(32'h39d3e749),
	.w3(32'hb9e702cc),
	.w4(32'h3a84cccb),
	.w5(32'hbb54c7e7),
	.w6(32'hbbc2c3a9),
	.w7(32'h3b351dc2),
	.w8(32'hbab9e971),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc425a69),
	.w1(32'hbc488e9d),
	.w2(32'hba6806c0),
	.w3(32'h3c522c1d),
	.w4(32'hbb92a328),
	.w5(32'hbb149e9e),
	.w6(32'h3931c9ff),
	.w7(32'hba6324e5),
	.w8(32'hbbcd2635),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6bc0),
	.w1(32'hbbbaa00f),
	.w2(32'hb9aa19cb),
	.w3(32'h38701c8e),
	.w4(32'h3ba18347),
	.w5(32'hba01b172),
	.w6(32'hbb5d5ee1),
	.w7(32'h3b725967),
	.w8(32'h3b388e1a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc7342),
	.w1(32'h3a6bd1d8),
	.w2(32'hba5ecdb1),
	.w3(32'hbb045a85),
	.w4(32'hba52beb2),
	.w5(32'hbc07e873),
	.w6(32'hbb62abde),
	.w7(32'hbc5b9ab3),
	.w8(32'hbac90dc3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54b472),
	.w1(32'hb5db549a),
	.w2(32'h3b47695e),
	.w3(32'hbb02ac9e),
	.w4(32'h3b82a095),
	.w5(32'hbb3bdadb),
	.w6(32'h3b54a6ba),
	.w7(32'h383e5647),
	.w8(32'hbaeddab9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b6de3),
	.w1(32'h3b1f9697),
	.w2(32'hb9f81876),
	.w3(32'hba4d9dc0),
	.w4(32'h39fb21d2),
	.w5(32'h3ccf98a2),
	.w6(32'h3b0c6cb1),
	.w7(32'h3b222277),
	.w8(32'hbb529239),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b8092),
	.w1(32'h3c32e1c3),
	.w2(32'h3b3e062c),
	.w3(32'hbc8b8da2),
	.w4(32'hba53f348),
	.w5(32'h3b02eda3),
	.w6(32'hbcb201dd),
	.w7(32'hbc23f18f),
	.w8(32'hbb2e3567),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb260d49),
	.w1(32'hbb248897),
	.w2(32'hbc04898a),
	.w3(32'h3b8ebced),
	.w4(32'h3bc405e2),
	.w5(32'h3a32cb5b),
	.w6(32'h39386c1f),
	.w7(32'hbab29557),
	.w8(32'h3b428c1d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5b829),
	.w1(32'hbb59ec35),
	.w2(32'h3ca02f6f),
	.w3(32'h3ab3680e),
	.w4(32'h3b97ca5f),
	.w5(32'h3a5f852e),
	.w6(32'h3afdd6fe),
	.w7(32'hbae72a38),
	.w8(32'hbb5aa7d9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30f8ed),
	.w1(32'h3b12059d),
	.w2(32'hba5bdf7c),
	.w3(32'h3c9bed3a),
	.w4(32'hbb4fb5fe),
	.w5(32'hbbbae5b8),
	.w6(32'hb9df8d1f),
	.w7(32'hbc5b75ee),
	.w8(32'hba96851a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b3090),
	.w1(32'hbc8081d0),
	.w2(32'hb8cc56dc),
	.w3(32'hbc73cece),
	.w4(32'hbc4021a4),
	.w5(32'h3bae2990),
	.w6(32'hba3aee9e),
	.w7(32'hb84d5041),
	.w8(32'h3a527ab7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba637f84),
	.w1(32'h3b0ee95e),
	.w2(32'hbb5e4454),
	.w3(32'hbb248e6e),
	.w4(32'h3b584b7b),
	.w5(32'hbbe4b937),
	.w6(32'hbb8e5c9a),
	.w7(32'hbb9cde64),
	.w8(32'hbc04f5c8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1262cc),
	.w1(32'hbaffc303),
	.w2(32'h3a91f951),
	.w3(32'h3be106d2),
	.w4(32'hbb8426d5),
	.w5(32'hbb693746),
	.w6(32'h3bc49210),
	.w7(32'h3b66c704),
	.w8(32'hbb0659f5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b82aa),
	.w1(32'hba9b70a0),
	.w2(32'hbc213ba6),
	.w3(32'h3b9883a3),
	.w4(32'h3c397fee),
	.w5(32'h3a24909d),
	.w6(32'hbb0abb41),
	.w7(32'h3b45bcd8),
	.w8(32'hbac16043),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7969ad),
	.w1(32'hbb4e5339),
	.w2(32'h39c9e6b2),
	.w3(32'hbb6fbd9e),
	.w4(32'h36de9934),
	.w5(32'hba1986ad),
	.w6(32'hba15a634),
	.w7(32'hbaba8d16),
	.w8(32'h3a5a2610),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60d9ba),
	.w1(32'hba8cbd00),
	.w2(32'h3b27927f),
	.w3(32'hba10aed5),
	.w4(32'hbb922e74),
	.w5(32'hbb3aaec9),
	.w6(32'hbba34a4a),
	.w7(32'hbc93a3f6),
	.w8(32'hba9da1d0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ea2ee),
	.w1(32'hb97fc032),
	.w2(32'hbb91c33e),
	.w3(32'hbb03706a),
	.w4(32'hbbe4c6ee),
	.w5(32'h3ac05d01),
	.w6(32'hbbdf0b91),
	.w7(32'h3a52d6f9),
	.w8(32'hbb9d62c4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32f8c9),
	.w1(32'h3b8f31b0),
	.w2(32'hba54f7a0),
	.w3(32'hbb97563e),
	.w4(32'hbb0005c6),
	.w5(32'h3b6bb83d),
	.w6(32'hbc1a7d4f),
	.w7(32'hbb83cc3c),
	.w8(32'hb9ac3f6b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9245c3),
	.w1(32'hba21233b),
	.w2(32'hbae928ae),
	.w3(32'hbb4192f5),
	.w4(32'h3b09791a),
	.w5(32'hbaeee101),
	.w6(32'hbc6ef943),
	.w7(32'hba750928),
	.w8(32'h3b1b8abb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23fdff),
	.w1(32'hba93625d),
	.w2(32'h3a174d06),
	.w3(32'h3aa8359e),
	.w4(32'h3a5670de),
	.w5(32'hba105e1b),
	.w6(32'h379c699d),
	.w7(32'h3acb56fa),
	.w8(32'h3a807697),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7af37e),
	.w1(32'hbc850419),
	.w2(32'hbb9c288c),
	.w3(32'hbb6fca15),
	.w4(32'h3bd9b5ca),
	.w5(32'h3b5fefa1),
	.w6(32'h399446ea),
	.w7(32'h3ce14021),
	.w8(32'hbc073ed4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac446a7),
	.w1(32'hba3b2901),
	.w2(32'h3b90bbde),
	.w3(32'hbb0ce661),
	.w4(32'hbc64d02c),
	.w5(32'h3b1c15ed),
	.w6(32'hbab3e098),
	.w7(32'hbb11477a),
	.w8(32'hbb5faa8c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a6cd54),
	.w1(32'h3b6a410d),
	.w2(32'hba562506),
	.w3(32'h3b3747b0),
	.w4(32'hba66de21),
	.w5(32'hba2f8702),
	.w6(32'hbc0c4bfa),
	.w7(32'hbafa63e4),
	.w8(32'h3adc4c84),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b62fd),
	.w1(32'h39c22cbf),
	.w2(32'h3b2e1832),
	.w3(32'hba0bfb30),
	.w4(32'hbb61f286),
	.w5(32'h3a962cd6),
	.w6(32'hbb13bca7),
	.w7(32'h3a4d5e5d),
	.w8(32'h3b47f036),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bd014),
	.w1(32'h3af06a6a),
	.w2(32'h3b28cdd3),
	.w3(32'hba46545d),
	.w4(32'h3a72c630),
	.w5(32'h3b864306),
	.w6(32'hbafe2b03),
	.w7(32'h3a8168d5),
	.w8(32'h3a2ab8a5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3706),
	.w1(32'hbb357fe1),
	.w2(32'hb87f0528),
	.w3(32'hbc083075),
	.w4(32'hbb9dd665),
	.w5(32'h3ab140dc),
	.w6(32'h3a903db3),
	.w7(32'hb9236faa),
	.w8(32'h3b86ac66),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874fc3),
	.w1(32'h3b6259ab),
	.w2(32'hbb576741),
	.w3(32'h3baf8511),
	.w4(32'hb9c6b9f8),
	.w5(32'hbb3a54f6),
	.w6(32'hbb960b87),
	.w7(32'hbb2eacc9),
	.w8(32'hba0ed3ad),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadf798),
	.w1(32'h3b03f595),
	.w2(32'hbc3045ef),
	.w3(32'h3aa5a65d),
	.w4(32'hbb0b674f),
	.w5(32'hbb4ac106),
	.w6(32'hb9305d05),
	.w7(32'h3a9e2ad0),
	.w8(32'hba0921f5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab8097),
	.w1(32'h38e10de6),
	.w2(32'hbc0f5a7a),
	.w3(32'hb9cb536a),
	.w4(32'h3b462272),
	.w5(32'hbaa1ca54),
	.w6(32'hbbd3861b),
	.w7(32'h3adba8f2),
	.w8(32'hbc2c8d92),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8063135),
	.w1(32'hb870f5e6),
	.w2(32'hba809038),
	.w3(32'h3af851fb),
	.w4(32'hbb14440d),
	.w5(32'hbb16d01a),
	.w6(32'hbc05154c),
	.w7(32'h3c8f5a34),
	.w8(32'hbba4fd74),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843313),
	.w1(32'hbb22802f),
	.w2(32'hbbb73b95),
	.w3(32'hbba1c04d),
	.w4(32'h3b45665b),
	.w5(32'hbc6d2dc4),
	.w6(32'hbb962885),
	.w7(32'hbb6b28a9),
	.w8(32'hbb3bf992),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccfdc0),
	.w1(32'hbbf1d619),
	.w2(32'h3a2986bd),
	.w3(32'h3b82f27b),
	.w4(32'hbb334fb8),
	.w5(32'hbb8bcf2c),
	.w6(32'h3b5d0af5),
	.w7(32'h3b93e4c6),
	.w8(32'hbbb7a1c3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc916eeb),
	.w1(32'hba178d10),
	.w2(32'h3b58af68),
	.w3(32'h38ca78af),
	.w4(32'hba8c324d),
	.w5(32'h39b8622f),
	.w6(32'hbc24528f),
	.w7(32'hbadb2ada),
	.w8(32'h3bb21655),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a222c19),
	.w1(32'h3a9adad3),
	.w2(32'h3a37290f),
	.w3(32'h3a3347c1),
	.w4(32'h3aeff804),
	.w5(32'h3b1df31f),
	.w6(32'h3b1b60cd),
	.w7(32'h3b120205),
	.w8(32'h39fba291),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975a8c2),
	.w1(32'hbb6c8e8a),
	.w2(32'hbc08114a),
	.w3(32'hbb6eddaf),
	.w4(32'h3a420d7e),
	.w5(32'h3c09c7b5),
	.w6(32'h3cce3498),
	.w7(32'hbbaebbc7),
	.w8(32'hbb9bf466),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39194d5f),
	.w1(32'hba6b9917),
	.w2(32'h3bab8f10),
	.w3(32'hb9a2cc53),
	.w4(32'hbb83450c),
	.w5(32'h3a695e77),
	.w6(32'h3af6d90c),
	.w7(32'h3b0b973f),
	.w8(32'h3986b123),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af16bda),
	.w1(32'h3c884ba9),
	.w2(32'h3afa4bb8),
	.w3(32'h3943643f),
	.w4(32'hbaa5c69f),
	.w5(32'h39b5e9ce),
	.w6(32'h3acf68ce),
	.w7(32'h3b136d79),
	.w8(32'hba227a33),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f323e3),
	.w1(32'hb9a3d3f9),
	.w2(32'hb99440f8),
	.w3(32'h3c9c7690),
	.w4(32'h3b0ace18),
	.w5(32'h3aab7ea7),
	.w6(32'hbb180cc1),
	.w7(32'h3cc100bc),
	.w8(32'h3984d0bb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc732516),
	.w1(32'hba7a51dd),
	.w2(32'hbb0851ba),
	.w3(32'h39dafe90),
	.w4(32'hbb0dc4f8),
	.w5(32'h3b72480f),
	.w6(32'hbb34b307),
	.w7(32'hbc756cc4),
	.w8(32'hbc40fd4e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade2379),
	.w1(32'h3b0b9214),
	.w2(32'hbbbf0e4b),
	.w3(32'hb9c9c51a),
	.w4(32'hb9ea9315),
	.w5(32'hbb64af8a),
	.w6(32'h3982d4fe),
	.w7(32'hbbf7bd49),
	.w8(32'hb9a90c05),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b569d1f),
	.w1(32'h39feda10),
	.w2(32'hbbcb22cf),
	.w3(32'h3b2371c0),
	.w4(32'h3b7fa005),
	.w5(32'hba1576b7),
	.w6(32'hbc0e6c82),
	.w7(32'h3b61a2f0),
	.w8(32'hbb8468cf),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970e49e),
	.w1(32'hbb10185f),
	.w2(32'hbb48ce4d),
	.w3(32'hbb896c38),
	.w4(32'h3ae7c839),
	.w5(32'hbb89dd86),
	.w6(32'hbb50139c),
	.w7(32'hbaa34d92),
	.w8(32'hbbb53518),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48090b),
	.w1(32'h39da54ce),
	.w2(32'hba11b3c1),
	.w3(32'hb8d5c528),
	.w4(32'h39ffa8bf),
	.w5(32'h38408291),
	.w6(32'hbb908bb5),
	.w7(32'h3b2e38b5),
	.w8(32'h3b0aea6f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b8d11),
	.w1(32'h3a5bfaf6),
	.w2(32'hbbc86e33),
	.w3(32'h3a8750ed),
	.w4(32'h3a86233f),
	.w5(32'hb9aa2616),
	.w6(32'h3ad0311e),
	.w7(32'h3b50181b),
	.w8(32'hbbe5abe1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085c4d),
	.w1(32'h3a974e89),
	.w2(32'hb9b20454),
	.w3(32'hba1cf3b2),
	.w4(32'h3a60328b),
	.w5(32'h3a8c5a1f),
	.w6(32'hbb1a0005),
	.w7(32'hbba93c2c),
	.w8(32'hbb246fb1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee49f7),
	.w1(32'h39d50748),
	.w2(32'h3b09a0ca),
	.w3(32'hba828b07),
	.w4(32'hba008c65),
	.w5(32'h3b7e16f6),
	.w6(32'h3a76d708),
	.w7(32'h38ae6358),
	.w8(32'h3a8f806b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a335766),
	.w1(32'h3ac10740),
	.w2(32'hbb608bff),
	.w3(32'hbab8358e),
	.w4(32'hbba4619c),
	.w5(32'hbaa9e019),
	.w6(32'hb9a0c8a6),
	.w7(32'hbbdd4bba),
	.w8(32'h3aaaf24b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff623e),
	.w1(32'h3c24ae16),
	.w2(32'h3b9cf490),
	.w3(32'hbba7da14),
	.w4(32'h3b937541),
	.w5(32'h3bd10ea0),
	.w6(32'hbc58cefe),
	.w7(32'hbb8b451e),
	.w8(32'hbb506aa4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b638fb7),
	.w1(32'h3b0433b7),
	.w2(32'h3b24289c),
	.w3(32'h3ba60de1),
	.w4(32'h3b844c4c),
	.w5(32'hbbb948fb),
	.w6(32'h3b134d0a),
	.w7(32'hba45f9fa),
	.w8(32'h3a14195e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c958090),
	.w1(32'hbbd3da26),
	.w2(32'hbad33bb4),
	.w3(32'hbb3eba69),
	.w4(32'hbbb189f0),
	.w5(32'hbb35897f),
	.w6(32'hbb1a3388),
	.w7(32'hba62fe03),
	.w8(32'hbbcc104d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2828f4),
	.w1(32'hba7a8325),
	.w2(32'hbc1e5cd1),
	.w3(32'h3b6cb10e),
	.w4(32'hbb46d7f9),
	.w5(32'hbadca675),
	.w6(32'h3b897387),
	.w7(32'h3abcb13c),
	.w8(32'hba02984c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c97de),
	.w1(32'hbb3463fa),
	.w2(32'hba6098bb),
	.w3(32'h3b23b2e8),
	.w4(32'h3c2ddfd6),
	.w5(32'hbc1f3660),
	.w6(32'h39f5ae13),
	.w7(32'h3a7246ff),
	.w8(32'hbc31e738),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552b76),
	.w1(32'h3abd4e32),
	.w2(32'hbb0e0dd2),
	.w3(32'h3c263a49),
	.w4(32'h3a7e8fc2),
	.w5(32'h3be9ceb8),
	.w6(32'hbbad6374),
	.w7(32'hb99959fd),
	.w8(32'hbb5b7e58),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdc4f6),
	.w1(32'hbb914dd6),
	.w2(32'hbc2fd803),
	.w3(32'h3adb168d),
	.w4(32'h3bad8c2b),
	.w5(32'hbafbdcc6),
	.w6(32'hbb32cddf),
	.w7(32'hbbc47d3e),
	.w8(32'hbba9c9ee),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d754),
	.w1(32'h3b9f4010),
	.w2(32'h38cac43c),
	.w3(32'hbab7c7c3),
	.w4(32'h39c2d4cd),
	.w5(32'hb9be4bf3),
	.w6(32'h3a336fad),
	.w7(32'hba42650b),
	.w8(32'h3b0ac25f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c355d),
	.w1(32'hbba974bd),
	.w2(32'hb927aa6d),
	.w3(32'hbb05d8dd),
	.w4(32'hbb85c3ec),
	.w5(32'hbbae2e30),
	.w6(32'hbb59a204),
	.w7(32'hbac70266),
	.w8(32'hbb799b79),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7bc79),
	.w1(32'hbb29e6da),
	.w2(32'hbaf93bfa),
	.w3(32'hbbe0d73a),
	.w4(32'h3c97e4e7),
	.w5(32'h3adcf777),
	.w6(32'hbb96c481),
	.w7(32'h3c3803a7),
	.w8(32'h3af684d2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8294c),
	.w1(32'hba0acd87),
	.w2(32'hbb85abb8),
	.w3(32'h3a5cbb75),
	.w4(32'h3af6ac11),
	.w5(32'hbb008864),
	.w6(32'h3a88849a),
	.w7(32'h3bfbf082),
	.w8(32'hbb1a331e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82c698),
	.w1(32'h3be17926),
	.w2(32'hbaa7c9bf),
	.w3(32'hbb7645bd),
	.w4(32'h3b9fd1d2),
	.w5(32'hba3a823f),
	.w6(32'hbba5c763),
	.w7(32'h38cc9cad),
	.w8(32'hbb10ba53),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1adab5),
	.w1(32'hbb2f0bb5),
	.w2(32'hbb111cd0),
	.w3(32'h3bcb1c85),
	.w4(32'h3b01164e),
	.w5(32'hbbc5c352),
	.w6(32'hbc53debc),
	.w7(32'hbb770566),
	.w8(32'hbc27dbf6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cc377),
	.w1(32'h3b65e226),
	.w2(32'hbb4ef67e),
	.w3(32'h3b42d7f6),
	.w4(32'hba8ab606),
	.w5(32'h3afe7c83),
	.w6(32'h3b1f4e81),
	.w7(32'hba870130),
	.w8(32'h3b362f02),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb845f7b),
	.w1(32'h3b791725),
	.w2(32'h3abd0d70),
	.w3(32'h3bd520ee),
	.w4(32'hb83ece44),
	.w5(32'h3b98f8d2),
	.w6(32'hb4583356),
	.w7(32'hbb6816e1),
	.w8(32'hbaa5d081),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2f7ce),
	.w1(32'hbb9aba00),
	.w2(32'h3d0a15ab),
	.w3(32'hba2d1bd3),
	.w4(32'hbb96eb2a),
	.w5(32'hb9852c3c),
	.w6(32'hbb80ce35),
	.w7(32'h3b3a87a3),
	.w8(32'hbbc81039),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139954),
	.w1(32'hbc04068f),
	.w2(32'h3bf0bdeb),
	.w3(32'hbc1efe9e),
	.w4(32'hbba8300a),
	.w5(32'hba72337f),
	.w6(32'hbb113f65),
	.w7(32'hb9a728ed),
	.w8(32'hbb16d4ea),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f5407),
	.w1(32'hbb1783ae),
	.w2(32'h3bceb4d4),
	.w3(32'hba46ee65),
	.w4(32'hbbbdc8ec),
	.w5(32'h3cd0bd27),
	.w6(32'hbadb723b),
	.w7(32'hbb11d42d),
	.w8(32'h3bfb9103),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33ad3e),
	.w1(32'hb9a299d2),
	.w2(32'h3a535ad8),
	.w3(32'h3a3b98c3),
	.w4(32'hba8a27db),
	.w5(32'hbb0076e3),
	.w6(32'h3af78859),
	.w7(32'h3c56008c),
	.w8(32'h39f68bee),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fdd38),
	.w1(32'hba9bb55e),
	.w2(32'hbc527774),
	.w3(32'h3b8e620e),
	.w4(32'hbaa986d9),
	.w5(32'hba61777c),
	.w6(32'hbc1cb5ec),
	.w7(32'hbadea6d2),
	.w8(32'hbbfeb57e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a209),
	.w1(32'hbc287206),
	.w2(32'h3c9021fd),
	.w3(32'h3b64708a),
	.w4(32'h3b45a08c),
	.w5(32'hbb6a0c53),
	.w6(32'h3bba28a8),
	.w7(32'h3aa8f8b6),
	.w8(32'hbafe5819),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ef11),
	.w1(32'h3ae8638a),
	.w2(32'h3b71fd8b),
	.w3(32'hbabc8b17),
	.w4(32'h3a949d89),
	.w5(32'h3a49dd5c),
	.w6(32'h3afd639a),
	.w7(32'h3ae449ae),
	.w8(32'h3afd2ea5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf649f),
	.w1(32'hbb2932ea),
	.w2(32'hba6e515c),
	.w3(32'h3b6ce542),
	.w4(32'h3a82dc83),
	.w5(32'hbb18ab91),
	.w6(32'hb936f482),
	.w7(32'hbb4400c8),
	.w8(32'h3c027c92),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3afb7b),
	.w1(32'hbad10c94),
	.w2(32'h3ad1274f),
	.w3(32'h3b820aa7),
	.w4(32'h3a663978),
	.w5(32'h388528d4),
	.w6(32'h3b48f1f3),
	.w7(32'hba6d7ea2),
	.w8(32'hba9cb3e7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fa660),
	.w1(32'hbb800e54),
	.w2(32'h3af0ef70),
	.w3(32'h37c53210),
	.w4(32'h39b2d0a8),
	.w5(32'h3b67df62),
	.w6(32'hb8f01f94),
	.w7(32'h3b5ea43e),
	.w8(32'hbaa83324),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac400e0),
	.w1(32'hbc80b4be),
	.w2(32'h3b530d31),
	.w3(32'h3af847bc),
	.w4(32'hbc8506bc),
	.w5(32'h3ac883aa),
	.w6(32'hba1fe64d),
	.w7(32'h3b67ef9a),
	.w8(32'h3bbba058),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28e1ba),
	.w1(32'h3a920f6c),
	.w2(32'hba4b7dc8),
	.w3(32'h3af122ff),
	.w4(32'h3bcf7bc5),
	.w5(32'h3b3d6db3),
	.w6(32'hbadb39c4),
	.w7(32'hbad8437c),
	.w8(32'hb982250e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd34da),
	.w1(32'h3b925edb),
	.w2(32'h3b94835c),
	.w3(32'hbb6e29b2),
	.w4(32'hbb740208),
	.w5(32'h3b8459c0),
	.w6(32'hba2da95c),
	.w7(32'hbbe87596),
	.w8(32'hbb7d1eba),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77160c),
	.w1(32'hbba75885),
	.w2(32'hba88d7f9),
	.w3(32'hbc2e0f8e),
	.w4(32'hbb617cdd),
	.w5(32'hba142d67),
	.w6(32'hbac80f45),
	.w7(32'hb93cc688),
	.w8(32'hbae18918),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aaae8),
	.w1(32'h3b378483),
	.w2(32'hbc19d24d),
	.w3(32'h3b0f4f38),
	.w4(32'h3b45af72),
	.w5(32'hba8bcc55),
	.w6(32'hbba3f244),
	.w7(32'hbb1708b1),
	.w8(32'hbba61512),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc345090),
	.w1(32'hba69bd4a),
	.w2(32'h3b5acd56),
	.w3(32'hbb918cf9),
	.w4(32'hbc40a663),
	.w5(32'hbad1cada),
	.w6(32'hbb45a6f9),
	.w7(32'hbbb5cc54),
	.w8(32'h3a41a432),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4253e0),
	.w1(32'h3c911b2b),
	.w2(32'h37a293fb),
	.w3(32'h3ae05cd5),
	.w4(32'h3a842518),
	.w5(32'h3ad61855),
	.w6(32'hbb55072c),
	.w7(32'hbad69d69),
	.w8(32'h39821187),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb04a5),
	.w1(32'h398bc3e6),
	.w2(32'hbb38512b),
	.w3(32'h3d0f0e7b),
	.w4(32'hba23675a),
	.w5(32'hbb352f84),
	.w6(32'h3b395ba0),
	.w7(32'hbc66e660),
	.w8(32'hbbc3f64f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0222d),
	.w1(32'hbc812577),
	.w2(32'hbabcb543),
	.w3(32'h390ccd5a),
	.w4(32'h3954dc43),
	.w5(32'h3b1b13f0),
	.w6(32'hbb093d27),
	.w7(32'h3bf900ec),
	.w8(32'hbba43abb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47c9ca),
	.w1(32'h3a8a5a22),
	.w2(32'hbb12f922),
	.w3(32'h3b03b985),
	.w4(32'hbb0df9ae),
	.w5(32'h3aff5736),
	.w6(32'h3a0362ae),
	.w7(32'h3be7279d),
	.w8(32'hbbe049f5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf00cc),
	.w1(32'hbb7c7450),
	.w2(32'h3b953b45),
	.w3(32'hbc0c2ea2),
	.w4(32'hbc787167),
	.w5(32'hbb00a077),
	.w6(32'hbbfd318d),
	.w7(32'hba1ea337),
	.w8(32'hbb90f423),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1504b1),
	.w1(32'h3bfbe067),
	.w2(32'hbb961fe2),
	.w3(32'hbb2943c0),
	.w4(32'hbbb06705),
	.w5(32'hb94ba7cb),
	.w6(32'hba5afebf),
	.w7(32'hbaf95204),
	.w8(32'hba41eecd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157f96),
	.w1(32'hbb9a061d),
	.w2(32'hbb288822),
	.w3(32'hba447b31),
	.w4(32'h3bafc88a),
	.w5(32'hb9fa055d),
	.w6(32'hbb961ada),
	.w7(32'hbc510c34),
	.w8(32'h3c016702),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3918b8),
	.w1(32'hbbec19cc),
	.w2(32'hbb863b89),
	.w3(32'hbc100bc6),
	.w4(32'hbbb68727),
	.w5(32'h3b09380e),
	.w6(32'h3a5e4093),
	.w7(32'hbae3ac7c),
	.w8(32'hbb46acd8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bdfd5),
	.w1(32'h3b6c9e9a),
	.w2(32'hbb97deec),
	.w3(32'h3c2275bc),
	.w4(32'hbc686f83),
	.w5(32'h3bf7b460),
	.w6(32'hbb2509af),
	.w7(32'h3aab873f),
	.w8(32'hbb900359),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4a7a),
	.w1(32'hbb66f984),
	.w2(32'hbbfe78a3),
	.w3(32'h3b77b563),
	.w4(32'h3b27c336),
	.w5(32'h3bc2fbc9),
	.w6(32'hbb41a388),
	.w7(32'hbb9bfd28),
	.w8(32'h3bc7e9a4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80faff),
	.w1(32'h3b408ff4),
	.w2(32'hbb4160dd),
	.w3(32'h3a93e071),
	.w4(32'h3a48164e),
	.w5(32'h3baf59ee),
	.w6(32'hbae5c2d8),
	.w7(32'hbc74ba3e),
	.w8(32'h3c86948a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3668b0),
	.w1(32'hba79db9a),
	.w2(32'h3810db65),
	.w3(32'h3c8b0501),
	.w4(32'hbbba3975),
	.w5(32'h3c1dc673),
	.w6(32'h3853334d),
	.w7(32'hbbc48380),
	.w8(32'h3999a9d2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99676a),
	.w1(32'h3b57cb95),
	.w2(32'h3bb86ab0),
	.w3(32'hbc0ad5d7),
	.w4(32'hbab20de5),
	.w5(32'h3b040894),
	.w6(32'hbbbf0637),
	.w7(32'hbc2eb7c2),
	.w8(32'h3ad5eb2c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a819e56),
	.w1(32'hbb3dea3e),
	.w2(32'hbc9e2c95),
	.w3(32'hbbaaa8f0),
	.w4(32'hbb91ba50),
	.w5(32'h3bb165d7),
	.w6(32'h3b7f894a),
	.w7(32'hbc55447f),
	.w8(32'hbbae01e2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb234ff0),
	.w1(32'hb989f06f),
	.w2(32'h3a243889),
	.w3(32'hba25d93b),
	.w4(32'hbb8b745c),
	.w5(32'h3a6cfd4b),
	.w6(32'hbb56f6a1),
	.w7(32'hbbf8b21c),
	.w8(32'hbbc22a88),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedb317),
	.w1(32'hbb883c55),
	.w2(32'hbc742a92),
	.w3(32'hbc457dcc),
	.w4(32'hbbf211eb),
	.w5(32'hbbc029bb),
	.w6(32'h397d2c10),
	.w7(32'h3b8dfa9c),
	.w8(32'hbb0026e5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2fef9),
	.w1(32'h3b911fc5),
	.w2(32'hbb1d663f),
	.w3(32'hbb25e536),
	.w4(32'hbc1c6418),
	.w5(32'hb8c2c4e1),
	.w6(32'hba1dd02b),
	.w7(32'hb8d3bafd),
	.w8(32'h3afc4a03),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd1662),
	.w1(32'h3c158bdd),
	.w2(32'h3c0ae1d5),
	.w3(32'hbaa14b85),
	.w4(32'h3c979363),
	.w5(32'h3c8749f1),
	.w6(32'h3a150a41),
	.w7(32'hba8737a2),
	.w8(32'hbb2b3edc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc454f8d),
	.w1(32'hb98df0d2),
	.w2(32'h3c8b7a5c),
	.w3(32'hbc33d400),
	.w4(32'h3cc0a621),
	.w5(32'h3cd2ebd9),
	.w6(32'hbbc26874),
	.w7(32'h3bd3911f),
	.w8(32'h3c7fe080),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f746f0),
	.w1(32'h3a923c4e),
	.w2(32'hbb8ae291),
	.w3(32'h3cc5caa6),
	.w4(32'h3ba71d55),
	.w5(32'hb8962b3f),
	.w6(32'hbb84fd19),
	.w7(32'hbc3f0fa2),
	.w8(32'hba69e761),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a9f69),
	.w1(32'hb9bf66d0),
	.w2(32'hba4d66d9),
	.w3(32'h3a069183),
	.w4(32'h3ae6e00f),
	.w5(32'hbc1e2f01),
	.w6(32'hbc055472),
	.w7(32'hbb384015),
	.w8(32'h3b016d52),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa37164),
	.w1(32'hba832700),
	.w2(32'h3aa416e7),
	.w3(32'hbc81480c),
	.w4(32'hbb85d06f),
	.w5(32'h3b00e09a),
	.w6(32'h38ace35b),
	.w7(32'hbac57d35),
	.w8(32'hbb091ea1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d8a3),
	.w1(32'hbbdafb5a),
	.w2(32'h3a903e62),
	.w3(32'hbb8a83e6),
	.w4(32'hbbd0f475),
	.w5(32'hbc2760a1),
	.w6(32'h3b5e3a66),
	.w7(32'h3ab2fe94),
	.w8(32'h3c32a701),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a782c),
	.w1(32'hbb3984c0),
	.w2(32'hba894805),
	.w3(32'hbb52d33f),
	.w4(32'hbb2c4fc2),
	.w5(32'h3a9b3d10),
	.w6(32'hbbbd5774),
	.w7(32'h3b0b1f06),
	.w8(32'h3b90d931),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a94d),
	.w1(32'h3b3d13f7),
	.w2(32'h39d9840d),
	.w3(32'h3aee8ccf),
	.w4(32'hbb105095),
	.w5(32'hbac7001c),
	.w6(32'hb9e3b88c),
	.w7(32'h3aaea575),
	.w8(32'h3ad4fc17),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd2efd),
	.w1(32'hbc69e65a),
	.w2(32'hbb66c898),
	.w3(32'h399f18af),
	.w4(32'hbc06329f),
	.w5(32'hbb06605f),
	.w6(32'h3abe500d),
	.w7(32'hbbe4be6d),
	.w8(32'h38e16361),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe859a),
	.w1(32'hbac4ec36),
	.w2(32'hbb776ecc),
	.w3(32'hb93d84a7),
	.w4(32'hbacd6008),
	.w5(32'hbbc9889e),
	.w6(32'hbb0c983d),
	.w7(32'hbab6805f),
	.w8(32'hbbb102b8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919415e),
	.w1(32'hbbe4230f),
	.w2(32'h3c398085),
	.w3(32'hbb4ffee2),
	.w4(32'h3c36be31),
	.w5(32'hbaefd720),
	.w6(32'hbbdfd879),
	.w7(32'hbabfe017),
	.w8(32'h3a9983cd),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb713b3),
	.w1(32'hbb88efe3),
	.w2(32'h3bcdafa7),
	.w3(32'hbbb83918),
	.w4(32'h3b9375b7),
	.w5(32'h3c36cf93),
	.w6(32'hbbdb9c57),
	.w7(32'hbc3c2793),
	.w8(32'hba94d9f7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ef4b),
	.w1(32'h3bc00f5b),
	.w2(32'hbaa88606),
	.w3(32'hbbdba402),
	.w4(32'hbae41a55),
	.w5(32'hb9d99a96),
	.w6(32'hbbab18b7),
	.w7(32'hbb407668),
	.w8(32'hbc867f86),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990a672),
	.w1(32'hbab26fdc),
	.w2(32'hbabd48f7),
	.w3(32'hbac73eac),
	.w4(32'hbbbbf2a6),
	.w5(32'hbd06dca5),
	.w6(32'h3a4decab),
	.w7(32'hbb8fc6c2),
	.w8(32'h3ba501bb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd185797),
	.w1(32'hbc174f72),
	.w2(32'hba8b7cc3),
	.w3(32'hbbacbe41),
	.w4(32'hbba286ce),
	.w5(32'h3ba83781),
	.w6(32'hbc8d9110),
	.w7(32'hbc2319f1),
	.w8(32'hbc2fe8ee),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e720e),
	.w1(32'hbafba141),
	.w2(32'h3aaaf26b),
	.w3(32'h3b21a885),
	.w4(32'h3b68bfee),
	.w5(32'hbc0956d9),
	.w6(32'h39493e23),
	.w7(32'h3b204fb0),
	.w8(32'h3b7a004e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ff31),
	.w1(32'h3a9ac1c4),
	.w2(32'h3b8b1ce3),
	.w3(32'h3b8e8ef9),
	.w4(32'h3cb36a4f),
	.w5(32'hbc304f4c),
	.w6(32'hbb076cfa),
	.w7(32'h3a9de86a),
	.w8(32'h3bd30ee8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b820d2),
	.w1(32'h3c088b2e),
	.w2(32'hbb80402f),
	.w3(32'h3bc1f03a),
	.w4(32'hbabb64cf),
	.w5(32'h3b5b2f43),
	.w6(32'hbb187458),
	.w7(32'hbadb6cec),
	.w8(32'h3bfda158),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0bb4a5),
	.w1(32'h3a5c74fd),
	.w2(32'hbbbad786),
	.w3(32'hbb223a8e),
	.w4(32'h3bfcc190),
	.w5(32'h3aa76a80),
	.w6(32'h3c00a5f3),
	.w7(32'hbaf94d06),
	.w8(32'hbb1bc2fc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4124),
	.w1(32'h3a5a48a0),
	.w2(32'hbb1d5071),
	.w3(32'h3b814eab),
	.w4(32'h3c506cee),
	.w5(32'hbc2cda27),
	.w6(32'h3acc3571),
	.w7(32'hbb092ec3),
	.w8(32'h3bcff760),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29445f),
	.w1(32'hbc60219c),
	.w2(32'hbb1ec559),
	.w3(32'hbbe06f73),
	.w4(32'hb89ea3e2),
	.w5(32'hbc517dd0),
	.w6(32'h3cfe17ed),
	.w7(32'h3d78a373),
	.w8(32'h389afbba),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a20e4),
	.w1(32'hbc4d8e2b),
	.w2(32'hbb269ed7),
	.w3(32'h3c35638f),
	.w4(32'hbc418963),
	.w5(32'hba51e1cf),
	.w6(32'hbbaabc0c),
	.w7(32'hbbd7687d),
	.w8(32'hbb2adf65),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61084b),
	.w1(32'h3c8c8671),
	.w2(32'h3aed0f30),
	.w3(32'hbb434c15),
	.w4(32'h3a572618),
	.w5(32'h3be167d0),
	.w6(32'h3a9b2cb0),
	.w7(32'h3b9a71cf),
	.w8(32'hba34f77b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2f6d30),
	.w1(32'hbc15d823),
	.w2(32'hbcb9fe8a),
	.w3(32'hbb274c77),
	.w4(32'h3b862035),
	.w5(32'hbc587b17),
	.w6(32'h3d376967),
	.w7(32'h3b844c9f),
	.w8(32'hbc909838),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f14e),
	.w1(32'h3bd1ebe8),
	.w2(32'hbb8e0c62),
	.w3(32'hbad835ad),
	.w4(32'hbab46475),
	.w5(32'h3c5ce09e),
	.w6(32'hbbf6b25a),
	.w7(32'hbba331cd),
	.w8(32'h3bd91b9c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9c4ded),
	.w1(32'h391d459d),
	.w2(32'hbba5f7b1),
	.w3(32'h39c7308a),
	.w4(32'h3c727eef),
	.w5(32'hbbfc60d9),
	.w6(32'hbbc59ff8),
	.w7(32'h3bc26375),
	.w8(32'hbbb0d789),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00ddc),
	.w1(32'hbc1a3232),
	.w2(32'hbbdfca2d),
	.w3(32'hbb364dd9),
	.w4(32'hbbbcb1b1),
	.w5(32'h398c8240),
	.w6(32'hbb9ed55b),
	.w7(32'hbb5b0a0f),
	.w8(32'hba461af5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102ce2),
	.w1(32'hbae8c017),
	.w2(32'hb8a10a9e),
	.w3(32'hbb708546),
	.w4(32'h3b7d760f),
	.w5(32'h3bdaf476),
	.w6(32'h3b7b185d),
	.w7(32'hb95f2ddd),
	.w8(32'h3c4bd479),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73406db),
	.w1(32'hba8e415b),
	.w2(32'hbbf1ac7d),
	.w3(32'hbb37ac2b),
	.w4(32'hbbd76d3f),
	.w5(32'hbbc0c6ae),
	.w6(32'h3b840937),
	.w7(32'hbc2e88d0),
	.w8(32'hba6d7cec),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f546),
	.w1(32'hbaaa55b0),
	.w2(32'h3c19cec3),
	.w3(32'h3d425a3e),
	.w4(32'hbb2e9d6e),
	.w5(32'hbba2bef8),
	.w6(32'h3b6111a2),
	.w7(32'hbc0a3359),
	.w8(32'hbcd7053c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a6a09),
	.w1(32'hbb2efa7a),
	.w2(32'hb8239bf8),
	.w3(32'hbb887b1d),
	.w4(32'h3b8a5cf9),
	.w5(32'hbbd05984),
	.w6(32'hbbf9f65f),
	.w7(32'h3ac334d5),
	.w8(32'hbb2e9593),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bf3bb),
	.w1(32'hbc1c68d4),
	.w2(32'hbaffb948),
	.w3(32'hbb2414c9),
	.w4(32'h3c1541c4),
	.w5(32'hbc16f623),
	.w6(32'hbc491d52),
	.w7(32'hbbfa9d27),
	.w8(32'h3c45bead),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1924e5),
	.w1(32'h3b7cdbf0),
	.w2(32'hbb0c8c01),
	.w3(32'h3c33f163),
	.w4(32'hbbd8480c),
	.w5(32'h3a563102),
	.w6(32'hbd044ee5),
	.w7(32'h3cabf7fd),
	.w8(32'hbc37a8ed),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad0586),
	.w1(32'hbaa97214),
	.w2(32'h3bff50eb),
	.w3(32'h3b004a84),
	.w4(32'hbb5211f1),
	.w5(32'h396a09cd),
	.w6(32'h3b0936ea),
	.w7(32'hbad8b33a),
	.w8(32'hb9d66cb1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07a3b),
	.w1(32'hbc47107b),
	.w2(32'h3c03e563),
	.w3(32'h3ac96985),
	.w4(32'h3cbf2855),
	.w5(32'hbb65cee5),
	.w6(32'hbbf39646),
	.w7(32'hba436b64),
	.w8(32'hbb16dfc5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718934),
	.w1(32'h3b40ac49),
	.w2(32'hbb5f1cdc),
	.w3(32'hbb69598c),
	.w4(32'hbaef6ce7),
	.w5(32'hbc0585d9),
	.w6(32'h39c6c5e0),
	.w7(32'hbb75b926),
	.w8(32'h39a80130),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c981625),
	.w1(32'hbc248877),
	.w2(32'hbc172f98),
	.w3(32'hbc00acf5),
	.w4(32'hbc88d4d6),
	.w5(32'h3b629d03),
	.w6(32'hbb982ce9),
	.w7(32'hbb393e30),
	.w8(32'hbb1467b6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c64e0),
	.w1(32'hba2ce05f),
	.w2(32'hbb0c2b3e),
	.w3(32'hbb594d36),
	.w4(32'hbaa6d536),
	.w5(32'hbca280a0),
	.w6(32'h3c265bc7),
	.w7(32'h3bf45ac9),
	.w8(32'hbbdb5480),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28fe0c),
	.w1(32'hb7590a89),
	.w2(32'h3ab76d5d),
	.w3(32'h38870d14),
	.w4(32'hb9550035),
	.w5(32'h399cc329),
	.w6(32'h3a0e98ae),
	.w7(32'hbb3a2487),
	.w8(32'hbb249e49),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab973a4),
	.w1(32'h3d16d019),
	.w2(32'h3b57b119),
	.w3(32'hbc38c2d4),
	.w4(32'hbb93d650),
	.w5(32'hbaa07539),
	.w6(32'hbb23dbab),
	.w7(32'hbc25d224),
	.w8(32'hbba39890),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule