module layer_8_featuremap_207(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13636a),
	.w1(32'h3c892574),
	.w2(32'h397d29f3),
	.w3(32'h3b016e21),
	.w4(32'h3c3103dc),
	.w5(32'h3be2a93b),
	.w6(32'h3c4daef1),
	.w7(32'hbc348e8a),
	.w8(32'h3caba82d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1e95c),
	.w1(32'hbb27c3a5),
	.w2(32'hb9d259f6),
	.w3(32'h3bf205bc),
	.w4(32'hbb404de1),
	.w5(32'hbb2b3dbc),
	.w6(32'hbb869032),
	.w7(32'hbaad5328),
	.w8(32'hba2a9945),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb703a64),
	.w1(32'h3c056d70),
	.w2(32'hbadcaf88),
	.w3(32'hbb9bd40a),
	.w4(32'h3c28c42b),
	.w5(32'h3af4c235),
	.w6(32'h3ba05055),
	.w7(32'hbb2271bf),
	.w8(32'h3c3b8dae),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca347e6),
	.w1(32'h3bc503c9),
	.w2(32'h3c8031be),
	.w3(32'h3cb2128e),
	.w4(32'h3b81df63),
	.w5(32'h3c0e14b5),
	.w6(32'h3b6209b4),
	.w7(32'h3c52bd5b),
	.w8(32'h3c86b862),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd26d5d),
	.w1(32'h3a660dc0),
	.w2(32'h3b219f8a),
	.w3(32'h3c8e9ad9),
	.w4(32'hbb0a592d),
	.w5(32'h3b334f2b),
	.w6(32'hbba4fbe0),
	.w7(32'hba316b21),
	.w8(32'hbba6af3c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a0808),
	.w1(32'h3a2b762d),
	.w2(32'hbc6ef8fb),
	.w3(32'hbb6ca401),
	.w4(32'hbb53213e),
	.w5(32'hbc811ea7),
	.w6(32'h3c0dbcf0),
	.w7(32'hbc77fc09),
	.w8(32'h3b97f4c9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b734191),
	.w1(32'hba30dd65),
	.w2(32'h3a206038),
	.w3(32'hbc0521ea),
	.w4(32'h3a88b878),
	.w5(32'h3a72f24b),
	.w6(32'h3a8e8240),
	.w7(32'h3ad62590),
	.w8(32'hbacaf2ed),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc66c),
	.w1(32'hbc389e0a),
	.w2(32'h3c91c805),
	.w3(32'hba0befed),
	.w4(32'hbc43ac3d),
	.w5(32'h3bcba66d),
	.w6(32'hbc8513f5),
	.w7(32'h3c39a720),
	.w8(32'h3c38f04c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c805025),
	.w1(32'h3aa7e10c),
	.w2(32'hb92bdc6b),
	.w3(32'h3b2017be),
	.w4(32'h39088746),
	.w5(32'h3b175f5a),
	.w6(32'hbb6e9363),
	.w7(32'hba13a904),
	.w8(32'hbc30a278),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cf170),
	.w1(32'h3b6f1b7c),
	.w2(32'hbc8ba9f2),
	.w3(32'hbc340ae9),
	.w4(32'h3c0db25a),
	.w5(32'hbc064eff),
	.w6(32'hb961bcfb),
	.w7(32'hbc010da9),
	.w8(32'h3c96f09b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ce94),
	.w1(32'h3b79e1d4),
	.w2(32'hbba731d4),
	.w3(32'h3a065489),
	.w4(32'h3c4b4721),
	.w5(32'hbb2443a7),
	.w6(32'hb95b6489),
	.w7(32'hbb2a9863),
	.w8(32'h3a363cc5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc981e2),
	.w1(32'h3b97e009),
	.w2(32'h3b7f16d0),
	.w3(32'hbb8bc42f),
	.w4(32'h3a87c7e4),
	.w5(32'h3aa5d3a3),
	.w6(32'h386216ca),
	.w7(32'h3aa1eb7b),
	.w8(32'h3b9cd402),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9bce),
	.w1(32'hbad7605b),
	.w2(32'hbb5edc73),
	.w3(32'hbb755498),
	.w4(32'h3a339932),
	.w5(32'h3970d43d),
	.w6(32'h3bd76344),
	.w7(32'h3b53386e),
	.w8(32'h3bb89090),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb960cb),
	.w1(32'h3b9c5c40),
	.w2(32'h3c2d4f04),
	.w3(32'hba9e589c),
	.w4(32'h3beba116),
	.w5(32'h3bd2de6a),
	.w6(32'h3b9d9a0c),
	.w7(32'h3af6fade),
	.w8(32'h3c5e816e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6d5e6),
	.w1(32'hbb265f46),
	.w2(32'hbbf42b7a),
	.w3(32'h3ca66109),
	.w4(32'hbac6aee1),
	.w5(32'hbbaef013),
	.w6(32'hba96e3c1),
	.w7(32'hbb514c9e),
	.w8(32'h3a80773e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995fda2),
	.w1(32'h3cb9f0cb),
	.w2(32'hbbaed7b6),
	.w3(32'h3af0cbe5),
	.w4(32'h3c871967),
	.w5(32'h3afbe6fc),
	.w6(32'h3c9db251),
	.w7(32'hbb9b318c),
	.w8(32'hbb9b93d7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb267b58),
	.w1(32'h3a693069),
	.w2(32'hbc07e6ad),
	.w3(32'hbc3d8de2),
	.w4(32'h3becb7c0),
	.w5(32'hbc4de3fa),
	.w6(32'h3c0d62ba),
	.w7(32'hbb91b330),
	.w8(32'h3bc0cd86),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c499545),
	.w1(32'h3c8d054f),
	.w2(32'h3cc29c98),
	.w3(32'h3a81edb9),
	.w4(32'h3c1458eb),
	.w5(32'h3c919d00),
	.w6(32'h3c709ad7),
	.w7(32'h3c8eec20),
	.w8(32'h3c48933e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08bce9),
	.w1(32'h3d16e29e),
	.w2(32'hbc7c1423),
	.w3(32'h3cb8d09b),
	.w4(32'h3d0937fd),
	.w5(32'hba0c6e92),
	.w6(32'hbae0ce06),
	.w7(32'hbc971de0),
	.w8(32'h3ccedbbd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3ac2b),
	.w1(32'h3b67c5db),
	.w2(32'hb99fcc96),
	.w3(32'h3c0db461),
	.w4(32'h3aea7382),
	.w5(32'hbabae48e),
	.w6(32'hbb823ae0),
	.w7(32'hbb8ecb08),
	.w8(32'hbaf8f416),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac5f80),
	.w1(32'hbc02da98),
	.w2(32'hbc550813),
	.w3(32'hbb94b1f5),
	.w4(32'h390d239e),
	.w5(32'hbb90fb3f),
	.w6(32'h39ae20fb),
	.w7(32'h3b0652c2),
	.w8(32'h3b23378e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc379a6e),
	.w1(32'hbc2db11b),
	.w2(32'hbcaa3ce7),
	.w3(32'hbb85a4d7),
	.w4(32'hbb0e1950),
	.w5(32'hbc3e0e66),
	.w6(32'hbb4d86d5),
	.w7(32'hbb777929),
	.w8(32'hbbbf97de),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc21437),
	.w1(32'h3ba65f5a),
	.w2(32'hbbf0e4c3),
	.w3(32'hbc60efc4),
	.w4(32'h3c2065db),
	.w5(32'hbbe000ad),
	.w6(32'hba3714b8),
	.w7(32'hbc593748),
	.w8(32'h3c2b5f75),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bc405),
	.w1(32'h3b99c5ff),
	.w2(32'hbb9861da),
	.w3(32'h3adaf0ee),
	.w4(32'h3c8438f8),
	.w5(32'hbae0e95b),
	.w6(32'h3b45927a),
	.w7(32'h3c4be770),
	.w8(32'h3afb3e8e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb39397),
	.w1(32'hbc1d0067),
	.w2(32'hbc060e43),
	.w3(32'h3b6192c2),
	.w4(32'h3ad85e1b),
	.w5(32'h3b5e7473),
	.w6(32'hbbcba3a5),
	.w7(32'h3a7f29e0),
	.w8(32'h3be4179f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbfd21),
	.w1(32'hbb8bc142),
	.w2(32'hbb881d7c),
	.w3(32'h3bd289ea),
	.w4(32'h3bee4d60),
	.w5(32'h3c749636),
	.w6(32'hbc652e04),
	.w7(32'hbb749244),
	.w8(32'h3a857c56),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12d56),
	.w1(32'hbc331a51),
	.w2(32'hbc92d411),
	.w3(32'hbaeccb63),
	.w4(32'hbba0e54b),
	.w5(32'hbcb09767),
	.w6(32'hbb7ec42a),
	.w7(32'hbbe456f9),
	.w8(32'hbb176206),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ecc43),
	.w1(32'h3c1ff25d),
	.w2(32'h3bcbbf6e),
	.w3(32'hbc72b33f),
	.w4(32'h3caea56e),
	.w5(32'h3c2ee45c),
	.w6(32'h3c9f0003),
	.w7(32'hbd20e619),
	.w8(32'hbc6ecccc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78730c),
	.w1(32'h3c52a8ca),
	.w2(32'h3bc16daa),
	.w3(32'hbbc13929),
	.w4(32'h3bf21efd),
	.w5(32'h3b5a1f9e),
	.w6(32'h3c2f6f13),
	.w7(32'h3aa84011),
	.w8(32'hbbc7e34d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc699108),
	.w1(32'h3869e4b1),
	.w2(32'h3b1d54fb),
	.w3(32'hbc641c64),
	.w4(32'hbbdf2911),
	.w5(32'h3769f6c5),
	.w6(32'hbae75d14),
	.w7(32'hba4edce8),
	.w8(32'hbbb2f398),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5a95),
	.w1(32'hbb873305),
	.w2(32'h39994313),
	.w3(32'hbc097299),
	.w4(32'hbbe0b70f),
	.w5(32'hbbd49e69),
	.w6(32'h38c90a00),
	.w7(32'hba0d2b08),
	.w8(32'h3c0e2eea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c094642),
	.w1(32'hbb2c6938),
	.w2(32'hbc72711a),
	.w3(32'h3ba68aa4),
	.w4(32'h3a8caec9),
	.w5(32'hbc001b32),
	.w6(32'hbbafc9dc),
	.w7(32'hbc5a3691),
	.w8(32'h3bfd1dd8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ed63b),
	.w1(32'hbc51dc63),
	.w2(32'hbc888069),
	.w3(32'h3bad2e12),
	.w4(32'hbc0f2554),
	.w5(32'hbc84adf3),
	.w6(32'hbc1ce922),
	.w7(32'hbc75e7a9),
	.w8(32'hbc1cd07d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa600),
	.w1(32'h3b79fc3a),
	.w2(32'h3b1be877),
	.w3(32'hbc378b7c),
	.w4(32'hbb328d9d),
	.w5(32'h3c16a326),
	.w6(32'h3c51e469),
	.w7(32'h3bb6e55e),
	.w8(32'h3c6e8ee2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b833a),
	.w1(32'hbb86d2e8),
	.w2(32'hbb9dab5b),
	.w3(32'h3c544d5a),
	.w4(32'hbc27876e),
	.w5(32'hbc24257e),
	.w6(32'hbba725c2),
	.w7(32'hbbce3b06),
	.w8(32'hbbbcaa99),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d11d),
	.w1(32'h3c574d43),
	.w2(32'h3b3a5912),
	.w3(32'h3970834d),
	.w4(32'h3be4f703),
	.w5(32'hbac8f27f),
	.w6(32'h3b85888b),
	.w7(32'hbc15ac82),
	.w8(32'h3b0532bf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11df3e),
	.w1(32'h3b569dbe),
	.w2(32'h3b44ed76),
	.w3(32'hbb1de392),
	.w4(32'h3b4464d7),
	.w5(32'h3ac3e48d),
	.w6(32'h3b968f19),
	.w7(32'h3b5955a2),
	.w8(32'h3a4b46e4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239ebe),
	.w1(32'hba82127f),
	.w2(32'h3b339843),
	.w3(32'hbb529f2b),
	.w4(32'hbaaf42b0),
	.w5(32'h3b072d5c),
	.w6(32'hbb72a65c),
	.w7(32'h3ab5c164),
	.w8(32'hbb1feb18),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c7e6),
	.w1(32'h3afd4294),
	.w2(32'h3bfd0674),
	.w3(32'h3aa020e1),
	.w4(32'h3b8e3e19),
	.w5(32'h3bcaf326),
	.w6(32'hbb7994b5),
	.w7(32'h3c078f10),
	.w8(32'h3b6cc246),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc759ed),
	.w1(32'h3c683f8b),
	.w2(32'h3b6a3a00),
	.w3(32'h3ab9e54a),
	.w4(32'h3c564849),
	.w5(32'hbabfdc42),
	.w6(32'h3c0d323c),
	.w7(32'h3c1e940e),
	.w8(32'h3c356e79),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5f92),
	.w1(32'h3b4b2c37),
	.w2(32'hb9b8efc6),
	.w3(32'h3c428090),
	.w4(32'h3b65d230),
	.w5(32'h3a95218e),
	.w6(32'hbc1b047f),
	.w7(32'hbc680620),
	.w8(32'h3bc53322),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80066a),
	.w1(32'h3bdce341),
	.w2(32'hbc2439e3),
	.w3(32'hbb3391f7),
	.w4(32'h3ba05aa8),
	.w5(32'hbc4cfb3b),
	.w6(32'h3b70e51a),
	.w7(32'hbc44103c),
	.w8(32'h3bb0eb76),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9614b0),
	.w1(32'hbc222358),
	.w2(32'h3af90794),
	.w3(32'hbaacc54b),
	.w4(32'hbbeca62a),
	.w5(32'hba982505),
	.w6(32'hbb601533),
	.w7(32'h39fb6fd6),
	.w8(32'hbb03b36e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b17d2),
	.w1(32'hbace3488),
	.w2(32'h3cfc242e),
	.w3(32'h3a983145),
	.w4(32'hbc2f6976),
	.w5(32'h3c979d86),
	.w6(32'h3a7a12dc),
	.w7(32'h3c1ca28c),
	.w8(32'h3c5c735d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca36cb),
	.w1(32'h3c6a5d37),
	.w2(32'hbcece4c4),
	.w3(32'h3c926b16),
	.w4(32'h3c76f14c),
	.w5(32'hbcb171f8),
	.w6(32'h3bd513fb),
	.w7(32'hbc669bae),
	.w8(32'h3c8549e5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b267e43),
	.w1(32'hbace5539),
	.w2(32'hbc084b82),
	.w3(32'h3b02b76a),
	.w4(32'hb8279ed0),
	.w5(32'hbb8163d0),
	.w6(32'hba23bcaa),
	.w7(32'hbb896670),
	.w8(32'hbb07bbba),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba78e8),
	.w1(32'h3b99b31b),
	.w2(32'hbb992938),
	.w3(32'hbb96cc8d),
	.w4(32'h3bc09aea),
	.w5(32'hbb317a31),
	.w6(32'h3b7122f9),
	.w7(32'h3a24e4bc),
	.w8(32'h3b97c458),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba966efb),
	.w1(32'h3c885451),
	.w2(32'hbae5958c),
	.w3(32'hb96bdd4a),
	.w4(32'h3c45909e),
	.w5(32'h3ac50f2b),
	.w6(32'h3b259707),
	.w7(32'hbb28420d),
	.w8(32'h3c588026),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155969),
	.w1(32'h3b818927),
	.w2(32'hbc3409b4),
	.w3(32'h3b83b729),
	.w4(32'hb9b2ce73),
	.w5(32'hbc563a77),
	.w6(32'h3b16e05e),
	.w7(32'hbb280dc0),
	.w8(32'h3b09c89f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c069c85),
	.w1(32'h3ca1be07),
	.w2(32'hbb4583d8),
	.w3(32'h3ab9ddf1),
	.w4(32'h3c795636),
	.w5(32'h3bf4b691),
	.w6(32'h3bc80115),
	.w7(32'hbc5b72fa),
	.w8(32'h3c342ba9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47d88d),
	.w1(32'hbc08fc6e),
	.w2(32'hbc13faf5),
	.w3(32'h3a1fc764),
	.w4(32'hbbf0b94d),
	.w5(32'hbc1141d3),
	.w6(32'hbc063165),
	.w7(32'hbc70fae2),
	.w8(32'hbb92e7a2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba842d37),
	.w1(32'h3c75c280),
	.w2(32'h3bd59f99),
	.w3(32'h3bab7909),
	.w4(32'h3ca4f17b),
	.w5(32'h3bdaa56d),
	.w6(32'h39ae8d96),
	.w7(32'hbad0bc6b),
	.w8(32'h3b9abce3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4bbf),
	.w1(32'h3b158864),
	.w2(32'h3b39808d),
	.w3(32'hbaf17d67),
	.w4(32'h3bb5c527),
	.w5(32'h3b4416fa),
	.w6(32'hbb2724ba),
	.w7(32'h3b3d3854),
	.w8(32'h3bda278a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba49dab),
	.w1(32'hbbb19072),
	.w2(32'h3cab4eea),
	.w3(32'h3bb4eb7a),
	.w4(32'hbbfb9785),
	.w5(32'h3c8cb42e),
	.w6(32'hbbaa0cfc),
	.w7(32'h3c444325),
	.w8(32'h3c174aa7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70c5da),
	.w1(32'hba3a24ea),
	.w2(32'h3c511958),
	.w3(32'h3c1a91e4),
	.w4(32'hbb870b1f),
	.w5(32'h3c3b0dce),
	.w6(32'hbc33486d),
	.w7(32'h3b9e708b),
	.w8(32'h3b2c10b5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b243ed7),
	.w1(32'h3b0a0667),
	.w2(32'h3cbfa207),
	.w3(32'hb860333e),
	.w4(32'hbbd0fa83),
	.w5(32'h3cbb499a),
	.w6(32'h372e4d68),
	.w7(32'h3a32f338),
	.w8(32'h3b5d6ac2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccea59),
	.w1(32'hbb8a7ff1),
	.w2(32'h3c4a2d29),
	.w3(32'h3c311aa9),
	.w4(32'hbbe31f4e),
	.w5(32'h39a1a0d6),
	.w6(32'h3a2e4912),
	.w7(32'hb9e7bda6),
	.w8(32'hbc6ef6e4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e7290),
	.w1(32'hbb995219),
	.w2(32'hbb9ca50b),
	.w3(32'hbbde4d6b),
	.w4(32'hba848fea),
	.w5(32'hbb4b7e2f),
	.w6(32'hb9516db3),
	.w7(32'h3a62acb2),
	.w8(32'h3a9d26b1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bf597),
	.w1(32'h3ab859bb),
	.w2(32'hbb86acbe),
	.w3(32'h38a2de20),
	.w4(32'h3ae9649c),
	.w5(32'hbb9f0667),
	.w6(32'h3b23af25),
	.w7(32'hbafbdb7e),
	.w8(32'hb915609b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05bd2),
	.w1(32'h3c1429fa),
	.w2(32'h3bc0b2e5),
	.w3(32'hbb4ac8d0),
	.w4(32'h3c0bc809),
	.w5(32'hbac14c0a),
	.w6(32'h3b8718db),
	.w7(32'h3baf7e84),
	.w8(32'h39641912),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d945c),
	.w1(32'hbc2ed152),
	.w2(32'hbb95816f),
	.w3(32'hbab0ef1f),
	.w4(32'h3b5989d8),
	.w5(32'hbc079c44),
	.w6(32'hbbb3a52d),
	.w7(32'hbb536b2f),
	.w8(32'h3adce630),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39875272),
	.w1(32'hba3adb63),
	.w2(32'h3a8921f2),
	.w3(32'h3ba4a6e8),
	.w4(32'h39c8398b),
	.w5(32'hba25f2dd),
	.w6(32'h39334270),
	.w7(32'h3bbb8ca4),
	.w8(32'h3b8967ba),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13819b),
	.w1(32'h3c2df961),
	.w2(32'h3cd750e4),
	.w3(32'h3bbce0b4),
	.w4(32'h3c2489aa),
	.w5(32'h3cf4399b),
	.w6(32'hbb608099),
	.w7(32'h3c36464d),
	.w8(32'h3c4a6bf3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69c9f4),
	.w1(32'hbae0366a),
	.w2(32'h38d95e04),
	.w3(32'h3bc07a34),
	.w4(32'hba824c66),
	.w5(32'hbb1eba72),
	.w6(32'hb9eb17e1),
	.w7(32'h3b8e04c9),
	.w8(32'h3b91baf8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8290c4),
	.w1(32'hbb9fa7a6),
	.w2(32'hbbf11d5d),
	.w3(32'hbb926a1b),
	.w4(32'hbb7e1b4e),
	.w5(32'hbbfd3270),
	.w6(32'hbb989719),
	.w7(32'hbbb22af6),
	.w8(32'h3a983edf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b056),
	.w1(32'h3c275564),
	.w2(32'h3b11aadf),
	.w3(32'hbbd0ac70),
	.w4(32'h3c8aae7a),
	.w5(32'hb9992798),
	.w6(32'h3b8c672c),
	.w7(32'h3b80ea4a),
	.w8(32'h3c8584bf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdf5ef),
	.w1(32'hbb880da0),
	.w2(32'hb937c844),
	.w3(32'h3be3d69c),
	.w4(32'h3bc0fa08),
	.w5(32'hbb603761),
	.w6(32'h3b655d4f),
	.w7(32'h3c1e1580),
	.w8(32'h3cd224c9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf164a1),
	.w1(32'h3b1fa453),
	.w2(32'hbbb7207d),
	.w3(32'h3c5742ab),
	.w4(32'h3bae5b11),
	.w5(32'h3b5fcd84),
	.w6(32'h3b11cc6b),
	.w7(32'hbb2a6f95),
	.w8(32'hb9c42bae),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b172ea1),
	.w1(32'hbb05bd3b),
	.w2(32'h3ba7f460),
	.w3(32'h39c8b312),
	.w4(32'hbafc2c03),
	.w5(32'hb99560bf),
	.w6(32'hba70752c),
	.w7(32'h3b845776),
	.w8(32'h3bb20eb7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79405d),
	.w1(32'h3ba8e1da),
	.w2(32'hbb9f057b),
	.w3(32'h3bcdd38b),
	.w4(32'h3bce427f),
	.w5(32'hbb53d455),
	.w6(32'hbb8453f9),
	.w7(32'hbc2fbdff),
	.w8(32'hba89f627),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f7630),
	.w1(32'h3bd64ec3),
	.w2(32'hbc0c2c18),
	.w3(32'hbb0ae937),
	.w4(32'h3be611a4),
	.w5(32'hbb97f641),
	.w6(32'hb9270d8b),
	.w7(32'hbc0dff2a),
	.w8(32'hbbc64c9f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2506c9),
	.w1(32'h3c29f8b1),
	.w2(32'hbbfe7f86),
	.w3(32'hbb831072),
	.w4(32'h3c18e445),
	.w5(32'hbb2979d9),
	.w6(32'hba916cef),
	.w7(32'hbb62beee),
	.w8(32'h3b6354c0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7cad8),
	.w1(32'h3c0c6054),
	.w2(32'hbc6a6739),
	.w3(32'h3c03878d),
	.w4(32'h3bceb8ed),
	.w5(32'hbb925707),
	.w6(32'h3bae7fd0),
	.w7(32'h3a489ea9),
	.w8(32'h3c336e5d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba10eaf),
	.w1(32'hbb322495),
	.w2(32'hbb300d2c),
	.w3(32'h3c10980b),
	.w4(32'hbabdd9c7),
	.w5(32'h3aae0030),
	.w6(32'hbbb4186c),
	.w7(32'hbb3f26c3),
	.w8(32'h3a28be66),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169dcc),
	.w1(32'h3b6cb192),
	.w2(32'hbc8805cf),
	.w3(32'h3b8314b7),
	.w4(32'h3ac8ceed),
	.w5(32'hbc349090),
	.w6(32'h3c2ac121),
	.w7(32'hbc1a119c),
	.w8(32'h39d7aedb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64f5cf),
	.w1(32'h3c37fd76),
	.w2(32'h3c40c917),
	.w3(32'hbaa2c38e),
	.w4(32'h3be9d50e),
	.w5(32'h3c228a1f),
	.w6(32'h3a42069f),
	.w7(32'h395b874b),
	.w8(32'h3c347d0d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5f7d5),
	.w1(32'hbc25afdf),
	.w2(32'hbb59f4b8),
	.w3(32'h3ca2ce3a),
	.w4(32'hbc29014f),
	.w5(32'hbb85bea1),
	.w6(32'hbbc956eb),
	.w7(32'hbbdacbc8),
	.w8(32'hbbea0cc3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe70f56),
	.w1(32'h3b37f6a5),
	.w2(32'h3c79c070),
	.w3(32'h3a1d21d7),
	.w4(32'h3b5dc317),
	.w5(32'h3c6469f1),
	.w6(32'hba804c8b),
	.w7(32'h3c12b7b3),
	.w8(32'h3b52e7dc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1d9a8),
	.w1(32'h3c6f64a0),
	.w2(32'hbbdf94bc),
	.w3(32'h3a6f96d7),
	.w4(32'h3caa365a),
	.w5(32'h3b1dd7da),
	.w6(32'h3be747bd),
	.w7(32'hbbc97624),
	.w8(32'h3b810292),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b55b),
	.w1(32'h3bde1030),
	.w2(32'h3c47316f),
	.w3(32'h3bd089ad),
	.w4(32'h3b582ae1),
	.w5(32'h3c814de2),
	.w6(32'h3c09bd80),
	.w7(32'hbb3c2733),
	.w8(32'hbb696fbf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0070f6),
	.w1(32'hbc2cbc4c),
	.w2(32'hbca63212),
	.w3(32'hbaf72722),
	.w4(32'hbbd2d6ef),
	.w5(32'hbc7f7cfa),
	.w6(32'hbb23a3ed),
	.w7(32'hbc33d7c2),
	.w8(32'hbb431196),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e1e7),
	.w1(32'h3bb4c37c),
	.w2(32'h3b41570d),
	.w3(32'hbbd29c5a),
	.w4(32'hb9ac2259),
	.w5(32'h3b147344),
	.w6(32'h3ac98102),
	.w7(32'h3ab4fc5f),
	.w8(32'h3c1b3e04),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdea03c),
	.w1(32'h3c2a8862),
	.w2(32'h3b56f467),
	.w3(32'h3bd252a5),
	.w4(32'h3b717887),
	.w5(32'h3c137c1f),
	.w6(32'hbc0d010b),
	.w7(32'hbc06073d),
	.w8(32'h3b94ebb2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3f32d),
	.w1(32'h3b569521),
	.w2(32'h3c89fca0),
	.w3(32'h3ce67293),
	.w4(32'h3b8fd7f7),
	.w5(32'h3c44307a),
	.w6(32'hbb26ffe4),
	.w7(32'h3ba17000),
	.w8(32'h3b995282),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e003d),
	.w1(32'h3b7a03e2),
	.w2(32'hbb8f2e95),
	.w3(32'hba9ac803),
	.w4(32'h3c416b06),
	.w5(32'h3bd738d5),
	.w6(32'hbc322a4c),
	.w7(32'hbc5b06bd),
	.w8(32'h3c16b458),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e97af),
	.w1(32'h3c1a0dd7),
	.w2(32'h3b828f0e),
	.w3(32'hba88b0f2),
	.w4(32'h3c1f3fb0),
	.w5(32'h3aee6b00),
	.w6(32'h3b2078d2),
	.w7(32'h3bed62e8),
	.w8(32'h3be2b7aa),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2491d9),
	.w1(32'h3b8b15e8),
	.w2(32'hb9ce6671),
	.w3(32'hbbc47a96),
	.w4(32'h3ba81e3d),
	.w5(32'hba0146e5),
	.w6(32'h3aea6052),
	.w7(32'h3a9be921),
	.w8(32'h3ba0cc45),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab42515),
	.w1(32'hbba28aab),
	.w2(32'hbbb49caf),
	.w3(32'h3a089dff),
	.w4(32'h3bffa9ae),
	.w5(32'h3a325d26),
	.w6(32'hbb4d04ca),
	.w7(32'hbc275a08),
	.w8(32'hbbcff74c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b84c9),
	.w1(32'h3af17426),
	.w2(32'h3a917a11),
	.w3(32'hbb14bc9b),
	.w4(32'hbb83d78b),
	.w5(32'hbb2d8420),
	.w6(32'h3b811d28),
	.w7(32'h3b842a22),
	.w8(32'h3bbe55e6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19efec),
	.w1(32'h3c06a6fa),
	.w2(32'h3b86638d),
	.w3(32'hb63c31aa),
	.w4(32'h3bfc843c),
	.w5(32'h3bae5e51),
	.w6(32'h3b36aaeb),
	.w7(32'hbabf0c05),
	.w8(32'h3cc1ce76),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0c637),
	.w1(32'h3a411ab3),
	.w2(32'hbb2d938a),
	.w3(32'h3ca625d4),
	.w4(32'h3b8c3176),
	.w5(32'hbbec6126),
	.w6(32'h3b76352f),
	.w7(32'h3add5352),
	.w8(32'h3bc5365a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73941e),
	.w1(32'h3bd286ae),
	.w2(32'h3bce5956),
	.w3(32'hbb4b98a5),
	.w4(32'h3bf24004),
	.w5(32'h3baec8d4),
	.w6(32'h3be518c0),
	.w7(32'h3bc06c4e),
	.w8(32'h3c4370a3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66b00c),
	.w1(32'hba2807ce),
	.w2(32'hbb72898d),
	.w3(32'h3c1d0040),
	.w4(32'h39adf070),
	.w5(32'hbae6d29c),
	.w6(32'h3b000792),
	.w7(32'h39b06abe),
	.w8(32'hbb74e111),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3710),
	.w1(32'hb91efb5f),
	.w2(32'hba14df1f),
	.w3(32'hbbfa0e55),
	.w4(32'h3b29a7a5),
	.w5(32'h3a2d8f3c),
	.w6(32'hbb5eb087),
	.w7(32'hbb0d941c),
	.w8(32'h3b869df9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6afc10),
	.w1(32'hbc6627e1),
	.w2(32'h3c917099),
	.w3(32'hbbb40035),
	.w4(32'hbc55ed38),
	.w5(32'h3c4897a0),
	.w6(32'hbc3f9238),
	.w7(32'h3bf09d72),
	.w8(32'h3c403105),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14f123),
	.w1(32'h3b6bcae3),
	.w2(32'h3b1a3abd),
	.w3(32'h3c1339e8),
	.w4(32'h3a619478),
	.w5(32'h3b19a12a),
	.w6(32'h39a43283),
	.w7(32'hba8c4c71),
	.w8(32'hb99c173b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd1121),
	.w1(32'h3b9a267a),
	.w2(32'h3bbd9345),
	.w3(32'hba7b8106),
	.w4(32'h3b0e6cca),
	.w5(32'h3c8383b6),
	.w6(32'hbb72be71),
	.w7(32'h3a7f5e32),
	.w8(32'h3ac230c2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c058d7c),
	.w1(32'hb88075c9),
	.w2(32'h3c96c6d8),
	.w3(32'h3c02c7cd),
	.w4(32'h3b492c20),
	.w5(32'h3ae64a18),
	.w6(32'h3b493772),
	.w7(32'h3b675619),
	.w8(32'h3c6ce7b5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd145c),
	.w1(32'h3b9c4aff),
	.w2(32'h3cb26b22),
	.w3(32'h3ba74d4b),
	.w4(32'h3bc93f9d),
	.w5(32'h3c4105aa),
	.w6(32'hbb900794),
	.w7(32'h3be7e3d6),
	.w8(32'h3a872f29),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0b4d9),
	.w1(32'hbc3e9200),
	.w2(32'h3ab7c1e1),
	.w3(32'hbb8671cc),
	.w4(32'hbbacc820),
	.w5(32'h3b62db5c),
	.w6(32'hbc4ae4ce),
	.w7(32'h3b3ba7a9),
	.w8(32'h3b2ef3b2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a908b6d),
	.w1(32'h3a450188),
	.w2(32'h3920be1e),
	.w3(32'hba7ae190),
	.w4(32'h3b411089),
	.w5(32'hbb395280),
	.w6(32'h3bf7d817),
	.w7(32'h3c49c636),
	.w8(32'h3b9303dd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd50f3e),
	.w1(32'hbcaae245),
	.w2(32'hbc908627),
	.w3(32'h3bc5a8c3),
	.w4(32'hbc8dc94e),
	.w5(32'hbc96ccb8),
	.w6(32'hbcaeea3e),
	.w7(32'hbc5a0fa5),
	.w8(32'hbb0072dc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc752e1f),
	.w1(32'h3c418d45),
	.w2(32'h3b00a558),
	.w3(32'hbc319f84),
	.w4(32'h3b627f30),
	.w5(32'h3b201016),
	.w6(32'h3c261918),
	.w7(32'h3a7a35ac),
	.w8(32'h3c60f9ce),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b84c7),
	.w1(32'hbb7cccbe),
	.w2(32'hbb6168e5),
	.w3(32'h3ca409b8),
	.w4(32'hbb2f91c9),
	.w5(32'h3b65675e),
	.w6(32'h3bc78a47),
	.w7(32'h3ca03d45),
	.w8(32'h3c24c66a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026993),
	.w1(32'h3cc8d177),
	.w2(32'hbc1482a7),
	.w3(32'h3ca44c77),
	.w4(32'h3c7dc0c0),
	.w5(32'hbc7860e8),
	.w6(32'h3c8c363f),
	.w7(32'h3a632b93),
	.w8(32'hbc20ebee),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13d0ae),
	.w1(32'hbb0167da),
	.w2(32'hbc3426f1),
	.w3(32'hbc325f7d),
	.w4(32'h3b299b0c),
	.w5(32'hbbfbe422),
	.w6(32'h3acc493a),
	.w7(32'hbbc41c1a),
	.w8(32'h3b52f1d1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856b0c),
	.w1(32'hbb29dd4b),
	.w2(32'hbb7dbd13),
	.w3(32'hbb6e165b),
	.w4(32'hbb1efced),
	.w5(32'h3a20b13c),
	.w6(32'hbbc7cc7c),
	.w7(32'hbac3a1a7),
	.w8(32'h3bf3b988),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba8b7),
	.w1(32'hbbcfa656),
	.w2(32'h3b20b17b),
	.w3(32'h3c196a3b),
	.w4(32'hbb02eaa5),
	.w5(32'h3a382ecf),
	.w6(32'hbb6623a2),
	.w7(32'h3b7cbebe),
	.w8(32'h3b57c3af),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c965a),
	.w1(32'h3bc6dc2c),
	.w2(32'h3c384aef),
	.w3(32'hbacf1926),
	.w4(32'h3ba1341c),
	.w5(32'h3c2495e0),
	.w6(32'h3b919c3b),
	.w7(32'h3bd5aaf2),
	.w8(32'h3b0d3ab5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836419),
	.w1(32'h3adce7da),
	.w2(32'h3a9d1901),
	.w3(32'h3a84b867),
	.w4(32'h3b2c4f35),
	.w5(32'h3b16bc78),
	.w6(32'hbba4a05e),
	.w7(32'hb92192fe),
	.w8(32'h3aa5b617),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7198bf),
	.w1(32'h3c7a4587),
	.w2(32'h3b51a37f),
	.w3(32'h3adf3b30),
	.w4(32'h3c3332a3),
	.w5(32'h3c1269ce),
	.w6(32'h3bd1dec6),
	.w7(32'hbad3d956),
	.w8(32'h3b221586),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d9a30),
	.w1(32'hbb0e4a5a),
	.w2(32'hbbe14ef6),
	.w3(32'h3c84d989),
	.w4(32'hba9ba4a0),
	.w5(32'hbb801f01),
	.w6(32'hbb0ff70d),
	.w7(32'hbbad9975),
	.w8(32'h3a5cc0a1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6b6f),
	.w1(32'hb9162988),
	.w2(32'h3c18fb40),
	.w3(32'hbb3076fa),
	.w4(32'h3c1c2deb),
	.w5(32'h3be9deb2),
	.w6(32'h3c6a4fab),
	.w7(32'h3c488f51),
	.w8(32'h3bc35827),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c308187),
	.w1(32'hbbbdb19f),
	.w2(32'hbc886c9f),
	.w3(32'h3bd4f946),
	.w4(32'hbb97aae2),
	.w5(32'hbb920aeb),
	.w6(32'h39a6f812),
	.w7(32'hbb1ee578),
	.w8(32'h3b940e8c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26b326),
	.w1(32'h3b8d5254),
	.w2(32'hbac96d1f),
	.w3(32'hbbbbfa5b),
	.w4(32'h3b96575c),
	.w5(32'h39bf8f1e),
	.w6(32'h3b08ea9d),
	.w7(32'hbae780f6),
	.w8(32'h3bc56dd3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd9b82),
	.w1(32'hbb331f68),
	.w2(32'h3ad7353a),
	.w3(32'h3b5ccb95),
	.w4(32'hbafc8137),
	.w5(32'hba6e69cc),
	.w6(32'hbb897826),
	.w7(32'hbac12e2f),
	.w8(32'hb9af99e0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2da4d9),
	.w1(32'h3a29a86e),
	.w2(32'hbc0d77fb),
	.w3(32'h3ae5260e),
	.w4(32'h3a37e5f7),
	.w5(32'hbba338e3),
	.w6(32'h3af7348b),
	.w7(32'hbc258397),
	.w8(32'hbaf0ff80),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1473d),
	.w1(32'h3bec52c2),
	.w2(32'h3c823b57),
	.w3(32'hbb8752ef),
	.w4(32'h3b68e701),
	.w5(32'h3c2d1267),
	.w6(32'h37c26c98),
	.w7(32'h3b756712),
	.w8(32'h3bedd381),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa33c3),
	.w1(32'hbc3864ba),
	.w2(32'hbc8ab770),
	.w3(32'h3bc44fd2),
	.w4(32'hbba4ea13),
	.w5(32'hbc36b1d8),
	.w6(32'hbbfb2144),
	.w7(32'hbc1ccecd),
	.w8(32'h3bdd3425),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e8592),
	.w1(32'h3bceed0e),
	.w2(32'hbbb4b2ca),
	.w3(32'hbb30a07f),
	.w4(32'h3b97fd03),
	.w5(32'hbbb1385f),
	.w6(32'h3c18b6da),
	.w7(32'hbac62576),
	.w8(32'h3ac5b571),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13be7e),
	.w1(32'h3b055ec3),
	.w2(32'hbb5439c6),
	.w3(32'h3a8627fc),
	.w4(32'hbc44a972),
	.w5(32'hbb499faf),
	.w6(32'h3ba00843),
	.w7(32'hbbfd6845),
	.w8(32'h3bd16b82),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61b4e2),
	.w1(32'h3b803487),
	.w2(32'hbc51bbb1),
	.w3(32'h3bf616f4),
	.w4(32'h3be0e791),
	.w5(32'hbc3e76f4),
	.w6(32'hb98757fc),
	.w7(32'hbc515d18),
	.w8(32'h3ba60f06),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5a402),
	.w1(32'hbb785bde),
	.w2(32'hbb8c5e67),
	.w3(32'hba236747),
	.w4(32'hbb8c2675),
	.w5(32'hbbaddf38),
	.w6(32'hbb4c7761),
	.w7(32'hbb76b1be),
	.w8(32'hbb20a631),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0167),
	.w1(32'h3bbbebab),
	.w2(32'h3c11081e),
	.w3(32'hbbdb480d),
	.w4(32'h3b805003),
	.w5(32'h3bd2418e),
	.w6(32'h3adfd5cd),
	.w7(32'h3bcf71fe),
	.w8(32'h3bb060b8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb48719),
	.w1(32'h3b9b3a0f),
	.w2(32'h3c6e5cbd),
	.w3(32'h3b83d980),
	.w4(32'hbb1d39af),
	.w5(32'h3be6ba90),
	.w6(32'h3b9a2bc1),
	.w7(32'h3c20a9d1),
	.w8(32'h3cda2911),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d136cc8),
	.w1(32'h3c196279),
	.w2(32'hbb157e95),
	.w3(32'h3ca80064),
	.w4(32'h3be623c7),
	.w5(32'hbb0c880b),
	.w6(32'h3c0442f8),
	.w7(32'h3b451c71),
	.w8(32'h3c3fe7b4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7833),
	.w1(32'h3a212919),
	.w2(32'hbb545d31),
	.w3(32'h3b8abbfa),
	.w4(32'hbadfec13),
	.w5(32'hbb8dc5d3),
	.w6(32'hbb31c79c),
	.w7(32'hbb62466a),
	.w8(32'hbb42dd56),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb8225),
	.w1(32'hbc91d35d),
	.w2(32'h3993c811),
	.w3(32'hbb2bc10b),
	.w4(32'hbbfd7f71),
	.w5(32'h3ba5b60d),
	.w6(32'hbbec2e6f),
	.w7(32'hbb8d5216),
	.w8(32'h3a53307a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule