module layer_8_featuremap_185(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb9a7d),
	.w1(32'hbc24403e),
	.w2(32'hbcce737d),
	.w3(32'hbc957b07),
	.w4(32'hbba61faf),
	.w5(32'hbc49e90f),
	.w6(32'hbb82de50),
	.w7(32'hbc25b2f6),
	.w8(32'h3c2664ca),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b40d8),
	.w1(32'hbb807d23),
	.w2(32'h3b14f932),
	.w3(32'h3b227abe),
	.w4(32'hbb90cea3),
	.w5(32'hbb0a3dd1),
	.w6(32'hba17a9c0),
	.w7(32'h3b088210),
	.w8(32'h3a3ba500),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29b64),
	.w1(32'h39ea4746),
	.w2(32'h3ba785cb),
	.w3(32'hbba099d6),
	.w4(32'hbbdb2b0c),
	.w5(32'h3ba9f849),
	.w6(32'hba92e10a),
	.w7(32'hbb860c4a),
	.w8(32'h3b611fb5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90596e),
	.w1(32'h3b5f8ad6),
	.w2(32'hbb8adaa6),
	.w3(32'h3b000597),
	.w4(32'hbbfc0819),
	.w5(32'hbb87ef41),
	.w6(32'h3ba6b3a9),
	.w7(32'hbb94bfd5),
	.w8(32'hbb3e32da),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fa006),
	.w1(32'h3ad52b0c),
	.w2(32'h3b601b0e),
	.w3(32'hbc0492c3),
	.w4(32'h3a6d4894),
	.w5(32'h3af0b474),
	.w6(32'hba151078),
	.w7(32'h3be540de),
	.w8(32'h3b0b7a06),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920918),
	.w1(32'hbc0bc77f),
	.w2(32'hb9d77c21),
	.w3(32'hbbdfbd35),
	.w4(32'hbb6ec7b4),
	.w5(32'h3c29e409),
	.w6(32'hbb82b001),
	.w7(32'h3b8d1040),
	.w8(32'hbb910c58),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9e3dc),
	.w1(32'h3bef4ac2),
	.w2(32'h3ae4b062),
	.w3(32'h3c65f179),
	.w4(32'h3ba395c7),
	.w5(32'h3b67b412),
	.w6(32'h3b5d1cfe),
	.w7(32'h3b597405),
	.w8(32'h3b1d9e7f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e439b),
	.w1(32'h3ca16bef),
	.w2(32'hbb4337ba),
	.w3(32'h3bbd52da),
	.w4(32'h3ba152fe),
	.w5(32'hbb723f2f),
	.w6(32'h3c0bd6ed),
	.w7(32'h3b9386c0),
	.w8(32'hbb46bb0b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ff8eb),
	.w1(32'h3c1f6cf1),
	.w2(32'hbb66f541),
	.w3(32'hbc132963),
	.w4(32'h3bb29c95),
	.w5(32'hbc05a14d),
	.w6(32'h3bca6ef6),
	.w7(32'h3b515236),
	.w8(32'h3b861edc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b8b82),
	.w1(32'hbc3d6bcd),
	.w2(32'hbc3f74cb),
	.w3(32'hbb5fd417),
	.w4(32'hbc6f7b5f),
	.w5(32'hbb3a83e2),
	.w6(32'hbba436b3),
	.w7(32'h3c3e951c),
	.w8(32'h3c54e712),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c949851),
	.w1(32'hbcc13663),
	.w2(32'h3c2a201b),
	.w3(32'h3bf71839),
	.w4(32'hbcefe52f),
	.w5(32'hbc5217b6),
	.w6(32'hbc38978a),
	.w7(32'h3b889e4f),
	.w8(32'hbb0de898),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc586b),
	.w1(32'hba0b320e),
	.w2(32'hbb8a3aaf),
	.w3(32'h3ba4cb32),
	.w4(32'hbbd0b662),
	.w5(32'hbb1ab7f5),
	.w6(32'hba8d27d6),
	.w7(32'h3ba0e942),
	.w8(32'h3ae94648),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02522e),
	.w1(32'hbbd30771),
	.w2(32'hbc2b224c),
	.w3(32'hb9825fdd),
	.w4(32'h3ac5c2bd),
	.w5(32'h3a8c65ab),
	.w6(32'hbb3d8884),
	.w7(32'hbb9c934d),
	.w8(32'h3bf1a9e7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05d795),
	.w1(32'h3aca9609),
	.w2(32'h3b89ae68),
	.w3(32'h398d9127),
	.w4(32'hbc10121c),
	.w5(32'h38c9e57d),
	.w6(32'hba820958),
	.w7(32'h3b83d25e),
	.w8(32'hbae7684e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd59c2),
	.w1(32'h3c013d17),
	.w2(32'hbb721b89),
	.w3(32'h399436bc),
	.w4(32'h3bad51e8),
	.w5(32'h3ae8e41f),
	.w6(32'h3b9bc3ac),
	.w7(32'hbb017424),
	.w8(32'hbb8ebfe7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccc329),
	.w1(32'hbc772920),
	.w2(32'hbbc8ce9c),
	.w3(32'h37fb63ec),
	.w4(32'hbc65e026),
	.w5(32'hbbabc9a5),
	.w6(32'hbc5d8baf),
	.w7(32'hbc168ab5),
	.w8(32'h3c262ba1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb30d26),
	.w1(32'hbbe5b21f),
	.w2(32'hba0becd4),
	.w3(32'h3ca12ee7),
	.w4(32'hbb0f7360),
	.w5(32'hbac61e74),
	.w6(32'h3ba92537),
	.w7(32'hbc1b2924),
	.w8(32'hbc1862ae),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4402ce),
	.w1(32'hbad4860c),
	.w2(32'hb98746ea),
	.w3(32'hbc04c316),
	.w4(32'hbb259078),
	.w5(32'hbb040976),
	.w6(32'hbc51da41),
	.w7(32'h3b1e189b),
	.w8(32'h3c0dccba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d651a87),
	.w1(32'hbc725d0f),
	.w2(32'hbd53d077),
	.w3(32'h3c9b0585),
	.w4(32'hbca784a1),
	.w5(32'hbd2e942c),
	.w6(32'hbb5487d8),
	.w7(32'hbd06d0e7),
	.w8(32'h3c8042b4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabe661),
	.w1(32'hbb88db0e),
	.w2(32'hbbfd0f55),
	.w3(32'h3c9a7373),
	.w4(32'h3b16e10e),
	.w5(32'h3b3de11a),
	.w6(32'h3b991c74),
	.w7(32'h3b21c532),
	.w8(32'h3b89220d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700abe),
	.w1(32'h3c8f1d81),
	.w2(32'hbb460827),
	.w3(32'h3b5a647e),
	.w4(32'h3c5949cf),
	.w5(32'hb9aa46af),
	.w6(32'h3c289161),
	.w7(32'hbab7dd1a),
	.w8(32'hbc1299ab),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64fd4),
	.w1(32'hbbf604cf),
	.w2(32'hbb0b84b6),
	.w3(32'h391f55bf),
	.w4(32'hbc190cb5),
	.w5(32'hbb311556),
	.w6(32'hbb1f21d7),
	.w7(32'hbc0e1bfd),
	.w8(32'hbbebceae),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89be44),
	.w1(32'hbcc9136b),
	.w2(32'hbc891428),
	.w3(32'h3ccbcd33),
	.w4(32'hbd0cea30),
	.w5(32'hbc25ba88),
	.w6(32'hbc82847f),
	.w7(32'hbcb0b06b),
	.w8(32'hbb89c1f8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1dffa0),
	.w1(32'hbba49fc0),
	.w2(32'hbc91fdbf),
	.w3(32'h3caa1563),
	.w4(32'hbb1eba2e),
	.w5(32'hbc0e89ba),
	.w6(32'hbb3383a3),
	.w7(32'hbba6cc29),
	.w8(32'hbc765c1d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79c54a),
	.w1(32'hbbd3e26d),
	.w2(32'hbbe42021),
	.w3(32'hbbcdc15f),
	.w4(32'hbbfe4145),
	.w5(32'h3a6e6d92),
	.w6(32'hba958c1d),
	.w7(32'hbb64a5ad),
	.w8(32'hbc16bab0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91eff),
	.w1(32'h3c2bf133),
	.w2(32'h3aba9dd4),
	.w3(32'h3b896005),
	.w4(32'h3a139f2b),
	.w5(32'h3ade0daa),
	.w6(32'h3c9c2a8d),
	.w7(32'h3beb4598),
	.w8(32'h3ba8969e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab5d7),
	.w1(32'hbc411a26),
	.w2(32'hbb2fa1a7),
	.w3(32'hbbef9252),
	.w4(32'hbc1f4ea3),
	.w5(32'hbb3fd9d2),
	.w6(32'hb9a2cdb3),
	.w7(32'h3b9005e0),
	.w8(32'h3b141aeb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9b66b0),
	.w1(32'h3d0b035e),
	.w2(32'hbd603bb0),
	.w3(32'h3d853913),
	.w4(32'h3cf13e1b),
	.w5(32'hbd8abb41),
	.w6(32'h3d6fa71b),
	.w7(32'h3cb536db),
	.w8(32'hbd378735),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb091e),
	.w1(32'h3a5567ea),
	.w2(32'h3b1594a1),
	.w3(32'hbc088397),
	.w4(32'hbaa48ea1),
	.w5(32'hbbb515aa),
	.w6(32'hbab842fe),
	.w7(32'hbbf24d8c),
	.w8(32'hbb990bc5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbbca3),
	.w1(32'h3a9c1a14),
	.w2(32'h3b6bf047),
	.w3(32'hbc2f7b97),
	.w4(32'h3ad21a50),
	.w5(32'h3c02a278),
	.w6(32'hb9cb8340),
	.w7(32'h3b73ac4e),
	.w8(32'hb9e47746),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1c829),
	.w1(32'h3c041b82),
	.w2(32'h3c17dd18),
	.w3(32'h3c1181f9),
	.w4(32'h3ba14f1a),
	.w5(32'h3a5c98f2),
	.w6(32'h3aa9a5c6),
	.w7(32'h3b9ce57f),
	.w8(32'h3af0e6b9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddfc8c),
	.w1(32'hbc83966b),
	.w2(32'hbc0c940f),
	.w3(32'hbbe3d20d),
	.w4(32'hbb711762),
	.w5(32'hbbfc0e48),
	.w6(32'hbb903ef4),
	.w7(32'hbb839f0f),
	.w8(32'hbb80b99d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d2ba7),
	.w1(32'hbba45e9c),
	.w2(32'h3ccc5fc8),
	.w3(32'h3c3d75c4),
	.w4(32'hbc1288ca),
	.w5(32'h3b8531ef),
	.w6(32'hbb71a5ac),
	.w7(32'h3c662065),
	.w8(32'hbafc6374),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a20d5),
	.w1(32'hba1f60b0),
	.w2(32'hbc025a22),
	.w3(32'hbb6df054),
	.w4(32'h3b2e2730),
	.w5(32'hbbafe2d6),
	.w6(32'h3a9d460b),
	.w7(32'hbb1ec22a),
	.w8(32'h3a984b36),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9651eb),
	.w1(32'h3bec9956),
	.w2(32'h3c1b15ed),
	.w3(32'hbca8c203),
	.w4(32'h3c1b6b8b),
	.w5(32'h3c9b04f3),
	.w6(32'h3ac629aa),
	.w7(32'h3c243e54),
	.w8(32'h3b1e8db5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d73a6),
	.w1(32'h3c4c0a9a),
	.w2(32'h39089af0),
	.w3(32'h3c5ed7fb),
	.w4(32'h3c090ff8),
	.w5(32'h3ae917a4),
	.w6(32'h3b67ec6a),
	.w7(32'h37ef2311),
	.w8(32'hbbfafb6d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6c223),
	.w1(32'h3bd6a530),
	.w2(32'h3b6c82a0),
	.w3(32'h3c45a23c),
	.w4(32'h3bb90bd2),
	.w5(32'h3b8922b6),
	.w6(32'h3b3ed45b),
	.w7(32'hbb0526ec),
	.w8(32'hbc1d8059),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12b986),
	.w1(32'h3c43ff9f),
	.w2(32'hbbcd743f),
	.w3(32'hbbd4d00f),
	.w4(32'h3bdc0ed4),
	.w5(32'hbba3549e),
	.w6(32'h3be60e79),
	.w7(32'hbb1f1222),
	.w8(32'hbbdbc411),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e1afe),
	.w1(32'hbbaa6fa8),
	.w2(32'hbc377aeb),
	.w3(32'hbc3e9c13),
	.w4(32'hbc1bca34),
	.w5(32'hbc31f0d6),
	.w6(32'hbb085ad8),
	.w7(32'hbc0c7bdd),
	.w8(32'hbb7770be),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fc53),
	.w1(32'h3c0d0217),
	.w2(32'h3a82f5d1),
	.w3(32'h3b6ece3b),
	.w4(32'h3b8de390),
	.w5(32'hbbf4180c),
	.w6(32'h3ac4dcfc),
	.w7(32'h3b99bc31),
	.w8(32'h3ad6edca),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa92aa),
	.w1(32'h3b181581),
	.w2(32'h3bae5690),
	.w3(32'h3b00d6e0),
	.w4(32'h3aef895c),
	.w5(32'h3c09c0ed),
	.w6(32'h3bb77797),
	.w7(32'h3bde1654),
	.w8(32'h3ca101a2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99b27d),
	.w1(32'hbbc2ca9f),
	.w2(32'hbc2fe8d3),
	.w3(32'hbb3ea917),
	.w4(32'hbbb1f4f3),
	.w5(32'hbc27425a),
	.w6(32'h3b89674b),
	.w7(32'hbbaedb5d),
	.w8(32'hb8f3cb0a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b99e7),
	.w1(32'hbbbbf457),
	.w2(32'h3c94434d),
	.w3(32'h3b1c693c),
	.w4(32'hbba13043),
	.w5(32'h3c48af3e),
	.w6(32'hbc335a99),
	.w7(32'hbaee5dc5),
	.w8(32'hbc4a1d04),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe0538),
	.w1(32'hbc997375),
	.w2(32'hbb45de40),
	.w3(32'hbc0b40bd),
	.w4(32'hbc4d95f8),
	.w5(32'hbc2bdde9),
	.w6(32'hbc3d12bb),
	.w7(32'hbbda33c1),
	.w8(32'h3b56fee9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d244137),
	.w1(32'hbbb66215),
	.w2(32'hbc4dfc11),
	.w3(32'h3cd84891),
	.w4(32'hbc8a1ec0),
	.w5(32'hbcafd0cd),
	.w6(32'h3c642cf4),
	.w7(32'hbc38c2bd),
	.w8(32'hbc5bded6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0c7e),
	.w1(32'hbbd8d377),
	.w2(32'hbc93ccad),
	.w3(32'hba294386),
	.w4(32'hbc4d1113),
	.w5(32'hbc46dcd1),
	.w6(32'h3b31da0c),
	.w7(32'hbbfb29ec),
	.w8(32'hbb2ab19a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b4d0f),
	.w1(32'hbc70ddb1),
	.w2(32'hbbddb6b6),
	.w3(32'hbb58607d),
	.w4(32'hbc677740),
	.w5(32'hb9e0689d),
	.w6(32'hbc1127bc),
	.w7(32'hbc478923),
	.w8(32'hbb5b504e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e5d3e),
	.w1(32'hbc701c38),
	.w2(32'hbcc18328),
	.w3(32'h3c73df18),
	.w4(32'hbc6622ff),
	.w5(32'hbcc67f13),
	.w6(32'hbb64a271),
	.w7(32'hbc93337b),
	.w8(32'hbc1e97ac),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52aade),
	.w1(32'hbc1506cc),
	.w2(32'h3b9c5974),
	.w3(32'h385f2d2f),
	.w4(32'hbae91403),
	.w5(32'h3c4069ea),
	.w6(32'hbbf84ada),
	.w7(32'hbc135ed2),
	.w8(32'hbbd2a6f7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c807fda),
	.w1(32'hbb088475),
	.w2(32'hbc3cae78),
	.w3(32'h3c0532ca),
	.w4(32'hbc01cb2d),
	.w5(32'hbcc0637e),
	.w6(32'h3a8b1087),
	.w7(32'h3b615529),
	.w8(32'h3c1d7e8e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e4671),
	.w1(32'hb9dd2c60),
	.w2(32'hbc1ef3d9),
	.w3(32'hbb62c6ce),
	.w4(32'h3a6f5122),
	.w5(32'hbba7ff32),
	.w6(32'hbc40d5ce),
	.w7(32'hbbfbd994),
	.w8(32'h3bf56d78),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0998a4),
	.w1(32'hbc236fc1),
	.w2(32'hbca091d4),
	.w3(32'h3c859c3d),
	.w4(32'hbbdd73c9),
	.w5(32'hbc93f32f),
	.w6(32'h3bc7fcc1),
	.w7(32'hbcb69df2),
	.w8(32'h3bab91fa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf83b1a),
	.w1(32'h3b8d3db1),
	.w2(32'hba0765e8),
	.w3(32'h3c1dbb99),
	.w4(32'h3b7e67d6),
	.w5(32'h39a64b59),
	.w6(32'h3bdba680),
	.w7(32'h3b4647db),
	.w8(32'h3b5e61c4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b477870),
	.w1(32'hbc3495f5),
	.w2(32'hbcaded89),
	.w3(32'h3b7e7d7f),
	.w4(32'hbc52844f),
	.w5(32'hbc896474),
	.w6(32'hbb5a2ea3),
	.w7(32'hbc5e5167),
	.w8(32'hbc1bac57),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc2dd3),
	.w1(32'h3bd2d1ce),
	.w2(32'h3beb61ad),
	.w3(32'hbb4cfd96),
	.w4(32'h3bbea3a1),
	.w5(32'hba1e8c3e),
	.w6(32'hbac21b2d),
	.w7(32'h3a85a02a),
	.w8(32'h3bf41779),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d12e646),
	.w1(32'hbbcd2ce6),
	.w2(32'hbd025b8b),
	.w3(32'h3c1e8343),
	.w4(32'hbc121788),
	.w5(32'hbd04faa8),
	.w6(32'hbc121810),
	.w7(32'h3af8aab3),
	.w8(32'h3b6656da),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7fecbd),
	.w1(32'h3bbc3cd2),
	.w2(32'h3ce6202a),
	.w3(32'h3c1cdee2),
	.w4(32'hbab9f767),
	.w5(32'h3c8ea138),
	.w6(32'hbbc3b24c),
	.w7(32'h3bb6aa77),
	.w8(32'hbc5dc49c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98ed2a),
	.w1(32'h3abd82d5),
	.w2(32'h3c06612d),
	.w3(32'hbc23c2bc),
	.w4(32'h3b59dba9),
	.w5(32'h3b864534),
	.w6(32'h3b2f6511),
	.w7(32'h39bddead),
	.w8(32'hbc35e664),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5da89),
	.w1(32'h3a73abf2),
	.w2(32'hbc28f7cc),
	.w3(32'h3ab72237),
	.w4(32'hbac5cced),
	.w5(32'hbc7a90a1),
	.w6(32'h3c0275cc),
	.w7(32'hbb87270e),
	.w8(32'hbc52dbff),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc948c6b),
	.w1(32'hbbe7d262),
	.w2(32'hbc4d93cb),
	.w3(32'hbc4889dc),
	.w4(32'hbc794051),
	.w5(32'hbbd335d2),
	.w6(32'hbb74a5f8),
	.w7(32'hbc922b2a),
	.w8(32'hbc1b1cca),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf338f7),
	.w1(32'h3ae883a5),
	.w2(32'hba90cda7),
	.w3(32'hb994a69d),
	.w4(32'hbb0bbb00),
	.w5(32'hbaa0a6b7),
	.w6(32'h3bb35714),
	.w7(32'h3bb3d0e5),
	.w8(32'h3b7f9bc5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8c9df),
	.w1(32'h3c122131),
	.w2(32'hbc334a22),
	.w3(32'h3b038c71),
	.w4(32'hbae82ad7),
	.w5(32'h39697ce5),
	.w6(32'h3c642812),
	.w7(32'hbb93f8d9),
	.w8(32'hbbf1c610),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6a551),
	.w1(32'h3a82e2cb),
	.w2(32'hbc0613b2),
	.w3(32'h3bc170ba),
	.w4(32'h3bc0d1c5),
	.w5(32'h3a632ce1),
	.w6(32'h3a8d193b),
	.w7(32'h3a6b3bf4),
	.w8(32'h3bb357dc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b39d0),
	.w1(32'hbb3c3a73),
	.w2(32'h3a85a00d),
	.w3(32'hbc09c94e),
	.w4(32'hbb83c1b8),
	.w5(32'hbbb691bb),
	.w6(32'hbb14f489),
	.w7(32'h3a258be7),
	.w8(32'hbafb7ca5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba506b80),
	.w1(32'hbb5dc8aa),
	.w2(32'hbae38562),
	.w3(32'hbc0f5c10),
	.w4(32'hba828869),
	.w5(32'hba988b40),
	.w6(32'hba272fa9),
	.w7(32'hbb85bfc6),
	.w8(32'hbbb5ef1e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f25e64),
	.w1(32'h3b1579bc),
	.w2(32'hbb309ccc),
	.w3(32'h39aa4822),
	.w4(32'hbb0b2ceb),
	.w5(32'hbbeccd5f),
	.w6(32'h3c6583f6),
	.w7(32'h3b872fa6),
	.w8(32'hba0aa5e2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd81f3e),
	.w1(32'hbc333f91),
	.w2(32'hbc706958),
	.w3(32'hbb2da185),
	.w4(32'hbbb8d7fc),
	.w5(32'hba395f2c),
	.w6(32'hbc5fec67),
	.w7(32'hbc5edc38),
	.w8(32'h3aedc8be),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e5c92),
	.w1(32'h3beb50e6),
	.w2(32'hbc1344ea),
	.w3(32'h3c6f163b),
	.w4(32'h3a209ea9),
	.w5(32'hbb018feb),
	.w6(32'hbb9d0317),
	.w7(32'hbb3614b9),
	.w8(32'h3c0851f8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5517f3),
	.w1(32'hbba1e46b),
	.w2(32'hbc348477),
	.w3(32'h3c49b153),
	.w4(32'hbbc7a5ae),
	.w5(32'hbc297add),
	.w6(32'hbbdde9b3),
	.w7(32'h3b5112c6),
	.w8(32'hbbe66383),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf1a4),
	.w1(32'h3ce3c70f),
	.w2(32'hbc983e8c),
	.w3(32'h3c9e7842),
	.w4(32'h3c13c9bd),
	.w5(32'hbcd35220),
	.w6(32'h3c9b4215),
	.w7(32'hbc99212b),
	.w8(32'hbd0fb71f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4d88),
	.w1(32'hbb2e477d),
	.w2(32'hbcc32cc8),
	.w3(32'h3bd33059),
	.w4(32'hba8275e3),
	.w5(32'hbc896172),
	.w6(32'h3becd464),
	.w7(32'hba4b0a14),
	.w8(32'h3c6ef95b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13a946),
	.w1(32'h3bf39b65),
	.w2(32'h3c857862),
	.w3(32'h3c8dfaa2),
	.w4(32'h3b0f7dc2),
	.w5(32'h3c08553b),
	.w6(32'h3c251bc7),
	.w7(32'h3b94b718),
	.w8(32'hbb9d05ae),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c164d),
	.w1(32'hbbe465ea),
	.w2(32'h3c0309a3),
	.w3(32'h3b07db06),
	.w4(32'hbb0a410f),
	.w5(32'h3c0abf48),
	.w6(32'hbbf4219c),
	.w7(32'hbb1e4a47),
	.w8(32'hbae69aa6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79c5b7),
	.w1(32'h3b804c18),
	.w2(32'h3c3e6b31),
	.w3(32'h3c2684f8),
	.w4(32'hbba3cc50),
	.w5(32'h3c0376c8),
	.w6(32'hbb85bd10),
	.w7(32'h3c645a36),
	.w8(32'hbb9e1bc9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03936e),
	.w1(32'hbb1e79f7),
	.w2(32'hbc0e044c),
	.w3(32'h3b27d111),
	.w4(32'hbb68431e),
	.w5(32'h3a74f644),
	.w6(32'h3a748fb9),
	.w7(32'hbadba3c2),
	.w8(32'h3ac7a5b7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0942d2),
	.w1(32'h3b85c520),
	.w2(32'h3cdc4aac),
	.w3(32'h3cadd282),
	.w4(32'hbb8f264b),
	.w5(32'h3ce2316d),
	.w6(32'hbbacc91f),
	.w7(32'h3c7adb4d),
	.w8(32'h3c429c87),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce8073),
	.w1(32'hba1fa704),
	.w2(32'h3c0d5b67),
	.w3(32'h3cdb4b3a),
	.w4(32'hbbbdd26d),
	.w5(32'hbb1241b2),
	.w6(32'hbb8f8eec),
	.w7(32'hbb6961f3),
	.w8(32'hbbcbc563),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c2172),
	.w1(32'h3c32d297),
	.w2(32'h3bf1482b),
	.w3(32'h3c212621),
	.w4(32'h3b65bc37),
	.w5(32'hba0bbd8c),
	.w6(32'h3ba2e93a),
	.w7(32'hbbaf4e56),
	.w8(32'h3bee06ce),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0eacfe),
	.w1(32'hbc967df5),
	.w2(32'hbcded4ab),
	.w3(32'h3bf4f86d),
	.w4(32'hbca899b4),
	.w5(32'hbcc4339e),
	.w6(32'hbba1b8d9),
	.w7(32'hbc1ebab4),
	.w8(32'h3c162715),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23c256),
	.w1(32'hbbc8605a),
	.w2(32'h3bda380c),
	.w3(32'h3b741fa3),
	.w4(32'hbc4a074d),
	.w5(32'hbb503c41),
	.w6(32'hbbdb2f3a),
	.w7(32'h3b8ba6f0),
	.w8(32'h3afd909d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c892226),
	.w1(32'h3c67abdc),
	.w2(32'h3c05477d),
	.w3(32'h3bf2e685),
	.w4(32'h3b98b704),
	.w5(32'h3bd10def),
	.w6(32'h3bfb84ec),
	.w7(32'h3b80eb55),
	.w8(32'hbba3105a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4356e),
	.w1(32'hbc61e6d9),
	.w2(32'hbb08cf17),
	.w3(32'h3a6a3244),
	.w4(32'h3a866f8a),
	.w5(32'hbb9495ea),
	.w6(32'h3c6a38b5),
	.w7(32'h3c0feb1a),
	.w8(32'hbc6fc7e4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba24f5e),
	.w1(32'hbc6e6b7e),
	.w2(32'hbb8374a0),
	.w3(32'h3b5d134e),
	.w4(32'hbc45c117),
	.w5(32'hbb0c6d97),
	.w6(32'hbb95e72c),
	.w7(32'hbc1d1dca),
	.w8(32'h3be3b4dc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0aca76),
	.w1(32'h3d04090d),
	.w2(32'h3c08356e),
	.w3(32'h3ca3e881),
	.w4(32'h3bd19284),
	.w5(32'h3c384bde),
	.w6(32'h3bc14b89),
	.w7(32'hbbb210b3),
	.w8(32'h3c59f3bd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ae91e),
	.w1(32'h3be5579a),
	.w2(32'hbc052406),
	.w3(32'h3c93e8e3),
	.w4(32'hbb58eece),
	.w5(32'hbc3e7d3d),
	.w6(32'h3c74a2d5),
	.w7(32'h3c39491a),
	.w8(32'h3c2392fb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af72c7e),
	.w1(32'hbc563bd7),
	.w2(32'h3b32689e),
	.w3(32'hb9eb7536),
	.w4(32'h3bb80dcc),
	.w5(32'h3a9dbb36),
	.w6(32'hbb97a5a4),
	.w7(32'hbc01bb7d),
	.w8(32'h3a8b8073),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf36bd),
	.w1(32'h39f37c34),
	.w2(32'h3aec93b4),
	.w3(32'h3c2e494e),
	.w4(32'h3a5d856e),
	.w5(32'hbb07f3e9),
	.w6(32'h3ad9d96c),
	.w7(32'h3c2184dd),
	.w8(32'h3c40e9c5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66262c),
	.w1(32'h3a72480f),
	.w2(32'h3bafa593),
	.w3(32'h39cb6f37),
	.w4(32'h3940b1e8),
	.w5(32'h3b8b60ff),
	.w6(32'h3bf8d027),
	.w7(32'h3b8d55c8),
	.w8(32'hba301a50),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab6096),
	.w1(32'h3b496748),
	.w2(32'h3a50ada3),
	.w3(32'hb9c1c77e),
	.w4(32'hbbbe421b),
	.w5(32'hbbb9a79d),
	.w6(32'hbb8e64cf),
	.w7(32'h3a8d5bac),
	.w8(32'hbacc083b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9c52e),
	.w1(32'hbbccd645),
	.w2(32'h3c54b854),
	.w3(32'hbbc885dc),
	.w4(32'hbc0033f6),
	.w5(32'h3b9195f1),
	.w6(32'hbc307581),
	.w7(32'hbb47a7f9),
	.w8(32'h3bc70d66),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8266fb),
	.w1(32'hbc3686f3),
	.w2(32'h3bf19626),
	.w3(32'h3b01d356),
	.w4(32'h3b9cd8fc),
	.w5(32'h3c1fcef5),
	.w6(32'hbbe1ed02),
	.w7(32'hbad10daa),
	.w8(32'hba0de0f1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c108469),
	.w1(32'h3c01218e),
	.w2(32'h3b64b464),
	.w3(32'h3c770a2a),
	.w4(32'h3baf1088),
	.w5(32'hba833ca9),
	.w6(32'h3b7fb1ec),
	.w7(32'h3bb64b8e),
	.w8(32'h3ad0f925),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9c056),
	.w1(32'h3b2c136f),
	.w2(32'h3c06caa2),
	.w3(32'hbc110ea7),
	.w4(32'h3b8491de),
	.w5(32'h3bb825ba),
	.w6(32'h3b45da05),
	.w7(32'h3bc0ae5e),
	.w8(32'h3b8ecf81),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b728482),
	.w1(32'hbc0603d9),
	.w2(32'hbad4748d),
	.w3(32'h3ae2c604),
	.w4(32'hbc162b5f),
	.w5(32'hbb440e50),
	.w6(32'hbb0727cd),
	.w7(32'hba50a118),
	.w8(32'h3b4297c5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c047c1f),
	.w1(32'hbc275b29),
	.w2(32'h3c8bb27d),
	.w3(32'h3b9c95e7),
	.w4(32'hbc200098),
	.w5(32'h3c20441f),
	.w6(32'hbc804d91),
	.w7(32'h3b889aa9),
	.w8(32'h3c8bb59d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d21ca59),
	.w1(32'h3c857660),
	.w2(32'hbbbabc00),
	.w3(32'h3cbd9a98),
	.w4(32'h3ba047ef),
	.w5(32'hbc60190c),
	.w6(32'h3c71d1ad),
	.w7(32'hbb6b9d7c),
	.w8(32'hbc0e3b53),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb727fd),
	.w1(32'h3c543937),
	.w2(32'h3cc52f06),
	.w3(32'hbb49e782),
	.w4(32'h3b23f00d),
	.w5(32'h3c8e5376),
	.w6(32'h3c294835),
	.w7(32'h3bbb0d5f),
	.w8(32'h3b44a992),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c9059),
	.w1(32'hbc6264bb),
	.w2(32'h3b6349bc),
	.w3(32'h3bb4c58b),
	.w4(32'hbc87bf30),
	.w5(32'hbbaf5b6b),
	.w6(32'hbc955da6),
	.w7(32'hbbc0cce2),
	.w8(32'h3b96f0cc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd8615),
	.w1(32'hbc88b079),
	.w2(32'hbba9b2a0),
	.w3(32'h3c8e69da),
	.w4(32'hbc672161),
	.w5(32'hbb3c0a1b),
	.w6(32'hbc42d4cb),
	.w7(32'hbcc0b25b),
	.w8(32'hbb4140b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85681c),
	.w1(32'hbcb97216),
	.w2(32'h3cec0d4d),
	.w3(32'h3c1c500b),
	.w4(32'hbc185918),
	.w5(32'h3d05b688),
	.w6(32'hbc7d2e6a),
	.w7(32'h3c18a603),
	.w8(32'hbb86b40f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35c641),
	.w1(32'h3b2f8489),
	.w2(32'h3b604548),
	.w3(32'h3c14b17b),
	.w4(32'h3c10abf8),
	.w5(32'h3b9214ff),
	.w6(32'h3b175751),
	.w7(32'h3c0af8af),
	.w8(32'h3bcd1b06),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b789ff6),
	.w1(32'h3891b170),
	.w2(32'hbc6876da),
	.w3(32'hbba9a8ea),
	.w4(32'h3a2bdb94),
	.w5(32'hbc406dd4),
	.w6(32'hbc2165d6),
	.w7(32'hbc36e988),
	.w8(32'hbc440ee3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95477e),
	.w1(32'h3babcc6b),
	.w2(32'h3c4b2bf1),
	.w3(32'hbc807d66),
	.w4(32'h3bc8ce94),
	.w5(32'hba80bb5e),
	.w6(32'h3c06802f),
	.w7(32'h3c15627c),
	.w8(32'hba724f95),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66198d),
	.w1(32'hbc32f37b),
	.w2(32'h3c6c803a),
	.w3(32'hbb0db31f),
	.w4(32'hba5f7eb9),
	.w5(32'h3a9356a1),
	.w6(32'hbb82fee7),
	.w7(32'h3ab39592),
	.w8(32'hbbe79297),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd82773),
	.w1(32'hbcb34e5b),
	.w2(32'h3b91dae4),
	.w3(32'hbbedc99f),
	.w4(32'hbc9fb8e0),
	.w5(32'h3b47155b),
	.w6(32'hbccce52f),
	.w7(32'hbbb1e031),
	.w8(32'h3a97e2b1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b1fc6),
	.w1(32'h3c2828c5),
	.w2(32'hbc4e6ec1),
	.w3(32'h3ca7e770),
	.w4(32'h3c18aa97),
	.w5(32'hbc098e8e),
	.w6(32'h3c60222a),
	.w7(32'hbb9651ce),
	.w8(32'hbc0739b1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aaa38),
	.w1(32'h3bc4990d),
	.w2(32'h3bab4d4d),
	.w3(32'h3bf0dd28),
	.w4(32'hbb876472),
	.w5(32'hbbbd4fb4),
	.w6(32'hbae2a830),
	.w7(32'h3bb2de44),
	.w8(32'h3bc6d2a4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ea46b),
	.w1(32'h3c0f7a94),
	.w2(32'h3c18149a),
	.w3(32'h3a213b18),
	.w4(32'h3be8c312),
	.w5(32'h3c57b16c),
	.w6(32'hba85c929),
	.w7(32'hbb1e42df),
	.w8(32'hbaaf1dfb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006231),
	.w1(32'h3c657e93),
	.w2(32'h39c24c99),
	.w3(32'hbac73306),
	.w4(32'h3c859678),
	.w5(32'h3be2f8d6),
	.w6(32'h3c4f9a28),
	.w7(32'h3be8d525),
	.w8(32'hbb190956),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1267d9),
	.w1(32'h3a5ee570),
	.w2(32'h3ac7d5ed),
	.w3(32'hbb3342d2),
	.w4(32'h3b23d6d1),
	.w5(32'h3a7b863d),
	.w6(32'h3a9ce927),
	.w7(32'h3a9ce272),
	.w8(32'h3a078722),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90f5db),
	.w1(32'h3a5783ec),
	.w2(32'h3beb63b0),
	.w3(32'h3b14ccfc),
	.w4(32'h3b1c77a1),
	.w5(32'h3c1b804b),
	.w6(32'h39bab43c),
	.w7(32'h3b2100d8),
	.w8(32'h3bbb8f16),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3b7e),
	.w1(32'hbb8e0a95),
	.w2(32'h3a3bb644),
	.w3(32'hbb39d130),
	.w4(32'hbb00ea67),
	.w5(32'h3b081801),
	.w6(32'hba8faa1e),
	.w7(32'h3917f46c),
	.w8(32'h3b5a2165),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4abe0),
	.w1(32'h3bab2999),
	.w2(32'h3bd9945c),
	.w3(32'hb9b6b9a5),
	.w4(32'hb8231724),
	.w5(32'h3c04faeb),
	.w6(32'h3a85e82d),
	.w7(32'h3b850d65),
	.w8(32'h3bc5488f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a5218),
	.w1(32'h3af47f95),
	.w2(32'h3bb674bd),
	.w3(32'h39868ac4),
	.w4(32'h3b715fac),
	.w5(32'h3b6ea76d),
	.w6(32'hbb81842c),
	.w7(32'hbc004d9e),
	.w8(32'hbc23902c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c176a02),
	.w1(32'hbb5d3aca),
	.w2(32'hbc2fa89c),
	.w3(32'h3ac4fff9),
	.w4(32'hbb8a3857),
	.w5(32'hbc614f5e),
	.w6(32'hbadcd028),
	.w7(32'hbb523340),
	.w8(32'h3a95146a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6225b6),
	.w1(32'hbb54551b),
	.w2(32'hba86a988),
	.w3(32'hbbe170e0),
	.w4(32'hba9bb676),
	.w5(32'hba9814de),
	.w6(32'hbaefb22a),
	.w7(32'hbb46b465),
	.w8(32'hbb4f5f46),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1679a5),
	.w1(32'hb89e618a),
	.w2(32'hbc4537b2),
	.w3(32'hbb11f02c),
	.w4(32'h3b969b60),
	.w5(32'hbc42ce8d),
	.w6(32'h3bf4f7fb),
	.w7(32'hbb849713),
	.w8(32'h3c16d16a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b753fff),
	.w1(32'h3bbce966),
	.w2(32'h3bc015df),
	.w3(32'h3c80e16d),
	.w4(32'h3b99ab48),
	.w5(32'h3b3ee34a),
	.w6(32'h3bac3b80),
	.w7(32'h3c19f25e),
	.w8(32'h3bf1bddf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ba15b),
	.w1(32'hbc5982cb),
	.w2(32'h3b16095f),
	.w3(32'hbb59259f),
	.w4(32'hbc09acfb),
	.w5(32'hbc216a6c),
	.w6(32'hba134365),
	.w7(32'h3c69a6a6),
	.w8(32'h3c02c605),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bf24d),
	.w1(32'hbb64d915),
	.w2(32'hbbdcd63d),
	.w3(32'h3824a233),
	.w4(32'hbb9164a3),
	.w5(32'hbc0af568),
	.w6(32'h3b6b8565),
	.w7(32'h3a8dadb2),
	.w8(32'hb9dd5b61),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbade79c),
	.w1(32'hbc7f7649),
	.w2(32'hbc6e61ef),
	.w3(32'h3b20f444),
	.w4(32'hbc81bd29),
	.w5(32'hbca3bae3),
	.w6(32'hbba80030),
	.w7(32'hbbc3690d),
	.w8(32'hba83781a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af94f84),
	.w1(32'hbc7d89e6),
	.w2(32'hb9225bc3),
	.w3(32'hbbf91216),
	.w4(32'hbc3e53f7),
	.w5(32'hbbc75ed8),
	.w6(32'hbc2f4f48),
	.w7(32'h3bbbaf3b),
	.w8(32'h3bebc663),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85d1d4),
	.w1(32'hbbbc68d6),
	.w2(32'h3bb07846),
	.w3(32'hba9a0e5a),
	.w4(32'hbb8a1e40),
	.w5(32'h3ac8d1d3),
	.w6(32'hbb742777),
	.w7(32'h3b9bc503),
	.w8(32'h3b73403e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0b90e),
	.w1(32'hbac6e06a),
	.w2(32'h3b32f758),
	.w3(32'hbb3864dc),
	.w4(32'h398cafcc),
	.w5(32'h3b5cb446),
	.w6(32'h3ac54575),
	.w7(32'h3bbbd788),
	.w8(32'h3b0770d0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b508f11),
	.w1(32'hbbf52fc5),
	.w2(32'hbc132d6d),
	.w3(32'h3ab393e7),
	.w4(32'hbbce66de),
	.w5(32'hbbac7bef),
	.w6(32'hbb7c6dd9),
	.w7(32'hbb99686e),
	.w8(32'hbaf1eb92),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90454e),
	.w1(32'hba194649),
	.w2(32'hbbd1308d),
	.w3(32'hbc296782),
	.w4(32'h3b139c43),
	.w5(32'hbb89c97a),
	.w6(32'hbb83d398),
	.w7(32'hb9cb2057),
	.w8(32'hbbf7ab5b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29968b),
	.w1(32'hbabe6aa8),
	.w2(32'hbab8aa72),
	.w3(32'h3b4a2ae8),
	.w4(32'hba771ca6),
	.w5(32'h39e4132f),
	.w6(32'h39a5a256),
	.w7(32'h3af16e4f),
	.w8(32'h3aac9424),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02484b),
	.w1(32'hbc4010df),
	.w2(32'hbc6461ec),
	.w3(32'h3c0c214d),
	.w4(32'hbc5d44c2),
	.w5(32'hbc827cd7),
	.w6(32'h3b69e5bf),
	.w7(32'hbbf30c48),
	.w8(32'hbb9c83ce),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule