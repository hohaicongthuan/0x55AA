module layer_6_featuremap_63(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf8862),
	.w1(32'h3bdb5cc1),
	.w2(32'hbad9a8ee),
	.w3(32'h3a9bd7f3),
	.w4(32'hba0fab40),
	.w5(32'h3a240728),
	.w6(32'h3b4096b0),
	.w7(32'hba76e12a),
	.w8(32'h3b8f2ce0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf4fde),
	.w1(32'h3b28ba5d),
	.w2(32'h3b24fd78),
	.w3(32'h3a935da9),
	.w4(32'hbaff94e0),
	.w5(32'h3a09d5da),
	.w6(32'h3baaaef7),
	.w7(32'hbb51a2b4),
	.w8(32'hbc6bc10c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26da7),
	.w1(32'hbc8df143),
	.w2(32'h3a22381b),
	.w3(32'h3b70037a),
	.w4(32'h3a688d3e),
	.w5(32'hbb95ae32),
	.w6(32'h3ab52e5d),
	.w7(32'hbb6de027),
	.w8(32'hbb2f6256),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58ad78),
	.w1(32'hbabd193d),
	.w2(32'h3b8db580),
	.w3(32'h3794ccdf),
	.w4(32'h3bc78379),
	.w5(32'h3b8eb4a1),
	.w6(32'hbb62964f),
	.w7(32'h3b872cc0),
	.w8(32'h39ac930b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9200f),
	.w1(32'hbb722a0e),
	.w2(32'hbc74dcb8),
	.w3(32'hbc8d4fc5),
	.w4(32'hbc9496ef),
	.w5(32'h3bb7f1b2),
	.w6(32'hbcd2b048),
	.w7(32'hbd224af0),
	.w8(32'hbcc6d08f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91a194),
	.w1(32'hbae9cb9e),
	.w2(32'hbb9c8d2b),
	.w3(32'hbbf4bc26),
	.w4(32'h38957cd2),
	.w5(32'h3c1bbf03),
	.w6(32'hbbdfaf22),
	.w7(32'hbb9a8ac3),
	.w8(32'h3c2ba0d7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819438),
	.w1(32'hbc1a9581),
	.w2(32'h3bcf5289),
	.w3(32'hbbb9b312),
	.w4(32'hbb7b6d01),
	.w5(32'hbc378b7b),
	.w6(32'hbb2d06d5),
	.w7(32'h3bfd007c),
	.w8(32'hbc03e173),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a782bf2),
	.w1(32'hbc88f40a),
	.w2(32'h3c170e33),
	.w3(32'h3c70bc6d),
	.w4(32'hbb2edd13),
	.w5(32'h3c288dc4),
	.w6(32'h3c5d4fc1),
	.w7(32'h3ccfed6f),
	.w8(32'h3c240a32),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2a37b),
	.w1(32'h3ccd4d3e),
	.w2(32'h3b1f2881),
	.w3(32'hbcb1d208),
	.w4(32'hbca3e45b),
	.w5(32'h3bb98410),
	.w6(32'hbc29d54a),
	.w7(32'hbd1594d7),
	.w8(32'hbd188621),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced7596),
	.w1(32'hb9eb7423),
	.w2(32'hba2deec6),
	.w3(32'hbb9917ce),
	.w4(32'h3aec918d),
	.w5(32'h3c07855a),
	.w6(32'hbb64a835),
	.w7(32'hbb31791a),
	.w8(32'h3ba079b9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a239074),
	.w1(32'hbc37d920),
	.w2(32'hbc3c160b),
	.w3(32'hba4f2e23),
	.w4(32'hbcb0c7b2),
	.w5(32'hbcda7375),
	.w6(32'hbc938b16),
	.w7(32'hbd17006d),
	.w8(32'hbce424d6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bcb4f),
	.w1(32'h3c691686),
	.w2(32'hbb022894),
	.w3(32'h3b938b3a),
	.w4(32'h3ab6852c),
	.w5(32'h3d08bd67),
	.w6(32'h3bc20cc2),
	.w7(32'hbb444fba),
	.w8(32'h3cd34c72),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabec59e),
	.w1(32'h388964a4),
	.w2(32'h3c1a0eec),
	.w3(32'hbb088f16),
	.w4(32'h3bd71320),
	.w5(32'hbb63ec59),
	.w6(32'h3a94ba49),
	.w7(32'h3c0bc6d4),
	.w8(32'hbbe39529),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52b9b5),
	.w1(32'h3c669f29),
	.w2(32'h39637a70),
	.w3(32'hbbc5155d),
	.w4(32'h3bdcff39),
	.w5(32'h3c209b83),
	.w6(32'hbb833542),
	.w7(32'hbd0feec0),
	.w8(32'hbc25d14a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca291a8),
	.w1(32'hba9572bf),
	.w2(32'h3a8708aa),
	.w3(32'hbaf764b4),
	.w4(32'hbb515001),
	.w5(32'h3974f861),
	.w6(32'h3a6ec5b7),
	.w7(32'h3b597b81),
	.w8(32'h3b8accc2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68621e),
	.w1(32'h3baaec0c),
	.w2(32'h3b7be8c3),
	.w3(32'h3a7b8b2b),
	.w4(32'h386029e4),
	.w5(32'hbb9da385),
	.w6(32'h3b2505a3),
	.w7(32'hb9ce5da2),
	.w8(32'hbbb0f62f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba890dc),
	.w1(32'h3cca5312),
	.w2(32'h3a194af2),
	.w3(32'hbc29945e),
	.w4(32'hbcbdb8ec),
	.w5(32'h3c1b3012),
	.w6(32'hbc02d5d8),
	.w7(32'hbd12c1af),
	.w8(32'hbb8879e8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8685dd),
	.w1(32'h3b71013a),
	.w2(32'h3bf07f55),
	.w3(32'hba2a97e5),
	.w4(32'h3b12e641),
	.w5(32'h3bd23309),
	.w6(32'h3ace6ba1),
	.w7(32'h3b5eb84a),
	.w8(32'h3b997ff7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04af83),
	.w1(32'hba0ed6ea),
	.w2(32'h3accf865),
	.w3(32'h3b2561f2),
	.w4(32'h3b6d9b68),
	.w5(32'h3b94c064),
	.w6(32'h3b5c4868),
	.w7(32'h3bb35317),
	.w8(32'h3c0cbe3b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb95e62),
	.w1(32'h3d2b4200),
	.w2(32'h3bb6355f),
	.w3(32'h3c39cce3),
	.w4(32'hbc24e7b8),
	.w5(32'h3d214c9c),
	.w6(32'h3d1dcdbd),
	.w7(32'hbc552471),
	.w8(32'h3c9352f9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeefcd9),
	.w1(32'h3b3bab7f),
	.w2(32'h3b8191c2),
	.w3(32'h3b522a3b),
	.w4(32'h3a5aa764),
	.w5(32'h3ad15194),
	.w6(32'h3b837fc4),
	.w7(32'h3bb05bdd),
	.w8(32'hba82e2ba),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898d58),
	.w1(32'h3bb5ec93),
	.w2(32'h3c0a1dfd),
	.w3(32'h3b6110ae),
	.w4(32'h3ba52d38),
	.w5(32'hbbc1dc39),
	.w6(32'h3b2daca7),
	.w7(32'h3b04cc1e),
	.w8(32'hbc44b400),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd680f),
	.w1(32'hbd33f35f),
	.w2(32'hbc35a5b6),
	.w3(32'hbc97ba52),
	.w4(32'h3cc6257b),
	.w5(32'h3cdafa4d),
	.w6(32'hbd05c353),
	.w7(32'h3c525b7a),
	.w8(32'h3d1d8eb1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5763d),
	.w1(32'h3cf9ad3d),
	.w2(32'h3d09ee68),
	.w3(32'hbb186a6e),
	.w4(32'h3cc1a1d9),
	.w5(32'hbc7c6c53),
	.w6(32'h3bd7422d),
	.w7(32'h3d162d12),
	.w8(32'h3b9faded),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f62c1),
	.w1(32'h3c8be8c0),
	.w2(32'hbb0cdfad),
	.w3(32'hbcd5cd3f),
	.w4(32'h3b22b0fd),
	.w5(32'h3b0e0e49),
	.w6(32'hbd1aedde),
	.w7(32'hbd3119d7),
	.w8(32'hbce11842),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb00d07),
	.w1(32'h3ca69d47),
	.w2(32'h3c334d99),
	.w3(32'hbb748264),
	.w4(32'h3c241686),
	.w5(32'h3cef6b94),
	.w6(32'hb9c2f6e8),
	.w7(32'hbac9fb1c),
	.w8(32'h3cd1796d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6db3cf),
	.w1(32'h3b64d732),
	.w2(32'h3bb365b9),
	.w3(32'h3b360c77),
	.w4(32'h3af5df63),
	.w5(32'hbb4e9470),
	.w6(32'h3b2d60dc),
	.w7(32'h3b8f87d5),
	.w8(32'h3c4dd023),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c1772),
	.w1(32'hbb9c9339),
	.w2(32'h3a7b0918),
	.w3(32'hbafc4309),
	.w4(32'hbbb48973),
	.w5(32'hbc264501),
	.w6(32'hb99f8bc3),
	.w7(32'h3a77a20a),
	.w8(32'hbc125fab),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a05b),
	.w1(32'h39a2498a),
	.w2(32'h39d48f25),
	.w3(32'h3b4e28da),
	.w4(32'h39b7bb10),
	.w5(32'hb99b1d2b),
	.w6(32'h3aa893ae),
	.w7(32'hba830c30),
	.w8(32'hba4182cd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc4e97),
	.w1(32'h3c925840),
	.w2(32'h3c0dec93),
	.w3(32'hbc8110bc),
	.w4(32'hbb989bbb),
	.w5(32'h3cc7e174),
	.w6(32'hb9e619bb),
	.w7(32'hbc74c877),
	.w8(32'hbc44b838),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47476a),
	.w1(32'hbcf09290),
	.w2(32'hbcc2f264),
	.w3(32'hbcb25c7c),
	.w4(32'h3c5357c5),
	.w5(32'h3c5ad84f),
	.w6(32'hbd0d2090),
	.w7(32'h3b62fd24),
	.w8(32'h3d2391ba),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb59c6b),
	.w1(32'hbc25f985),
	.w2(32'hbc61856f),
	.w3(32'hbcfeb447),
	.w4(32'hbcf10536),
	.w5(32'hbc61ae22),
	.w6(32'hbcee7acb),
	.w7(32'hbd15c61f),
	.w8(32'hbc71593d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b21f),
	.w1(32'h3d168422),
	.w2(32'h3ccfce6d),
	.w3(32'h3c439697),
	.w4(32'hbc89ade8),
	.w5(32'hbb866350),
	.w6(32'h3d1a2c4a),
	.w7(32'h3c0d316f),
	.w8(32'hbcd9a3b9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e8c6),
	.w1(32'h3ca0d0e0),
	.w2(32'hbcc16f8b),
	.w3(32'hbc8d35f2),
	.w4(32'hbc947c04),
	.w5(32'h3cd183b7),
	.w6(32'hbc003de3),
	.w7(32'hbd415259),
	.w8(32'hbb8225ee),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc976d4),
	.w1(32'h3ba9f914),
	.w2(32'hbae1d1b0),
	.w3(32'hba1f85d6),
	.w4(32'h3a4ccb17),
	.w5(32'h3bfa7acb),
	.w6(32'hbb48e171),
	.w7(32'hbbc28d60),
	.w8(32'h3b93378d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dc6e4),
	.w1(32'hbc21e280),
	.w2(32'h3cb6c008),
	.w3(32'h3beb058a),
	.w4(32'h3bad8f3e),
	.w5(32'hbb4b73df),
	.w6(32'h3bafad85),
	.w7(32'h3cabbad2),
	.w8(32'h3c0bb637),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe8017),
	.w1(32'h3b4f8272),
	.w2(32'hbbbc766a),
	.w3(32'hbb146df3),
	.w4(32'h3ac1dd13),
	.w5(32'h3c027d7c),
	.w6(32'hbbdc1a71),
	.w7(32'hbbc2ea0c),
	.w8(32'h3c16aa42),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fab905),
	.w1(32'hba812905),
	.w2(32'hbb4e9bca),
	.w3(32'hbb58af15),
	.w4(32'hbb5f4654),
	.w5(32'hbb1619e9),
	.w6(32'hbb6186c3),
	.w7(32'hbb96146c),
	.w8(32'hbb8aedc2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb638263),
	.w1(32'hbb9c4a11),
	.w2(32'h3b30d88a),
	.w3(32'h3b7defa5),
	.w4(32'h3bdcd831),
	.w5(32'h3b1cbe52),
	.w6(32'hbabe7c3a),
	.w7(32'hbc0f4329),
	.w8(32'hb919dcef),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa006af),
	.w1(32'h3d2de5df),
	.w2(32'h3d2ef06b),
	.w3(32'hbc8a0a0f),
	.w4(32'hbcc1e7b2),
	.w5(32'hbc8e6b66),
	.w6(32'h3c892e80),
	.w7(32'hbb69c517),
	.w8(32'hbd40cf9f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48c835),
	.w1(32'hbcc8199d),
	.w2(32'hbd74eecd),
	.w3(32'hbca738d0),
	.w4(32'hbbad9830),
	.w5(32'h3cd64f18),
	.w6(32'hbd336c0d),
	.w7(32'hbd699ac8),
	.w8(32'h3bebc5dd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2b080),
	.w1(32'h3b643bc5),
	.w2(32'h3c093d63),
	.w3(32'h3b987baf),
	.w4(32'h3bf2d983),
	.w5(32'h3b6bd1e5),
	.w6(32'h3bbd6dbc),
	.w7(32'h3c303ccf),
	.w8(32'h3b9804f7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878b7e),
	.w1(32'h3bf47a83),
	.w2(32'h3bb48917),
	.w3(32'h3bd49ffa),
	.w4(32'h3c159834),
	.w5(32'h3c997f3f),
	.w6(32'h3bd0685e),
	.w7(32'h3b821fb7),
	.w8(32'h3c992be3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c531134),
	.w1(32'h3c074ef0),
	.w2(32'h3bc59103),
	.w3(32'h3bcc88de),
	.w4(32'h3a687ac0),
	.w5(32'hbb3da2a9),
	.w6(32'h3befe190),
	.w7(32'h3ba5d56b),
	.w8(32'h3bf63dea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1964a),
	.w1(32'h3c28cf6d),
	.w2(32'h3c3302e6),
	.w3(32'h3b9b0898),
	.w4(32'h3b4b64e0),
	.w5(32'h3b3d03bb),
	.w6(32'h3bba1679),
	.w7(32'h3b3007bb),
	.w8(32'h39e8cc30),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b16ab),
	.w1(32'hbc4d93c1),
	.w2(32'hbc0829c5),
	.w3(32'hbc7d4cf4),
	.w4(32'hbcdfd59d),
	.w5(32'hbc886f4a),
	.w6(32'hbb850381),
	.w7(32'hbd05d423),
	.w8(32'hbcac4f9a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94b4c2),
	.w1(32'hbc1cdc42),
	.w2(32'h3ba72bee),
	.w3(32'hbb82dbc3),
	.w4(32'hba8afcc0),
	.w5(32'hba54be2f),
	.w6(32'h3c00415b),
	.w7(32'h3c1c0839),
	.w8(32'hbbbf0850),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf0279),
	.w1(32'h3b89eb04),
	.w2(32'hbc4d02b8),
	.w3(32'hbcd55489),
	.w4(32'hbcee1129),
	.w5(32'h3c3a0794),
	.w6(32'hbbe95465),
	.w7(32'hbd46e87c),
	.w8(32'hbc4237ff),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbc956),
	.w1(32'hbb9ecb3a),
	.w2(32'hbbc038e2),
	.w3(32'hbc0a823c),
	.w4(32'hbbd8978f),
	.w5(32'hbba6d044),
	.w6(32'hbc2ca1cf),
	.w7(32'hbc0a8449),
	.w8(32'hbbd511e8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004d6b),
	.w1(32'hbc88d50d),
	.w2(32'h3bed586d),
	.w3(32'hbc06b092),
	.w4(32'h3c194663),
	.w5(32'h3adff617),
	.w6(32'hbc636c52),
	.w7(32'h3c27e245),
	.w8(32'h3c9bcb24),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdb8a5),
	.w1(32'h3b859019),
	.w2(32'h3c4262aa),
	.w3(32'hbad69526),
	.w4(32'h3b7adc67),
	.w5(32'h3a8f9e89),
	.w6(32'hbb83ed70),
	.w7(32'h3b891a6b),
	.w8(32'hbbe08fe6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc995ba),
	.w1(32'hb9e5bf55),
	.w2(32'h3c5d3d21),
	.w3(32'h3c20f7bf),
	.w4(32'h3c2c21c2),
	.w5(32'h3bcb1db5),
	.w6(32'h3bda7b6e),
	.w7(32'h3c326c36),
	.w8(32'h3bf74583),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c153dce),
	.w1(32'h3a9416fe),
	.w2(32'h3cbd9986),
	.w3(32'hbbe84ca1),
	.w4(32'h3ae1de76),
	.w5(32'h3b6b4b87),
	.w6(32'hbbdfab90),
	.w7(32'h3bce0b6d),
	.w8(32'h3ba9a418),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be21564),
	.w1(32'hbc53b72a),
	.w2(32'h3a563b3e),
	.w3(32'hbc245c67),
	.w4(32'hbc7dd27d),
	.w5(32'hbce96c97),
	.w6(32'hbc2fb111),
	.w7(32'hbba7f325),
	.w8(32'hbca94a26),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b058ce1),
	.w1(32'h3b481326),
	.w2(32'h3c4bd76a),
	.w3(32'h3b00ab2f),
	.w4(32'h3b8f19ef),
	.w5(32'h3a9ba5a8),
	.w6(32'h3bd67536),
	.w7(32'h3c40d70a),
	.w8(32'hbb8531ed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302b58),
	.w1(32'hbc3d714e),
	.w2(32'h3a2d9309),
	.w3(32'hbbc69f77),
	.w4(32'hbc2bad08),
	.w5(32'h3b87a354),
	.w6(32'hbbba68e9),
	.w7(32'hbc8679bc),
	.w8(32'hbc755a76),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad103),
	.w1(32'hba98104e),
	.w2(32'h3b4db84b),
	.w3(32'h3997ba50),
	.w4(32'hbb23be35),
	.w5(32'hbb8f44ac),
	.w6(32'h3a4961d1),
	.w7(32'h3b5cc6ee),
	.w8(32'hbbf17c0f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b847852),
	.w1(32'h3b9515f2),
	.w2(32'hbc8064e9),
	.w3(32'hbb2de3dc),
	.w4(32'hbb2205b5),
	.w5(32'hbb860b5e),
	.w6(32'hbc96834b),
	.w7(32'hbb4c64ca),
	.w8(32'hbaf8b821),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b3425),
	.w1(32'hbb9ff77a),
	.w2(32'hbbde5bd0),
	.w3(32'hbbd560c1),
	.w4(32'hbbaf020c),
	.w5(32'hbbb63152),
	.w6(32'hbc048359),
	.w7(32'hbc03009c),
	.w8(32'hbb9dc2cd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40d045),
	.w1(32'h3aede561),
	.w2(32'h3b6ca1e8),
	.w3(32'h3a33f176),
	.w4(32'h3b91bf18),
	.w5(32'h3bab2ba1),
	.w6(32'hbc89e943),
	.w7(32'h3ba73ab1),
	.w8(32'hba678721),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e728f),
	.w1(32'hbc338c0b),
	.w2(32'hbb788aab),
	.w3(32'hbc8fde98),
	.w4(32'hbbc48722),
	.w5(32'hbb7e4400),
	.w6(32'hbc80c547),
	.w7(32'hbbf2d56e),
	.w8(32'hbb3eadd2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47fd0f),
	.w1(32'hbbb61189),
	.w2(32'hbc006b23),
	.w3(32'hbc820861),
	.w4(32'hbd09f56b),
	.w5(32'h3bc0cf62),
	.w6(32'hbcbf7937),
	.w7(32'hbcdf4b83),
	.w8(32'hbd1efa40),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf29b69),
	.w1(32'hbcbcfc58),
	.w2(32'hbc623b61),
	.w3(32'hbcaa93d0),
	.w4(32'hbc841add),
	.w5(32'h38f806dd),
	.w6(32'hbd1ec972),
	.w7(32'hbca1085f),
	.w8(32'hbc696a4f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bc53e),
	.w1(32'h3bdc5655),
	.w2(32'h3bddeaca),
	.w3(32'hb9e82704),
	.w4(32'h38b7fb34),
	.w5(32'h3a970b50),
	.w6(32'h3a7ddcef),
	.w7(32'h3ac33401),
	.w8(32'h3c3c2d84),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule