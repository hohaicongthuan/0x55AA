module layer_10_featuremap_4(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc375e4),
	.w1(32'hbbc261ed),
	.w2(32'h3b80c824),
	.w3(32'h3c132e4a),
	.w4(32'h3b5fa7ae),
	.w5(32'hbb627e92),
	.w6(32'h3ba60fdc),
	.w7(32'h39f92993),
	.w8(32'hbc8fc78f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178792),
	.w1(32'h3a89757e),
	.w2(32'hbc637071),
	.w3(32'hbc38f2ab),
	.w4(32'h3c30e0cb),
	.w5(32'h3b76b563),
	.w6(32'hbcb34bbc),
	.w7(32'hbb6ea20d),
	.w8(32'hba10ed81),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d40d9),
	.w1(32'hbc298db2),
	.w2(32'h3c567337),
	.w3(32'h3b5ff860),
	.w4(32'hbb112306),
	.w5(32'h3c663d21),
	.w6(32'h3b5804a6),
	.w7(32'h3b815807),
	.w8(32'h3c228778),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c15c1),
	.w1(32'h3c328162),
	.w2(32'h3c16f286),
	.w3(32'h3c760241),
	.w4(32'h3c64a65f),
	.w5(32'hbb920268),
	.w6(32'h3c8d01ca),
	.w7(32'h3cb1dfaa),
	.w8(32'h3bc65c72),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbcd26),
	.w1(32'h3a4935e0),
	.w2(32'hbc4fecee),
	.w3(32'hbb7559a2),
	.w4(32'hbc1926e3),
	.w5(32'hbcd98887),
	.w6(32'h3b3dacda),
	.w7(32'h3a6c942a),
	.w8(32'hbbaaaaf0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4da4b),
	.w1(32'h3adf80b2),
	.w2(32'hbb96c581),
	.w3(32'hb9c63499),
	.w4(32'h3c0c341c),
	.w5(32'hbb1f89a0),
	.w6(32'h3bd9863e),
	.w7(32'h3c256102),
	.w8(32'hba4c4d44),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd35b46),
	.w1(32'h3bc80078),
	.w2(32'hbcb3e6ff),
	.w3(32'h3c0d176e),
	.w4(32'hbc0a0e03),
	.w5(32'hbc6c3c6f),
	.w6(32'hbb983f73),
	.w7(32'hbbe35114),
	.w8(32'hbceabf6d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd723acf),
	.w1(32'hbd70cc35),
	.w2(32'hbd288fe5),
	.w3(32'hbd0e257c),
	.w4(32'hbd372b92),
	.w5(32'hbd143476),
	.w6(32'hbd392366),
	.w7(32'hbd87ae8b),
	.w8(32'hbc3d102a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aea45),
	.w1(32'h3b5e540c),
	.w2(32'hbc815840),
	.w3(32'h3c051fc8),
	.w4(32'hbbb5c287),
	.w5(32'hbc2c27c6),
	.w6(32'h3bbf8010),
	.w7(32'hbb9b5864),
	.w8(32'hbc395328),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5a2e3),
	.w1(32'hbb0929ec),
	.w2(32'hbca75a91),
	.w3(32'h3c612063),
	.w4(32'hbb83d6e5),
	.w5(32'hbc483a62),
	.w6(32'hbc88731e),
	.w7(32'hbcade630),
	.w8(32'hbd12c692),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab843c3),
	.w1(32'h38a863e5),
	.w2(32'h3c174f0b),
	.w3(32'h3ad6b4d9),
	.w4(32'h3b1ff063),
	.w5(32'h3c42c100),
	.w6(32'h3b45e3cb),
	.w7(32'h3a59a713),
	.w8(32'h3c3a363a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfcd777),
	.w1(32'h3d04b80a),
	.w2(32'hbc4adbff),
	.w3(32'h3c941419),
	.w4(32'h3c9248dd),
	.w5(32'hbc2363b5),
	.w6(32'h3c4018a3),
	.w7(32'h3c88390c),
	.w8(32'hbca8945e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08813b),
	.w1(32'h3be39e1b),
	.w2(32'hbcc4d8a7),
	.w3(32'h3ce70f41),
	.w4(32'h3b49c715),
	.w5(32'hbc929cab),
	.w6(32'hbbfac13a),
	.w7(32'hbc5e5dc0),
	.w8(32'hbd0d80f0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68aaef),
	.w1(32'hb9fe66bb),
	.w2(32'hbcb1758a),
	.w3(32'h3c80b981),
	.w4(32'h3b3abacd),
	.w5(32'hbc9dae78),
	.w6(32'h3c0079ee),
	.w7(32'hbb87c814),
	.w8(32'hbc3bc84d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059db9),
	.w1(32'h3b579572),
	.w2(32'hbbbfea6c),
	.w3(32'hbb505aac),
	.w4(32'h3a409350),
	.w5(32'h3bddbbe3),
	.w6(32'hbb7878ad),
	.w7(32'hbbba8ed9),
	.w8(32'hbb875f38),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd002f6),
	.w1(32'hbcb6435d),
	.w2(32'hbc733efd),
	.w3(32'h3b3ba9a2),
	.w4(32'h3ad73638),
	.w5(32'h3bd59a18),
	.w6(32'hbc99f750),
	.w7(32'hbc803327),
	.w8(32'hbcc46ffd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c8543),
	.w1(32'h3a7effba),
	.w2(32'h3b29b6ad),
	.w3(32'h3b12bd28),
	.w4(32'h3aeb6d51),
	.w5(32'h3bf68191),
	.w6(32'h3b8caf3b),
	.w7(32'h3b21aaed),
	.w8(32'h38af378f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc842d36),
	.w1(32'hbbd7e2f8),
	.w2(32'hbd0efdcb),
	.w3(32'hbb9ebbab),
	.w4(32'hbc5479fb),
	.w5(32'hbce6103b),
	.w6(32'hbd181720),
	.w7(32'hbc974970),
	.w8(32'hbd1a4a74),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ebc20),
	.w1(32'hbab32fe3),
	.w2(32'hbc7e597d),
	.w3(32'h3c3618c8),
	.w4(32'hba8bb202),
	.w5(32'hbc6feaa1),
	.w6(32'hbbf31fa9),
	.w7(32'hbc499328),
	.w8(32'hbca59acb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01462f),
	.w1(32'h3b0832e4),
	.w2(32'h3ae1a6c8),
	.w3(32'hbb9954db),
	.w4(32'hbbd6a767),
	.w5(32'h3aa9f8fb),
	.w6(32'h3b61c491),
	.w7(32'hbae4728b),
	.w8(32'h3baf3617),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918a205),
	.w1(32'h3a5dd75c),
	.w2(32'hbbcd0171),
	.w3(32'h3b92eae7),
	.w4(32'h3acbdb69),
	.w5(32'hbc2b8ea8),
	.w6(32'h3bc191b3),
	.w7(32'h3b9610c6),
	.w8(32'hbb64043c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812c2d),
	.w1(32'h3c4aace9),
	.w2(32'hbc3001e4),
	.w3(32'hbc9d5ee2),
	.w4(32'hbc6a3832),
	.w5(32'hbbdf588c),
	.w6(32'hbb796a11),
	.w7(32'hbc67c0b4),
	.w8(32'h39ee588e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1a41a),
	.w1(32'hbd217874),
	.w2(32'hbd1bef1c),
	.w3(32'h3c7129a1),
	.w4(32'h398ca0fd),
	.w5(32'hbc924de1),
	.w6(32'hbd91b776),
	.w7(32'hbd389a92),
	.w8(32'hbd95ce7a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e78a8),
	.w1(32'h3c1cb3bb),
	.w2(32'hbc1e46a8),
	.w3(32'h3c98c51e),
	.w4(32'h3c58726d),
	.w5(32'hbb9e2d05),
	.w6(32'hbbefd189),
	.w7(32'hbc44608a),
	.w8(32'hbcd393bc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3a5ff),
	.w1(32'h3c112d61),
	.w2(32'hba783032),
	.w3(32'h3cdc0346),
	.w4(32'h3c6f7208),
	.w5(32'h3c471da2),
	.w6(32'h3ca07a58),
	.w7(32'hbc6cee37),
	.w8(32'hbcd159b9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc104ce),
	.w1(32'hbbfca82e),
	.w2(32'h3c140dfe),
	.w3(32'h3c204e74),
	.w4(32'h3ab69927),
	.w5(32'h3afbba92),
	.w6(32'hba3412db),
	.w7(32'h39c7309a),
	.w8(32'h3c2a9472),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb661bf),
	.w1(32'h3b7342c0),
	.w2(32'h3b4e495f),
	.w3(32'h3ba1108a),
	.w4(32'hbac5bfe5),
	.w5(32'h3bf7f918),
	.w6(32'hba9ba530),
	.w7(32'hbb6a1d58),
	.w8(32'h3b221756),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e3ba317),
	.w1(32'hbd0a9196),
	.w2(32'hbd1ed7cd),
	.w3(32'h3e17bfe3),
	.w4(32'hbd7b0208),
	.w5(32'hbd422a29),
	.w6(32'h3e221947),
	.w7(32'hbd520fff),
	.w8(32'hbcbe99b8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4d51),
	.w1(32'h3b7bc9f1),
	.w2(32'hbc4d6036),
	.w3(32'h3cc108f2),
	.w4(32'h3c69d02c),
	.w5(32'hbbeae074),
	.w6(32'h3cbbe7f5),
	.w7(32'h3c58ff61),
	.w8(32'hbb3edbcb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e1871fd),
	.w1(32'h3b329602),
	.w2(32'hbc6d4a57),
	.w3(32'h3dd286d9),
	.w4(32'hbca85a6e),
	.w5(32'hbcf84688),
	.w6(32'h3db2ac81),
	.w7(32'hbcb37d77),
	.w8(32'hbd069e9a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993e5ec),
	.w1(32'hbb0d1e42),
	.w2(32'hbba69e01),
	.w3(32'h3b569235),
	.w4(32'h3b1e0597),
	.w5(32'hbc59dadc),
	.w6(32'hba78eece),
	.w7(32'hbace7d05),
	.w8(32'hbc735ffb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60b9d0),
	.w1(32'h3b869200),
	.w2(32'hbc108056),
	.w3(32'hbc3d3a79),
	.w4(32'hbb7b1a27),
	.w5(32'hbcc43b8c),
	.w6(32'hbc42d80e),
	.w7(32'hbbcc5578),
	.w8(32'hbc4d589f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b56e1),
	.w1(32'h3a68a64b),
	.w2(32'hbc7203c6),
	.w3(32'hbc7c5908),
	.w4(32'hbb94dd6a),
	.w5(32'hbb6d9a55),
	.w6(32'hbcfc45ec),
	.w7(32'hbcf62ca4),
	.w8(32'hbc9a638b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff63b6),
	.w1(32'hbbdd850b),
	.w2(32'h3b3c23ca),
	.w3(32'h3b50881e),
	.w4(32'h3ae77fa3),
	.w5(32'hbab7eb71),
	.w6(32'hbb5930ca),
	.w7(32'hbc1d417d),
	.w8(32'hbc89af2a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a519d),
	.w1(32'hbbc0bd6d),
	.w2(32'h38de8edc),
	.w3(32'hbc3ded76),
	.w4(32'h3b8a3f78),
	.w5(32'hba4ab9f4),
	.w6(32'hbc674c24),
	.w7(32'hbaadce89),
	.w8(32'hbb2ece53),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb495a1),
	.w1(32'hbc17201f),
	.w2(32'hbbe5d5fc),
	.w3(32'hbadd9c49),
	.w4(32'hbbec14ea),
	.w5(32'hbc8787de),
	.w6(32'hbc403036),
	.w7(32'hbbb45b8c),
	.w8(32'hbc27e083),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd82879f),
	.w1(32'h3c795be5),
	.w2(32'hbd4d7497),
	.w3(32'hbbd56904),
	.w4(32'h3d04ce79),
	.w5(32'h3b6ae493),
	.w6(32'hbd5c5660),
	.w7(32'h3d316f4d),
	.w8(32'hbc8141bd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9ba6fe),
	.w1(32'h3bc69292),
	.w2(32'hbd34d95b),
	.w3(32'h3d8ff2a5),
	.w4(32'h3cd3c2d5),
	.w5(32'hbd19c75b),
	.w6(32'h3d8dea6d),
	.w7(32'hbb393e0d),
	.w8(32'hbd36c047),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e221dfa),
	.w1(32'h3c8580aa),
	.w2(32'hbd3f67a6),
	.w3(32'h3de30b02),
	.w4(32'hbca8dc2b),
	.w5(32'hbd7041be),
	.w6(32'h3dfa5279),
	.w7(32'hbb1aeffc),
	.w8(32'hbd791b75),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92a572),
	.w1(32'hbc108c10),
	.w2(32'h3bdcaddd),
	.w3(32'hbc96079d),
	.w4(32'hbba55255),
	.w5(32'h3bbbd187),
	.w6(32'hbc6599c7),
	.w7(32'hbc3046e5),
	.w8(32'h3a5c3313),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e13a),
	.w1(32'hbada6078),
	.w2(32'hbbc5da62),
	.w3(32'h3ba3d046),
	.w4(32'hbb8a9b74),
	.w5(32'hbc50f830),
	.w6(32'h3bec8eab),
	.w7(32'hbb2736c2),
	.w8(32'hbc3c601f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cb8a5),
	.w1(32'h3c10371f),
	.w2(32'hbc2831b2),
	.w3(32'hbcb8bc59),
	.w4(32'hbbb766ef),
	.w5(32'h3a10fc34),
	.w6(32'hbccc45c1),
	.w7(32'hbc83c12e),
	.w8(32'h3c08a6ae),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c606c93),
	.w1(32'h3c31f166),
	.w2(32'hbc4c9039),
	.w3(32'h3bbfe69c),
	.w4(32'h3c212d29),
	.w5(32'hbc32e06f),
	.w6(32'h3c0c420e),
	.w7(32'h3b690fcc),
	.w8(32'hbb3f3fa4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f4a4a),
	.w1(32'hbcf71061),
	.w2(32'hbd0acdcf),
	.w3(32'h3c1460ab),
	.w4(32'hbc8639eb),
	.w5(32'hbd3b7634),
	.w6(32'hbc751e84),
	.w7(32'hbcddf711),
	.w8(32'hbd91c8b2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75d411),
	.w1(32'hbbb9f754),
	.w2(32'hbcc13c13),
	.w3(32'h3c8cff59),
	.w4(32'h3c7539e0),
	.w5(32'hbcc36e1c),
	.w6(32'h3bdc8b3c),
	.w7(32'hbbfa2b86),
	.w8(32'hbd337639),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e385f),
	.w1(32'hbbf13715),
	.w2(32'hbc710eb5),
	.w3(32'h3bddeb07),
	.w4(32'hbc811dc8),
	.w5(32'h3b8880e4),
	.w6(32'hbd112c18),
	.w7(32'hbd2160d0),
	.w8(32'hbc8f6b95),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2eed),
	.w1(32'h3b589d8a),
	.w2(32'hbc867b87),
	.w3(32'hbb5139ed),
	.w4(32'h3bf419f0),
	.w5(32'hbbb012e3),
	.w6(32'hbc26cfd3),
	.w7(32'hbcabf093),
	.w8(32'hbca3b376),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31df9d),
	.w1(32'h3a805554),
	.w2(32'hbd1eca63),
	.w3(32'h3c198c53),
	.w4(32'h3b17f964),
	.w5(32'hbd479057),
	.w6(32'hbce4500b),
	.w7(32'hbcca66a8),
	.w8(32'hbd5ae1f0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f703),
	.w1(32'h3bb6dfb9),
	.w2(32'h3b64fd95),
	.w3(32'hbb1045d2),
	.w4(32'h3bd09cce),
	.w5(32'h3b60e6c6),
	.w6(32'h3b025fd1),
	.w7(32'h3c1d056a),
	.w8(32'h3bc8e2d3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0f23a),
	.w1(32'hbb5b0650),
	.w2(32'h3c0a14d6),
	.w3(32'h3c158697),
	.w4(32'hbb77c58f),
	.w5(32'h3c12fb76),
	.w6(32'h3c1287db),
	.w7(32'hbbdf51e1),
	.w8(32'h3ad54676),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c767ef3),
	.w1(32'hba87c186),
	.w2(32'hbbd4f409),
	.w3(32'h3c8557f3),
	.w4(32'h3c1073cc),
	.w5(32'hbc482d08),
	.w6(32'h3bae1cca),
	.w7(32'h3c3aff6b),
	.w8(32'hbba29fc1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab20816),
	.w1(32'hbc9be64e),
	.w2(32'hbba651ce),
	.w3(32'hbc44307f),
	.w4(32'hbc45445b),
	.w5(32'hbad9eadb),
	.w6(32'hbcae650b),
	.w7(32'hbc8f36d5),
	.w8(32'hbce91a8b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b003453),
	.w1(32'hba4470df),
	.w2(32'hbbc1d10f),
	.w3(32'h3c510b0a),
	.w4(32'h3b54c438),
	.w5(32'hbb1e064f),
	.w6(32'h3b7c9c24),
	.w7(32'hbadef2e8),
	.w8(32'hbbbe6d46),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18496d),
	.w1(32'hbbcad4ac),
	.w2(32'hbc98c043),
	.w3(32'hbbbf8e1c),
	.w4(32'hbbe5b148),
	.w5(32'hbcdf80e6),
	.w6(32'hbd032e84),
	.w7(32'hbcfa7f1e),
	.w8(32'hbd56d96e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c50f7),
	.w1(32'hbcbb2242),
	.w2(32'hbbb051ef),
	.w3(32'h3c71a9eb),
	.w4(32'hbc8d2ecf),
	.w5(32'hbcf03850),
	.w6(32'hbae9d67b),
	.w7(32'hbb491b02),
	.w8(32'hbcb47ca4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb34872),
	.w1(32'hbbaf4965),
	.w2(32'hbcc18250),
	.w3(32'hbc9e6660),
	.w4(32'hbb84e270),
	.w5(32'hbc7000fb),
	.w6(32'hbc0b99a5),
	.w7(32'hbc1633a0),
	.w8(32'hbc444c77),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81b64b),
	.w1(32'hbc46f95c),
	.w2(32'h3bb43bbb),
	.w3(32'hbc828344),
	.w4(32'hbcacd7aa),
	.w5(32'h3c29dbc2),
	.w6(32'hbca35121),
	.w7(32'hbc7ee30c),
	.w8(32'h3bfa0f08),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1de2be),
	.w1(32'hbb902ca3),
	.w2(32'h3b5e1814),
	.w3(32'h3c5bef9d),
	.w4(32'hbac2e20f),
	.w5(32'hba305d0c),
	.w6(32'h3c4299f8),
	.w7(32'hbaf584d4),
	.w8(32'hbbb20363),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15805b),
	.w1(32'hbb4bcd40),
	.w2(32'hbbb1ba6e),
	.w3(32'h3b44f901),
	.w4(32'hbb336fab),
	.w5(32'h3a01b97c),
	.w6(32'h3b73e4fb),
	.w7(32'h3a402773),
	.w8(32'hbb254d48),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2603a8),
	.w1(32'hb98bbda5),
	.w2(32'hbbfaae5c),
	.w3(32'h3be4d340),
	.w4(32'h3b25ef70),
	.w5(32'hbc07ddef),
	.w6(32'h3ba0fe21),
	.w7(32'h3c0a7070),
	.w8(32'hbc27577f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2885),
	.w1(32'hbbe83176),
	.w2(32'hbc8bf8b5),
	.w3(32'h3c511aa3),
	.w4(32'h3b48a242),
	.w5(32'hbc9a87c4),
	.w6(32'hbc609da6),
	.w7(32'hbc0d06b8),
	.w8(32'hbc887ce3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61fdf7),
	.w1(32'hbc2605d1),
	.w2(32'hbc6f2803),
	.w3(32'h3c8aba5d),
	.w4(32'hbc4405d4),
	.w5(32'hbc963876),
	.w6(32'hba4de94d),
	.w7(32'hbc22937f),
	.w8(32'hbc6f9500),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9212),
	.w1(32'hbc17f291),
	.w2(32'hbb43fe47),
	.w3(32'hba6c5b09),
	.w4(32'hbc04928c),
	.w5(32'h3a16c951),
	.w6(32'hbb5d4e0e),
	.w7(32'hbbda8d4d),
	.w8(32'hbbacb842),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa9d5e),
	.w1(32'hbadf5fdc),
	.w2(32'hbc2a4d86),
	.w3(32'hbb4b1f63),
	.w4(32'hbb081190),
	.w5(32'hb7ba04c6),
	.w6(32'hbc120cbd),
	.w7(32'hbb750fa2),
	.w8(32'h3a746c39),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11d44b),
	.w1(32'hbbb95cf8),
	.w2(32'hbb18ab21),
	.w3(32'h3c3ba6b9),
	.w4(32'h3b059af9),
	.w5(32'hbb8a34bc),
	.w6(32'h3c5175ff),
	.w7(32'h3bd828f4),
	.w8(32'hbb0c72f9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a701686),
	.w1(32'hbad3c740),
	.w2(32'hbb3d6d14),
	.w3(32'hbb3749bf),
	.w4(32'hb9b419e0),
	.w5(32'hb9bf8360),
	.w6(32'hbaaa530b),
	.w7(32'hb91a2b9d),
	.w8(32'h3b11d3f7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257d75),
	.w1(32'hbb2fc1cf),
	.w2(32'hbc29194c),
	.w3(32'h3c61e41e),
	.w4(32'h3bc1d0bc),
	.w5(32'hbb95f382),
	.w6(32'hbbe76dad),
	.w7(32'hbca7cb6d),
	.w8(32'hbd2159a6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87e0d2),
	.w1(32'h3c298a82),
	.w2(32'hbab5ef23),
	.w3(32'h3c14179a),
	.w4(32'h3c96ff96),
	.w5(32'hbc10f94e),
	.w6(32'hbd3bd858),
	.w7(32'hbcfac660),
	.w8(32'hbd24c805),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc852ea2),
	.w1(32'hbcbdee47),
	.w2(32'hbcfe2329),
	.w3(32'hbc1e4f38),
	.w4(32'hbc941731),
	.w5(32'hbcf9dd32),
	.w6(32'hbd2b37c6),
	.w7(32'hbd1903ec),
	.w8(32'hbd3948e4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d803139),
	.w1(32'h3beb3d72),
	.w2(32'hbcccdeec),
	.w3(32'h3d046a78),
	.w4(32'hb848f742),
	.w5(32'h3a8385e7),
	.w6(32'h3c62c054),
	.w7(32'hbd2f17c4),
	.w8(32'hbd314023),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39ac70),
	.w1(32'h3c0684bd),
	.w2(32'h3b08f17d),
	.w3(32'h3c3da8d3),
	.w4(32'h3c3efd16),
	.w5(32'h3b135042),
	.w6(32'h3c35a060),
	.w7(32'h3c4542c1),
	.w8(32'h3af4f076),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff693),
	.w1(32'h3be46ffe),
	.w2(32'hbba072e4),
	.w3(32'h3b9cd7e1),
	.w4(32'h3c596d43),
	.w5(32'hba190cae),
	.w6(32'h3bb283e7),
	.w7(32'h3c46a712),
	.w8(32'h3bd17586),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58814c),
	.w1(32'h3a510192),
	.w2(32'h39b731ce),
	.w3(32'h3c8e3890),
	.w4(32'h3c810243),
	.w5(32'h3b2892a6),
	.w6(32'h3b285431),
	.w7(32'h3b8f9b08),
	.w8(32'h3c1b5a52),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd5bc6),
	.w1(32'hbb2fc852),
	.w2(32'hbc415ca2),
	.w3(32'h3be20ab5),
	.w4(32'hba540a5d),
	.w5(32'hbc2c95dc),
	.w6(32'h3b5a4e92),
	.w7(32'hbbb18475),
	.w8(32'hbc5edb1f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e82b1),
	.w1(32'hbb92ce6f),
	.w2(32'hbc10b20b),
	.w3(32'hbbab0001),
	.w4(32'hbb17b93e),
	.w5(32'h3afedb33),
	.w6(32'hbb11bb59),
	.w7(32'hba53a956),
	.w8(32'hba12dd82),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd9de5),
	.w1(32'hbcd8c7a7),
	.w2(32'hbbaa518c),
	.w3(32'h3993e4eb),
	.w4(32'hbcad8a4b),
	.w5(32'hbb8d01dd),
	.w6(32'hbb6eb439),
	.w7(32'hbcdf67e6),
	.w8(32'hbcab78b4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc195a40),
	.w1(32'hbc177f9c),
	.w2(32'hbc79efa4),
	.w3(32'h3c35a9f5),
	.w4(32'hbc0ad9d3),
	.w5(32'hbc9b1f15),
	.w6(32'hbc0bd818),
	.w7(32'hbb9c0646),
	.w8(32'hbcc68902),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c955edc),
	.w1(32'hbb59247d),
	.w2(32'hbc68637a),
	.w3(32'h3cc83f40),
	.w4(32'h3c1be9c3),
	.w5(32'hbac29969),
	.w6(32'h3c1b1d08),
	.w7(32'h3abfd7dd),
	.w8(32'hbc0fe6a2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a0e6d),
	.w1(32'h3b857700),
	.w2(32'hbc01469a),
	.w3(32'hbca37aa4),
	.w4(32'hbc2da147),
	.w5(32'hb9c9a5d9),
	.w6(32'hbccc7a18),
	.w7(32'hbcaa01a3),
	.w8(32'hbc44551d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb79240),
	.w1(32'h3bb6f3cf),
	.w2(32'hbb06f789),
	.w3(32'h3cad5af4),
	.w4(32'h3c56b172),
	.w5(32'h3c279fd4),
	.w6(32'hbb4bff96),
	.w7(32'hbc8b7f23),
	.w8(32'hbc469109),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9246c),
	.w1(32'hbc115814),
	.w2(32'hbc1a923a),
	.w3(32'h3abf505f),
	.w4(32'hbbf2a820),
	.w5(32'h39ffef79),
	.w6(32'h3bcddde6),
	.w7(32'hbbf2b5ac),
	.w8(32'hbc342684),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84b199),
	.w1(32'hbc2c1f0e),
	.w2(32'hbc67ae39),
	.w3(32'h3bfa33e0),
	.w4(32'hbc12cbfa),
	.w5(32'h3b60606e),
	.w6(32'hbc31f32e),
	.w7(32'hbc9f9745),
	.w8(32'hbc273450),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bb653),
	.w1(32'h3c057c51),
	.w2(32'hbb6edfce),
	.w3(32'h3c6fcf94),
	.w4(32'h3c795fd2),
	.w5(32'hbb8c1672),
	.w6(32'h3c4dc651),
	.w7(32'h3c9450af),
	.w8(32'hbafa03ed),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eb566),
	.w1(32'h3a8d662b),
	.w2(32'hba9ddf8e),
	.w3(32'h39ef6d3d),
	.w4(32'hb99ca82c),
	.w5(32'h3bd0ce15),
	.w6(32'hbbab1876),
	.w7(32'hbb43adab),
	.w8(32'h3c44ec52),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49633b),
	.w1(32'h3c3ebae9),
	.w2(32'hbb0ea04b),
	.w3(32'h3c6a58f4),
	.w4(32'h3c5a085e),
	.w5(32'h3bfd53c4),
	.w6(32'h3bd3d537),
	.w7(32'h3b7cd406),
	.w8(32'hbc39d593),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd153d6),
	.w1(32'hb9e83ef1),
	.w2(32'hb9ac2077),
	.w3(32'hbab6c22e),
	.w4(32'h3bc60dbe),
	.w5(32'hbb1b58e4),
	.w6(32'hbb9ac7ef),
	.w7(32'hb8a05750),
	.w8(32'hb9f8f6d4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28de57),
	.w1(32'h3b224f19),
	.w2(32'hbc127ab9),
	.w3(32'hbcba0059),
	.w4(32'h3bbe9c2b),
	.w5(32'hbb950393),
	.w6(32'hbcb132d9),
	.w7(32'hbc3a4e45),
	.w8(32'hbc7b0576),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad22166),
	.w1(32'h3bb5de62),
	.w2(32'h3bd66a70),
	.w3(32'hbb4a2d7d),
	.w4(32'h3a1e7a50),
	.w5(32'h3b0f3105),
	.w6(32'hbb787d26),
	.w7(32'h3b192637),
	.w8(32'hbba312cc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a717),
	.w1(32'hbc1c6044),
	.w2(32'h3c594adf),
	.w3(32'hbbab1252),
	.w4(32'h3bb4026f),
	.w5(32'h38aedc8b),
	.w6(32'hbca0edbc),
	.w7(32'hbc8384cc),
	.w8(32'hbc936331),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac08a8),
	.w1(32'hbc70fcbd),
	.w2(32'hbcfda186),
	.w3(32'hbcfc7503),
	.w4(32'hbc21034e),
	.w5(32'hbd012340),
	.w6(32'hbd6245fb),
	.w7(32'hbcbc838f),
	.w8(32'hbd504fb2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d87337e),
	.w1(32'h3bda3ecd),
	.w2(32'hbc4e490b),
	.w3(32'h3d77f408),
	.w4(32'hbb40f868),
	.w5(32'hbd0c7935),
	.w6(32'h3d81b7cf),
	.w7(32'h3b338e0c),
	.w8(32'hbd0aedb1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9232cb),
	.w1(32'h3ab0f12b),
	.w2(32'h3b604a2c),
	.w3(32'h3c696244),
	.w4(32'h3c652918),
	.w5(32'h3c1ed08c),
	.w6(32'hbd12925c),
	.w7(32'h3aa06912),
	.w8(32'hbcd03212),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8cb00),
	.w1(32'h3b2d6cc5),
	.w2(32'hbc35e607),
	.w3(32'h3c616d21),
	.w4(32'hbba75931),
	.w5(32'hbcee50d5),
	.w6(32'h3c12db82),
	.w7(32'hbba20f17),
	.w8(32'hbcc16438),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86252c),
	.w1(32'hbb15cfc3),
	.w2(32'hbcae2820),
	.w3(32'hbc255dfa),
	.w4(32'h3c44f434),
	.w5(32'h3ac081dd),
	.w6(32'hbd294a02),
	.w7(32'hbca00d83),
	.w8(32'hbcfc3d78),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc253fa8),
	.w1(32'hbc6f58ed),
	.w2(32'h3c2adda5),
	.w3(32'hbb87d5e9),
	.w4(32'hbc9c2792),
	.w5(32'h3ca90060),
	.w6(32'hbc4daf43),
	.w7(32'hbcd3f3f9),
	.w8(32'hbc8c735f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e663a),
	.w1(32'h3b20016b),
	.w2(32'hbc85f223),
	.w3(32'h3d8e0158),
	.w4(32'hba98d410),
	.w5(32'hbc90a72f),
	.w6(32'h3d7ea328),
	.w7(32'hbc93d457),
	.w8(32'hbcdb2fa1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79de92),
	.w1(32'hbc80b4b8),
	.w2(32'hbb8d302d),
	.w3(32'h3b7cb1d1),
	.w4(32'hbc8bd92e),
	.w5(32'h393cc0d8),
	.w6(32'h3b66d2e0),
	.w7(32'hbc47afa7),
	.w8(32'h3b12cfd8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86566c),
	.w1(32'hbb9fbb24),
	.w2(32'hbc583697),
	.w3(32'h3cc4b81b),
	.w4(32'hb9f87900),
	.w5(32'hbcabebf1),
	.w6(32'hbca4855c),
	.w7(32'hbcbd6277),
	.w8(32'hbd605e5d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4615eb),
	.w1(32'hbc0b699b),
	.w2(32'hbcc94f13),
	.w3(32'h3c314c96),
	.w4(32'hbc2cba7c),
	.w5(32'hbc5e9b8e),
	.w6(32'hbca1456a),
	.w7(32'hbd0e9adc),
	.w8(32'hbd33b218),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd13743b),
	.w1(32'hbac1a2aa),
	.w2(32'hbd508bc9),
	.w3(32'hbc8faa44),
	.w4(32'h3ba128cb),
	.w5(32'hbc77d1cb),
	.w6(32'hbdb441af),
	.w7(32'hbc341008),
	.w8(32'hbc95d01e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d25c895),
	.w1(32'hbb8223ef),
	.w2(32'hbd1bdb63),
	.w3(32'h3cc3ba99),
	.w4(32'hbbaf2142),
	.w5(32'hbca880c7),
	.w6(32'h3cdb86dc),
	.w7(32'hbbe2e386),
	.w8(32'hbcebbb61),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3a258),
	.w1(32'h3be453f6),
	.w2(32'hbc2bce09),
	.w3(32'h3cdc1d0c),
	.w4(32'h3bbed4c4),
	.w5(32'h3b81b8e9),
	.w6(32'h3aeb3353),
	.w7(32'hbc3d44b7),
	.w8(32'hbbe9a7b2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda4ade),
	.w1(32'h3c816d6c),
	.w2(32'hbcedb644),
	.w3(32'hbc2c4f3d),
	.w4(32'h3bfc5420),
	.w5(32'h3b240ac1),
	.w6(32'hbd1a21e5),
	.w7(32'h3c1eea86),
	.w8(32'hbcc6311e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c3073),
	.w1(32'h3b323125),
	.w2(32'hbc1b35f7),
	.w3(32'hba2951d3),
	.w4(32'h3b5b8e33),
	.w5(32'hb80b1c7c),
	.w6(32'hbbc2090a),
	.w7(32'h3a3f24cc),
	.w8(32'hbb8754f7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdbc5fed),
	.w1(32'hbbbfe51d),
	.w2(32'hbd537bad),
	.w3(32'hbd6338af),
	.w4(32'h3c680caf),
	.w5(32'hbce7f9ce),
	.w6(32'hbd920866),
	.w7(32'hbc4b034c),
	.w8(32'hbcd0fa95),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a5460),
	.w1(32'h3ca61ca6),
	.w2(32'hbc944b32),
	.w3(32'h3c5fc29c),
	.w4(32'h3c1b38ae),
	.w5(32'hbcaefef4),
	.w6(32'h3be35ae5),
	.w7(32'hbbf855a2),
	.w8(32'hbca127f5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc6002),
	.w1(32'h3c088172),
	.w2(32'hbbdd2b23),
	.w3(32'h3beb5f35),
	.w4(32'h3c35c093),
	.w5(32'h3b9c5f2a),
	.w6(32'h3c2f50ac),
	.w7(32'h3c1a9849),
	.w8(32'h3c173061),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fb16a),
	.w1(32'hbc34d601),
	.w2(32'hbbe07537),
	.w3(32'hbc7c61b4),
	.w4(32'hbc268ea8),
	.w5(32'h3b3efa6c),
	.w6(32'hbc8a23ff),
	.w7(32'hbc4336e6),
	.w8(32'hbb1518bd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8c0a0),
	.w1(32'h3bf451a0),
	.w2(32'hbc8a1dcd),
	.w3(32'h3cf274be),
	.w4(32'h3c6bc06e),
	.w5(32'hbcb9ead4),
	.w6(32'h3b218a33),
	.w7(32'hba87f3f9),
	.w8(32'hbce906bf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee3db9),
	.w1(32'h3c88d6cb),
	.w2(32'hbbeb83ba),
	.w3(32'h3c38b172),
	.w4(32'hbb1e68ec),
	.w5(32'h3bb04e67),
	.w6(32'h3b680649),
	.w7(32'hbc4db41b),
	.w8(32'h3ae7bdc4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d25f26e),
	.w1(32'h3a698780),
	.w2(32'hbcb7e047),
	.w3(32'h3d55f64e),
	.w4(32'h3c12782b),
	.w5(32'hbc41e07a),
	.w6(32'h3d7cb98f),
	.w7(32'h3bbaece4),
	.w8(32'hbc9177d1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0368c3),
	.w1(32'hba22d6c4),
	.w2(32'hbc1bd693),
	.w3(32'h3aeb530f),
	.w4(32'h3c477500),
	.w5(32'hbc58ae77),
	.w6(32'hbc094a36),
	.w7(32'hbadec1d7),
	.w8(32'hbca5c5a5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7004ea),
	.w1(32'h3c494948),
	.w2(32'hbb1ddcf2),
	.w3(32'hbc44fc99),
	.w4(32'hbbab07d1),
	.w5(32'hbc217086),
	.w6(32'hbd6124d5),
	.w7(32'hbcb700a0),
	.w8(32'hbc482a1b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1be856),
	.w1(32'hbb809a6e),
	.w2(32'hbcb1d0cd),
	.w3(32'hbc99b32f),
	.w4(32'h3ac9cf8f),
	.w5(32'hbbd6e539),
	.w6(32'hbd43d531),
	.w7(32'hbcf03ebb),
	.w8(32'hbccadb4b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a40d),
	.w1(32'hbc07e038),
	.w2(32'hba2aa8e0),
	.w3(32'hbc39e2a0),
	.w4(32'hbc948dbc),
	.w5(32'h3bb3a088),
	.w6(32'hbc8a8f3a),
	.w7(32'hbcc8be9e),
	.w8(32'hbbb30ac3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e02562),
	.w1(32'h3b8f760b),
	.w2(32'hbc1dbc75),
	.w3(32'h3bcae945),
	.w4(32'h3be941b9),
	.w5(32'hbb576436),
	.w6(32'h3b8f6a7d),
	.w7(32'h3ba0e85f),
	.w8(32'hbb0511cd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31b233),
	.w1(32'hbb3cafee),
	.w2(32'h3b16e32a),
	.w3(32'hbb402570),
	.w4(32'hbb8fd9b0),
	.w5(32'h3bb87366),
	.w6(32'hbb60f3a5),
	.w7(32'hbb9a084c),
	.w8(32'h3b349d82),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad90514),
	.w1(32'h3bac3b1e),
	.w2(32'hbc4b2b0d),
	.w3(32'hba03de58),
	.w4(32'h3b4f504b),
	.w5(32'hbc9e1428),
	.w6(32'hb8efa865),
	.w7(32'h39ed0891),
	.w8(32'hbbeabc71),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51be5e),
	.w1(32'hbc619f0d),
	.w2(32'hbb79a9e6),
	.w3(32'hbcac3233),
	.w4(32'hbc72a329),
	.w5(32'hbbdf6ebf),
	.w6(32'hbc2b6cf6),
	.w7(32'h3b077c98),
	.w8(32'hbb8cdd76),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c852613),
	.w1(32'hbb903007),
	.w2(32'hbbd07fd5),
	.w3(32'h3cabdb6e),
	.w4(32'hbac9fbe0),
	.w5(32'hbb07d6e3),
	.w6(32'h3c60cb4b),
	.w7(32'hbc53ba70),
	.w8(32'hbcbe58d6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222063),
	.w1(32'hbc1c4160),
	.w2(32'hba8bfdcc),
	.w3(32'h3b3d19d5),
	.w4(32'hbc021d97),
	.w5(32'hbb5cb0a7),
	.w6(32'h3baf483f),
	.w7(32'hbc2e93ac),
	.w8(32'hbaefe9d9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4431a6),
	.w1(32'h3b163e2e),
	.w2(32'hbc6312a1),
	.w3(32'h3acfd073),
	.w4(32'hbbf8d132),
	.w5(32'hbba2ca63),
	.w6(32'hbc2b3367),
	.w7(32'hbc1de837),
	.w8(32'hbc30a189),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d04208a),
	.w1(32'h3a5fa7c9),
	.w2(32'hbc49fa77),
	.w3(32'h3d251bfa),
	.w4(32'h3c13e8e1),
	.w5(32'hbc32d751),
	.w6(32'h3d19c953),
	.w7(32'hbb8dbb9f),
	.w8(32'hbcdbe27b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f87f),
	.w1(32'h3a78ef11),
	.w2(32'hbaaf08ec),
	.w3(32'hbc5b121f),
	.w4(32'hbb7b3645),
	.w5(32'h3990e5fb),
	.w6(32'hbbd13b55),
	.w7(32'h3b427d49),
	.w8(32'h396c4bc5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae41eb),
	.w1(32'hbac74dd1),
	.w2(32'hba8f51f4),
	.w3(32'h3afb3b93),
	.w4(32'h3b6bad7f),
	.w5(32'hbb334577),
	.w6(32'h3aa33de7),
	.w7(32'h3a7e2035),
	.w8(32'hbc6284a4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b21d),
	.w1(32'hbbd0dc9d),
	.w2(32'hbb89b5a4),
	.w3(32'hbc58ce03),
	.w4(32'hbad9cf86),
	.w5(32'hba36fafd),
	.w6(32'hbc070ec2),
	.w7(32'h3c86a63d),
	.w8(32'hbbbf78a9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5135c),
	.w1(32'h3bc716a0),
	.w2(32'h3b2bf18a),
	.w3(32'h3baf1e5d),
	.w4(32'h3c405005),
	.w5(32'hbb8a601b),
	.w6(32'hbb130c4a),
	.w7(32'h3b66aff8),
	.w8(32'hbbb3861a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8b631),
	.w1(32'hbc1cfc3e),
	.w2(32'hbb8c87cb),
	.w3(32'hbc40f66c),
	.w4(32'hbb78275a),
	.w5(32'hbbf9e18b),
	.w6(32'hbd1b116a),
	.w7(32'hbd01ba9e),
	.w8(32'hbcb81727),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07f23),
	.w1(32'hbc0dd029),
	.w2(32'hbcd91097),
	.w3(32'hbc67fe97),
	.w4(32'hbc4be607),
	.w5(32'hbbb0ef18),
	.w6(32'hbd04477a),
	.w7(32'hbcd14f40),
	.w8(32'hbceebc69),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd002231),
	.w1(32'hbb89a90d),
	.w2(32'h37b3f78d),
	.w3(32'hbc3a38b9),
	.w4(32'hbc66f6e7),
	.w5(32'hbbab97e7),
	.w6(32'hbc4ece70),
	.w7(32'hbc87e745),
	.w8(32'hbb218f18),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b6cdb),
	.w1(32'h3aae355c),
	.w2(32'hbc139a82),
	.w3(32'hbcc59fb8),
	.w4(32'h3b5e4044),
	.w5(32'hbb1704b2),
	.w6(32'hbcccb27f),
	.w7(32'h3b071b98),
	.w8(32'h3b1044d3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beebb2d),
	.w1(32'h3b609e53),
	.w2(32'hbbbc1720),
	.w3(32'h3ce6c84c),
	.w4(32'h3c7f9629),
	.w5(32'hbc5f3bbb),
	.w6(32'h3c78b1f3),
	.w7(32'h3b6712f4),
	.w8(32'hbc86cda7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ec043),
	.w1(32'hbc9799da),
	.w2(32'hbc1cdca9),
	.w3(32'hbc477863),
	.w4(32'hbb8550cc),
	.w5(32'hbb8c57f5),
	.w6(32'hbb4e6ef4),
	.w7(32'hbc4bcb8e),
	.w8(32'hbbfa221a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03e0dc),
	.w1(32'hbc4a2357),
	.w2(32'hbcb855d3),
	.w3(32'hbcbcf755),
	.w4(32'hbc64fc6f),
	.w5(32'hbc4d6d27),
	.w6(32'hbc8ad2ad),
	.w7(32'hbca9de9a),
	.w8(32'hbc9a7fbb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d9af6),
	.w1(32'hbc972254),
	.w2(32'hbce3a27d),
	.w3(32'h3b801e95),
	.w4(32'hbccc75d9),
	.w5(32'hbcd16ec6),
	.w6(32'hbcab9096),
	.w7(32'hbd15c398),
	.w8(32'hbd51a0c6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc96dee),
	.w1(32'h3c0e8025),
	.w2(32'hb9ef44b1),
	.w3(32'hbb0f128a),
	.w4(32'h3c8c70fc),
	.w5(32'h38de3da4),
	.w6(32'h3bbb301e),
	.w7(32'h3b7049b7),
	.w8(32'hbc28398a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9368746),
	.w1(32'hbb13f870),
	.w2(32'hbc4fe0e8),
	.w3(32'hbbe3ea66),
	.w4(32'h3bf9fb8b),
	.w5(32'hb98a8b90),
	.w6(32'hbd07053b),
	.w7(32'hbc5c696b),
	.w8(32'hbc61f4e2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacb9f4),
	.w1(32'hbcd554a9),
	.w2(32'hbc84cf47),
	.w3(32'hb9841554),
	.w4(32'hbca61c26),
	.w5(32'hbc4dd9fc),
	.w6(32'hbc8fc30f),
	.w7(32'hbcf3f57e),
	.w8(32'hbcd89459),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c109b),
	.w1(32'hbb28dbe0),
	.w2(32'h3b0f828e),
	.w3(32'hbc1e6b39),
	.w4(32'h3b893887),
	.w5(32'h3c909897),
	.w6(32'hbceab013),
	.w7(32'hbc89bbfe),
	.w8(32'hbb2391be),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96f979),
	.w1(32'hbb26e29f),
	.w2(32'hbc23fd1c),
	.w3(32'h3cc165c3),
	.w4(32'h3b75284e),
	.w5(32'hbbf87f02),
	.w6(32'h3b69d2db),
	.w7(32'hbc5bc4a2),
	.w8(32'hbc8f08ed),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9009904),
	.w1(32'hbaa6cf7e),
	.w2(32'h3b853407),
	.w3(32'h3a8ba9cb),
	.w4(32'h3ac2c182),
	.w5(32'h3c18529f),
	.w6(32'hbb3f53b7),
	.w7(32'hbabd9c40),
	.w8(32'hbb087653),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e0e943d),
	.w1(32'hbc3ae359),
	.w2(32'hbc4c22a2),
	.w3(32'h3ddb877f),
	.w4(32'hbcff922d),
	.w5(32'hbd74b734),
	.w6(32'h3ddfc4ba),
	.w7(32'hbd135b81),
	.w8(32'hbd79fb8a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68c7a),
	.w1(32'hbc03e507),
	.w2(32'hbc4ff26c),
	.w3(32'hbcb5b329),
	.w4(32'hbc89a6e8),
	.w5(32'hba9580a6),
	.w6(32'hbcdede71),
	.w7(32'hbc7e0ff9),
	.w8(32'hba6393ee),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d36cc),
	.w1(32'h3b529df6),
	.w2(32'hbada1282),
	.w3(32'h3aeb080b),
	.w4(32'h3b66b878),
	.w5(32'hb87d2977),
	.w6(32'h3a483441),
	.w7(32'h3a985e9c),
	.w8(32'h39f2609a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10cf6a),
	.w1(32'hbb034457),
	.w2(32'hbbfee5da),
	.w3(32'hb92e9a0c),
	.w4(32'hba672c73),
	.w5(32'hbbb17687),
	.w6(32'hb9c68388),
	.w7(32'hb8ae71eb),
	.w8(32'hbbfbd9e3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcf827),
	.w1(32'h3b8b3364),
	.w2(32'hbb2124dc),
	.w3(32'hba8de90d),
	.w4(32'h3bd179b2),
	.w5(32'hbba732a7),
	.w6(32'hbb94bb71),
	.w7(32'hbbdc9ae5),
	.w8(32'hbb786543),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167ba9),
	.w1(32'hbb7b1b9a),
	.w2(32'hbce7d430),
	.w3(32'hba431a9a),
	.w4(32'h3c3b3563),
	.w5(32'hbc86ec6d),
	.w6(32'hbb186374),
	.w7(32'h3b3d4bdf),
	.w8(32'hbc75f36b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7c1a5),
	.w1(32'h3c95781d),
	.w2(32'hbc0f1399),
	.w3(32'h3ad65ea9),
	.w4(32'h3a78f6c8),
	.w5(32'hbc3b8969),
	.w6(32'hbcc98bf5),
	.w7(32'hbd1d876b),
	.w8(32'hbcc8c218),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19cfeb),
	.w1(32'h3b2f0572),
	.w2(32'hbbbd7900),
	.w3(32'h3b1a3a5d),
	.w4(32'h3b6f4a02),
	.w5(32'h3bc7161b),
	.w6(32'h3afb3f93),
	.w7(32'h3a83c04a),
	.w8(32'h3c3eacd3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c0961),
	.w1(32'h3b760724),
	.w2(32'hbcd22048),
	.w3(32'h3d0d1bc7),
	.w4(32'h3b32c43b),
	.w5(32'hbca09d57),
	.w6(32'h3b14804c),
	.w7(32'hbcaf29af),
	.w8(32'hbd0ce0f5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce54d6),
	.w1(32'h3bde12fc),
	.w2(32'hbbc14108),
	.w3(32'h3bccee82),
	.w4(32'h3ba9ec60),
	.w5(32'h37d23ac6),
	.w6(32'hbb604f72),
	.w7(32'hbbf45bd1),
	.w8(32'hbc1ed1b6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cb0d4),
	.w1(32'hbbe324e7),
	.w2(32'hbbe6738f),
	.w3(32'hb9fdede1),
	.w4(32'hbbfec476),
	.w5(32'h3bb25707),
	.w6(32'hbc71fb34),
	.w7(32'hbc4817b0),
	.w8(32'hbc45a455),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dcbfbfd),
	.w1(32'hbce318be),
	.w2(32'hbd0a6674),
	.w3(32'h3dbea475),
	.w4(32'hbcc7aca8),
	.w5(32'hbcd154d0),
	.w6(32'h3dc82261),
	.w7(32'hbce11c7b),
	.w8(32'hbd0fde88),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3a04),
	.w1(32'h3bd3a7fe),
	.w2(32'h3b9991cd),
	.w3(32'hbc731718),
	.w4(32'hbbe49321),
	.w5(32'h3c013f9d),
	.w6(32'hbc4f1810),
	.w7(32'hbc8e1c9f),
	.w8(32'h3bc5c43a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b7832),
	.w1(32'h3b0da007),
	.w2(32'h3a9eebea),
	.w3(32'h3c83c371),
	.w4(32'h3c44359a),
	.w5(32'h390ed937),
	.w6(32'h3ca04922),
	.w7(32'h3c7ae82a),
	.w8(32'h3abdb292),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd76503),
	.w1(32'h3be95b32),
	.w2(32'h3b68c8eb),
	.w3(32'h3ca72ce8),
	.w4(32'h3b864954),
	.w5(32'h3b9e2265),
	.w6(32'h3c846a9b),
	.w7(32'hbb10091d),
	.w8(32'hbbb93ff2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70cc24),
	.w1(32'hbbe6704c),
	.w2(32'h39867578),
	.w3(32'h3be7d13b),
	.w4(32'hbb6d7cb1),
	.w5(32'hbb73dc6f),
	.w6(32'hbb983d13),
	.w7(32'hbbb11799),
	.w8(32'hbbf7482b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c224332),
	.w1(32'hbb1a61ad),
	.w2(32'hbc194321),
	.w3(32'h3c1df8f5),
	.w4(32'h3c1a75a5),
	.w5(32'hbc07ba31),
	.w6(32'h3c3152f3),
	.w7(32'h3bd57074),
	.w8(32'hbc28b5af),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19cfe1),
	.w1(32'h3a3a7215),
	.w2(32'hbbd347f8),
	.w3(32'hbb343e98),
	.w4(32'hba8d5af7),
	.w5(32'hbbbc50b8),
	.w6(32'hbc1bbb41),
	.w7(32'hbbcada90),
	.w8(32'hbc1b0d39),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b823b95),
	.w1(32'h3b535027),
	.w2(32'h3b972de6),
	.w3(32'h3b069ce8),
	.w4(32'hbb1f681c),
	.w5(32'h3b63edad),
	.w6(32'hbb3c44ac),
	.w7(32'hbbad6df4),
	.w8(32'hbb13ada6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6b960),
	.w1(32'hbbf1470c),
	.w2(32'hbc856fdc),
	.w3(32'h3c266fd7),
	.w4(32'h3c482795),
	.w5(32'hbad92e89),
	.w6(32'hbc627acf),
	.w7(32'hbc05b05a),
	.w8(32'hbc83c31b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c356460),
	.w1(32'h3c4bd474),
	.w2(32'hbb93c057),
	.w3(32'h3b68dea7),
	.w4(32'h3b56d60b),
	.w5(32'hbbf17a58),
	.w6(32'h3ba83174),
	.w7(32'h3aeb7b21),
	.w8(32'hbc3eafb1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d13ffa9),
	.w1(32'hbc09c27a),
	.w2(32'hbb73d375),
	.w3(32'h3ca08076),
	.w4(32'hbc64ff2e),
	.w5(32'hbc2dd325),
	.w6(32'h3c7c3b49),
	.w7(32'hbc5f7cc0),
	.w8(32'hbc968a55),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e8287),
	.w1(32'h3b639308),
	.w2(32'h3b21b093),
	.w3(32'h399c87c2),
	.w4(32'h3b0a116f),
	.w5(32'h3c110f99),
	.w6(32'h39ccf0f2),
	.w7(32'h3ab8dbb8),
	.w8(32'h3be81725),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3b61e),
	.w1(32'h3c5fecf7),
	.w2(32'h3a2295e6),
	.w3(32'h3ca71525),
	.w4(32'h3b959dff),
	.w5(32'hbc9ef2ee),
	.w6(32'h3befe3c0),
	.w7(32'hbb4fd6eb),
	.w8(32'hbcc94912),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03630b),
	.w1(32'h3c26670f),
	.w2(32'h3bb75db4),
	.w3(32'hbbb5f124),
	.w4(32'h3c08e0d4),
	.w5(32'hb9821e90),
	.w6(32'hbb7165f5),
	.w7(32'h3a552605),
	.w8(32'h3bc2a7e0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7fe4e),
	.w1(32'hbb08717f),
	.w2(32'h3b5dc9a9),
	.w3(32'hbb316acf),
	.w4(32'h3aadeb94),
	.w5(32'h3aaa2e0f),
	.w6(32'h3bbaab91),
	.w7(32'h3c49be92),
	.w8(32'hbc4ec50d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f7ce6),
	.w1(32'hbc4543ed),
	.w2(32'hbbb043d5),
	.w3(32'h3cc36699),
	.w4(32'h3c0fb90a),
	.w5(32'h3aefe89d),
	.w6(32'h3b3ff08d),
	.w7(32'h3bd0b283),
	.w8(32'hbb303a6a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25547f),
	.w1(32'h3bfdbe67),
	.w2(32'hbcc602f9),
	.w3(32'h3bfab160),
	.w4(32'h3b86eb35),
	.w5(32'hbcbf77fa),
	.w6(32'hbd1326dc),
	.w7(32'hbbec2ae2),
	.w8(32'hbd0e9946),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c981c8f),
	.w1(32'h3cd31191),
	.w2(32'h3aebd516),
	.w3(32'h3c0c9386),
	.w4(32'h3cad9d74),
	.w5(32'hbba03c77),
	.w6(32'hbbcc6238),
	.w7(32'h390af9de),
	.w8(32'h39778df9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc61054),
	.w1(32'h3b53b8e9),
	.w2(32'hba950528),
	.w3(32'h3c964989),
	.w4(32'h3c0d6142),
	.w5(32'h3a604234),
	.w6(32'h3c8df954),
	.w7(32'hbb4cfb61),
	.w8(32'hbc4d0800),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafc605),
	.w1(32'hbb3fa7a3),
	.w2(32'hbb4810c9),
	.w3(32'h3cbf17d3),
	.w4(32'hbbb89524),
	.w5(32'hbc25f6a8),
	.w6(32'h3cae7b65),
	.w7(32'hbc2962e5),
	.w8(32'hbc63365f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf99b79),
	.w1(32'hbc8274d4),
	.w2(32'hbbf61c0f),
	.w3(32'h3c4d4384),
	.w4(32'hbcbb6a12),
	.w5(32'hbca36341),
	.w6(32'hbc8ee9d1),
	.w7(32'hbce3a56d),
	.w8(32'hbd3aadbd),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd431d3),
	.w1(32'hbaa834cf),
	.w2(32'hbca1bc18),
	.w3(32'hbb003bdc),
	.w4(32'h3a98e360),
	.w5(32'hbc5cc90e),
	.w6(32'hbc67440c),
	.w7(32'hbc284800),
	.w8(32'hbcaf4889),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bc3de),
	.w1(32'hbc424d46),
	.w2(32'hbc39a2d1),
	.w3(32'hbc3b410e),
	.w4(32'hbc265628),
	.w5(32'hbc1faf76),
	.w6(32'hbcb4c1da),
	.w7(32'hbcba68cc),
	.w8(32'hbd0082d8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed30a3),
	.w1(32'hbbbe2dbf),
	.w2(32'hbaa56466),
	.w3(32'h3b09000d),
	.w4(32'h3b248d66),
	.w5(32'hbba16395),
	.w6(32'hbbe2217d),
	.w7(32'hbba89456),
	.w8(32'hbbd9957d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3765ca),
	.w1(32'hba9215ad),
	.w2(32'hbbc2ee8c),
	.w3(32'h3b7eb29b),
	.w4(32'h3bbc5aeb),
	.w5(32'hbbba53a0),
	.w6(32'hbbb2acce),
	.w7(32'hbc46cf14),
	.w8(32'hbc4c8101),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23be78),
	.w1(32'h3c4eaa57),
	.w2(32'h3a4b5d73),
	.w3(32'h3b8e32df),
	.w4(32'h3cc41028),
	.w5(32'h3b4343cb),
	.w6(32'hbc716188),
	.w7(32'hbbf4031e),
	.w8(32'h3b67c02b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4ca6d),
	.w1(32'hbc0d4474),
	.w2(32'hbaf3ff56),
	.w3(32'hb9e2a11b),
	.w4(32'h3aa22187),
	.w5(32'hbb319289),
	.w6(32'h3bb3950d),
	.w7(32'hbb97f1bc),
	.w8(32'hbc1577f6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d4104),
	.w1(32'h3b784e0e),
	.w2(32'h3ba6eb2d),
	.w3(32'hbbb49a9c),
	.w4(32'hbbb53369),
	.w5(32'h3b87db25),
	.w6(32'hbc2c7fda),
	.w7(32'hbc1b3b11),
	.w8(32'h3b5265d6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc455cdb),
	.w1(32'hbbc93bb2),
	.w2(32'hbc4ee52b),
	.w3(32'hbb55f414),
	.w4(32'h3aa63d11),
	.w5(32'hbc0997c8),
	.w6(32'hbc42d31e),
	.w7(32'hbc576f73),
	.w8(32'hbcf33d39),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34fce4),
	.w1(32'h3bf4fa25),
	.w2(32'hbc1c1c02),
	.w3(32'h3ae42048),
	.w4(32'h3b702325),
	.w5(32'hbc480927),
	.w6(32'hbbd13adc),
	.w7(32'hba8658eb),
	.w8(32'hbc7a36e6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba744d5c),
	.w1(32'h3c076e90),
	.w2(32'h3ab234b2),
	.w3(32'hbc67e947),
	.w4(32'hbacee617),
	.w5(32'hbabddbb0),
	.w6(32'hbc829113),
	.w7(32'hbc401b3c),
	.w8(32'hbbe5816d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe4ba1),
	.w1(32'hbaa650ba),
	.w2(32'hbc101a30),
	.w3(32'h3c647ea8),
	.w4(32'h3c33a494),
	.w5(32'hba2630a9),
	.w6(32'h3c5c19f3),
	.w7(32'hbbc3d793),
	.w8(32'hbbefd2e2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205d9b),
	.w1(32'h3cc2fc1c),
	.w2(32'hbc8e2542),
	.w3(32'hbc812f39),
	.w4(32'h3cb8064d),
	.w5(32'hbc8305b0),
	.w6(32'hbcf18b18),
	.w7(32'h3bdb03d0),
	.w8(32'hbc702055),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ecdf5),
	.w1(32'hbcc3565c),
	.w2(32'hbc909c00),
	.w3(32'hbcebaf59),
	.w4(32'hbc91c862),
	.w5(32'hbbef7508),
	.w6(32'hbce4d2bc),
	.w7(32'hbc5b1ed1),
	.w8(32'hbc58e5f6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb114473),
	.w1(32'hb9cb5e2a),
	.w2(32'hbb3d35b9),
	.w3(32'hbb9f8669),
	.w4(32'h376c1a8b),
	.w5(32'h3aa82509),
	.w6(32'hbb7c153d),
	.w7(32'hbb07f868),
	.w8(32'h3af9e9e5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b03e),
	.w1(32'hbc8be576),
	.w2(32'hbd425edf),
	.w3(32'h3b9c8e81),
	.w4(32'hbc4b62c4),
	.w5(32'hbd4cec54),
	.w6(32'hbd556989),
	.w7(32'hbce234af),
	.w8(32'hbd900e9a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d723d8a),
	.w1(32'hba0c6057),
	.w2(32'hbb3301bd),
	.w3(32'h3d53284c),
	.w4(32'hbbde4735),
	.w5(32'h39ebb2b2),
	.w6(32'h3d5542e5),
	.w7(32'hbc91b6cc),
	.w8(32'hbc2620de),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13a25),
	.w1(32'h3b40b6ab),
	.w2(32'h3b84c2f1),
	.w3(32'h3be9d3e3),
	.w4(32'h3bbd37c6),
	.w5(32'hbc0ea29b),
	.w6(32'h3b8b8279),
	.w7(32'hbc170e1f),
	.w8(32'hbc1eeea6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f39bb),
	.w1(32'hba5aace0),
	.w2(32'hba752e7d),
	.w3(32'hbbabd23c),
	.w4(32'h3996b1c5),
	.w5(32'hbac3e762),
	.w6(32'hbaf3f326),
	.w7(32'hbbbee33f),
	.w8(32'h3b24fcea),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bbecd),
	.w1(32'hb7af5a34),
	.w2(32'hb99c5d66),
	.w3(32'hbb4d719b),
	.w4(32'h3a8ccf7f),
	.w5(32'h3bbccb4d),
	.w6(32'hbba29155),
	.w7(32'hbafdd473),
	.w8(32'h3bc213c7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14d325),
	.w1(32'hbb50625d),
	.w2(32'hba64d725),
	.w3(32'h3c0ad7f8),
	.w4(32'h3b6633fa),
	.w5(32'hbaa4875c),
	.w6(32'h3c053a11),
	.w7(32'h3b894c96),
	.w8(32'h3aea9e8f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff1cbe),
	.w1(32'h3bc478de),
	.w2(32'hbb216088),
	.w3(32'hbabfb262),
	.w4(32'h3993352a),
	.w5(32'hba2b81e8),
	.w6(32'hbbbc2312),
	.w7(32'hbb3665fe),
	.w8(32'hbb7e3632),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cde51),
	.w1(32'hbbe36a06),
	.w2(32'hbbd8cc37),
	.w3(32'h3ba9d321),
	.w4(32'hba476403),
	.w5(32'hbaf273f8),
	.w6(32'hbc4b51b7),
	.w7(32'hbc72a986),
	.w8(32'hbc37bfc3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9c27),
	.w1(32'h3b70e6f3),
	.w2(32'hbaefce71),
	.w3(32'h3a8100a2),
	.w4(32'h3c35b782),
	.w5(32'h3c49fe13),
	.w6(32'h3b2f86eb),
	.w7(32'hbab702d2),
	.w8(32'hbbd96b65),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88f62d),
	.w1(32'hba9a76e9),
	.w2(32'h3b2d75c6),
	.w3(32'h3be76472),
	.w4(32'hbb1759ff),
	.w5(32'h38e59a20),
	.w6(32'h3aced482),
	.w7(32'hba1d687d),
	.w8(32'h3921ba7e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8344c9),
	.w1(32'h3bb63b68),
	.w2(32'hbc0cef60),
	.w3(32'h3c60de4b),
	.w4(32'h3a883920),
	.w5(32'hbc3c5716),
	.w6(32'hbc94f5d0),
	.w7(32'hbc90c03b),
	.w8(32'hbd2c6da3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76facb),
	.w1(32'hbbc54f35),
	.w2(32'hbc56c23b),
	.w3(32'h3cabe4b6),
	.w4(32'h3b76ee91),
	.w5(32'hbc7c6175),
	.w6(32'hb9595a99),
	.w7(32'hbb02bd72),
	.w8(32'hbb90da90),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac37a9),
	.w1(32'hbb563d90),
	.w2(32'hbb59e053),
	.w3(32'hbb3d0856),
	.w4(32'hbb42a863),
	.w5(32'h3bfa2850),
	.w6(32'h3a06eac3),
	.w7(32'h3ac33c7a),
	.w8(32'h3bac1916),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5351e9),
	.w1(32'hbbf312d1),
	.w2(32'hbc8ae0c7),
	.w3(32'hbbf6997a),
	.w4(32'hbb4cbefd),
	.w5(32'hbc9e804d),
	.w6(32'hbb492104),
	.w7(32'hbadd9e86),
	.w8(32'hbbf9797e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0909e),
	.w1(32'h3cb8a0ca),
	.w2(32'h3a9de553),
	.w3(32'hbbbe25c8),
	.w4(32'h3cb0ba95),
	.w5(32'hbbaecc1d),
	.w6(32'hbc8c4203),
	.w7(32'hbad8b1ab),
	.w8(32'hbbc67518),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe4603),
	.w1(32'h3cd22ab0),
	.w2(32'hbcbd9081),
	.w3(32'h3cb36eff),
	.w4(32'h3cc6c7d3),
	.w5(32'hbcdd7fa2),
	.w6(32'hba4bd4a0),
	.w7(32'hba1c1d1e),
	.w8(32'hbd1e2a73),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e61a8),
	.w1(32'h3cbb45bf),
	.w2(32'hbc2baead),
	.w3(32'hbbc4913e),
	.w4(32'h3cfefcf4),
	.w5(32'h3bcf4b33),
	.w6(32'hbc26f215),
	.w7(32'h3adb1c62),
	.w8(32'hbbafcaf2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1faae2),
	.w1(32'h3ab03a98),
	.w2(32'hbb68f079),
	.w3(32'h3c0c66c0),
	.w4(32'h3b09459e),
	.w5(32'h3b34ca39),
	.w6(32'h3a28b38d),
	.w7(32'hbb283f6e),
	.w8(32'hbc1d0bda),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c373de7),
	.w1(32'h3bd45cf7),
	.w2(32'hbc28998b),
	.w3(32'h3be2d179),
	.w4(32'h3b77fffa),
	.w5(32'hbc99ad30),
	.w6(32'h3b8f7562),
	.w7(32'h3b08cabd),
	.w8(32'hbc8b9bf4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce372d7),
	.w1(32'h3c49e0e4),
	.w2(32'hbc9f3033),
	.w3(32'h3c5677b4),
	.w4(32'h3c206154),
	.w5(32'hbb7e9b63),
	.w6(32'h3c1e0b30),
	.w7(32'hbc85c690),
	.w8(32'hbcb66a31),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d800f),
	.w1(32'hbb2c3ea7),
	.w2(32'hbbf2125d),
	.w3(32'hba90c40f),
	.w4(32'hbb3e0ec3),
	.w5(32'hbbba97f7),
	.w6(32'hbc784c00),
	.w7(32'hbc373c01),
	.w8(32'hbc9f02c1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cecd1bb),
	.w1(32'h3c867270),
	.w2(32'hbc3aa851),
	.w3(32'h3c87ed1d),
	.w4(32'h3b5ae222),
	.w5(32'hbc5d6851),
	.w6(32'hbc9f8457),
	.w7(32'hbcea7fb5),
	.w8(32'hbd06eb84),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810d97),
	.w1(32'hbb13b585),
	.w2(32'h3b238fe1),
	.w3(32'hbb0f3fd1),
	.w4(32'hbb890097),
	.w5(32'h3ad7d3a8),
	.w6(32'h3964889c),
	.w7(32'hbb1471c8),
	.w8(32'hbb89dc58),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd8fd),
	.w1(32'h3b8411f4),
	.w2(32'h3b34685c),
	.w3(32'hbaa6060d),
	.w4(32'hbac19835),
	.w5(32'h3b86b6a8),
	.w6(32'hbbb60c15),
	.w7(32'hbba5d4d0),
	.w8(32'h3bd1dee4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cd621),
	.w1(32'h3ca4fc8b),
	.w2(32'hbc205db7),
	.w3(32'h3c2f96b9),
	.w4(32'h3ca70cec),
	.w5(32'h3adbb0f5),
	.w6(32'hbd002c70),
	.w7(32'hbc571c6b),
	.w8(32'hbbf8dcdb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5b71b),
	.w1(32'hbbcd98ff),
	.w2(32'hbca51a82),
	.w3(32'h3c6f03b0),
	.w4(32'h3bf7f095),
	.w5(32'hbc610840),
	.w6(32'hbd160ef5),
	.w7(32'hbcefb4cb),
	.w8(32'hbd0388ef),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bd1a7),
	.w1(32'h3aad9382),
	.w2(32'hbb9cb9cb),
	.w3(32'h39d4af63),
	.w4(32'h3c3a4cba),
	.w5(32'h3b879985),
	.w6(32'hbc6d4c33),
	.w7(32'hbc0289fe),
	.w8(32'hbc5bb684),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7481fc),
	.w1(32'h3abd24be),
	.w2(32'h3c36f3af),
	.w3(32'hbb7fc9bd),
	.w4(32'hbc46250d),
	.w5(32'hbb86a33d),
	.w6(32'hbbf69664),
	.w7(32'hbc9a1352),
	.w8(32'hbcb06142),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57513b),
	.w1(32'hbb8a3f7d),
	.w2(32'h3903a88c),
	.w3(32'hbb97b570),
	.w4(32'hba619812),
	.w5(32'hba350564),
	.w6(32'hbbe51db4),
	.w7(32'hbb81f4a7),
	.w8(32'hb89dfb10),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad96dd),
	.w1(32'hbbc6eba8),
	.w2(32'hbb500891),
	.w3(32'hbb1782d7),
	.w4(32'hbbb9ecd0),
	.w5(32'hbc22a908),
	.w6(32'hbb3de106),
	.w7(32'hbae28991),
	.w8(32'hbb9c94a8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a757545),
	.w1(32'h3c10a665),
	.w2(32'hbbf72644),
	.w3(32'hbc24286e),
	.w4(32'hbb35a015),
	.w5(32'hbcdffc83),
	.w6(32'hbd0edeb5),
	.w7(32'h3b8c3ba3),
	.w8(32'hbca69289),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80a009),
	.w1(32'h3a03e433),
	.w2(32'hbbb3aac0),
	.w3(32'hbb13bab5),
	.w4(32'hbcc5c870),
	.w5(32'hbaca86ab),
	.w6(32'hbd0f98d6),
	.w7(32'hbd0d42ca),
	.w8(32'hbc9bd69e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf8658),
	.w1(32'hbcde9052),
	.w2(32'hbc8be0bd),
	.w3(32'hbac3022f),
	.w4(32'hbcc53184),
	.w5(32'hbc5e6ca4),
	.w6(32'hbc984806),
	.w7(32'h3b0690e1),
	.w8(32'hbcabe5e3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1f1ca9),
	.w1(32'h3c583697),
	.w2(32'h39e129d6),
	.w3(32'h3cc6b037),
	.w4(32'h3be7bf26),
	.w5(32'hbb8eb311),
	.w6(32'h3cb4dbcf),
	.w7(32'h3b2c39d3),
	.w8(32'hbc858018),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5fe6),
	.w1(32'hbba9f6e8),
	.w2(32'hbca2541c),
	.w3(32'h3c82e2c0),
	.w4(32'hba545f60),
	.w5(32'hbc0445f2),
	.w6(32'h3ca30d11),
	.w7(32'hbbf35f7f),
	.w8(32'hbc8ef16a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87465a),
	.w1(32'hbc31ecb1),
	.w2(32'h3ba70ba4),
	.w3(32'h3a6a1818),
	.w4(32'hbb3c12ff),
	.w5(32'h3c1ac4f0),
	.w6(32'h3b88544c),
	.w7(32'hbb71cf89),
	.w8(32'h3bc73455),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd54e4),
	.w1(32'hbc31c6a9),
	.w2(32'hbc3277ba),
	.w3(32'hba8e050a),
	.w4(32'hbc83a2fc),
	.w5(32'hbc506bd1),
	.w6(32'h3bbb3f95),
	.w7(32'hb8ae084c),
	.w8(32'hbc949514),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17e4b9),
	.w1(32'h3d391cdb),
	.w2(32'h3c78926f),
	.w3(32'h3c47de88),
	.w4(32'h3cd28d72),
	.w5(32'h3b80edd2),
	.w6(32'hbc825e67),
	.w7(32'hbc3881d1),
	.w8(32'h3ab9398b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba046e09),
	.w1(32'h39970cde),
	.w2(32'h3b4763f5),
	.w3(32'hb9c4000d),
	.w4(32'h3a0a6ee8),
	.w5(32'h3bcd566b),
	.w6(32'h394c8c23),
	.w7(32'h3b8db847),
	.w8(32'h3ac0a40d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111e80),
	.w1(32'h3c7d6160),
	.w2(32'hba91aa00),
	.w3(32'hbbdb86e9),
	.w4(32'h3c086a06),
	.w5(32'hbb9916f6),
	.w6(32'hbba0346e),
	.w7(32'hbbe6272c),
	.w8(32'hbc6e2050),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab608),
	.w1(32'hbc943fb8),
	.w2(32'hba694f3e),
	.w3(32'hbb730346),
	.w4(32'hbaf18976),
	.w5(32'hbb091c5e),
	.w6(32'hbd29404a),
	.w7(32'hbd0a5008),
	.w8(32'hbcbcd13a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b0631),
	.w1(32'h3bdb4149),
	.w2(32'hbb845e58),
	.w3(32'h3c044d63),
	.w4(32'h3bf9b06d),
	.w5(32'h3b9c9a3b),
	.w6(32'hbb61b1bf),
	.w7(32'hba24badd),
	.w8(32'hbbae1bbb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89ded6),
	.w1(32'h3bc4726c),
	.w2(32'hbbc052a5),
	.w3(32'h3b22f5f6),
	.w4(32'hbb3802b2),
	.w5(32'hbbf915ea),
	.w6(32'h3c007544),
	.w7(32'hbb020f10),
	.w8(32'hba96a3b6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb82cd),
	.w1(32'h3c4e7fbb),
	.w2(32'hbd20349b),
	.w3(32'hbc8286d2),
	.w4(32'h3ba52de7),
	.w5(32'hbcc50f66),
	.w6(32'hbd863aa8),
	.w7(32'hbc6102fb),
	.w8(32'hbd13fa04),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b411a7b),
	.w1(32'hbbd35885),
	.w2(32'hbb4cc9db),
	.w3(32'h3b96ffbb),
	.w4(32'hbbe750c7),
	.w5(32'hbb39e3fa),
	.w6(32'hbcbda2b7),
	.w7(32'hbcae575a),
	.w8(32'hbc567dbe),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4492bb),
	.w1(32'hbb89adf5),
	.w2(32'hbb83573a),
	.w3(32'hbb613e47),
	.w4(32'hbb4f24ab),
	.w5(32'hbbc7c2d0),
	.w6(32'hb99962f3),
	.w7(32'h3afe659f),
	.w8(32'hbb4c1562),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4998ca),
	.w1(32'h3ac2ff8a),
	.w2(32'hbc33fada),
	.w3(32'hbb6cca99),
	.w4(32'hbaea0ec6),
	.w5(32'hbc337ffa),
	.w6(32'hbc99eafa),
	.w7(32'hbc8056e8),
	.w8(32'hbcba25b6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b465f),
	.w1(32'h3c17bc1c),
	.w2(32'hb9db69c1),
	.w3(32'hbaea4661),
	.w4(32'h3c243396),
	.w5(32'hbb5a7b23),
	.w6(32'hbbb69c1d),
	.w7(32'h3b9a237d),
	.w8(32'hbc0611af),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f247c9),
	.w1(32'h3be4782d),
	.w2(32'hb9487438),
	.w3(32'hba036f93),
	.w4(32'h3c0907d4),
	.w5(32'h3b86419a),
	.w6(32'hbc54df67),
	.w7(32'hbb9ad785),
	.w8(32'h3b8dd4d9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeba522),
	.w1(32'hbb2a4464),
	.w2(32'hbad8e669),
	.w3(32'h3be0d683),
	.w4(32'h3a83f361),
	.w5(32'hbba3ddef),
	.w6(32'hba0c3ec6),
	.w7(32'h392f10e3),
	.w8(32'hbb3ae0f1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8769ed),
	.w1(32'h3c1dedfd),
	.w2(32'h3a69e93d),
	.w3(32'h39dc80ad),
	.w4(32'h3b79d07e),
	.w5(32'hbb87b461),
	.w6(32'hbbab7e53),
	.w7(32'hbb9b3d02),
	.w8(32'hb900bb3f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f03d),
	.w1(32'h3c25c6ce),
	.w2(32'hbaa47d21),
	.w3(32'hbb16e23e),
	.w4(32'hbb2bc2e0),
	.w5(32'hbc50f8d1),
	.w6(32'h3961cce7),
	.w7(32'hbbc84b85),
	.w8(32'hbc00e596),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08e3eb),
	.w1(32'h3bcdc980),
	.w2(32'hbbf5211c),
	.w3(32'hbb29ad99),
	.w4(32'hbb958c2b),
	.w5(32'hbc8eec8c),
	.w6(32'hbcb1ab31),
	.w7(32'hbcf9f8ed),
	.w8(32'hbd3144d5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c14e1),
	.w1(32'h3c4f2943),
	.w2(32'hbca9b7e0),
	.w3(32'hbbb75db2),
	.w4(32'h3ba29ae9),
	.w5(32'hbc45fd2b),
	.w6(32'hbcc4a1d8),
	.w7(32'hbcd4ac90),
	.w8(32'hbca097da),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbad8f9),
	.w1(32'h3bda4531),
	.w2(32'hbc5b5c1e),
	.w3(32'h3ca0cab1),
	.w4(32'hbaf8130e),
	.w5(32'hbc89b372),
	.w6(32'hbbf35fac),
	.w7(32'hbc9738f8),
	.w8(32'hbd18dac5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae178c6),
	.w1(32'h3adea59f),
	.w2(32'hbb5fd13c),
	.w3(32'hbbcd38d1),
	.w4(32'h3bedfb0c),
	.w5(32'hba8a51dd),
	.w6(32'hbbd89d6d),
	.w7(32'hbba65f56),
	.w8(32'hbbb8357d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b62b7),
	.w1(32'hb9d983fe),
	.w2(32'hbc27a237),
	.w3(32'h3a338e79),
	.w4(32'h3b402cb6),
	.w5(32'hbc3add5c),
	.w6(32'hbbc3640f),
	.w7(32'hbb939f50),
	.w8(32'h3b4904aa),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb674674),
	.w1(32'h3b31fb7f),
	.w2(32'hbc1d553e),
	.w3(32'hbcad8082),
	.w4(32'hbcb53fad),
	.w5(32'hba574021),
	.w6(32'hbb2e9661),
	.w7(32'hbc195a10),
	.w8(32'h37b50229),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f5a91),
	.w1(32'hba13a188),
	.w2(32'h3c0c42e4),
	.w3(32'h3be6e56e),
	.w4(32'h3c57c534),
	.w5(32'h3c00e862),
	.w6(32'h3b83ee33),
	.w7(32'h3bee5cc0),
	.w8(32'h3bded80e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde0005),
	.w1(32'hbc864718),
	.w2(32'hbc2c2621),
	.w3(32'h3a91b205),
	.w4(32'hbbd81a2c),
	.w5(32'hbbcb6922),
	.w6(32'hbbbe666c),
	.w7(32'hbc6a920b),
	.w8(32'hbc3b5cb9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d11e9),
	.w1(32'hbb06dacf),
	.w2(32'hbb7540c0),
	.w3(32'h3b6ddf5b),
	.w4(32'hba953a70),
	.w5(32'h3a544b47),
	.w6(32'h3bbba1f3),
	.w7(32'hbaf5275a),
	.w8(32'h38d64b05),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba999ff6),
	.w1(32'hbad18265),
	.w2(32'hbb4f2391),
	.w3(32'h3bd1ec80),
	.w4(32'hbbb51fba),
	.w5(32'hbc0e9126),
	.w6(32'h3a3a8686),
	.w7(32'h3b309913),
	.w8(32'hbbc72287),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebe5fb),
	.w1(32'hbb814dcd),
	.w2(32'hbca38b07),
	.w3(32'hbc350bbe),
	.w4(32'hbadbebda),
	.w5(32'hbc72af81),
	.w6(32'hbbbf8a9b),
	.w7(32'hbb9fd29c),
	.w8(32'hbc25c551),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23311d),
	.w1(32'h3af97056),
	.w2(32'hba6727d5),
	.w3(32'hbaecd888),
	.w4(32'hba8ad070),
	.w5(32'hbc33f219),
	.w6(32'hbb24b56c),
	.w7(32'h3a246a80),
	.w8(32'hbbe80ba0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb44486),
	.w1(32'h3cacfbd6),
	.w2(32'hbbde2412),
	.w3(32'hbb50071b),
	.w4(32'h3c1220a6),
	.w5(32'hbb99f069),
	.w6(32'hbc36f39f),
	.w7(32'hbab29b17),
	.w8(32'hbc076c28),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed35ef),
	.w1(32'h3b614d73),
	.w2(32'hbbb505a9),
	.w3(32'h3b82c299),
	.w4(32'h3ba2fc71),
	.w5(32'hbb879777),
	.w6(32'hbb03371e),
	.w7(32'h3ade03e0),
	.w8(32'hbb95d251),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823176),
	.w1(32'hbc0e3082),
	.w2(32'hbc83da0d),
	.w3(32'hbbd865da),
	.w4(32'hbc4d5b0e),
	.w5(32'h3c54f7f9),
	.w6(32'hbcb0bb70),
	.w7(32'hbcd594b9),
	.w8(32'hbc439978),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02576b),
	.w1(32'hba35f8ac),
	.w2(32'h3aee0808),
	.w3(32'h3ae8abba),
	.w4(32'h3a5b631f),
	.w5(32'h3b849686),
	.w6(32'h3b839a6a),
	.w7(32'h3ad9904a),
	.w8(32'h3bccf780),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e02ac),
	.w1(32'h3ca6b35d),
	.w2(32'h3c12cbbc),
	.w3(32'hbc856dd1),
	.w4(32'h3bdaacfa),
	.w5(32'h3c021ce2),
	.w6(32'hbcde3b8e),
	.w7(32'h3b0d5f27),
	.w8(32'h3c2c7489),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule