module layer_6_featuremap_14(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb796f62f),
	.w1(32'hb76ef4ce),
	.w2(32'hb829a666),
	.w3(32'hb66c3717),
	.w4(32'h35940fff),
	.w5(32'hb75b2e6b),
	.w6(32'hb6201c86),
	.w7(32'hb6c99cad),
	.w8(32'hb7be3070),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8257c9a),
	.w1(32'hb7dc6cab),
	.w2(32'hb8bdd026),
	.w3(32'hb6c03334),
	.w4(32'h359c0bb5),
	.w5(32'hb885aafc),
	.w6(32'hb717666b),
	.w7(32'hb653c9e2),
	.w8(32'hb889e7f0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c79bd3),
	.w1(32'hb74e036e),
	.w2(32'h36ad4cf7),
	.w3(32'hb7f00778),
	.w4(32'hb7cba14c),
	.w5(32'hb724a2e0),
	.w6(32'h36655ee8),
	.w7(32'h38145d38),
	.w8(32'h384efb0d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a38880),
	.w1(32'h395e89b8),
	.w2(32'h38dea8a7),
	.w3(32'h3991781e),
	.w4(32'h39216f5a),
	.w5(32'h38fd32ce),
	.w6(32'h39585627),
	.w7(32'h3915139e),
	.w8(32'h38c12945),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894c607),
	.w1(32'h381a22f8),
	.w2(32'h36488e7b),
	.w3(32'h3866f7cb),
	.w4(32'h37e26780),
	.w5(32'h37b04ebf),
	.w6(32'h378a56ba),
	.w7(32'h37807d56),
	.w8(32'h37fb5154),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f0001),
	.w1(32'h383930e7),
	.w2(32'h382f7125),
	.w3(32'h388be3c6),
	.w4(32'h383da60d),
	.w5(32'h384e3a38),
	.w6(32'h387ee268),
	.w7(32'h384fecd7),
	.w8(32'h382e4552),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3889e977),
	.w1(32'h38aa6566),
	.w2(32'h3a6ba23b),
	.w3(32'hb991061c),
	.w4(32'hb9912d0d),
	.w5(32'h3a21f686),
	.w6(32'hb9a2286d),
	.w7(32'hb9ab57c8),
	.w8(32'h3a0af80f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912fd28),
	.w1(32'h386b5c49),
	.w2(32'h38cfb8af),
	.w3(32'h38d78408),
	.w4(32'h381bce19),
	.w5(32'h38b1b191),
	.w6(32'h393099f0),
	.w7(32'h388f85c9),
	.w8(32'h38dfbf53),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a76ab),
	.w1(32'h3703269b),
	.w2(32'h37b4a9d2),
	.w3(32'hb7f46423),
	.w4(32'hb723fe72),
	.w5(32'h386fa32a),
	.w6(32'hb8338d59),
	.w7(32'hb78e5381),
	.w8(32'h38927928),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da18cf),
	.w1(32'h38da00e6),
	.w2(32'h398c39e7),
	.w3(32'hb6b8c2fb),
	.w4(32'hb7bd5671),
	.w5(32'h3990885e),
	.w6(32'h3817b269),
	.w7(32'h380f8565),
	.w8(32'h3993ca22),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381746e7),
	.w1(32'h3898a78a),
	.w2(32'h38c9bed7),
	.w3(32'h389521bd),
	.w4(32'h390ec587),
	.w5(32'h390b4354),
	.w6(32'h38c273cd),
	.w7(32'h3934649d),
	.w8(32'h393e4738),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c16a9d),
	.w1(32'hb6b31a79),
	.w2(32'h39008b95),
	.w3(32'hb7b82586),
	.w4(32'hb81c0384),
	.w5(32'h38b3bee1),
	.w6(32'hb7b22a4a),
	.w7(32'hb86ad54b),
	.w8(32'h38d1a999),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84130a5),
	.w1(32'hb7e2e579),
	.w2(32'hb76fb9a5),
	.w3(32'hb7f3fad4),
	.w4(32'hb63015a5),
	.w5(32'hb66234c0),
	.w6(32'hb74bc99c),
	.w7(32'hb7aa991d),
	.w8(32'hb7506e7b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911e6ce),
	.w1(32'hb893bb40),
	.w2(32'h3a098210),
	.w3(32'hb980e910),
	.w4(32'hb932ee1f),
	.w5(32'h3a1f9f51),
	.w6(32'hb9f186c4),
	.w7(32'hb996ac59),
	.w8(32'h39eb64ce),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c6550),
	.w1(32'hb878c981),
	.w2(32'h387ec1fb),
	.w3(32'hb8d2e232),
	.w4(32'hb8c87f5b),
	.w5(32'h386360c7),
	.w6(32'hb8af23b3),
	.w7(32'hb8bb2043),
	.w8(32'h3881c990),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d66a28),
	.w1(32'hb789bfbb),
	.w2(32'h39479f0b),
	.w3(32'h3779c613),
	.w4(32'hb815ed9e),
	.w5(32'h392bef9b),
	.w6(32'h3870446f),
	.w7(32'h37dc28f6),
	.w8(32'h39906563),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d334d),
	.w1(32'hb944a052),
	.w2(32'h3923b77c),
	.w3(32'hb93f4c86),
	.w4(32'hb99ae3f6),
	.w5(32'h392cc8f3),
	.w6(32'hb89f1209),
	.w7(32'hb774fe08),
	.w8(32'h39d8e639),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b57410),
	.w1(32'hb64aa531),
	.w2(32'hb7555ae5),
	.w3(32'h370ad310),
	.w4(32'hb58a5c3f),
	.w5(32'hb731d36d),
	.w6(32'h3730b29f),
	.w7(32'h36b30809),
	.w8(32'hb6fdaed2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eba244),
	.w1(32'h398315a6),
	.w2(32'h38d72fb0),
	.w3(32'h39a5e96b),
	.w4(32'h38af9f2d),
	.w5(32'h3804da9c),
	.w6(32'h398bb676),
	.w7(32'h3893d3ee),
	.w8(32'h3883ed26),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f64e1),
	.w1(32'h38557295),
	.w2(32'hb890f9f0),
	.w3(32'h385fa297),
	.w4(32'h372caaae),
	.w5(32'h38c55e7e),
	.w6(32'h38df6cee),
	.w7(32'h3900af66),
	.w8(32'h38e0a8a7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d6ebdd),
	.w1(32'h37ea5aa0),
	.w2(32'h37a083f0),
	.w3(32'h379a80d5),
	.w4(32'h37c638bf),
	.w5(32'h36cfbc29),
	.w6(32'h3799a046),
	.w7(32'h380eccf6),
	.w8(32'h37029106),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0c67a),
	.w1(32'h395e27db),
	.w2(32'h38e0fb41),
	.w3(32'h39b53179),
	.w4(32'h397bc671),
	.w5(32'h3985980c),
	.w6(32'h39c7d87a),
	.w7(32'h39a09120),
	.w8(32'h39936efc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee7351),
	.w1(32'hb8c42d14),
	.w2(32'h3994af70),
	.w3(32'hb976a350),
	.w4(32'hb95f08d6),
	.w5(32'hb68baa18),
	.w6(32'hb8fcffe4),
	.w7(32'hb8f3e97f),
	.w8(32'h3838bc75),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38687f46),
	.w1(32'h390c69fb),
	.w2(32'h38f21e99),
	.w3(32'h39092364),
	.w4(32'h390643ec),
	.w5(32'h392e5b8d),
	.w6(32'h397f8c68),
	.w7(32'h398dd30b),
	.w8(32'h398a916f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f5277),
	.w1(32'h39883574),
	.w2(32'h38f63945),
	.w3(32'h39908c12),
	.w4(32'hb54eae1a),
	.w5(32'hb89ca16f),
	.w6(32'h39913557),
	.w7(32'h38961fc2),
	.w8(32'h37500d0b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44bd05),
	.w1(32'h3a1d2b8f),
	.w2(32'h3a3b9856),
	.w3(32'h39f3fdae),
	.w4(32'h399cc50d),
	.w5(32'h3a3bd4da),
	.w6(32'h39612976),
	.w7(32'h392b5fb9),
	.w8(32'h3a0ff8e2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38739ecd),
	.w1(32'h383929df),
	.w2(32'h38b3451f),
	.w3(32'h38d43f9f),
	.w4(32'h38c69a43),
	.w5(32'h391ee7bb),
	.w6(32'h3898b955),
	.w7(32'h3859cbc2),
	.w8(32'h38ac0707),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372adf84),
	.w1(32'hb90d6197),
	.w2(32'h384e96af),
	.w3(32'h37d2194c),
	.w4(32'hb90364a6),
	.w5(32'h38614d3f),
	.w6(32'h37c307cd),
	.w7(32'hb90a56e6),
	.w8(32'h3842925f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70eda1d),
	.w1(32'h3767d5fe),
	.w2(32'h38751976),
	.w3(32'h37e45e17),
	.w4(32'h3857a397),
	.w5(32'h380e7f69),
	.w6(32'h37f3d12a),
	.w7(32'h3846ed39),
	.w8(32'h38419f75),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fb07a),
	.w1(32'h3a617016),
	.w2(32'h3a4bf379),
	.w3(32'h3a46240c),
	.w4(32'h3a05036e),
	.w5(32'h3a467afc),
	.w6(32'h39cf928e),
	.w7(32'h398ed8e2),
	.w8(32'h3a05ce40),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aab2b0),
	.w1(32'hbad91fbd),
	.w2(32'hb963d1b7),
	.w3(32'hb6895139),
	.w4(32'hba457ecc),
	.w5(32'hba991141),
	.w6(32'hbafbd314),
	.w7(32'hb7bdf4cb),
	.w8(32'h3abcd612),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a8fbc),
	.w1(32'hbb98fda5),
	.w2(32'hbb926fd6),
	.w3(32'hba5f1a4e),
	.w4(32'hbb4b4d41),
	.w5(32'hbb49a77b),
	.w6(32'hbb9d568a),
	.w7(32'hbb7cb02e),
	.w8(32'hbac3dc99),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb311308),
	.w1(32'hb7d4a888),
	.w2(32'hbb1de129),
	.w3(32'hbb13d53a),
	.w4(32'h3b6c986a),
	.w5(32'h3b39a74f),
	.w6(32'hbb6a3fa5),
	.w7(32'hbb91943d),
	.w8(32'hbb308bef),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8d3da),
	.w1(32'hbb7ee0ec),
	.w2(32'hbb23df01),
	.w3(32'h3b5fd633),
	.w4(32'hbb39570e),
	.w5(32'hbaf8a24c),
	.w6(32'hbbba3a1f),
	.w7(32'hbb94b14c),
	.w8(32'hbb3e9fc0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c772e),
	.w1(32'h3a8311e0),
	.w2(32'h3abce5f8),
	.w3(32'hb9f7c6f9),
	.w4(32'h39f1e687),
	.w5(32'h3a583a81),
	.w6(32'h3a082e85),
	.w7(32'h3a10b3ee),
	.w8(32'hbb0db626),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43fc8f),
	.w1(32'hbb0e4085),
	.w2(32'hbbaa22d0),
	.w3(32'hba802868),
	.w4(32'hbad22c63),
	.w5(32'hbb712c25),
	.w6(32'h3908a606),
	.w7(32'hbad4cc5f),
	.w8(32'hb9e6c14b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d5b94),
	.w1(32'hbb8b2530),
	.w2(32'hbb5e025b),
	.w3(32'hba746d2d),
	.w4(32'hbb897e7a),
	.w5(32'hbb6933eb),
	.w6(32'hbb871574),
	.w7(32'hbb764b5c),
	.w8(32'hbb827f54),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb719966),
	.w1(32'hbaa5084f),
	.w2(32'hb96c6b2d),
	.w3(32'hbb84068e),
	.w4(32'hbb483de7),
	.w5(32'hba708348),
	.w6(32'hbaf91721),
	.w7(32'hbb234e6d),
	.w8(32'hbb17d84f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9854705),
	.w1(32'hb96a37e2),
	.w2(32'hba257baa),
	.w3(32'hba0e1d16),
	.w4(32'h38a4c194),
	.w5(32'hb9954d05),
	.w6(32'h3a0f98c9),
	.w7(32'h39b93eb5),
	.w8(32'h3a95ae35),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3988ad),
	.w1(32'hbaf895a1),
	.w2(32'hbb3f1ff8),
	.w3(32'h3a537976),
	.w4(32'hbb57a32c),
	.w5(32'hbb4e5a9a),
	.w6(32'hbb2f7dbe),
	.w7(32'hbb58c021),
	.w8(32'hbb0d936d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b2720),
	.w1(32'hbb6480c4),
	.w2(32'hbb54add8),
	.w3(32'hbb2726f6),
	.w4(32'hbb5bd944),
	.w5(32'hbb5f4899),
	.w6(32'hbb6ad25b),
	.w7(32'hbb63b455),
	.w8(32'hbb5c6af0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c0b74),
	.w1(32'hb96d9d03),
	.w2(32'hb90e23ca),
	.w3(32'hbb5b1f18),
	.w4(32'hb95a03d7),
	.w5(32'hb89a3068),
	.w6(32'hb862546b),
	.w7(32'hb73be478),
	.w8(32'h39a1422f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fadc8),
	.w1(32'h3ade5353),
	.w2(32'h3b1e11ad),
	.w3(32'hb899e930),
	.w4(32'h3a9f4c48),
	.w5(32'h3ac1c58c),
	.w6(32'hb939ce66),
	.w7(32'h39f6cfbb),
	.w8(32'hbaad3f4b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a0258),
	.w1(32'hbb9550ac),
	.w2(32'hbb46bb1c),
	.w3(32'h38cd15b2),
	.w4(32'hbbe341c9),
	.w5(32'hbb050558),
	.w6(32'hbb70b52a),
	.w7(32'hbb7e7260),
	.w8(32'hbb915cb2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9426f),
	.w1(32'hb9cbe18c),
	.w2(32'h3a902557),
	.w3(32'h3a8075fa),
	.w4(32'h39c40708),
	.w5(32'h3afe7793),
	.w6(32'hb949ba28),
	.w7(32'h3a6bcb6d),
	.w8(32'hba53927c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0af93),
	.w1(32'h3b4bc5c1),
	.w2(32'h3b384ea5),
	.w3(32'hb98aa799),
	.w4(32'h3b3b201d),
	.w5(32'h3b19aa76),
	.w6(32'h3b81302e),
	.w7(32'h3b88b664),
	.w8(32'h3b7c8112),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ee571),
	.w1(32'hbb03a4e5),
	.w2(32'hbaca7d34),
	.w3(32'h3a9eb787),
	.w4(32'hbab79d66),
	.w5(32'h3a1755bb),
	.w6(32'hbb297327),
	.w7(32'hbb169fb9),
	.w8(32'hbab8fdc1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131e00),
	.w1(32'hb87f1bff),
	.w2(32'h3ab3ebe8),
	.w3(32'h3abb9701),
	.w4(32'h3a8f7d0a),
	.w5(32'h3af97949),
	.w6(32'hbad8f1f6),
	.w7(32'h3996b0b5),
	.w8(32'h3a442332),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a60414),
	.w1(32'hbb638456),
	.w2(32'hbba9d246),
	.w3(32'hb8b2633b),
	.w4(32'hbb5bfd94),
	.w5(32'hbb859fa7),
	.w6(32'hbb096c6e),
	.w7(32'hbb092a97),
	.w8(32'hbab4a66e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63a3aa),
	.w1(32'h3be17d47),
	.w2(32'h3b6c663b),
	.w3(32'hbaec104f),
	.w4(32'h3ba8ad24),
	.w5(32'h3b199b8d),
	.w6(32'h3be43d10),
	.w7(32'h3b464f5d),
	.w8(32'hbb608714),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907211),
	.w1(32'hbb6cc5a3),
	.w2(32'hbb676a56),
	.w3(32'hbba4b0f2),
	.w4(32'hbb5f9aeb),
	.w5(32'hbb656e04),
	.w6(32'hbb78a62b),
	.w7(32'hbb78fb93),
	.w8(32'hbb640faf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72fdd1),
	.w1(32'hbb42d51b),
	.w2(32'hba4b1192),
	.w3(32'hbb7ba68f),
	.w4(32'hbb43dc1d),
	.w5(32'hba298a28),
	.w6(32'hbb3d2d9a),
	.w7(32'hba9113f1),
	.w8(32'hbaf02323),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f03b3),
	.w1(32'h3751073e),
	.w2(32'hb84eafb3),
	.w3(32'hbb176bb0),
	.w4(32'h382a5447),
	.w5(32'h3a1d7573),
	.w6(32'hb9c7cd07),
	.w7(32'hba8298b0),
	.w8(32'hba2b8fb2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fc2e0),
	.w1(32'hbb9ff879),
	.w2(32'hbb9fa51c),
	.w3(32'hb81452ab),
	.w4(32'hbba9722f),
	.w5(32'hbba7407a),
	.w6(32'hbb9c9648),
	.w7(32'hbba8b306),
	.w8(32'hbbb3e538),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac393d),
	.w1(32'h3a56cfff),
	.w2(32'hb9187479),
	.w3(32'hbbaf914b),
	.w4(32'h3aee5955),
	.w5(32'h3a92d6f4),
	.w6(32'hba66cf6b),
	.w7(32'hbb0072ab),
	.w8(32'hbb27b45f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6e10),
	.w1(32'hba6378a0),
	.w2(32'hbabdf346),
	.w3(32'hb919ddc0),
	.w4(32'hbae9d9a3),
	.w5(32'hbb3998a1),
	.w6(32'hbb13ed84),
	.w7(32'hbaca8c3e),
	.w8(32'hba870949),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8acf67),
	.w1(32'hb9bb3c54),
	.w2(32'hbb0d5868),
	.w3(32'hbadc1115),
	.w4(32'h3aca5bde),
	.w5(32'h3ab5104b),
	.w6(32'hb90455fa),
	.w7(32'hba9b0ec1),
	.w8(32'h3b0bc43c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cac21),
	.w1(32'h3a7bd5df),
	.w2(32'h3a08033e),
	.w3(32'h3a5e8822),
	.w4(32'h3b47f5a3),
	.w5(32'h3b0c59df),
	.w6(32'h3ad7b5c6),
	.w7(32'h3b0220bb),
	.w8(32'h3b83a486),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b744c6a),
	.w1(32'hbb272670),
	.w2(32'hbb168d9c),
	.w3(32'h3b754cc1),
	.w4(32'hbb200c8b),
	.w5(32'hbb196701),
	.w6(32'hba8bf977),
	.w7(32'hb99166c4),
	.w8(32'hb9d9199a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bb61e),
	.w1(32'hba941523),
	.w2(32'hb963941b),
	.w3(32'hbad16e6c),
	.w4(32'hb9bf3fe8),
	.w5(32'h3adcec27),
	.w6(32'hbab1f6cb),
	.w7(32'hbaefe304),
	.w8(32'hba10997f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac271cd),
	.w1(32'h3a857969),
	.w2(32'h3b4efead),
	.w3(32'h3b197ed2),
	.w4(32'hba4b33a2),
	.w5(32'h3ac455cc),
	.w6(32'h3adba81d),
	.w7(32'h3af52c5f),
	.w8(32'h3a668196),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd29a4),
	.w1(32'hba64efdf),
	.w2(32'hbac8fcd2),
	.w3(32'h384b5991),
	.w4(32'hba955bc7),
	.w5(32'hbab87999),
	.w6(32'hb66a0be8),
	.w7(32'hba793b0d),
	.w8(32'hb8ce2bbc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa86a14),
	.w1(32'h3ab7f275),
	.w2(32'h3a917c36),
	.w3(32'h3a92bb27),
	.w4(32'h3a8b595f),
	.w5(32'h3a52cc6f),
	.w6(32'h3a1a0e1e),
	.w7(32'h39b94fce),
	.w8(32'h39bc8c03),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41e367),
	.w1(32'h39eaf715),
	.w2(32'h3991437b),
	.w3(32'h3a004ed7),
	.w4(32'h3965a5c7),
	.w5(32'h39a48e58),
	.w6(32'h39c54d25),
	.w7(32'h39674dcb),
	.w8(32'h39a2df09),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule