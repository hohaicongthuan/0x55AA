module layer_8_featuremap_198(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9379f2),
	.w1(32'h3b80d30f),
	.w2(32'h3ccbd2d0),
	.w3(32'h3c0796c7),
	.w4(32'hbbe136ac),
	.w5(32'h3b0f0dfb),
	.w6(32'h39cc404d),
	.w7(32'h3caf75c0),
	.w8(32'h3cb91f09),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca09f1b),
	.w1(32'hbb4ecb5b),
	.w2(32'h3a8d30f3),
	.w3(32'h3ae6fe81),
	.w4(32'h38c9d1c0),
	.w5(32'h3a8d979b),
	.w6(32'hb6f38dfb),
	.w7(32'h3a0c0374),
	.w8(32'h3aa94ec7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882c0c4),
	.w1(32'h3be1962c),
	.w2(32'h3b6c4805),
	.w3(32'h3b98a525),
	.w4(32'h3b9bd04e),
	.w5(32'h3be3702e),
	.w6(32'hbac884bc),
	.w7(32'h39a8e349),
	.w8(32'hb9887556),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b991e62),
	.w1(32'hbc18eee4),
	.w2(32'hbc9c178f),
	.w3(32'hba3ef7f0),
	.w4(32'h3bb1011b),
	.w5(32'h39edf858),
	.w6(32'hbc2ce19d),
	.w7(32'hbb89a43a),
	.w8(32'hbbd56207),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07cd92),
	.w1(32'h3b93afd3),
	.w2(32'hbb611aa8),
	.w3(32'hbc278581),
	.w4(32'h3c42ec19),
	.w5(32'h3b622d4d),
	.w6(32'h3a374c78),
	.w7(32'hbb8a1756),
	.w8(32'hbbc3b9d1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe61f58),
	.w1(32'hbc17383c),
	.w2(32'hbbe62a9f),
	.w3(32'h3b815be3),
	.w4(32'hbc581ab0),
	.w5(32'hbbba2cc3),
	.w6(32'h3b5ded7f),
	.w7(32'hbc0ae0e3),
	.w8(32'hbc982fde),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b31ee),
	.w1(32'h3b8d8163),
	.w2(32'hbb53cc3c),
	.w3(32'hbbfe1b9b),
	.w4(32'h3c637610),
	.w5(32'h3be59f95),
	.w6(32'hb98e1de3),
	.w7(32'hbc09901d),
	.w8(32'hbbfab8c8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9860d7),
	.w1(32'h3c69b11b),
	.w2(32'h3cb8d22e),
	.w3(32'h3b61d97c),
	.w4(32'h3b3286d1),
	.w5(32'h3bdf3643),
	.w6(32'h3c9ead67),
	.w7(32'h3cfa3896),
	.w8(32'h3cb4f25c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9401),
	.w1(32'h3976d140),
	.w2(32'hbc7da41a),
	.w3(32'hbb27f91a),
	.w4(32'hbadb6ee8),
	.w5(32'hbc91e5fa),
	.w6(32'h3c8b14bc),
	.w7(32'h3aa70953),
	.w8(32'hb9ae7b0c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c1b3),
	.w1(32'h3c98887e),
	.w2(32'h3c840358),
	.w3(32'hbb612bee),
	.w4(32'h3bf9e78d),
	.w5(32'h3ba6a76c),
	.w6(32'h3c20eb6c),
	.w7(32'h3cb410f0),
	.w8(32'h3c58a54f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b7f6c),
	.w1(32'h3bd87473),
	.w2(32'hbbf9a1ee),
	.w3(32'h3c256da4),
	.w4(32'h3c101c20),
	.w5(32'h3b5f8a96),
	.w6(32'hba562732),
	.w7(32'hba26dbbd),
	.w8(32'h3ad1c064),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bd3fa),
	.w1(32'hbc43df8e),
	.w2(32'hbc4c9667),
	.w3(32'h3be7d6af),
	.w4(32'hbbf7486a),
	.w5(32'hbc0d008e),
	.w6(32'hbc030679),
	.w7(32'hbc3b2695),
	.w8(32'hbc02edf9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc674f70),
	.w1(32'hba6e9dc9),
	.w2(32'h3a95537f),
	.w3(32'hbc596970),
	.w4(32'hbb6fb36c),
	.w5(32'hba53e37a),
	.w6(32'h3b1ecb78),
	.w7(32'hbb13a15f),
	.w8(32'h3af0cf52),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db04d),
	.w1(32'h3c8dde3f),
	.w2(32'h3cb82a3e),
	.w3(32'hbb9bb151),
	.w4(32'h3c5119e0),
	.w5(32'h3cc16d22),
	.w6(32'h3bf105b7),
	.w7(32'h3bf3a5c6),
	.w8(32'hb9a7cf77),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43d31b),
	.w1(32'h3c040367),
	.w2(32'h39cee47f),
	.w3(32'h3c4aea99),
	.w4(32'h3bd9de1e),
	.w5(32'h3b21bb25),
	.w6(32'h3ba8065b),
	.w7(32'hbb8f8ba2),
	.w8(32'hbb337521),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba074338),
	.w1(32'hb8919bba),
	.w2(32'h3bf022fa),
	.w3(32'hbac9df8c),
	.w4(32'h3c092b47),
	.w5(32'h3bd8f953),
	.w6(32'hbac2d59a),
	.w7(32'h3c01278b),
	.w8(32'h3c778679),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c977acb),
	.w1(32'hb8fc8ae4),
	.w2(32'hbb942088),
	.w3(32'hba5daa43),
	.w4(32'hbb314f62),
	.w5(32'hbc1122b0),
	.w6(32'hbb87db3e),
	.w7(32'hbc133b8a),
	.w8(32'hbc08f2ee),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec4cbd),
	.w1(32'h3b332d2d),
	.w2(32'h3b2f5795),
	.w3(32'hbae02f0d),
	.w4(32'h3c92eb22),
	.w5(32'h3cf15717),
	.w6(32'hba5ab172),
	.w7(32'hbbdcdca7),
	.w8(32'h3a8aeb87),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad1035),
	.w1(32'h3cbbb520),
	.w2(32'h3c101dd0),
	.w3(32'h3d025184),
	.w4(32'h3c8b5bc6),
	.w5(32'h3c8a38f9),
	.w6(32'h3c70fa7e),
	.w7(32'h3b850fae),
	.w8(32'h3ba5ee3a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c320eb6),
	.w1(32'h3b8a2bf8),
	.w2(32'hbab540e0),
	.w3(32'h3cae6b1b),
	.w4(32'hbaaa940f),
	.w5(32'hbb51d911),
	.w6(32'h3b20e23e),
	.w7(32'hbb8c9339),
	.w8(32'hbb9624bb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0e092),
	.w1(32'hbc3b7b8e),
	.w2(32'hbcb98ca1),
	.w3(32'hbc73e453),
	.w4(32'hbac5d510),
	.w5(32'hbb97db86),
	.w6(32'hbbfcbad1),
	.w7(32'hbc71a388),
	.w8(32'hbc84968e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc730c76),
	.w1(32'h3b1f6fd5),
	.w2(32'h3c4150a1),
	.w3(32'hba517155),
	.w4(32'h3b805823),
	.w5(32'h3c381442),
	.w6(32'h3bd0a85c),
	.w7(32'hbb0f83ae),
	.w8(32'hbaf7be2f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98b588),
	.w1(32'h3ccd6216),
	.w2(32'h3c79030d),
	.w3(32'h3c38da15),
	.w4(32'h3cf747ac),
	.w5(32'h3c5d42db),
	.w6(32'hbb153076),
	.w7(32'h3c21a4fc),
	.w8(32'h3b128136),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440cc2),
	.w1(32'h3b8c2fe5),
	.w2(32'h3bcc58d4),
	.w3(32'hbb8a3815),
	.w4(32'h3ae01b55),
	.w5(32'h3c3a03db),
	.w6(32'hbba16b0c),
	.w7(32'hbb8d6e58),
	.w8(32'hbc1de949),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad807ae),
	.w1(32'hbaedec9b),
	.w2(32'hbc80a2de),
	.w3(32'h3ac1f110),
	.w4(32'h3cb7994b),
	.w5(32'h3c2cb0b2),
	.w6(32'hbbd7ccaa),
	.w7(32'hbc2bcd8a),
	.w8(32'hbb9b5c29),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b4cb7),
	.w1(32'h3d0416bd),
	.w2(32'h3d55443f),
	.w3(32'h3c0d6b8a),
	.w4(32'h3cb85ae0),
	.w5(32'h3d0fffd6),
	.w6(32'h3c251c7e),
	.w7(32'h3cc54e41),
	.w8(32'h3c44b009),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82954c),
	.w1(32'hbc8910b8),
	.w2(32'hbcab8014),
	.w3(32'h3c97bec9),
	.w4(32'hbc45d744),
	.w5(32'hbbfe620f),
	.w6(32'hbc2777cb),
	.w7(32'hbc8e6084),
	.w8(32'hbc810334),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4ad89f),
	.w1(32'hbc86287d),
	.w2(32'hbc2cc747),
	.w3(32'hbcc3178a),
	.w4(32'hbb4b2c80),
	.w5(32'hbc6e91f0),
	.w6(32'hbd4a2591),
	.w7(32'hbc948972),
	.w8(32'hbb9052e4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe0c77),
	.w1(32'h3b9c613a),
	.w2(32'hbbd12288),
	.w3(32'h3a55b085),
	.w4(32'h3a860d1d),
	.w5(32'hbc0db404),
	.w6(32'h3b678b9c),
	.w7(32'hbc059d4e),
	.w8(32'hbb00309b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf48ff1),
	.w1(32'h375ede72),
	.w2(32'h395729dc),
	.w3(32'hbc8d5093),
	.w4(32'h3c536d22),
	.w5(32'h3c057c98),
	.w6(32'hbba94867),
	.w7(32'hbb7e7736),
	.w8(32'hbbc3e516),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cf1fb),
	.w1(32'h3c0b82d6),
	.w2(32'hbae2fc0e),
	.w3(32'h3c109568),
	.w4(32'h3abba54d),
	.w5(32'hbc4b9f1b),
	.w6(32'h3b86b437),
	.w7(32'hbc120b74),
	.w8(32'hbbf21493),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c975),
	.w1(32'h3b0f9e71),
	.w2(32'h3ba75c6e),
	.w3(32'hbc8b98c0),
	.w4(32'hbbd52c5b),
	.w5(32'h3a1702b1),
	.w6(32'h3c43f711),
	.w7(32'h3b914639),
	.w8(32'hbb1491ee),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994b2bc),
	.w1(32'hbb1480c6),
	.w2(32'hbc24df0b),
	.w3(32'hba92aaca),
	.w4(32'hbba3b141),
	.w5(32'h3a02ab3a),
	.w6(32'h3b24d8df),
	.w7(32'hbb991038),
	.w8(32'hbbc7592e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407a32),
	.w1(32'hbb7754b7),
	.w2(32'hbb9f59ee),
	.w3(32'h3b344367),
	.w4(32'h3c2260e5),
	.w5(32'hbb23ed98),
	.w6(32'hbbdc53a9),
	.w7(32'hbb4bff9c),
	.w8(32'h3bec6c39),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bfbcf),
	.w1(32'hbc22789a),
	.w2(32'hbb939a55),
	.w3(32'h3ac2fb10),
	.w4(32'hbc77c11b),
	.w5(32'hbc6f133a),
	.w6(32'hbb0e8cb1),
	.w7(32'h3aafd2cf),
	.w8(32'h3b7608c8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18c932),
	.w1(32'h3bd22d44),
	.w2(32'h3a908b7b),
	.w3(32'hbc906a35),
	.w4(32'h3c0f7d77),
	.w5(32'h3b172dee),
	.w6(32'hba4e1e9a),
	.w7(32'hbb8fc530),
	.w8(32'hba884286),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba334fe),
	.w1(32'h3a9417ea),
	.w2(32'hbbceba1a),
	.w3(32'h3becdf98),
	.w4(32'hbb1b0cbf),
	.w5(32'hbbdecc65),
	.w6(32'h3bde9ae8),
	.w7(32'h3b54e110),
	.w8(32'h3b7060b0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e168),
	.w1(32'h3c009382),
	.w2(32'hbb01bedb),
	.w3(32'hbbd4fd25),
	.w4(32'h3b064dcf),
	.w5(32'hbbe98d7a),
	.w6(32'h3c77034c),
	.w7(32'h3c215d81),
	.w8(32'h3c44a523),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f227),
	.w1(32'h3c839a2e),
	.w2(32'h3c95d6b3),
	.w3(32'hbb8d0b1a),
	.w4(32'h3cb6996d),
	.w5(32'h3d06d82d),
	.w6(32'hba198ce9),
	.w7(32'hbc12af01),
	.w8(32'hbc583f2f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945b9e),
	.w1(32'h3c08fae3),
	.w2(32'h3c1f048b),
	.w3(32'h3c845619),
	.w4(32'h3c239d26),
	.w5(32'h3c377008),
	.w6(32'h3c286b3b),
	.w7(32'h3b947b12),
	.w8(32'h3a320d1b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9176),
	.w1(32'hbbdc5cd7),
	.w2(32'hbbda3ccc),
	.w3(32'h3c36315d),
	.w4(32'hbc80e221),
	.w5(32'hbca3e9f0),
	.w6(32'hba3b5f00),
	.w7(32'h3bf1a30d),
	.w8(32'h3c820b41),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab677d),
	.w1(32'hbbfdd706),
	.w2(32'hbc503ed9),
	.w3(32'hbc9d5ff7),
	.w4(32'hbc0550cb),
	.w5(32'hbbfd70bf),
	.w6(32'hbb3c4ade),
	.w7(32'hbc137d53),
	.w8(32'h3b059a69),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9de637),
	.w1(32'h3aace0de),
	.w2(32'hbb89ce60),
	.w3(32'hb9f934fe),
	.w4(32'h3b9c1c19),
	.w5(32'h3c21cfa3),
	.w6(32'h3bcf95ad),
	.w7(32'hba35fb12),
	.w8(32'h39bd3dd5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f87cf),
	.w1(32'h3be8c1ea),
	.w2(32'h3c550544),
	.w3(32'h3b3e761b),
	.w4(32'h3cc1a5d9),
	.w5(32'h3d40c895),
	.w6(32'hbc1abbe8),
	.w7(32'hbc3660eb),
	.w8(32'hbb5473ba),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c900661),
	.w1(32'h3bbfac81),
	.w2(32'hbb3d22ee),
	.w3(32'h3d1d4f50),
	.w4(32'hbc4d021d),
	.w5(32'hbd0a24e2),
	.w6(32'h3c34531d),
	.w7(32'h3bfe097e),
	.w8(32'h3c663009),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc291265),
	.w1(32'h3b80ffeb),
	.w2(32'hbaec41a1),
	.w3(32'hbce04545),
	.w4(32'hb81b5e7c),
	.w5(32'hbbeb6a29),
	.w6(32'h39af55e4),
	.w7(32'hbbce2b8b),
	.w8(32'hbba1b3eb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34ec6c),
	.w1(32'h3b04608a),
	.w2(32'hbc08ddaa),
	.w3(32'hbbe7b7f2),
	.w4(32'h3cf3a283),
	.w5(32'h3d1129f0),
	.w6(32'hbcc1a6ec),
	.w7(32'hbd349ff3),
	.w8(32'hbd3b44aa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92100e),
	.w1(32'h3c3fdf68),
	.w2(32'h3c2c2dda),
	.w3(32'h3c78a755),
	.w4(32'h3c6d14ae),
	.w5(32'h3c6cf9a5),
	.w6(32'h3bee7904),
	.w7(32'h3ba1f032),
	.w8(32'h3a68269b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd35ca),
	.w1(32'h3c39cebc),
	.w2(32'h3c960cf0),
	.w3(32'h3c2967ef),
	.w4(32'h3c07dc95),
	.w5(32'h3ca25b36),
	.w6(32'h3988e33d),
	.w7(32'h3b63345c),
	.w8(32'h3b6ac0db),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfba52f),
	.w1(32'h3c5a547b),
	.w2(32'h3c9dc510),
	.w3(32'h3c430c14),
	.w4(32'h3c927108),
	.w5(32'h3cec9f8d),
	.w6(32'h3bdf8616),
	.w7(32'hbb0a8904),
	.w8(32'hbbd3527f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca176a),
	.w1(32'hbbdd0d03),
	.w2(32'hbbdd02af),
	.w3(32'h3c747a89),
	.w4(32'hbbbfb632),
	.w5(32'hbbd34bcc),
	.w6(32'hbb5ee554),
	.w7(32'hbc29ae41),
	.w8(32'hbb326133),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2d3e),
	.w1(32'h3928de24),
	.w2(32'hbae4dfbb),
	.w3(32'h3baa47fe),
	.w4(32'h3c0941b8),
	.w5(32'h3c37f7da),
	.w6(32'hbbdac6f5),
	.w7(32'hbabe89df),
	.w8(32'hbc1c8852),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1efb4b),
	.w1(32'h3976725b),
	.w2(32'hbbca64c1),
	.w3(32'h3c732300),
	.w4(32'h3bd036b9),
	.w5(32'hbb0a657b),
	.w6(32'hbb21b9dd),
	.w7(32'hbbaad9d5),
	.w8(32'hbaaae4b3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b421dc3),
	.w1(32'h3ba86be0),
	.w2(32'h3b538c73),
	.w3(32'h3bb9c526),
	.w4(32'h3b4beecb),
	.w5(32'h3adb337f),
	.w6(32'h3b361670),
	.w7(32'hbb19594e),
	.w8(32'h3bb9fda7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a067062),
	.w1(32'h3c65d8bb),
	.w2(32'h3c5d802c),
	.w3(32'h3b4361c4),
	.w4(32'h3c5de092),
	.w5(32'h3cd5df93),
	.w6(32'h3c0b1081),
	.w7(32'hbb7d32e0),
	.w8(32'hbb92def1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec1524),
	.w1(32'hba3cfc6c),
	.w2(32'h3c1cccdb),
	.w3(32'h3c962cab),
	.w4(32'h3c42f00d),
	.w5(32'h3cb07eae),
	.w6(32'hbb134baa),
	.w7(32'hbc2450aa),
	.w8(32'h38fadbf8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c700a94),
	.w1(32'h3c48f832),
	.w2(32'h3c245a78),
	.w3(32'h3c9fc269),
	.w4(32'h3c8a940c),
	.w5(32'h3c98a060),
	.w6(32'hbb7f7ef9),
	.w7(32'hb9ed0d2f),
	.w8(32'hbb8a06b4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb271135),
	.w1(32'hbb7f8821),
	.w2(32'hbb819492),
	.w3(32'h3b044035),
	.w4(32'h3b81b4f7),
	.w5(32'h3b31fcda),
	.w6(32'hbb4ad227),
	.w7(32'h3a835e26),
	.w8(32'h3b492599),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d2152),
	.w1(32'h39b44d5f),
	.w2(32'hbb0031b1),
	.w3(32'h3c21a035),
	.w4(32'h3bc1bd5f),
	.w5(32'h383eb1a4),
	.w6(32'hbbd26997),
	.w7(32'hbc0b41e9),
	.w8(32'hbc0af0ae),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c55e),
	.w1(32'h3bdf3b7f),
	.w2(32'h39a13eb7),
	.w3(32'h3a9b01e5),
	.w4(32'h3c1f4e7c),
	.w5(32'h3c2a3995),
	.w6(32'hbb64f67c),
	.w7(32'hbc057933),
	.w8(32'hbc142514),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81451f),
	.w1(32'h3ad2d106),
	.w2(32'hbba4b767),
	.w3(32'hbadf19ff),
	.w4(32'h3c10a2f2),
	.w5(32'hbbbdffec),
	.w6(32'h3b75d2ae),
	.w7(32'hbb73aaa2),
	.w8(32'hbbf62009),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9117),
	.w1(32'h3b241e6b),
	.w2(32'hbc41297d),
	.w3(32'hbc050a41),
	.w4(32'hbc8f6818),
	.w5(32'hbcf1ff99),
	.w6(32'h3c8b6702),
	.w7(32'h3bbee982),
	.w8(32'h3b42112f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c0697),
	.w1(32'h3bedb128),
	.w2(32'hbbf5a570),
	.w3(32'hbc82166b),
	.w4(32'hbc7d1296),
	.w5(32'hbd12b070),
	.w6(32'h3d004415),
	.w7(32'h3d1387ed),
	.w8(32'h3d282613),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b653f),
	.w1(32'hbb77a009),
	.w2(32'hba810b41),
	.w3(32'hbc331a87),
	.w4(32'h39eb66cb),
	.w5(32'h3ae3b90d),
	.w6(32'hbba994bb),
	.w7(32'hbb63cf4d),
	.w8(32'hbb9fd58f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b3da5),
	.w1(32'hbabab29e),
	.w2(32'hbbb20e2f),
	.w3(32'hbb837c77),
	.w4(32'hbbb76287),
	.w5(32'hbc22ecf8),
	.w6(32'h3b321d95),
	.w7(32'hbadc440c),
	.w8(32'hbb5311cf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce95fd),
	.w1(32'h3bcf1a6a),
	.w2(32'h3bee13c8),
	.w3(32'hbc2b5bfc),
	.w4(32'h3c0be31e),
	.w5(32'h3c3dcf33),
	.w6(32'h3a1350df),
	.w7(32'h3a7b170b),
	.w8(32'hbb8f02c3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c091),
	.w1(32'hbca6c9c4),
	.w2(32'hbd05a9cd),
	.w3(32'h3c359a98),
	.w4(32'hbca7034c),
	.w5(32'hbce9307d),
	.w6(32'hbc0f31b8),
	.w7(32'hbc681a41),
	.w8(32'hbc12fad3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1c841),
	.w1(32'hbb9d7b94),
	.w2(32'hbb8fda4a),
	.w3(32'hbcbe50cf),
	.w4(32'h3b91ff97),
	.w5(32'h3c51e118),
	.w6(32'hbc7eec9d),
	.w7(32'hbcbdbcdc),
	.w8(32'hbc9d96b0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d67f9),
	.w1(32'h3b63a3d5),
	.w2(32'h3bda52a6),
	.w3(32'h3bdc4bb6),
	.w4(32'h3ba2cb67),
	.w5(32'h3c20dd8e),
	.w6(32'hbba0ad9e),
	.w7(32'hbb94caa2),
	.w8(32'h3b7b3706),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c291641),
	.w1(32'h3c996be8),
	.w2(32'h3bf772f2),
	.w3(32'h3c923e35),
	.w4(32'h3cadd4ea),
	.w5(32'h3c736416),
	.w6(32'hbc015b34),
	.w7(32'h3bb160e8),
	.w8(32'h3b58f073),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c7777),
	.w1(32'h3ba489f8),
	.w2(32'hbc283f28),
	.w3(32'hbbd7b003),
	.w4(32'h3c17a88e),
	.w5(32'h3a660b8e),
	.w6(32'h3c5f665a),
	.w7(32'hbab7b415),
	.w8(32'hbb566e9c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d19a9),
	.w1(32'h3c5333ff),
	.w2(32'h3c2ada09),
	.w3(32'hbb892f13),
	.w4(32'h3bf77f4f),
	.w5(32'h3c317d37),
	.w6(32'h3b853c37),
	.w7(32'hb9861e88),
	.w8(32'hbb10eae3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd82b5),
	.w1(32'h3c768d02),
	.w2(32'h3c6fb4f7),
	.w3(32'h3b939a8f),
	.w4(32'h3c8b91a4),
	.w5(32'h3c8f69eb),
	.w6(32'h3bbe515f),
	.w7(32'hbafd7c29),
	.w8(32'h3c07bc9b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ccc78),
	.w1(32'h3b3a2611),
	.w2(32'hbbc6cac1),
	.w3(32'h3c496d09),
	.w4(32'h3bc2d2b3),
	.w5(32'hbbb2eb03),
	.w6(32'h3b462460),
	.w7(32'hbb1aa61d),
	.w8(32'h3b92c25b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39944201),
	.w1(32'h3b2cde0f),
	.w2(32'hbbb6d329),
	.w3(32'hb9a13261),
	.w4(32'h3b0f456f),
	.w5(32'h3b64ba48),
	.w6(32'hbba2d9cf),
	.w7(32'hbbf373ae),
	.w8(32'hbb241e5f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf43d31),
	.w1(32'h3b45a090),
	.w2(32'h3ba3fd6e),
	.w3(32'hbbaa6794),
	.w4(32'h3c81e27e),
	.w5(32'h3ce89f30),
	.w6(32'hbc54d394),
	.w7(32'hbc1028de),
	.w8(32'hbc1417cb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd868cc),
	.w1(32'h3a13bf04),
	.w2(32'hbbbde0e0),
	.w3(32'h3c4f1925),
	.w4(32'h3c3c74da),
	.w5(32'h3c4f8c4d),
	.w6(32'hbb9eea9a),
	.w7(32'hbb96eab4),
	.w8(32'hbaaaf1f1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7f3c3),
	.w1(32'h3ba29fca),
	.w2(32'h3b1d997a),
	.w3(32'hbb8b1a90),
	.w4(32'h3c5d5e89),
	.w5(32'h3c905a5e),
	.w6(32'hbbeec2b5),
	.w7(32'hbb82b2fd),
	.w8(32'h3a3c70f1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb247156),
	.w1(32'hbb629082),
	.w2(32'hbb86164c),
	.w3(32'h3bb810ee),
	.w4(32'h3c24f0b0),
	.w5(32'h3c44a544),
	.w6(32'h374cc446),
	.w7(32'h3b542b5a),
	.w8(32'h3ba85e6b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f301),
	.w1(32'hbaf99ba8),
	.w2(32'h3c22e6ca),
	.w3(32'h3abfad63),
	.w4(32'h3c6eaa3e),
	.w5(32'h3cee840a),
	.w6(32'hbc8457f7),
	.w7(32'hbc087ad8),
	.w8(32'hbb1295e2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb2d6),
	.w1(32'h3c174d59),
	.w2(32'h3c00ed9e),
	.w3(32'h3c3d44d8),
	.w4(32'h3c34582c),
	.w5(32'h3c3720ad),
	.w6(32'h3c046a7f),
	.w7(32'hbb1c02d4),
	.w8(32'hbb98aadf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8af4b1),
	.w1(32'h3c01137a),
	.w2(32'h3c306d7f),
	.w3(32'h3b535a6f),
	.w4(32'h3c5c9c5c),
	.w5(32'h3c7e8d3d),
	.w6(32'h39182842),
	.w7(32'h39eab579),
	.w8(32'h3c1436b5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a34e4),
	.w1(32'hbbe40339),
	.w2(32'hbc30dcbe),
	.w3(32'h3c12be5e),
	.w4(32'h3bd922ad),
	.w5(32'hbba4f191),
	.w6(32'hbb598d89),
	.w7(32'hbba1da89),
	.w8(32'hbc1869eb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e617c),
	.w1(32'hbbba1504),
	.w2(32'hbc7aaf8f),
	.w3(32'hbb5d52cc),
	.w4(32'hbb669053),
	.w5(32'hbbd6a99b),
	.w6(32'hba65d9e2),
	.w7(32'hbc3dabc2),
	.w8(32'hbb8e6601),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80cba8),
	.w1(32'h3c992507),
	.w2(32'h3c68f465),
	.w3(32'hbc3ceafe),
	.w4(32'h3c4443c4),
	.w5(32'h3b76e1b1),
	.w6(32'h3b739cd0),
	.w7(32'h3ba88536),
	.w8(32'hbb540833),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda8256),
	.w1(32'h37f417d7),
	.w2(32'hbc74bfd9),
	.w3(32'h3ba31dce),
	.w4(32'hbb75bffd),
	.w5(32'hbbef884e),
	.w6(32'hbc3bef58),
	.w7(32'hbc8bf551),
	.w8(32'hbc216ed3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94f7fe),
	.w1(32'h3ba21661),
	.w2(32'h3bd6d79a),
	.w3(32'hbc51ca3a),
	.w4(32'h3bb2ea96),
	.w5(32'h3c16a0b4),
	.w6(32'h3b24c0f4),
	.w7(32'h3aea31ec),
	.w8(32'hb80144d3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad65307),
	.w1(32'h3ba7394a),
	.w2(32'hbbc0adcd),
	.w3(32'h3c3e3c88),
	.w4(32'h3cbbd8bd),
	.w5(32'h3c6b817b),
	.w6(32'h3bfc5490),
	.w7(32'h3bcbba66),
	.w8(32'h3a1a5d75),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe94000),
	.w1(32'hbb382cf7),
	.w2(32'hbae307b9),
	.w3(32'h3bf8adde),
	.w4(32'h3c11b181),
	.w5(32'h3c1ceaf7),
	.w6(32'hba8a0d0f),
	.w7(32'hbba89a9a),
	.w8(32'hbbb4eff5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd902ea),
	.w1(32'h3c3e6837),
	.w2(32'h3c82c2c6),
	.w3(32'h3bd8e80e),
	.w4(32'h3c7cabfe),
	.w5(32'h3c8fcbfe),
	.w6(32'h3b924a34),
	.w7(32'h3b2e2af5),
	.w8(32'hbb8a5ca2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1122ac),
	.w1(32'h3c111b55),
	.w2(32'h3b08d010),
	.w3(32'hbacd2a2e),
	.w4(32'h3c93d346),
	.w5(32'h3cb88815),
	.w6(32'h3b260b38),
	.w7(32'h3aaeb7bc),
	.w8(32'h3a98399a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a1bd2),
	.w1(32'hbb53f4f5),
	.w2(32'hbbac5332),
	.w3(32'h3bfcfd81),
	.w4(32'h3bbd8702),
	.w5(32'hba73d6a4),
	.w6(32'h3ab4ac32),
	.w7(32'hbbd6299b),
	.w8(32'h3ac548ca),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1f5ce),
	.w1(32'hba9fbe12),
	.w2(32'h39bb9f17),
	.w3(32'h3b2a4da3),
	.w4(32'h39fcae9a),
	.w5(32'h3a0f8da4),
	.w6(32'h3b664895),
	.w7(32'h3a77c16c),
	.w8(32'h3b63cfd3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e32a8),
	.w1(32'h3b3fd66a),
	.w2(32'h3a8ebd10),
	.w3(32'hba9b632b),
	.w4(32'h3c20750a),
	.w5(32'h3c3a6ea4),
	.w6(32'hbb86809c),
	.w7(32'hbbe473fb),
	.w8(32'hbc0c2c6d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d7c5),
	.w1(32'h3c0cfbc6),
	.w2(32'h3c481da5),
	.w3(32'h3c1501fc),
	.w4(32'h3c5fc6af),
	.w5(32'h3d14c7a0),
	.w6(32'hbad6a71f),
	.w7(32'hbb8aef29),
	.w8(32'hbc08778d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16da88),
	.w1(32'hbb61e25e),
	.w2(32'hbb2256a2),
	.w3(32'h3ca26d96),
	.w4(32'hba18c268),
	.w5(32'hbb12a9f5),
	.w6(32'hbb75c18d),
	.w7(32'hbb6238af),
	.w8(32'h3b39923c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba881421),
	.w1(32'h3bb3f7e3),
	.w2(32'hbb36e803),
	.w3(32'hbb7559c8),
	.w4(32'h3bbe7199),
	.w5(32'h3c2744a4),
	.w6(32'hbc48503a),
	.w7(32'hbc46af3f),
	.w8(32'hbc11d9c2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7e2f),
	.w1(32'h3c20a8a3),
	.w2(32'h3c84ca1a),
	.w3(32'h3a8ca6d2),
	.w4(32'h3c8c17c0),
	.w5(32'h3cfe852c),
	.w6(32'h3b89aadc),
	.w7(32'hbb06930a),
	.w8(32'hbba8e784),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdba61),
	.w1(32'h3c5bebd1),
	.w2(32'h3ca1ece5),
	.w3(32'h3ca1eda8),
	.w4(32'h3d043fc8),
	.w5(32'h3d5cd9d3),
	.w6(32'hba37f147),
	.w7(32'hbc1002df),
	.w8(32'hbbd95db3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf102b7),
	.w1(32'hbc4529bd),
	.w2(32'hbc9a5f22),
	.w3(32'h3cc7d35d),
	.w4(32'hbc41592e),
	.w5(32'hbc6bc8cf),
	.w6(32'hbbca6535),
	.w7(32'hbc5b5d5c),
	.w8(32'hbb84bca8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb81377),
	.w1(32'hbca7ad89),
	.w2(32'hbd14f81b),
	.w3(32'hbc806467),
	.w4(32'hbc854016),
	.w5(32'hbcee1824),
	.w6(32'hbc473a22),
	.w7(32'hbcd647a5),
	.w8(32'hbc8aec35),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced1a96),
	.w1(32'hbc6ed471),
	.w2(32'hbc801797),
	.w3(32'hbca70461),
	.w4(32'hbcdc2195),
	.w5(32'hbd0184e1),
	.w6(32'h3c58df47),
	.w7(32'h3c985b87),
	.w8(32'h3c9366cd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d60f),
	.w1(32'h3bc89ce0),
	.w2(32'h3b82f874),
	.w3(32'hbc126775),
	.w4(32'h3c2611ec),
	.w5(32'hb996dfed),
	.w6(32'h3982084b),
	.w7(32'hba595751),
	.w8(32'h3ab9988e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854bdd),
	.w1(32'h3bc3d7e5),
	.w2(32'h3c420eb1),
	.w3(32'hbb93bef4),
	.w4(32'h3c618549),
	.w5(32'h3c9b3855),
	.w6(32'hbba04fac),
	.w7(32'h3a426a65),
	.w8(32'hbb8ae75b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55dc14),
	.w1(32'hbbb9dfc2),
	.w2(32'h3b746685),
	.w3(32'h3c5c526c),
	.w4(32'h3c400892),
	.w5(32'h3c846d0d),
	.w6(32'hbca277b4),
	.w7(32'h3b7add62),
	.w8(32'h3bfef330),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1143e5),
	.w1(32'h3c0645c9),
	.w2(32'h3b151b50),
	.w3(32'h3bd4e180),
	.w4(32'h3c210f3a),
	.w5(32'h3b98a2ea),
	.w6(32'hbb883d2d),
	.w7(32'hbc1eef7f),
	.w8(32'hb9fb8ac2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d253c),
	.w1(32'h3c04eb3d),
	.w2(32'h3ac41da5),
	.w3(32'h3be38fa4),
	.w4(32'h3cbf6360),
	.w5(32'h3ca33b6b),
	.w6(32'h3a827860),
	.w7(32'hbb4f8627),
	.w8(32'hbc030469),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9f57e),
	.w1(32'h3a39645b),
	.w2(32'hbaa38861),
	.w3(32'h3c4e1b9c),
	.w4(32'hbae160cf),
	.w5(32'h3ba8af25),
	.w6(32'h3b889660),
	.w7(32'hbb252ee8),
	.w8(32'h3a6a7e33),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaee23c),
	.w1(32'hbb96f674),
	.w2(32'hbc54f1a8),
	.w3(32'h3b961494),
	.w4(32'hbc5be521),
	.w5(32'hbccf9232),
	.w6(32'h3c76a7dd),
	.w7(32'h3bed0fe4),
	.w8(32'h3c1536ea),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3fe1),
	.w1(32'h3ab80d1d),
	.w2(32'h3a373a9d),
	.w3(32'hbc647af1),
	.w4(32'h3b7d16c4),
	.w5(32'h3af116bf),
	.w6(32'h3a747d96),
	.w7(32'h3b6f5500),
	.w8(32'h3b7cfc8c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79166f),
	.w1(32'h3b8672ca),
	.w2(32'h3c0d62f8),
	.w3(32'h3bd0a67e),
	.w4(32'h3b743898),
	.w5(32'h3c4b8a76),
	.w6(32'h3b4926ab),
	.w7(32'hb93ab06a),
	.w8(32'h3abb03ea),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ec1d4),
	.w1(32'hbacdbcc1),
	.w2(32'hbba028a8),
	.w3(32'h3c1441b8),
	.w4(32'hbb1b64b1),
	.w5(32'hbbdd36d5),
	.w6(32'h3a3746ca),
	.w7(32'hbb1bf08e),
	.w8(32'hbbc57f3a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfae1e0),
	.w1(32'h3cc5d9db),
	.w2(32'h3cf72700),
	.w3(32'hbc03e5d9),
	.w4(32'h3c89952c),
	.w5(32'h3d1b2b66),
	.w6(32'h3ca02ff7),
	.w7(32'h3cdf0ef4),
	.w8(32'h3ca1c5a7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb22115),
	.w1(32'h3b746564),
	.w2(32'h39f41592),
	.w3(32'h3c959801),
	.w4(32'h3c6342aa),
	.w5(32'h3ba12430),
	.w6(32'h398c97de),
	.w7(32'hbb49a0d0),
	.w8(32'hbbd06230),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf68d),
	.w1(32'hbb6b61c5),
	.w2(32'hbbc386a0),
	.w3(32'h3b330dd5),
	.w4(32'hbb90df92),
	.w5(32'hbb0e606e),
	.w6(32'hb96bef29),
	.w7(32'hbb90de6a),
	.w8(32'hbb2e6024),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ac05),
	.w1(32'hbb431530),
	.w2(32'hbb627341),
	.w3(32'hbb8d6c9d),
	.w4(32'hbacdd241),
	.w5(32'hbb69e645),
	.w6(32'hbb483def),
	.w7(32'hb9ae1729),
	.w8(32'h39c67c2c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed5cbe),
	.w1(32'hbabbe39d),
	.w2(32'hbb5e5908),
	.w3(32'hba391f68),
	.w4(32'hbbb8349a),
	.w5(32'hbc3b3f60),
	.w6(32'h3b5a60cd),
	.w7(32'hbb846d47),
	.w8(32'h3baec2ff),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2c292),
	.w1(32'h3c87fbe3),
	.w2(32'h3c94444f),
	.w3(32'hbbbf5241),
	.w4(32'h3c8142cc),
	.w5(32'h3c5a3ddd),
	.w6(32'h3c8038cf),
	.w7(32'h3c8e77cb),
	.w8(32'h3c807bd7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ca59b),
	.w1(32'hbb63091e),
	.w2(32'h3c287e7a),
	.w3(32'h3c1f704d),
	.w4(32'h3aa7058a),
	.w5(32'h3bba1a66),
	.w6(32'h3a8389d1),
	.w7(32'h3b8b6be8),
	.w8(32'h3b5daa03),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad64692),
	.w1(32'h3c06d03f),
	.w2(32'h3ba1ef42),
	.w3(32'h3a01d271),
	.w4(32'h3c44fa97),
	.w5(32'h3c1ec3a5),
	.w6(32'hbaf900a6),
	.w7(32'hbaf45784),
	.w8(32'hbb0f4476),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30bc37),
	.w1(32'hbb6a7d1c),
	.w2(32'h3b163336),
	.w3(32'h3bbfa39b),
	.w4(32'h3c07c18a),
	.w5(32'h3c0b9fcc),
	.w6(32'hbbbab777),
	.w7(32'hbbc675bd),
	.w8(32'h3a208926),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d0fc3),
	.w1(32'h3a0b5f0b),
	.w2(32'h3c092402),
	.w3(32'h3c4ef22c),
	.w4(32'h3a923105),
	.w5(32'h3ad5d681),
	.w6(32'hbb204e3b),
	.w7(32'h3bc4712c),
	.w8(32'h3a9b5f54),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9de335),
	.w1(32'hbbb72a8d),
	.w2(32'hbc0b7251),
	.w3(32'hbc6ae57a),
	.w4(32'h3ab91979),
	.w5(32'hbb574933),
	.w6(32'hbbaaec78),
	.w7(32'hbbbd5d52),
	.w8(32'hbbde9bdb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaec5b),
	.w1(32'h3ca7d443),
	.w2(32'h3cb8e209),
	.w3(32'hbb5204be),
	.w4(32'h3c27fbe3),
	.w5(32'h3c91af87),
	.w6(32'h3c6d019b),
	.w7(32'h3c98e190),
	.w8(32'h3c35a2bf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5762c3),
	.w1(32'h3c5321bd),
	.w2(32'h3c17bfe5),
	.w3(32'h3c0be65a),
	.w4(32'h3cb57b3b),
	.w5(32'h3c2b8f65),
	.w6(32'h3bbf7430),
	.w7(32'h3a908643),
	.w8(32'h3b98f0a8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24104b),
	.w1(32'h3acec5aa),
	.w2(32'h3c0d084c),
	.w3(32'h3b0e1545),
	.w4(32'h3c2d7599),
	.w5(32'h3c7349cc),
	.w6(32'h39512f91),
	.w7(32'h3a87b06e),
	.w8(32'hb6ed70e0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5efad),
	.w1(32'h3b2f9d3c),
	.w2(32'hbb9dd95b),
	.w3(32'h3bb5c063),
	.w4(32'hb8e819d4),
	.w5(32'hbb81283f),
	.w6(32'h3951ceb2),
	.w7(32'hba6dde23),
	.w8(32'h3a66e532),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc34be),
	.w1(32'h3b8f9ba8),
	.w2(32'h3999d252),
	.w3(32'h39014768),
	.w4(32'h3bf1d1d9),
	.w5(32'h394117c9),
	.w6(32'hbbc10354),
	.w7(32'hbc0ce52d),
	.w8(32'hba9b0ed3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule