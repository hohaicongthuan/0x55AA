module layer_10_featuremap_498(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd005e),
	.w1(32'hbb0e3aac),
	.w2(32'hb90cab83),
	.w3(32'hba47425d),
	.w4(32'hb9be6c58),
	.w5(32'hb8964977),
	.w6(32'h3b033596),
	.w7(32'hbb4a24c8),
	.w8(32'hbb136ff5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd049c),
	.w1(32'hbb6f7ed2),
	.w2(32'hbbab723a),
	.w3(32'hbc11de04),
	.w4(32'h3b0dd8ac),
	.w5(32'hbbaf5a4f),
	.w6(32'hbc06d0c7),
	.w7(32'h3b6e6314),
	.w8(32'hbaa5f780),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b778a87),
	.w1(32'hbb8922cc),
	.w2(32'h3bb65823),
	.w3(32'hbaa64664),
	.w4(32'hba1981d1),
	.w5(32'hba9bc332),
	.w6(32'hb8dc4b47),
	.w7(32'h3b0a0a75),
	.w8(32'hbbbb0811),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96256d6),
	.w1(32'hbac5ebd7),
	.w2(32'h3bc7defd),
	.w3(32'h3b5ef577),
	.w4(32'h3c329b97),
	.w5(32'hbb8c3bde),
	.w6(32'h3aaa377c),
	.w7(32'hba79f6e2),
	.w8(32'h3af3f04a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa74b6),
	.w1(32'h3a8df627),
	.w2(32'hbaa46800),
	.w3(32'hb95957d5),
	.w4(32'hbadaf30f),
	.w5(32'hb8a75d6d),
	.w6(32'hb99b3bc9),
	.w7(32'hbb913fc7),
	.w8(32'hbbacc705),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb181fab),
	.w1(32'hbb6e3e67),
	.w2(32'hbb66724e),
	.w3(32'hba706c40),
	.w4(32'hbb7f217c),
	.w5(32'hb9f22fdb),
	.w6(32'hbba34481),
	.w7(32'hbb1c4bc5),
	.w8(32'h3afac198),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc157861),
	.w1(32'h383bb122),
	.w2(32'h3b9c115a),
	.w3(32'hbb59481a),
	.w4(32'h3aa97b58),
	.w5(32'h3b2032dc),
	.w6(32'h3bbea2cc),
	.w7(32'hba44c718),
	.w8(32'hbba22673),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8ecf5),
	.w1(32'h3ba39235),
	.w2(32'h3c0f25c4),
	.w3(32'h3cbae81e),
	.w4(32'h3c3830f5),
	.w5(32'h3b7bafda),
	.w6(32'h3c868da0),
	.w7(32'h3c916789),
	.w8(32'h3c0a694b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5da3ea),
	.w1(32'h3a9431d6),
	.w2(32'h3badd8d3),
	.w3(32'hbb7d9cff),
	.w4(32'h3b6d8d8e),
	.w5(32'hbb280d79),
	.w6(32'h3857efea),
	.w7(32'h3ae641e0),
	.w8(32'h3a6357ed),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51173a),
	.w1(32'h3c08ae1b),
	.w2(32'h3ab90d09),
	.w3(32'hbbd1923d),
	.w4(32'h3aba32bc),
	.w5(32'hbbc404f5),
	.w6(32'h392d7182),
	.w7(32'h3acad23a),
	.w8(32'hbb0ce2b5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ab8e2),
	.w1(32'h3b84334d),
	.w2(32'h3b872977),
	.w3(32'h3abf26d7),
	.w4(32'hbb012d11),
	.w5(32'hbbbcae5e),
	.w6(32'hbb593199),
	.w7(32'h3a6d17b7),
	.w8(32'hba83254d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f5c7a),
	.w1(32'hbb8b34a0),
	.w2(32'h3b8a32fe),
	.w3(32'h39b7d199),
	.w4(32'hbb997985),
	.w5(32'h3b64224f),
	.w6(32'hbab8ba54),
	.w7(32'hbb98659a),
	.w8(32'hbb2e0006),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67aeb8),
	.w1(32'h3c222927),
	.w2(32'h3bb5e611),
	.w3(32'h3b88b90b),
	.w4(32'h3c32bb53),
	.w5(32'hbb991710),
	.w6(32'h3af5faeb),
	.w7(32'h3c0403dc),
	.w8(32'h3b902529),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a373927),
	.w1(32'h3bc6bba9),
	.w2(32'h3b3972f4),
	.w3(32'hbbad8b11),
	.w4(32'h3c044894),
	.w5(32'h3b43172b),
	.w6(32'hbbbd1571),
	.w7(32'h3bb26e56),
	.w8(32'h3a9aa300),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011e50),
	.w1(32'hbb02ce3a),
	.w2(32'h3bce22bd),
	.w3(32'h3b954d58),
	.w4(32'hbb9d69ad),
	.w5(32'hba8c9da7),
	.w6(32'h3a63a73f),
	.w7(32'hbbcb65b7),
	.w8(32'hbb0a04e8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207c23),
	.w1(32'hba89250d),
	.w2(32'h3a913e55),
	.w3(32'h3c316378),
	.w4(32'hbb4d3e08),
	.w5(32'h3b2cf5ef),
	.w6(32'h3c2f7901),
	.w7(32'h3b94580a),
	.w8(32'h3c0e4cd9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b058d9a),
	.w1(32'hba6830d7),
	.w2(32'h3ba5fdde),
	.w3(32'h3b8d4535),
	.w4(32'hbb45b82f),
	.w5(32'hbad85115),
	.w6(32'h3b42d868),
	.w7(32'hbaf57b61),
	.w8(32'hbb6cb312),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8a570),
	.w1(32'h3cbd19de),
	.w2(32'h3ccdaa19),
	.w3(32'h3d03f0da),
	.w4(32'h3cd33516),
	.w5(32'h3c84f903),
	.w6(32'h3cab03f3),
	.w7(32'h3cce01d5),
	.w8(32'h3c670dda),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ecab6),
	.w1(32'h3c03c2fb),
	.w2(32'h3c1e314c),
	.w3(32'h3c358ac8),
	.w4(32'h3c4f8f30),
	.w5(32'h3b51006c),
	.w6(32'h3c4b5070),
	.w7(32'h3c0b5bb4),
	.w8(32'h3acdd380),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6fc50),
	.w1(32'h3ab73b28),
	.w2(32'h3c26d1fb),
	.w3(32'h3ab314bb),
	.w4(32'h3b030e2b),
	.w5(32'h3b15333a),
	.w6(32'hbb6cafe4),
	.w7(32'h3b06814c),
	.w8(32'h3bd59924),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a396fa5),
	.w1(32'h3ad3eae4),
	.w2(32'hba806b8b),
	.w3(32'h39ce0020),
	.w4(32'h39224cb9),
	.w5(32'hbad323fb),
	.w6(32'h3a433a63),
	.w7(32'h3a924176),
	.w8(32'hb91ef737),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c161),
	.w1(32'hbb7e490e),
	.w2(32'hbbe0587c),
	.w3(32'h3a803971),
	.w4(32'hbbfe8397),
	.w5(32'h3a828c44),
	.w6(32'h3b615979),
	.w7(32'hbb02c244),
	.w8(32'h3a9987b2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc62a5),
	.w1(32'h3cd9846f),
	.w2(32'h3d106a07),
	.w3(32'h3cf00d58),
	.w4(32'h3cae79b7),
	.w5(32'h3c8a9227),
	.w6(32'h3d0169eb),
	.w7(32'h3cccce30),
	.w8(32'h3cad9b31),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6957f),
	.w1(32'hbbc2d136),
	.w2(32'hbc11b43a),
	.w3(32'hbbd1acc8),
	.w4(32'hbc18199d),
	.w5(32'hbc106d8a),
	.w6(32'hbbbb0cc9),
	.w7(32'hbb8d74c0),
	.w8(32'hbb8aa12d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8958ce4),
	.w1(32'hbbc901e3),
	.w2(32'hbc3247f7),
	.w3(32'hbc165e43),
	.w4(32'hbbd66c55),
	.w5(32'hbc055ac2),
	.w6(32'h3a91f633),
	.w7(32'h3b9f5016),
	.w8(32'h3bb3638d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7291a0),
	.w1(32'hbbe19a28),
	.w2(32'hbbb4df94),
	.w3(32'h3b9c9dd5),
	.w4(32'h390c696e),
	.w5(32'h3c410dab),
	.w6(32'hbb43d471),
	.w7(32'h3b128f0d),
	.w8(32'h3b9ca1fd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ada1),
	.w1(32'hbb51d194),
	.w2(32'hbb989a2d),
	.w3(32'hba749047),
	.w4(32'hbbabe4b8),
	.w5(32'hbb662849),
	.w6(32'h3bb0aeeb),
	.w7(32'hbb882f96),
	.w8(32'hbbc33982),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf3f82),
	.w1(32'hbba239c1),
	.w2(32'hbbbbf1ff),
	.w3(32'hbbb59a96),
	.w4(32'hbbff9cca),
	.w5(32'hbb933893),
	.w6(32'hbb485532),
	.w7(32'hba7b489d),
	.w8(32'h3bc98b24),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24b93b),
	.w1(32'h3b34bf41),
	.w2(32'h3b64b9c5),
	.w3(32'hba8f50ad),
	.w4(32'hbab4a9c2),
	.w5(32'hbc16e0f7),
	.w6(32'hb9a8686a),
	.w7(32'hbc00974c),
	.w8(32'hbb1e894c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf70c1),
	.w1(32'hbb804854),
	.w2(32'hbbce8a27),
	.w3(32'hbbff6d49),
	.w4(32'hbc4914eb),
	.w5(32'hbb64eb1a),
	.w6(32'hbc307919),
	.w7(32'hbbffdfae),
	.w8(32'hbc04df4c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e8499),
	.w1(32'h3a5eeed5),
	.w2(32'h3b9102c8),
	.w3(32'hba205583),
	.w4(32'hb9b34798),
	.w5(32'h3936adb7),
	.w6(32'hbb924eec),
	.w7(32'h3830f4d9),
	.w8(32'hbb313f6f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7557e4),
	.w1(32'hbad7dfff),
	.w2(32'h3a7b12d6),
	.w3(32'h39d78ba0),
	.w4(32'hbb498928),
	.w5(32'hbbcd2830),
	.w6(32'hbb258f43),
	.w7(32'hba386869),
	.w8(32'hba98afdd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae17ea),
	.w1(32'hbb6bc00d),
	.w2(32'hbba01b3d),
	.w3(32'hba2e32dc),
	.w4(32'hbaa2ffc2),
	.w5(32'hbb920ac2),
	.w6(32'h38a1e41f),
	.w7(32'h3923b1a9),
	.w8(32'h3b04bc1b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64ab9e),
	.w1(32'hbb1ac822),
	.w2(32'hbb316dce),
	.w3(32'hbaf13a9d),
	.w4(32'hbb3f9071),
	.w5(32'hbb924ae7),
	.w6(32'hbb103c56),
	.w7(32'h3a8b0982),
	.w8(32'hb8ae88c2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399376f2),
	.w1(32'hbb906dbb),
	.w2(32'hbc717e22),
	.w3(32'hba69301d),
	.w4(32'h3abfc3d4),
	.w5(32'hb99b762b),
	.w6(32'hb9b20757),
	.w7(32'h3bf1da73),
	.w8(32'h3c240256),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbfa63),
	.w1(32'hbb6b174a),
	.w2(32'h3a715080),
	.w3(32'h3b72f202),
	.w4(32'h3bce44f5),
	.w5(32'h3bb3f4a0),
	.w6(32'h3bec335c),
	.w7(32'h3a9091a8),
	.w8(32'h3a301d46),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a3fd),
	.w1(32'h3c6d94a9),
	.w2(32'h3c58e29c),
	.w3(32'h3bae58ec),
	.w4(32'h3c5f9123),
	.w5(32'h3a781d85),
	.w6(32'h3c0af550),
	.w7(32'h3c5e3915),
	.w8(32'h3c191d37),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ab3a1),
	.w1(32'hbca6cdea),
	.w2(32'hbc7775d6),
	.w3(32'hbcb14cd0),
	.w4(32'hbcb7c152),
	.w5(32'hbca31939),
	.w6(32'hbc617485),
	.w7(32'hbc47c469),
	.w8(32'hbbe106a5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257731),
	.w1(32'hbc7683db),
	.w2(32'hbc599125),
	.w3(32'hbc9d251d),
	.w4(32'hbc8dbb04),
	.w5(32'hbc5884eb),
	.w6(32'hbca6aac2),
	.w7(32'hbc474d2e),
	.w8(32'hbace2156),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc173),
	.w1(32'hbc1a41d6),
	.w2(32'hbbaf4374),
	.w3(32'hbbdca111),
	.w4(32'hbab798d5),
	.w5(32'hbbc0530f),
	.w6(32'hbb303edd),
	.w7(32'hbb1016c0),
	.w8(32'h3ac7e070),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0de0b3),
	.w1(32'h3b83f850),
	.w2(32'hba292ee8),
	.w3(32'hbb72f863),
	.w4(32'hbaea825d),
	.w5(32'h3b595379),
	.w6(32'hbbc7e841),
	.w7(32'hbbd3e2b1),
	.w8(32'h397076ff),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85ed06),
	.w1(32'h3a9689a6),
	.w2(32'h3b0c610c),
	.w3(32'h3b85cce3),
	.w4(32'h3a5b36cd),
	.w5(32'h3aaabd67),
	.w6(32'h39c6b9c0),
	.w7(32'hbb6b5ecc),
	.w8(32'hbb676a5a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97c47a),
	.w1(32'h391848fc),
	.w2(32'h3b6c4dee),
	.w3(32'hbb0b2cf9),
	.w4(32'h3b4372ab),
	.w5(32'hbc08c0aa),
	.w6(32'hbb1eed61),
	.w7(32'hbbbd8a49),
	.w8(32'hbbe16d15),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ce9d1),
	.w1(32'hb9e48411),
	.w2(32'hbb9c921d),
	.w3(32'h3bc083b8),
	.w4(32'h3b95de77),
	.w5(32'h3ba297e8),
	.w6(32'h3aa0a640),
	.w7(32'h3be20584),
	.w8(32'h3b8de147),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac787f1),
	.w1(32'hba0dcda2),
	.w2(32'hbb8cfd40),
	.w3(32'hbb30da60),
	.w4(32'hbb7b0727),
	.w5(32'hbbbab93f),
	.w6(32'hbb46564c),
	.w7(32'hbbb4fd18),
	.w8(32'hbb8faca1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3999d),
	.w1(32'hbb4b0f4c),
	.w2(32'hbc13a8ab),
	.w3(32'hbbc701f5),
	.w4(32'hbc2ef668),
	.w5(32'hbae3f896),
	.w6(32'hbb05323a),
	.w7(32'hbba20d65),
	.w8(32'hba8ed94e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36d2b1),
	.w1(32'h3b74bbcd),
	.w2(32'h3ba48089),
	.w3(32'h3b81750b),
	.w4(32'h3adaa691),
	.w5(32'hbc0767a5),
	.w6(32'h3c3b8499),
	.w7(32'h3ba338ea),
	.w8(32'h3aed59d0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea421b),
	.w1(32'h3d155ff1),
	.w2(32'h3cf46d25),
	.w3(32'h3cfa3528),
	.w4(32'h3d204091),
	.w5(32'h3c8ee915),
	.w6(32'h3ced1f67),
	.w7(32'h3d10963e),
	.w8(32'h3ca6ecca),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad15438),
	.w1(32'hbaa90b07),
	.w2(32'h3b58d41a),
	.w3(32'hbad2ec47),
	.w4(32'hbacb979b),
	.w5(32'h3b8cd620),
	.w6(32'hbac32c5b),
	.w7(32'hbb880a6f),
	.w8(32'h3a93b7f2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae56ddf),
	.w1(32'hbaf3dee5),
	.w2(32'h3a712e0b),
	.w3(32'h3c115e3d),
	.w4(32'hbb975a83),
	.w5(32'h3ba5e2a4),
	.w6(32'h3bb07248),
	.w7(32'hbaf0fc65),
	.w8(32'h3b3c74cc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc17e2c),
	.w1(32'hba0e4794),
	.w2(32'h3a7ccca1),
	.w3(32'h3c2c4515),
	.w4(32'hbb0a887f),
	.w5(32'hbb83661c),
	.w6(32'h3ac0fb33),
	.w7(32'hba99ea05),
	.w8(32'hba430615),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1f6b8),
	.w1(32'h3aa699ce),
	.w2(32'hbb0b7c7f),
	.w3(32'h3a060ab4),
	.w4(32'h3ac2c7fb),
	.w5(32'hb9eedc3a),
	.w6(32'h3beb1322),
	.w7(32'h3be00bd3),
	.w8(32'h3b5158a8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bcfc4),
	.w1(32'hbb5c030c),
	.w2(32'hbb86684d),
	.w3(32'hba39187e),
	.w4(32'hba88f0e8),
	.w5(32'hbbb569a4),
	.w6(32'hb908af30),
	.w7(32'h39f9fe75),
	.w8(32'h3a92c90f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29b971),
	.w1(32'h3c04a30e),
	.w2(32'h3b6dae5f),
	.w3(32'h3c80f3b3),
	.w4(32'h3c87e953),
	.w5(32'h3aa83f18),
	.w6(32'h3c91c1a6),
	.w7(32'h3cbe93c9),
	.w8(32'h3c940288),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcede7),
	.w1(32'h3ba478fe),
	.w2(32'h3b5e8be7),
	.w3(32'hbb5cf67f),
	.w4(32'h3ba32577),
	.w5(32'hb98f4fbd),
	.w6(32'h3ad9cecf),
	.w7(32'h3abf5898),
	.w8(32'h3b6165d1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70a15d),
	.w1(32'h3bbd3835),
	.w2(32'hba990f01),
	.w3(32'hbbb3daf9),
	.w4(32'h3c1f56cd),
	.w5(32'hbc1092ab),
	.w6(32'hbbda6c5f),
	.w7(32'h3c05cb7b),
	.w8(32'h3b04cc65),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8d77c),
	.w1(32'hb9c1c139),
	.w2(32'h3ad262d6),
	.w3(32'hbba5ac05),
	.w4(32'hbb591426),
	.w5(32'h3aab3b77),
	.w6(32'hbafaf824),
	.w7(32'hbb9298d3),
	.w8(32'hbb1a12e8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd6953),
	.w1(32'hbb84494b),
	.w2(32'hbb6ad2c6),
	.w3(32'h3aea4704),
	.w4(32'hba198f4f),
	.w5(32'h3ba029f6),
	.w6(32'hbb0b160c),
	.w7(32'h3a720618),
	.w8(32'hbab6cd6a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7e1e3),
	.w1(32'hbbffb399),
	.w2(32'hbb18f091),
	.w3(32'hbb8a6a00),
	.w4(32'h39b45fcb),
	.w5(32'hbab84b66),
	.w6(32'h39f88d60),
	.w7(32'hbb2ec870),
	.w8(32'hbb14ace4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970429d),
	.w1(32'hbb1da695),
	.w2(32'h394b9282),
	.w3(32'hba0f0ee2),
	.w4(32'h3a2f5da3),
	.w5(32'hbba0738e),
	.w6(32'hbac7ba78),
	.w7(32'h38ad7893),
	.w8(32'h392c0954),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24cd54),
	.w1(32'h3bc3fd1e),
	.w2(32'h3b98b3e7),
	.w3(32'h3c1271d1),
	.w4(32'h3b1e48dd),
	.w5(32'h3a7b13a2),
	.w6(32'h3bd71e34),
	.w7(32'h3bbebd3f),
	.w8(32'h3b60b6c3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a9544),
	.w1(32'h3c3db095),
	.w2(32'h3c4d22db),
	.w3(32'h3c3b663c),
	.w4(32'h3bac940e),
	.w5(32'h3b9c1c72),
	.w6(32'h3c0c632d),
	.w7(32'h3b6b6bab),
	.w8(32'h3bdeba2e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4fd7a),
	.w1(32'h3a860762),
	.w2(32'hbb2c834f),
	.w3(32'h3bba417e),
	.w4(32'h3be9099d),
	.w5(32'hbc2350e3),
	.w6(32'h3b44ff97),
	.w7(32'h3ae888b7),
	.w8(32'hbaf21451),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7dab4),
	.w1(32'hba7c2ae1),
	.w2(32'h3a19cbd8),
	.w3(32'hbbb3244f),
	.w4(32'hbb5fb1af),
	.w5(32'hbb17f373),
	.w6(32'hbc04c2e9),
	.w7(32'hbb8b5506),
	.w8(32'hbb1619f7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c58cb),
	.w1(32'hbba044a0),
	.w2(32'hbae696bf),
	.w3(32'h3a86f137),
	.w4(32'hba558a19),
	.w5(32'h397b6102),
	.w6(32'h39339642),
	.w7(32'h3a992f96),
	.w8(32'h3bae6f15),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af065),
	.w1(32'h3b7e9800),
	.w2(32'h3b93919b),
	.w3(32'h3b8035b7),
	.w4(32'h3b93a8eb),
	.w5(32'h3bcb2524),
	.w6(32'h3baf0ec0),
	.w7(32'hbadacc2a),
	.w8(32'h3a7cb398),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f7c67),
	.w1(32'hbb0f8085),
	.w2(32'hbbf6648c),
	.w3(32'h3bd439c6),
	.w4(32'hbbdbc447),
	.w5(32'hbc049063),
	.w6(32'h3c683dda),
	.w7(32'h3b76bb99),
	.w8(32'hbb6bfe8f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb915a),
	.w1(32'hb9fdf2a5),
	.w2(32'hbb7b6101),
	.w3(32'hbc248ea6),
	.w4(32'hbacfe7d5),
	.w5(32'hbb4b852a),
	.w6(32'hbbf84999),
	.w7(32'h3b727988),
	.w8(32'h3a635591),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96138c),
	.w1(32'h3c54b9ba),
	.w2(32'h3be1af60),
	.w3(32'h3c3959bb),
	.w4(32'h3bfd04b1),
	.w5(32'h3b9a2037),
	.w6(32'h3c4d413d),
	.w7(32'h3c17f376),
	.w8(32'h3c390fe2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92d70),
	.w1(32'hbc298b0e),
	.w2(32'h3aad37f0),
	.w3(32'hbc883927),
	.w4(32'hbc9df603),
	.w5(32'h3cca359d),
	.w6(32'hbc2902d3),
	.w7(32'hbb46690a),
	.w8(32'h3c925731),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dca07),
	.w1(32'hbbb3eca1),
	.w2(32'hbb096633),
	.w3(32'h3b927fb6),
	.w4(32'hbbf589e0),
	.w5(32'hbc0ade7d),
	.w6(32'h3c0a742e),
	.w7(32'hbb07bdb4),
	.w8(32'hbb8468ff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e774e),
	.w1(32'hbbd9e230),
	.w2(32'hbb2541c3),
	.w3(32'h39e6952b),
	.w4(32'hbb743299),
	.w5(32'hbb7ed5db),
	.w6(32'hbaaee2f7),
	.w7(32'hbc21cc07),
	.w8(32'hbc2116aa),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4bdad),
	.w1(32'hbace4075),
	.w2(32'h3b946c01),
	.w3(32'hb851ca62),
	.w4(32'hbbea03df),
	.w5(32'h3ccc8d0a),
	.w6(32'hbab6262f),
	.w7(32'hbb943cd3),
	.w8(32'h3c52cce2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c211ea),
	.w1(32'hbb041cc0),
	.w2(32'h3b7f53fe),
	.w3(32'hbb93226a),
	.w4(32'h3a6f6880),
	.w5(32'h3bd985ec),
	.w6(32'h3bb68d9d),
	.w7(32'h3a418a69),
	.w8(32'h3b846d42),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f3fc),
	.w1(32'hbc409b51),
	.w2(32'hbc00afee),
	.w3(32'hbb0ba1e3),
	.w4(32'h3b72d358),
	.w5(32'hbad7e3e4),
	.w6(32'h3aa91940),
	.w7(32'hbbff14ef),
	.w8(32'hbbb703bc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf99bf),
	.w1(32'h3c923492),
	.w2(32'h3c4f46ea),
	.w3(32'h3c8b9a9e),
	.w4(32'h3c490115),
	.w5(32'h3b954dc6),
	.w6(32'h3c426a00),
	.w7(32'h3c10a390),
	.w8(32'h3bd1a94b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab7ce8),
	.w1(32'h3c2e261c),
	.w2(32'h3c1e7045),
	.w3(32'h3c968dd3),
	.w4(32'h3ca98d9a),
	.w5(32'h3beba6cd),
	.w6(32'h3ce1b471),
	.w7(32'h3c2c2d30),
	.w8(32'h3be6d624),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9515a2),
	.w1(32'hbbfc9061),
	.w2(32'hbbd002a4),
	.w3(32'h3b4bb497),
	.w4(32'hbc5db338),
	.w5(32'hbbbcef34),
	.w6(32'h3b70922f),
	.w7(32'hbc435366),
	.w8(32'hbc10f2a9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b953d52),
	.w1(32'hbbaa09c6),
	.w2(32'hbb05c0a4),
	.w3(32'h3ac9e3ed),
	.w4(32'hbb83cffc),
	.w5(32'hbb041a8d),
	.w6(32'hbba58978),
	.w7(32'hbb0e9beb),
	.w8(32'h3b9dd4b8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d80ea5),
	.w1(32'hbaa3b493),
	.w2(32'hbc1514a8),
	.w3(32'h3ac24e32),
	.w4(32'hbb288303),
	.w5(32'hbb461a42),
	.w6(32'h3a8f4402),
	.w7(32'h3bc5b6e4),
	.w8(32'h3c315184),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd31c4),
	.w1(32'h3be489b8),
	.w2(32'hba648e57),
	.w3(32'hbc12149e),
	.w4(32'h3b9aa966),
	.w5(32'hbba3abfb),
	.w6(32'h3a309e50),
	.w7(32'h3bce11fc),
	.w8(32'hba582958),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c778bd8),
	.w1(32'h3c7bc347),
	.w2(32'h3c4364b5),
	.w3(32'h3cda4051),
	.w4(32'h3c3ff588),
	.w5(32'h3b4b7948),
	.w6(32'h3c80310b),
	.w7(32'h3c5e1749),
	.w8(32'h3c243dcc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f9535),
	.w1(32'h3b0a4617),
	.w2(32'hba85ff2c),
	.w3(32'hba60e78f),
	.w4(32'hbbb48f63),
	.w5(32'hbc1fce7c),
	.w6(32'hb998b800),
	.w7(32'hbab88841),
	.w8(32'h3ab6767e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f8ea5),
	.w1(32'hbb289697),
	.w2(32'hba727b0d),
	.w3(32'hbbc3524d),
	.w4(32'hbb9f5695),
	.w5(32'h3ac76682),
	.w6(32'h3b28a0cb),
	.w7(32'h3b794f59),
	.w8(32'h3c1598a5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1f045),
	.w1(32'hbbdd6f0b),
	.w2(32'h3a05d62a),
	.w3(32'hbb9e85a4),
	.w4(32'hbb8e05f9),
	.w5(32'h3c1c202d),
	.w6(32'hbb145497),
	.w7(32'hbc11790c),
	.w8(32'h3b09fdab),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8109d),
	.w1(32'hbc070d51),
	.w2(32'hbc3975d5),
	.w3(32'hbb450603),
	.w4(32'hbc244213),
	.w5(32'hbc69b800),
	.w6(32'h3b3968d9),
	.w7(32'h3b60fc8f),
	.w8(32'h3c81f29c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd53ec),
	.w1(32'hbc976924),
	.w2(32'hbc412096),
	.w3(32'hbc258c1f),
	.w4(32'hbc6d976f),
	.w5(32'h3bc46b0b),
	.w6(32'h3bd9ca58),
	.w7(32'hbbd2019b),
	.w8(32'hbb1f6e9a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ed57a),
	.w1(32'h3ae74964),
	.w2(32'hbb46733f),
	.w3(32'h3bbcecf6),
	.w4(32'h3b3407f3),
	.w5(32'hbc02dfd8),
	.w6(32'h3c099b8d),
	.w7(32'h3b33bbc1),
	.w8(32'h3c3e09e6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081d20),
	.w1(32'hbab65097),
	.w2(32'hbbdd46c1),
	.w3(32'hbb9a0068),
	.w4(32'hbc37cef8),
	.w5(32'hbbed65c4),
	.w6(32'h3b98b1ea),
	.w7(32'hbc13e87d),
	.w8(32'h3b42c562),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0476ab),
	.w1(32'h3cdfaec3),
	.w2(32'h3c852fa5),
	.w3(32'h3d2a8024),
	.w4(32'h3ce62c91),
	.w5(32'h3c115da3),
	.w6(32'h3d3831eb),
	.w7(32'h3cf0ba25),
	.w8(32'h3c139eec),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d06c),
	.w1(32'hbb0d8532),
	.w2(32'h3ac9bb11),
	.w3(32'hba534873),
	.w4(32'hba8c78c9),
	.w5(32'h3c560c42),
	.w6(32'hbbfb0aba),
	.w7(32'h391bb9fe),
	.w8(32'h3c6a0c39),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5534),
	.w1(32'h3c7bb56a),
	.w2(32'h3ac38df4),
	.w3(32'h3baab912),
	.w4(32'h3bd2b09d),
	.w5(32'hbbba1826),
	.w6(32'h3c6db768),
	.w7(32'h3c32446a),
	.w8(32'h3b5dc5bf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d7feb),
	.w1(32'hbb18a199),
	.w2(32'hbb0698d8),
	.w3(32'hbab3c715),
	.w4(32'hbbc4ea6a),
	.w5(32'hbc4cc689),
	.w6(32'hbc32c59d),
	.w7(32'h3b0bdfe5),
	.w8(32'h39c94e0a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5873),
	.w1(32'h3c2676fc),
	.w2(32'h3b07735f),
	.w3(32'h3b41cfdd),
	.w4(32'h3bca7c18),
	.w5(32'hb96df681),
	.w6(32'h3bb588e9),
	.w7(32'h3c44deb9),
	.w8(32'h3c432082),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba732c4b),
	.w1(32'hbbcc6e53),
	.w2(32'hbb04336e),
	.w3(32'hbbf97d68),
	.w4(32'hbc6df956),
	.w5(32'hbbbb99ea),
	.w6(32'hbaebfcc3),
	.w7(32'hbc375d54),
	.w8(32'h3b36eed0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7f429),
	.w1(32'hbc422c54),
	.w2(32'hbada081e),
	.w3(32'hbc5023e8),
	.w4(32'hbc17da25),
	.w5(32'h3cece773),
	.w6(32'hbb1742a9),
	.w7(32'hbc01254a),
	.w8(32'hbb88d9a7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0902f9),
	.w1(32'hba1d6805),
	.w2(32'hbb8e7de7),
	.w3(32'h3b28553a),
	.w4(32'hbb1c9fdc),
	.w5(32'hbbb90bd3),
	.w6(32'hbbc4ff54),
	.w7(32'h3b66f718),
	.w8(32'h3b893d2d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a995dad),
	.w1(32'h3ba78d19),
	.w2(32'h3c43c28e),
	.w3(32'hbac0a946),
	.w4(32'hba92554d),
	.w5(32'h3c348ae1),
	.w6(32'h3c1afacc),
	.w7(32'h3bef1950),
	.w8(32'h3bcc940c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e0547),
	.w1(32'hba99a19f),
	.w2(32'hbc46767f),
	.w3(32'hbc61e165),
	.w4(32'hbc28c518),
	.w5(32'hbbd23109),
	.w6(32'hbbc77cb3),
	.w7(32'h3b4aefb3),
	.w8(32'hba05d2ba),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c50f),
	.w1(32'h3cadea5d),
	.w2(32'h3c1d24d1),
	.w3(32'h3c8e54e8),
	.w4(32'h3d0c371a),
	.w5(32'h3c84e77c),
	.w6(32'h3c87b475),
	.w7(32'h3cbe1ff0),
	.w8(32'h3b84baa9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ff5c),
	.w1(32'hbcaf9a47),
	.w2(32'hbc8be02c),
	.w3(32'hbc8d7050),
	.w4(32'hbd0c223a),
	.w5(32'hbcc4562a),
	.w6(32'hbc96e01e),
	.w7(32'hbcbaeaa7),
	.w8(32'hbb767fac),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a926304),
	.w1(32'hbbc802f4),
	.w2(32'hbba2f61c),
	.w3(32'hbc7da1bc),
	.w4(32'hbbe4fd17),
	.w5(32'h3b56bce9),
	.w6(32'hbbc545b3),
	.w7(32'hbb6d5548),
	.w8(32'hbb87e908),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be00b83),
	.w1(32'h3c5e0518),
	.w2(32'h3b9f7064),
	.w3(32'hbb8862d1),
	.w4(32'hbb0a4c86),
	.w5(32'h39e5bd07),
	.w6(32'h3c1f8b5c),
	.w7(32'h3a7febfd),
	.w8(32'h3ba3fe81),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad43bed),
	.w1(32'hbb38b7d3),
	.w2(32'h3c4cb2ef),
	.w3(32'hb9d8ecce),
	.w4(32'hba7c0334),
	.w5(32'h3cd965e5),
	.w6(32'h3a79839f),
	.w7(32'hbb045f8b),
	.w8(32'h3c63d2a4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd45e8c),
	.w1(32'h3d08e315),
	.w2(32'h3d040d7f),
	.w3(32'h3cf75984),
	.w4(32'h3cb72a5c),
	.w5(32'h3c0375b9),
	.w6(32'h3d1fdd64),
	.w7(32'h3c836aaa),
	.w8(32'h3c948781),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0706),
	.w1(32'h3a9a5bcc),
	.w2(32'hbb94350d),
	.w3(32'hbbef3011),
	.w4(32'hbb6005e9),
	.w5(32'h3a8515b8),
	.w6(32'hbae5d439),
	.w7(32'hb91b3e0a),
	.w8(32'h3a77ae8a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab725d),
	.w1(32'h3be6bd30),
	.w2(32'hbb9b90dc),
	.w3(32'hbb60850f),
	.w4(32'h3a5ba5ff),
	.w5(32'hbc5825e4),
	.w6(32'h3b2fb000),
	.w7(32'h3ba08a00),
	.w8(32'h3b4b6e1a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07fcd9),
	.w1(32'h3b2bfd12),
	.w2(32'h3c0d548e),
	.w3(32'h3b190843),
	.w4(32'hbb584b88),
	.w5(32'h3bf5b768),
	.w6(32'hbb461491),
	.w7(32'h3bcf5a21),
	.w8(32'hba6a1b95),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964270),
	.w1(32'h39a426b1),
	.w2(32'h3b30a550),
	.w3(32'h3c6045f5),
	.w4(32'hba9019a3),
	.w5(32'h3c0b55df),
	.w6(32'h3c038e19),
	.w7(32'h3b736dd9),
	.w8(32'hbbf212a9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb220814),
	.w1(32'hbbf1f1a6),
	.w2(32'hbbb8aad4),
	.w3(32'hbbc4ee5d),
	.w4(32'hbc316336),
	.w5(32'h3c0b391b),
	.w6(32'hbbd825a5),
	.w7(32'hbc439fd9),
	.w8(32'hbaced4d2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91694),
	.w1(32'hba171c4a),
	.w2(32'h3a0b6308),
	.w3(32'hbb6a1340),
	.w4(32'hbb2d1519),
	.w5(32'hbaeb9376),
	.w6(32'h3b361a7c),
	.w7(32'h3c17845c),
	.w8(32'h3c14b956),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec7dc7),
	.w1(32'hbb1bda14),
	.w2(32'hba134e65),
	.w3(32'h3b69e024),
	.w4(32'hbbd1221c),
	.w5(32'hbbfc486c),
	.w6(32'hbbc215f7),
	.w7(32'h3bdb55a9),
	.w8(32'h3a8d862a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cda8e),
	.w1(32'h3bc4e339),
	.w2(32'h3bf453d6),
	.w3(32'hba326c55),
	.w4(32'h3c0e9c3c),
	.w5(32'h3b1f0f8d),
	.w6(32'h3b3d4a01),
	.w7(32'hb9abc8a6),
	.w8(32'hbbbd8548),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67e965),
	.w1(32'h3ae2fb87),
	.w2(32'hba0c9391),
	.w3(32'h3b9cc45a),
	.w4(32'hbb12fbde),
	.w5(32'h3be9cac3),
	.w6(32'h3bbd14d9),
	.w7(32'hbb515c12),
	.w8(32'h3af40c00),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b442f62),
	.w1(32'h3a6381ca),
	.w2(32'h3b9c50dc),
	.w3(32'h3bec0a8c),
	.w4(32'hbacc4a9e),
	.w5(32'h3bf6ae23),
	.w6(32'hbc001ab2),
	.w7(32'h3a20e0e7),
	.w8(32'hbad9bf40),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87138),
	.w1(32'hbbffa198),
	.w2(32'hba51eaac),
	.w3(32'hbc11d96c),
	.w4(32'hbc32c340),
	.w5(32'h3bae9fe5),
	.w6(32'hb8db5bc1),
	.w7(32'hbb9d3373),
	.w8(32'hbb4b55af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fdd9c),
	.w1(32'h3bba346e),
	.w2(32'hbaedad6a),
	.w3(32'h3a5e6b7d),
	.w4(32'h3c01eb96),
	.w5(32'h3bbd2631),
	.w6(32'hb852a22a),
	.w7(32'h3b38ae4b),
	.w8(32'h3ba1da5d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf791b),
	.w1(32'h3b1c7d8e),
	.w2(32'h3b3f62aa),
	.w3(32'hbc01d3eb),
	.w4(32'h3b86df4e),
	.w5(32'hbc29f9de),
	.w6(32'hb97fa206),
	.w7(32'h3a9e10ad),
	.w8(32'hbbd5da67),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e5092),
	.w1(32'hbaffb995),
	.w2(32'h3b589558),
	.w3(32'hbc26232b),
	.w4(32'hbbc24d3c),
	.w5(32'hbbab44b0),
	.w6(32'hbb845ff1),
	.w7(32'hbbef10c5),
	.w8(32'hbc345a9b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22c2c4),
	.w1(32'hbbd38e9b),
	.w2(32'hbaeac263),
	.w3(32'h381bb8a6),
	.w4(32'hbc60c519),
	.w5(32'h3caed7c8),
	.w6(32'hbb06b48d),
	.w7(32'hbbf17696),
	.w8(32'hb9854ccb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4ee04),
	.w1(32'h3aa9b95b),
	.w2(32'h3b0cb356),
	.w3(32'h3ada8f8d),
	.w4(32'hbb82b3dd),
	.w5(32'h3c014836),
	.w6(32'h3b0756fb),
	.w7(32'hbb13673c),
	.w8(32'h3bbfb859),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf196d6),
	.w1(32'h3c330f04),
	.w2(32'hba551501),
	.w3(32'h3c63872a),
	.w4(32'h3b8941ff),
	.w5(32'h3b970672),
	.w6(32'h3c816dcf),
	.w7(32'h3c3bde07),
	.w8(32'h3c02e601),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb8066),
	.w1(32'hbc2324e3),
	.w2(32'hbb9db650),
	.w3(32'h3c7e33a7),
	.w4(32'hbc9634ad),
	.w5(32'hbc0827f3),
	.w6(32'hbc19bc09),
	.w7(32'hbb86f54f),
	.w8(32'h3babb1b2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964ccaa),
	.w1(32'h3bd45a06),
	.w2(32'hbba2b0d2),
	.w3(32'h3a75c250),
	.w4(32'h3c09ff99),
	.w5(32'hbc0abf6f),
	.w6(32'h3ba4d67a),
	.w7(32'h3c589dd3),
	.w8(32'h3b282947),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a763929),
	.w1(32'h3b788ab0),
	.w2(32'h397ef9d5),
	.w3(32'h3ad75bd7),
	.w4(32'h3b99f2da),
	.w5(32'hbc03865f),
	.w6(32'h3c208b25),
	.w7(32'hbb9d9117),
	.w8(32'hbbde70ec),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fa5e2),
	.w1(32'hbb8e7f12),
	.w2(32'h3ad93814),
	.w3(32'h3af92d8e),
	.w4(32'h3b02a244),
	.w5(32'hbb67916c),
	.w6(32'h3baa6fc6),
	.w7(32'hbaf43fb6),
	.w8(32'h3b9010fc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6f6b6),
	.w1(32'hba13bea7),
	.w2(32'hbc115620),
	.w3(32'hbc1b78f1),
	.w4(32'h3a2f7780),
	.w5(32'hbc4f6e99),
	.w6(32'hbbb2c255),
	.w7(32'h3b4e6685),
	.w8(32'h3b51f09e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad38f56),
	.w1(32'hbc534a65),
	.w2(32'hbc2c4917),
	.w3(32'hbc7c2ed0),
	.w4(32'hbb77b526),
	.w5(32'h3ac9f0dc),
	.w6(32'h3c0314d2),
	.w7(32'hbb83ef72),
	.w8(32'h3ae033b5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c8f3),
	.w1(32'hbbf1e317),
	.w2(32'hbb161e81),
	.w3(32'h3b2d6a97),
	.w4(32'hbc022e6e),
	.w5(32'h3bfb8aa3),
	.w6(32'h3bc555b8),
	.w7(32'hbc241575),
	.w8(32'hbbef59af),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908fb0c),
	.w1(32'h3b89f3ae),
	.w2(32'h3b98b739),
	.w3(32'h3bf57b38),
	.w4(32'h3b03781b),
	.w5(32'h3ba6bbc5),
	.w6(32'hbb091eca),
	.w7(32'h3ade6c65),
	.w8(32'h3b22b2b1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8155),
	.w1(32'h3b645272),
	.w2(32'h3af5b78d),
	.w3(32'hb9e6ee18),
	.w4(32'h3ba67fdd),
	.w5(32'h3c4fee55),
	.w6(32'h3bf66d8a),
	.w7(32'hba9b09a4),
	.w8(32'h3c5677a4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba737cc),
	.w1(32'hbb8b65f9),
	.w2(32'hbb8218ad),
	.w3(32'hbb51f642),
	.w4(32'hbbc3305c),
	.w5(32'h3afd85b6),
	.w6(32'h3bcc0224),
	.w7(32'hbbcd3b2d),
	.w8(32'hbc3739a9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c018f5c),
	.w1(32'h3b7da549),
	.w2(32'hbabe58f5),
	.w3(32'hb8fcd61e),
	.w4(32'h3bb271c9),
	.w5(32'h3b971ec9),
	.w6(32'hbbe65808),
	.w7(32'h3b0d5742),
	.w8(32'hb90dfa40),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242b31),
	.w1(32'hb9f5671c),
	.w2(32'h3c108521),
	.w3(32'hbb178049),
	.w4(32'hbb8d3e17),
	.w5(32'hbc54d2fc),
	.w6(32'h3a434a8f),
	.w7(32'h3b8cfdcb),
	.w8(32'hbb01fc1c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c231498),
	.w1(32'h3af6f32d),
	.w2(32'h3b6b5424),
	.w3(32'h3b7b1c5c),
	.w4(32'h3bd9a437),
	.w5(32'h389d2b86),
	.w6(32'h3c7b419e),
	.w7(32'h3bf45542),
	.w8(32'h3b964961),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77de57),
	.w1(32'hbbb5596f),
	.w2(32'hbb591f19),
	.w3(32'hbb954997),
	.w4(32'hbb43d822),
	.w5(32'hbc3710dd),
	.w6(32'hbbb88f91),
	.w7(32'h3b1b07ab),
	.w8(32'hbbf678c0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c013818),
	.w1(32'hbb498199),
	.w2(32'h3b6b0830),
	.w3(32'hbbc6d8a4),
	.w4(32'hbbe0a396),
	.w5(32'h3ce40bb7),
	.w6(32'h3ba3630c),
	.w7(32'hba52f38b),
	.w8(32'h3bd9446f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8376bd),
	.w1(32'h3c81bc79),
	.w2(32'h3b8c263a),
	.w3(32'h3c7d449d),
	.w4(32'h3c4299d3),
	.w5(32'hbac7a9d2),
	.w6(32'h3c86090d),
	.w7(32'h3b9a8c95),
	.w8(32'hbb1a2633),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ad56),
	.w1(32'h3b4e8541),
	.w2(32'hbb9fe2f7),
	.w3(32'hba9ca71a),
	.w4(32'hbbb4a9e2),
	.w5(32'hba764c90),
	.w6(32'h3ab80ca4),
	.w7(32'hbb5720a9),
	.w8(32'hbbf1a63e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b3d0),
	.w1(32'hbb0cadd8),
	.w2(32'hbbc0df40),
	.w3(32'h3b8b22ee),
	.w4(32'hbbacb77c),
	.w5(32'hbc15bbc8),
	.w6(32'h3b82c53d),
	.w7(32'hbb46b17c),
	.w8(32'hbb58783a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac82b00),
	.w1(32'hbbd6a298),
	.w2(32'hbc01cca6),
	.w3(32'hb9101403),
	.w4(32'hbc27cf09),
	.w5(32'hbc128c61),
	.w6(32'h3b8a331a),
	.w7(32'hbaf5ec62),
	.w8(32'h3830d7d0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39341d),
	.w1(32'hbbdec88b),
	.w2(32'h3ace518e),
	.w3(32'hbc7e1ba4),
	.w4(32'hbc42ef75),
	.w5(32'h3c2ed1ab),
	.w6(32'hbc161025),
	.w7(32'hbc843167),
	.w8(32'h3bd87e4e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6b4b),
	.w1(32'hbb1d7c2d),
	.w2(32'h3b417fe4),
	.w3(32'hbba98722),
	.w4(32'hbb18a6b6),
	.w5(32'h3bfa6a9a),
	.w6(32'h3b77e142),
	.w7(32'hba472706),
	.w8(32'h3bd667c4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822118),
	.w1(32'h3a00d4b4),
	.w2(32'hbac0feec),
	.w3(32'h37fc6499),
	.w4(32'hbac591b8),
	.w5(32'hbb78f28f),
	.w6(32'h3b3b5e7d),
	.w7(32'h3ac3f2ae),
	.w8(32'hbb2317fc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbe1f5),
	.w1(32'hbb47c716),
	.w2(32'hba25bf96),
	.w3(32'h3b4e598e),
	.w4(32'hbbda5a71),
	.w5(32'hbb3e9970),
	.w6(32'hbb2f194f),
	.w7(32'hbbd16b60),
	.w8(32'hbb9db9ec),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52c4bb),
	.w1(32'hbb999947),
	.w2(32'h3b35b0fa),
	.w3(32'h3b52d254),
	.w4(32'h3a85889d),
	.w5(32'h3c1915cf),
	.w6(32'hbadc743a),
	.w7(32'hbbbf20de),
	.w8(32'hbabdce2c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42d4e0),
	.w1(32'hbc23faf3),
	.w2(32'hbab60d1c),
	.w3(32'hbc403a6e),
	.w4(32'hbc85bfa0),
	.w5(32'h3a4461e4),
	.w6(32'hbba70334),
	.w7(32'hbbb71e12),
	.w8(32'hbade01f0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d78bb),
	.w1(32'hba6d6678),
	.w2(32'h3bc81fc7),
	.w3(32'h3bb25eed),
	.w4(32'h3b355eea),
	.w5(32'h3bf1270b),
	.w6(32'h3c223e79),
	.w7(32'hbbe279c1),
	.w8(32'hbb0bf469),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc310317),
	.w1(32'h3c66666b),
	.w2(32'hb914b96f),
	.w3(32'hbc054ca3),
	.w4(32'h3c0b8607),
	.w5(32'hbc12b4ee),
	.w6(32'h3bdb2a11),
	.w7(32'h3bd0e8a5),
	.w8(32'h3c077e5b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7278a5),
	.w1(32'h3a6a8166),
	.w2(32'h3b092d06),
	.w3(32'hbba97155),
	.w4(32'hbb84b8e5),
	.w5(32'hbc399291),
	.w6(32'h3b5c1e63),
	.w7(32'h3a444d34),
	.w8(32'h3bbdd9f2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374a9d),
	.w1(32'hbb6f8808),
	.w2(32'hbbac3c8e),
	.w3(32'hbca2c792),
	.w4(32'hbbaaa55d),
	.w5(32'h3b99b388),
	.w6(32'hbbd56c37),
	.w7(32'h3b88bb27),
	.w8(32'h3bccb613),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca34ffc),
	.w1(32'h3c3fec16),
	.w2(32'h3bf829c1),
	.w3(32'hbaed82d2),
	.w4(32'h3c1b406a),
	.w5(32'h3b8aca2f),
	.w6(32'h3c236b7a),
	.w7(32'h3c6190b5),
	.w8(32'h3be3c08d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc3c2d),
	.w1(32'h3bda6a2b),
	.w2(32'h3c610d7d),
	.w3(32'hbb93c314),
	.w4(32'h3c363a23),
	.w5(32'h3c8ed92c),
	.w6(32'hbc2cea99),
	.w7(32'h3c90b449),
	.w8(32'h3cac5772),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32d591),
	.w1(32'h3bb3e755),
	.w2(32'hbacf863e),
	.w3(32'hbc73709e),
	.w4(32'h3ab2ec1a),
	.w5(32'hbc3b6f87),
	.w6(32'hbb750882),
	.w7(32'h3c158f2c),
	.w8(32'h3bad679c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57c229),
	.w1(32'hbb35e571),
	.w2(32'h3a0cd2dc),
	.w3(32'hbc2f1660),
	.w4(32'hbb9ebc39),
	.w5(32'hbbcca801),
	.w6(32'hbc8deb8b),
	.w7(32'hbbc16fb9),
	.w8(32'hbad097b1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c080452),
	.w1(32'hba16605a),
	.w2(32'hbaacbb2c),
	.w3(32'hbc0ba299),
	.w4(32'hbb728753),
	.w5(32'h3c8fe785),
	.w6(32'hba0e84e0),
	.w7(32'h3b5e53b4),
	.w8(32'h3ba12369),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b8db),
	.w1(32'hbc943a24),
	.w2(32'hba83d99e),
	.w3(32'hbc0f3144),
	.w4(32'hbcbda7dd),
	.w5(32'hbbe02126),
	.w6(32'hbbcd5370),
	.w7(32'hbc36334c),
	.w8(32'hba0861b1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21a005),
	.w1(32'hba9d7e7c),
	.w2(32'hbc2cdcf6),
	.w3(32'hbbe31f36),
	.w4(32'hbb05759b),
	.w5(32'hbcc588fe),
	.w6(32'h3a08de03),
	.w7(32'h3b85e303),
	.w8(32'hbc236bd1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8453910),
	.w1(32'hbb3ddb09),
	.w2(32'hbba1afc1),
	.w3(32'hbbe340eb),
	.w4(32'h3c185d64),
	.w5(32'hba8864c8),
	.w6(32'h3aeb2784),
	.w7(32'hbb3b4053),
	.w8(32'hb78d932b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61f6e8),
	.w1(32'hbb3095cf),
	.w2(32'h3b568dc7),
	.w3(32'h3b0276f7),
	.w4(32'hbb586214),
	.w5(32'h3c7c6451),
	.w6(32'h3bc179df),
	.w7(32'hbb4de618),
	.w8(32'h3bc54710),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ac26d),
	.w1(32'hbb4972f5),
	.w2(32'hbb7c9025),
	.w3(32'h3b78fcf3),
	.w4(32'hbbe12fae),
	.w5(32'h3b957b0c),
	.w6(32'h3b2e0cbe),
	.w7(32'hbac1668c),
	.w8(32'hba9cbe25),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a0db4),
	.w1(32'h3a94d470),
	.w2(32'hbc29a8b2),
	.w3(32'h3b317e04),
	.w4(32'hbac9183b),
	.w5(32'h39f77739),
	.w6(32'hba52ccd8),
	.w7(32'hb93c7100),
	.w8(32'hbba5221f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39153386),
	.w1(32'h3c1cdff7),
	.w2(32'h3acbce4f),
	.w3(32'hbb89b644),
	.w4(32'h3b8237b9),
	.w5(32'hbc1c08da),
	.w6(32'hbbac962d),
	.w7(32'h3c161ba2),
	.w8(32'hbbe8e2eb),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3ff3),
	.w1(32'hbbdfcbd7),
	.w2(32'h3aa1a65d),
	.w3(32'hbc27dcfb),
	.w4(32'hbb979bad),
	.w5(32'h3c8005a4),
	.w6(32'h39f089f8),
	.w7(32'hbba5f348),
	.w8(32'hbb4cced5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6982eb),
	.w1(32'hbc374272),
	.w2(32'h3a060bea),
	.w3(32'h3be53056),
	.w4(32'hbc39f64d),
	.w5(32'h3c196bcf),
	.w6(32'hb846b0e9),
	.w7(32'hbc2051fa),
	.w8(32'hbabb41c7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c82ea5),
	.w1(32'h3b42c51f),
	.w2(32'h3c12ec32),
	.w3(32'h3b139aee),
	.w4(32'hbab0f1c5),
	.w5(32'h3c5f5374),
	.w6(32'h3b9b1a79),
	.w7(32'hba4b86eb),
	.w8(32'h3b98e46e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6fec7),
	.w1(32'hbc0dab21),
	.w2(32'hbbef46e7),
	.w3(32'hbaab8158),
	.w4(32'hbc0b4264),
	.w5(32'h3c9ee531),
	.w6(32'h3b061058),
	.w7(32'hbc0c0ca6),
	.w8(32'hbc28b98e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ada9),
	.w1(32'hbc14e762),
	.w2(32'hbb912abb),
	.w3(32'hbb530748),
	.w4(32'hbc5eba10),
	.w5(32'h3a37de76),
	.w6(32'hbc5bb5cc),
	.w7(32'hbc117f08),
	.w8(32'hbb3f5979),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36b5ec),
	.w1(32'hbac76eac),
	.w2(32'h3b2c4bbc),
	.w3(32'h3c3d06f0),
	.w4(32'h3b85f5cb),
	.w5(32'hbb1fa697),
	.w6(32'h3c7b1bdb),
	.w7(32'h3b8ed301),
	.w8(32'h3c05c78f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc0a29),
	.w1(32'h3ab98071),
	.w2(32'h3be381b0),
	.w3(32'h37bd4f4b),
	.w4(32'hbaf2a852),
	.w5(32'hb98536ba),
	.w6(32'h3bbdca3c),
	.w7(32'h3aabb868),
	.w8(32'h3b890039),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba380cc),
	.w1(32'hbbbe646a),
	.w2(32'hba4c6937),
	.w3(32'hbb01f04d),
	.w4(32'hbc16e56b),
	.w5(32'h3c5fad46),
	.w6(32'h3b577f10),
	.w7(32'hbbcf0c8d),
	.w8(32'h39735ede),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04db91),
	.w1(32'hbbf7be36),
	.w2(32'hbc15e1f3),
	.w3(32'hbb611dcf),
	.w4(32'hbc19a51e),
	.w5(32'hbbd635cd),
	.w6(32'hbbb8c4da),
	.w7(32'hbc412c06),
	.w8(32'hbc593426),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04417c),
	.w1(32'hbb95fbbb),
	.w2(32'h3ad499df),
	.w3(32'h3c0a9fa6),
	.w4(32'hbbd2a47d),
	.w5(32'h3c370530),
	.w6(32'h3a57ff80),
	.w7(32'h3abb1e5a),
	.w8(32'h3a1e50d4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec9c7b),
	.w1(32'h3a79bd44),
	.w2(32'hbba71af7),
	.w3(32'hbb0c87f5),
	.w4(32'h3a434856),
	.w5(32'hbb7d5a27),
	.w6(32'h3b8e68ba),
	.w7(32'h3bf44662),
	.w8(32'hbb370861),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c099a25),
	.w1(32'h3b2cc4a2),
	.w2(32'hbba0286c),
	.w3(32'h3c7b3913),
	.w4(32'h3bc2c8b5),
	.w5(32'h3adeab3b),
	.w6(32'h3bebc131),
	.w7(32'h3c40fe2c),
	.w8(32'h3c62e41e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd57d4e),
	.w1(32'hbb991cb1),
	.w2(32'h3b9999bf),
	.w3(32'h3be87538),
	.w4(32'hbbf9fc8c),
	.w5(32'h3c88ac39),
	.w6(32'h3b425307),
	.w7(32'hbb89c087),
	.w8(32'hbb7448ef),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f7c6a),
	.w1(32'hbab86fe1),
	.w2(32'hbb2a72f2),
	.w3(32'h3c27e19e),
	.w4(32'h3b9cd7ab),
	.w5(32'hbbfda88f),
	.w6(32'h3a5d491f),
	.w7(32'h3c20b5de),
	.w8(32'h3b8489cc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94dbe6),
	.w1(32'h3b0dcddc),
	.w2(32'hbaee6510),
	.w3(32'hbb927eb3),
	.w4(32'h3ae8aa8e),
	.w5(32'hbc102a04),
	.w6(32'hbb148922),
	.w7(32'h3b8cda0f),
	.w8(32'hbaabeb20),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e085e8),
	.w1(32'h3a81232c),
	.w2(32'h39912942),
	.w3(32'h3c16e682),
	.w4(32'hbaac6418),
	.w5(32'hbbde9553),
	.w6(32'h3bcbc406),
	.w7(32'h39ef17b5),
	.w8(32'hbb0b29bf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a37a6),
	.w1(32'h3accd62a),
	.w2(32'hbb52a017),
	.w3(32'h3b80d144),
	.w4(32'hba8f4472),
	.w5(32'h3b848a3b),
	.w6(32'h3bb13f63),
	.w7(32'hbb6ab8af),
	.w8(32'hbbd071b6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be15fbf),
	.w1(32'h3b8ee34a),
	.w2(32'h3b5ae9d3),
	.w3(32'hb892f68b),
	.w4(32'hbb4a6c0e),
	.w5(32'hbbc4ffaf),
	.w6(32'h3c1681de),
	.w7(32'h3bfc469f),
	.w8(32'h3a479e93),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd71a9),
	.w1(32'h3b8f943d),
	.w2(32'h3b94e780),
	.w3(32'hbbd01075),
	.w4(32'h3a889570),
	.w5(32'h38abd24c),
	.w6(32'h3939ec0f),
	.w7(32'h3bffc4b0),
	.w8(32'h3b0c5db1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87c2a7),
	.w1(32'hb9c0154d),
	.w2(32'hba58d1e1),
	.w3(32'hbbf0ada8),
	.w4(32'hbafecdd7),
	.w5(32'h3c122a6b),
	.w6(32'h3b0cb032),
	.w7(32'h399c34c0),
	.w8(32'hbb877dc2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab19b1b),
	.w1(32'hb9f3d59c),
	.w2(32'h3b540df5),
	.w3(32'hba9ae931),
	.w4(32'hb9cd261e),
	.w5(32'h3cb7abc5),
	.w6(32'h3bdb2eda),
	.w7(32'h3b457047),
	.w8(32'h3be5bba1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f82f2),
	.w1(32'h3be7563e),
	.w2(32'hbb13087b),
	.w3(32'hbb370267),
	.w4(32'h3bdf3faa),
	.w5(32'hbc046d72),
	.w6(32'hbbc2188b),
	.w7(32'h3c1f71bc),
	.w8(32'hb9691208),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84c810),
	.w1(32'hbb99b6dd),
	.w2(32'h3a080287),
	.w3(32'h3bc98cb3),
	.w4(32'hbc9d792a),
	.w5(32'hbc2b3106),
	.w6(32'h3b1f6fb4),
	.w7(32'hbc0b145d),
	.w8(32'hb9287011),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2d746),
	.w1(32'hbacb32df),
	.w2(32'hbb9d3401),
	.w3(32'hbade577c),
	.w4(32'hbbf3e407),
	.w5(32'hbbcb64ac),
	.w6(32'hbba45c18),
	.w7(32'hbb22c68e),
	.w8(32'hbbc01b36),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b17d9),
	.w1(32'h3cae3db6),
	.w2(32'h3c4bbc9c),
	.w3(32'h3bbf3de3),
	.w4(32'h3cabf39c),
	.w5(32'h3cbf87a5),
	.w6(32'h3c0f71f9),
	.w7(32'h3c83c056),
	.w8(32'hba7fee09),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6795b7),
	.w1(32'hbc0f22a9),
	.w2(32'hbc975b93),
	.w3(32'hbc98de5e),
	.w4(32'hbc2868dd),
	.w5(32'hbc680c05),
	.w6(32'h3b1af20d),
	.w7(32'hba920779),
	.w8(32'h3ba63084),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc678930),
	.w1(32'h3a324699),
	.w2(32'hbba8ae00),
	.w3(32'h3c371469),
	.w4(32'h3acd535b),
	.w5(32'h3c283c20),
	.w6(32'hbbf4a14f),
	.w7(32'hb98b1067),
	.w8(32'h3ac4753d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ccb6f),
	.w1(32'h3ba4231f),
	.w2(32'hbb15b812),
	.w3(32'hbb12457e),
	.w4(32'h3c092f82),
	.w5(32'h3c70cd17),
	.w6(32'h3add4490),
	.w7(32'h3bb581f5),
	.w8(32'hbb8c3adb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ce5f1),
	.w1(32'h39d512f2),
	.w2(32'hbbb74f85),
	.w3(32'h37e7d051),
	.w4(32'hbb7c0fca),
	.w5(32'hbc09255f),
	.w6(32'hb8b9924e),
	.w7(32'hbb74cb9c),
	.w8(32'hbbdc4fae),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae14bac),
	.w1(32'h3b319a35),
	.w2(32'hbb16b4b4),
	.w3(32'h3b3392e7),
	.w4(32'h3ba2f721),
	.w5(32'hbc0dfa1f),
	.w6(32'h3a4a9e1f),
	.w7(32'h398ae6d4),
	.w8(32'hbbec9ac9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71ae31),
	.w1(32'hb9361a57),
	.w2(32'h3984be51),
	.w3(32'h3ac55abd),
	.w4(32'h3a2fda2c),
	.w5(32'h3c299b95),
	.w6(32'hbb6d51da),
	.w7(32'h3b8a785b),
	.w8(32'hbb6820a5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac851f4),
	.w1(32'h3b9f6fe2),
	.w2(32'h3b3033b2),
	.w3(32'h3bf58191),
	.w4(32'h3bef5edc),
	.w5(32'hbb0ac6d5),
	.w6(32'hba72dd32),
	.w7(32'h3c08ce00),
	.w8(32'h3c359d75),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad5573),
	.w1(32'h3b0bce3a),
	.w2(32'hbbd21f07),
	.w3(32'hbba452f1),
	.w4(32'h3b815597),
	.w5(32'hbb94510d),
	.w6(32'h3c54b3ca),
	.w7(32'h3c6ec06a),
	.w8(32'h3ab71190),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f6556),
	.w1(32'hbb9a9922),
	.w2(32'h3b8281ab),
	.w3(32'hbbd7be22),
	.w4(32'hbc0954e5),
	.w5(32'h3cb5187b),
	.w6(32'hbb91d5ef),
	.w7(32'hbaab37fa),
	.w8(32'h39b89a11),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18e195),
	.w1(32'hbb2f505f),
	.w2(32'h3c0fa629),
	.w3(32'hbb3f75fe),
	.w4(32'h3b8b4a71),
	.w5(32'h3cf9b872),
	.w6(32'hbaf3a5cb),
	.w7(32'h3b4e6000),
	.w8(32'h3ca7d1d2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13afbe),
	.w1(32'h3c2ea86f),
	.w2(32'h3be82fa7),
	.w3(32'h3ca0e4ea),
	.w4(32'h3c4d2caf),
	.w5(32'h3a45d592),
	.w6(32'h3c2691e5),
	.w7(32'h3bd7a7d6),
	.w8(32'hbc1196c1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae166f2),
	.w1(32'hbbc961a6),
	.w2(32'h3a4fad35),
	.w3(32'hbc6f1eab),
	.w4(32'hbb271c8a),
	.w5(32'hbb6f03d8),
	.w6(32'hbca99769),
	.w7(32'h3c81ca9c),
	.w8(32'h3b0db8ab),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c236e8d),
	.w1(32'h3c333984),
	.w2(32'h3b279dd4),
	.w3(32'h3bbe8063),
	.w4(32'h3c7307c2),
	.w5(32'h3c078847),
	.w6(32'hbbd97e39),
	.w7(32'h3c2e8763),
	.w8(32'h3b5b4492),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28482a),
	.w1(32'hbafeda32),
	.w2(32'hbc1f6598),
	.w3(32'h3c1d4608),
	.w4(32'hbc253cb4),
	.w5(32'hbc8aa555),
	.w6(32'h3c4f37a2),
	.w7(32'hbc219e5c),
	.w8(32'hbc2918c5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95570f),
	.w1(32'hba973c52),
	.w2(32'h3c018d69),
	.w3(32'hbb9f3cb9),
	.w4(32'hbb9cf52d),
	.w5(32'hbc0302b8),
	.w6(32'h3b49f4dd),
	.w7(32'h3b72ec41),
	.w8(32'h3bda797b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0072b),
	.w1(32'hbb21b732),
	.w2(32'hbb617591),
	.w3(32'hbc5f8a8b),
	.w4(32'hbc4feaf8),
	.w5(32'hbc241691),
	.w6(32'hbc199896),
	.w7(32'hbc252465),
	.w8(32'hbc331ded),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bfddf),
	.w1(32'h3b9b0f85),
	.w2(32'hbb8be1d8),
	.w3(32'hbb8879d5),
	.w4(32'h3c51f24d),
	.w5(32'hbb8fb7ec),
	.w6(32'hbb8bf60a),
	.w7(32'h3c1cc2b4),
	.w8(32'h3b7b2409),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2da135),
	.w1(32'h3ab4ceb8),
	.w2(32'hbb856ea6),
	.w3(32'hbc2799b2),
	.w4(32'h3bad1afb),
	.w5(32'h3a3752d0),
	.w6(32'hbbf5fbf7),
	.w7(32'hbb7f31dc),
	.w8(32'h3c02975b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0632ce),
	.w1(32'hbb2819dd),
	.w2(32'h3bbc87d3),
	.w3(32'hbb686129),
	.w4(32'hbb5acdae),
	.w5(32'h3c17aae7),
	.w6(32'hbb5f696f),
	.w7(32'hbbfd4e7c),
	.w8(32'h3b6a1f77),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde35b1),
	.w1(32'h3c5b37e9),
	.w2(32'hbbb5b212),
	.w3(32'h3c0ca22a),
	.w4(32'h3c452fec),
	.w5(32'h397f3c3d),
	.w6(32'h3c10a780),
	.w7(32'h3b3f01f0),
	.w8(32'h3c035212),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70cb15),
	.w1(32'h3bacb636),
	.w2(32'h3b1bd5a9),
	.w3(32'h3b7916b0),
	.w4(32'h3a6d7342),
	.w5(32'h3bbc2be0),
	.w6(32'h3c5fb006),
	.w7(32'h3c413bde),
	.w8(32'h3c36ac70),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c455c75),
	.w1(32'h3c038e16),
	.w2(32'hbbe36a49),
	.w3(32'h3cba15fe),
	.w4(32'h3a570c49),
	.w5(32'hbc2e9deb),
	.w6(32'h3c9b0a7f),
	.w7(32'h3bc436f8),
	.w8(32'hbbb623b4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b063494),
	.w1(32'hbaa7a567),
	.w2(32'hba912da3),
	.w3(32'hbb97e3b5),
	.w4(32'hbbe41bab),
	.w5(32'h38cebea1),
	.w6(32'h3b1b4f63),
	.w7(32'hbb4c685e),
	.w8(32'hbc13210c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac56885),
	.w1(32'h394969dd),
	.w2(32'hbc0c14ac),
	.w3(32'h3aa2fde4),
	.w4(32'hbba22621),
	.w5(32'h378193cf),
	.w6(32'hbbc1003c),
	.w7(32'hbc059396),
	.w8(32'hbbfba170),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78b74d),
	.w1(32'h3c5f7f54),
	.w2(32'hbabc8f48),
	.w3(32'h3bb14bdf),
	.w4(32'h3abac1e7),
	.w5(32'hbb72b362),
	.w6(32'h3c6b8c7d),
	.w7(32'h3cb8377b),
	.w8(32'h3bf6197f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e67c7),
	.w1(32'hbbe87a81),
	.w2(32'hbc5fc177),
	.w3(32'hbc845969),
	.w4(32'hbb97f59d),
	.w5(32'hbb6caac9),
	.w6(32'hbbdbe772),
	.w7(32'hbb13e346),
	.w8(32'hbb8f8a59),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0118fb),
	.w1(32'h3c239c30),
	.w2(32'h3a787738),
	.w3(32'hba0d5b80),
	.w4(32'h3c06f656),
	.w5(32'h3cae04b7),
	.w6(32'h3c34c568),
	.w7(32'hbaa4f67b),
	.w8(32'h3c6cae46),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178b8a),
	.w1(32'h3a9056cd),
	.w2(32'hbc31b4b5),
	.w3(32'hbb74f4ab),
	.w4(32'hbbadc0e8),
	.w5(32'hbc3a77cd),
	.w6(32'h3b5e136f),
	.w7(32'hbc7a0119),
	.w8(32'h3b2f7d35),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ce7e4),
	.w1(32'h3b10efda),
	.w2(32'h3b07e021),
	.w3(32'hbc68408d),
	.w4(32'h3c16f483),
	.w5(32'hbb22099c),
	.w6(32'h3a84d9c5),
	.w7(32'hbbc31bfd),
	.w8(32'h3a12a67b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc492c35),
	.w1(32'h3bc130ad),
	.w2(32'h3c2622d4),
	.w3(32'hbc4bd5c2),
	.w4(32'h3c76a500),
	.w5(32'h3cc3ba53),
	.w6(32'hbbf415e3),
	.w7(32'h3ba88d7c),
	.w8(32'h3c23cc5f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75ee24),
	.w1(32'h3caadd0a),
	.w2(32'h3c343274),
	.w3(32'h3c4fa8a1),
	.w4(32'h3cc6d976),
	.w5(32'h3c661928),
	.w6(32'h3c89841c),
	.w7(32'h3cde39a0),
	.w8(32'h3c043079),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b134e21),
	.w1(32'h3c90c5b7),
	.w2(32'h3c57e6ba),
	.w3(32'hba8ddcf5),
	.w4(32'h3c40e314),
	.w5(32'h3c612db3),
	.w6(32'h3bece595),
	.w7(32'h3c248ad0),
	.w8(32'h3c61814c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48f6f),
	.w1(32'hbc088988),
	.w2(32'hba8cca3e),
	.w3(32'h3a13e343),
	.w4(32'hbc860c3d),
	.w5(32'hbb51de1a),
	.w6(32'h3ba23cd4),
	.w7(32'hbbf3ecaf),
	.w8(32'h3a878624),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c547fd8),
	.w1(32'hbbc34350),
	.w2(32'hbb311bee),
	.w3(32'h3c0584fb),
	.w4(32'hbc10e8bc),
	.w5(32'hba79ddc2),
	.w6(32'h3b5c7b59),
	.w7(32'hbb03044e),
	.w8(32'h3b4c1bcc),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb4c18),
	.w1(32'h3b6f80c6),
	.w2(32'hbb12bd76),
	.w3(32'h3b1f3375),
	.w4(32'h3c6a0463),
	.w5(32'h3a51de67),
	.w6(32'h3b6a2844),
	.w7(32'hbbdb6bdb),
	.w8(32'h3bd72adf),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a70b1),
	.w1(32'h3c0a0cf8),
	.w2(32'h39ca3095),
	.w3(32'hbc0dc66b),
	.w4(32'h3c041243),
	.w5(32'hba93cfeb),
	.w6(32'h3bc09c4e),
	.w7(32'h3a562d6b),
	.w8(32'hbb97bb4e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38636c),
	.w1(32'hba026d0b),
	.w2(32'hbc65259a),
	.w3(32'hbc1a7922),
	.w4(32'hbc4c3a3b),
	.w5(32'hbc9748fc),
	.w6(32'hbc018794),
	.w7(32'hbc10e110),
	.w8(32'hbc4a58b2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65d34a),
	.w1(32'h3bab3ad2),
	.w2(32'h3af79974),
	.w3(32'hbcec9a83),
	.w4(32'h3c023715),
	.w5(32'h3bcf3c71),
	.w6(32'hbbfb8f75),
	.w7(32'h3c08423b),
	.w8(32'hba1f8705),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9193b),
	.w1(32'hbacfd4c5),
	.w2(32'h3c06d2f7),
	.w3(32'hb997e8be),
	.w4(32'h3b63ebb7),
	.w5(32'h3b88e660),
	.w6(32'hbbb229be),
	.w7(32'h3ba12046),
	.w8(32'h3b85ea8c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2600b4),
	.w1(32'hbb4f5c3e),
	.w2(32'h3c086d83),
	.w3(32'h3b37f852),
	.w4(32'hbc26b058),
	.w5(32'h3c0ffa54),
	.w6(32'h3a95561d),
	.w7(32'h3b1e5e38),
	.w8(32'h3b796af5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8483),
	.w1(32'h3b64e79d),
	.w2(32'hbaddb7ab),
	.w3(32'h3c459703),
	.w4(32'h3bc39525),
	.w5(32'hbbaa922b),
	.w6(32'hbb8a775a),
	.w7(32'hbb6c647c),
	.w8(32'h3b6f10d3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28e526),
	.w1(32'hbc47f5b8),
	.w2(32'hbc4c2e84),
	.w3(32'hbc07ea4e),
	.w4(32'hbcb8ad4d),
	.w5(32'hbc1eebc9),
	.w6(32'hbba2544a),
	.w7(32'hbb17fa8f),
	.w8(32'hbc10c123),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03e9bf),
	.w1(32'h3bc86fb6),
	.w2(32'h3c0d2719),
	.w3(32'h3b5c6c21),
	.w4(32'h3c238a6f),
	.w5(32'h3b7ddecf),
	.w6(32'h3c1fdadd),
	.w7(32'h3c4759c6),
	.w8(32'hbc090a41),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b201c7d),
	.w1(32'h39300ac7),
	.w2(32'h3bb0d997),
	.w3(32'h3ba32812),
	.w4(32'hbb48c659),
	.w5(32'h3ca5de68),
	.w6(32'h3884f035),
	.w7(32'h3b413d79),
	.w8(32'h3c521ab9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05cc5),
	.w1(32'h3b14f5c0),
	.w2(32'h3b020cbf),
	.w3(32'hbaf17503),
	.w4(32'h3bbae07d),
	.w5(32'h3ac89410),
	.w6(32'h3aa4e3fd),
	.w7(32'h3be219c4),
	.w8(32'h3b4d0353),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1570c3),
	.w1(32'h3c22506e),
	.w2(32'hbb04ea9d),
	.w3(32'h3c160241),
	.w4(32'h3b86a582),
	.w5(32'hbbbe2797),
	.w6(32'hb94922b9),
	.w7(32'h3c4e229d),
	.w8(32'h3b3189c5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39560ea1),
	.w1(32'h3b7ef606),
	.w2(32'hbbd91ce3),
	.w3(32'hbb12d3b0),
	.w4(32'h3c3a4e88),
	.w5(32'h3ac618f6),
	.w6(32'h3b64ee0d),
	.w7(32'h3b52e9e7),
	.w8(32'hbb33899d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c23fb),
	.w1(32'hbbd5059b),
	.w2(32'h3c799644),
	.w3(32'hba83ba8f),
	.w4(32'hbc21c763),
	.w5(32'h3c7f9b69),
	.w6(32'h3a74b7fc),
	.w7(32'hbb8737a9),
	.w8(32'h3b7bb2cd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b2d72),
	.w1(32'hbc1ab826),
	.w2(32'hbbefc7fd),
	.w3(32'h3c8aae83),
	.w4(32'hbc93928c),
	.w5(32'hbc72acc0),
	.w6(32'h3bb66e90),
	.w7(32'hbb5f220d),
	.w8(32'hbc1d9764),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780176),
	.w1(32'hbc0bb4d6),
	.w2(32'hbc25db1f),
	.w3(32'hbb5fd886),
	.w4(32'hbb378906),
	.w5(32'hbbe3925f),
	.w6(32'hbc2e12d5),
	.w7(32'h3ba2480a),
	.w8(32'h3b2b6274),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e42f),
	.w1(32'h3b21df26),
	.w2(32'hbba95dc3),
	.w3(32'h3a2818e7),
	.w4(32'hbc1c0374),
	.w5(32'h3ac0ca64),
	.w6(32'hbb05da5b),
	.w7(32'h3aa6755b),
	.w8(32'h3b1b816b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb851c),
	.w1(32'h3bb585b4),
	.w2(32'hbbceebb9),
	.w3(32'h3c377ece),
	.w4(32'h3b74164e),
	.w5(32'hbb762456),
	.w6(32'h3c6fb1bb),
	.w7(32'h3c3d6ccd),
	.w8(32'h3ab60d88),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbae5fd),
	.w1(32'hbaf4f484),
	.w2(32'hbc1e3846),
	.w3(32'h3b03adba),
	.w4(32'hbc0693fb),
	.w5(32'hbcc1af8c),
	.w6(32'hbb65c395),
	.w7(32'h3b291796),
	.w8(32'hbbec783d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d28ec),
	.w1(32'h3b7fb351),
	.w2(32'hbb744881),
	.w3(32'h3b02b490),
	.w4(32'hbb122f8c),
	.w5(32'h39fe4d50),
	.w6(32'h3c8bbef2),
	.w7(32'h3bcd0e93),
	.w8(32'hbbd63dd9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ef036),
	.w1(32'hbb8f5146),
	.w2(32'h3c4eb0a0),
	.w3(32'hbafe1c00),
	.w4(32'hbb8cb33a),
	.w5(32'h3c993b06),
	.w6(32'hbbd367f3),
	.w7(32'hbbf28e19),
	.w8(32'h3c5a23c1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4351e9),
	.w1(32'h3a892b3f),
	.w2(32'hbaf583ac),
	.w3(32'h3c3ded9b),
	.w4(32'hbabf57ee),
	.w5(32'hb93a8d70),
	.w6(32'h3c87a993),
	.w7(32'h3aadfd42),
	.w8(32'hbab1c70e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bd8b6),
	.w1(32'hbb822310),
	.w2(32'hbba71f13),
	.w3(32'h3b517d10),
	.w4(32'h382ed6db),
	.w5(32'hbc484bb1),
	.w6(32'h39f98ce0),
	.w7(32'h3a779609),
	.w8(32'hbb21fca8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f3b08),
	.w1(32'h3bac6dab),
	.w2(32'hbb6d3f25),
	.w3(32'hbc7bd703),
	.w4(32'h3be36516),
	.w5(32'hbb79a3f4),
	.w6(32'hba3aa42f),
	.w7(32'h3c07b567),
	.w8(32'hbbd3fcf9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3ffbc),
	.w1(32'hbafc8bc7),
	.w2(32'h3bd2ea53),
	.w3(32'h3a912552),
	.w4(32'hbb4be8e4),
	.w5(32'hbbceb129),
	.w6(32'hbb941476),
	.w7(32'hb98745dd),
	.w8(32'h3baf7465),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b8461),
	.w1(32'hbafef53c),
	.w2(32'h3bb0f7ce),
	.w3(32'hbc3c041b),
	.w4(32'hbb10acc1),
	.w5(32'h3ced55e1),
	.w6(32'h3a8f8b19),
	.w7(32'hbbea2f19),
	.w8(32'h3b5961a6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb731134),
	.w1(32'h39ce4ce0),
	.w2(32'h37628ee7),
	.w3(32'h3b840c40),
	.w4(32'h3c450452),
	.w5(32'h3bacf8db),
	.w6(32'hbc005b98),
	.w7(32'h3bd82842),
	.w8(32'h3b8ec15c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1febb1),
	.w1(32'hba2f5c81),
	.w2(32'h3accfff4),
	.w3(32'hbbdb7206),
	.w4(32'hbbcb8691),
	.w5(32'h3bd79063),
	.w6(32'hbbb4bc61),
	.w7(32'hba8afd87),
	.w8(32'h3c4153c4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc60070),
	.w1(32'h3c166943),
	.w2(32'hbb3e18b9),
	.w3(32'h3c5936e8),
	.w4(32'h3b731c66),
	.w5(32'hbc33c6f0),
	.w6(32'h3b6f4ac4),
	.w7(32'hbb7788b5),
	.w8(32'hbc11b5cb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb27a1),
	.w1(32'hbc75b898),
	.w2(32'hbc60682f),
	.w3(32'hbc8594c7),
	.w4(32'hbd0ddc03),
	.w5(32'hbce76308),
	.w6(32'hbb4a8419),
	.w7(32'hbb28d62f),
	.w8(32'hbc2788dc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbca94),
	.w1(32'hbc6d4298),
	.w2(32'hbbebf1cd),
	.w3(32'hbbc3374c),
	.w4(32'hbc761442),
	.w5(32'hbca5aeb4),
	.w6(32'h3a85d2c5),
	.w7(32'h3c6f9f03),
	.w8(32'hbb9a5269),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ee136),
	.w1(32'hb98f53b5),
	.w2(32'h3c0f6c6b),
	.w3(32'h3c23dcb6),
	.w4(32'h3a2f15a5),
	.w5(32'h3c20f3ef),
	.w6(32'h3bc04631),
	.w7(32'h3c60116e),
	.w8(32'h3b818f57),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46d563),
	.w1(32'hbbe1236b),
	.w2(32'hbb8ca15c),
	.w3(32'hbba3e2e2),
	.w4(32'h3aa35693),
	.w5(32'hbc2615ac),
	.w6(32'hbadc9a24),
	.w7(32'hbbfbd34d),
	.w8(32'hbbc086c9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0925fe),
	.w1(32'h3c40fb29),
	.w2(32'h3b76fc54),
	.w3(32'hbc59af65),
	.w4(32'h3bdf633c),
	.w5(32'hbac610a1),
	.w6(32'hbb33217d),
	.w7(32'h3bc00b20),
	.w8(32'h3b57b966),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule