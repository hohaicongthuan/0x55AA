module layer_10_featuremap_116(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb603aa21),
	.w1(32'h3601bcf0),
	.w2(32'hb68d9624),
	.w3(32'h3367e74b),
	.w4(32'h3743b77b),
	.w5(32'h3518f512),
	.w6(32'hb72b176b),
	.w7(32'hb6426982),
	.w8(32'h36c08bd0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fb4d9),
	.w1(32'h39b957f4),
	.w2(32'h398eded6),
	.w3(32'h39589684),
	.w4(32'h3996b6bf),
	.w5(32'h394a0cf8),
	.w6(32'hb7a01da2),
	.w7(32'h386a012a),
	.w8(32'h3844e8e4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34e2fcc4),
	.w1(32'h36d7bbb0),
	.w2(32'h370c66cb),
	.w3(32'h368a46cf),
	.w4(32'h37068faf),
	.w5(32'h37268305),
	.w6(32'h36812ef7),
	.w7(32'h364e2b43),
	.w8(32'h367e70b9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ef18b0),
	.w1(32'hb702213f),
	.w2(32'hb7cfc4b6),
	.w3(32'h35573a5a),
	.w4(32'h3696aae3),
	.w5(32'h3743c416),
	.w6(32'hb7426177),
	.w7(32'hb711b541),
	.w8(32'hb68e2fdf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b806df),
	.w1(32'h372714dc),
	.w2(32'hb5dbbb5e),
	.w3(32'h3727b9f0),
	.w4(32'h36fba916),
	.w5(32'h36d434b9),
	.w6(32'h3766512e),
	.w7(32'h375e254c),
	.w8(32'h3656a01f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36010428),
	.w1(32'h36a55d90),
	.w2(32'h36b9b9c6),
	.w3(32'h362038ed),
	.w4(32'h368fad17),
	.w5(32'h36eadaad),
	.w6(32'h36bebd3c),
	.w7(32'h370990cf),
	.w8(32'h36ba0623),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9182845),
	.w1(32'hb9ce9d6f),
	.w2(32'hba2d3fb7),
	.w3(32'hb95da84d),
	.w4(32'hb93f5196),
	.w5(32'hb98d6e84),
	.w6(32'hb75e68c0),
	.w7(32'h37c8b71f),
	.w8(32'hb8af5817),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f47f26),
	.w1(32'hba09e6a5),
	.w2(32'hba13a33c),
	.w3(32'h38ab5cd9),
	.w4(32'hb8a14333),
	.w5(32'hba126bac),
	.w6(32'hb9bd8f5d),
	.w7(32'h3901af55),
	.w8(32'hb92f4312),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38164b1c),
	.w1(32'h37854afd),
	.w2(32'hb84d1207),
	.w3(32'h3829e009),
	.w4(32'h381b5414),
	.w5(32'hb8130d47),
	.w6(32'h37de973a),
	.w7(32'h383f2b41),
	.w8(32'h37f9caac),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983ef48),
	.w1(32'hb98bb2d4),
	.w2(32'hb9d6265b),
	.w3(32'hb9d455bc),
	.w4(32'hb9b96025),
	.w5(32'hb9b0e529),
	.w6(32'hb89cf8b6),
	.w7(32'h38a74325),
	.w8(32'h38c9b9d9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3836d224),
	.w1(32'h3837e3bb),
	.w2(32'hb7f01316),
	.w3(32'hb72ba1e8),
	.w4(32'hb8a0b49b),
	.w5(32'hb7708f02),
	.w6(32'hb8d4440e),
	.w7(32'hb91c5e9e),
	.w8(32'h3782046b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c71fe),
	.w1(32'hb9bcefd8),
	.w2(32'hba0866ca),
	.w3(32'hb957edf8),
	.w4(32'hb9db10b4),
	.w5(32'hb7adee8c),
	.w6(32'hb9889827),
	.w7(32'hb926f11b),
	.w8(32'h3915a391),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e84b3),
	.w1(32'hba20c3d8),
	.w2(32'hba08b33a),
	.w3(32'hba11c3e5),
	.w4(32'hba0fc00f),
	.w5(32'hba0f6e1a),
	.w6(32'hb9757662),
	.w7(32'h37882621),
	.w8(32'h37d6d377),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389602e7),
	.w1(32'h38d0bf88),
	.w2(32'h38b49172),
	.w3(32'hb7d56b7f),
	.w4(32'hb7d6700b),
	.w5(32'h378cc12f),
	.w6(32'h38134046),
	.w7(32'h3811d941),
	.w8(32'h38bf8291),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b1a51),
	.w1(32'h3916961b),
	.w2(32'h37d59124),
	.w3(32'h392fcf56),
	.w4(32'h3940f3b4),
	.w5(32'h38f3668c),
	.w6(32'h36e56804),
	.w7(32'h391e9880),
	.w8(32'h38f3f0ed),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5c9cf),
	.w1(32'h39032796),
	.w2(32'h3900887e),
	.w3(32'hb9889297),
	.w4(32'hb8b96ad1),
	.w5(32'hb9c7f4a9),
	.w6(32'hb954bce7),
	.w7(32'h38921b6d),
	.w8(32'hb70573d5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3852559d),
	.w1(32'h36a66b5d),
	.w2(32'hb6eb6b5c),
	.w3(32'h3704350a),
	.w4(32'hb88078d4),
	.w5(32'hb888938e),
	.w6(32'hb80b3252),
	.w7(32'hb843e9ae),
	.w8(32'hb7ae4b5c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04af31),
	.w1(32'hba450ab8),
	.w2(32'hba67fece),
	.w3(32'hb9e2a09a),
	.w4(32'hb98d4d5e),
	.w5(32'hba1b446b),
	.w6(32'hb8deaae3),
	.w7(32'hb89e1d68),
	.w8(32'hb98e477a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfeb1e),
	.w1(32'hb9cad64c),
	.w2(32'hb9fc992c),
	.w3(32'hb9a63e1b),
	.w4(32'hb9830001),
	.w5(32'hb9bbae47),
	.w6(32'hb8bc2653),
	.w7(32'h38508221),
	.w8(32'hb839516d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a5b052),
	.w1(32'h35b52b60),
	.w2(32'h367837a2),
	.w3(32'h367ee77f),
	.w4(32'hb6b59cb3),
	.w5(32'hb4e7a7b2),
	.w6(32'hb714983f),
	.w7(32'h36e3a781),
	.w8(32'h359f04ad),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6efe53c),
	.w1(32'hb62f5f33),
	.w2(32'hb70262dc),
	.w3(32'hb68e8f78),
	.w4(32'hb5e9ac96),
	.w5(32'h35e57d4b),
	.w6(32'hb4907f38),
	.w7(32'h36706fae),
	.w8(32'h35dbd88b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e66261),
	.w1(32'h3803429d),
	.w2(32'h381426e2),
	.w3(32'h388d7db8),
	.w4(32'h37c87286),
	.w5(32'h37d560e8),
	.w6(32'h36f76faf),
	.w7(32'hb50600dc),
	.w8(32'h379ffb9c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb5586),
	.w1(32'hb92c5536),
	.w2(32'hb9838a50),
	.w3(32'hba7494e7),
	.w4(32'hb92270cc),
	.w5(32'hba041997),
	.w6(32'hb9c2f4ca),
	.w7(32'h39bd1bd1),
	.w8(32'hb9230582),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f23817),
	.w1(32'hb94284bd),
	.w2(32'hb9729dc2),
	.w3(32'hb960f923),
	.w4(32'hb9408974),
	.w5(32'hb9132d5e),
	.w6(32'hb880c95d),
	.w7(32'h36279f29),
	.w8(32'h384fed0e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f0b89),
	.w1(32'h3a086fc2),
	.w2(32'h39c91efb),
	.w3(32'h394b7b6d),
	.w4(32'h3a3058fa),
	.w5(32'h39ff2f22),
	.w6(32'hb7a9ab8b),
	.w7(32'h398f2614),
	.w8(32'h396baea2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f5cdd),
	.w1(32'h37333b13),
	.w2(32'hb7c9498a),
	.w3(32'h3825c9c0),
	.w4(32'h36d40f90),
	.w5(32'hb78b587b),
	.w6(32'h37bfb8be),
	.w7(32'h37ee72e1),
	.w8(32'h37098955),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61e06f4),
	.w1(32'hb6ff9867),
	.w2(32'h363b980d),
	.w3(32'h36fa7475),
	.w4(32'h367fd3b0),
	.w5(32'h376340ef),
	.w6(32'hb69d9cfd),
	.w7(32'h34e51f04),
	.w8(32'h369329b1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a69185),
	.w1(32'hb904fbcc),
	.w2(32'hb8ea6838),
	.w3(32'h392628c9),
	.w4(32'h39534de5),
	.w5(32'h37d1f3db),
	.w6(32'hb9c57cb5),
	.w7(32'hb96a7446),
	.w8(32'hba294d9a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4bbe9),
	.w1(32'hb88cf560),
	.w2(32'hb748b928),
	.w3(32'hb8a9efed),
	.w4(32'hb8a7e1a0),
	.w5(32'h38158def),
	.w6(32'hb93a5600),
	.w7(32'hb8fb7bdb),
	.w8(32'hb824ef97),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd914d),
	.w1(32'h393afca9),
	.w2(32'h37948e4a),
	.w3(32'h39f9eb2b),
	.w4(32'h3a142b3a),
	.w5(32'h399861e5),
	.w6(32'hb84f769a),
	.w7(32'h38350f33),
	.w8(32'hb54bde34),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb52e3a2a),
	.w1(32'hb608441e),
	.w2(32'h36362761),
	.w3(32'hb70af3d5),
	.w4(32'hb6d64ef8),
	.w5(32'h356f8807),
	.w6(32'hb6fb1e85),
	.w7(32'h357b1ee5),
	.w8(32'h3690631b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3601b1cb),
	.w1(32'h36dc87c1),
	.w2(32'hb75d0c20),
	.w3(32'h375c5900),
	.w4(32'hb73fd71b),
	.w5(32'hb822c818),
	.w6(32'hb79830ce),
	.w7(32'hb7b7c932),
	.w8(32'hb7cbe3f7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91328c5),
	.w1(32'hb92f8616),
	.w2(32'hb9657654),
	.w3(32'hb9816507),
	.w4(32'hb9898a6b),
	.w5(32'hb958b7d6),
	.w6(32'hb9032b74),
	.w7(32'hb8738348),
	.w8(32'hb844ce1c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892946c),
	.w1(32'h3934a863),
	.w2(32'h391b004d),
	.w3(32'h38f431e0),
	.w4(32'h39344813),
	.w5(32'h39178c5a),
	.w6(32'h37b21b75),
	.w7(32'h380af10b),
	.w8(32'h389b5886),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84875d2),
	.w1(32'hb848a522),
	.w2(32'hb7f97453),
	.w3(32'hb8ae091d),
	.w4(32'hb8ab0b46),
	.w5(32'h370f9f2b),
	.w6(32'hb8613f2e),
	.w7(32'hb87b585e),
	.w8(32'hb85a03f5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911d4d6),
	.w1(32'hb99ab6b4),
	.w2(32'hb9b7fed8),
	.w3(32'hb92bc22d),
	.w4(32'hb8fcad50),
	.w5(32'hb925ae83),
	.w6(32'hb861f0a2),
	.w7(32'hb81c4710),
	.w8(32'hb8800274),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acca3b),
	.w1(32'h3a64892b),
	.w2(32'h38e8bf56),
	.w3(32'h3a05ec09),
	.w4(32'h3907c364),
	.w5(32'hb81d26c7),
	.w6(32'h38e72f93),
	.w7(32'h39a0d931),
	.w8(32'h3a36d898),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d60a2),
	.w1(32'h38af7728),
	.w2(32'h39781fd9),
	.w3(32'h395a53d4),
	.w4(32'h39fb54f8),
	.w5(32'h3a2ac95a),
	.w6(32'hb94d45ce),
	.w7(32'h39408794),
	.w8(32'h390e1d2d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae49de),
	.w1(32'h39d2ca0f),
	.w2(32'h3a699d48),
	.w3(32'h3a074b67),
	.w4(32'h3a491363),
	.w5(32'h3a5e3d71),
	.w6(32'h355ce3d9),
	.w7(32'h394040c4),
	.w8(32'h39ab31d9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38667e37),
	.w1(32'h38aaf241),
	.w2(32'h37830ada),
	.w3(32'h38e32603),
	.w4(32'h38df00cc),
	.w5(32'h388381db),
	.w6(32'hb7a47fef),
	.w7(32'h37c8ac4a),
	.w8(32'h38425c24),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4c998),
	.w1(32'hb80ccec4),
	.w2(32'hb74bf368),
	.w3(32'h384e1756),
	.w4(32'hb7b6cf56),
	.w5(32'hb7160fb0),
	.w6(32'hb744b13f),
	.w7(32'hb783b080),
	.w8(32'hb6d2f00a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fa8888),
	.w1(32'hb88e1668),
	.w2(32'h37b35d55),
	.w3(32'hb6d3fe39),
	.w4(32'hb7c6e45b),
	.w5(32'hb60cd024),
	.w6(32'h3818d968),
	.w7(32'h37e9bd25),
	.w8(32'hb7e76133),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38992015),
	.w1(32'h38b01e8e),
	.w2(32'h3924bf27),
	.w3(32'h390f1a8d),
	.w4(32'h386d84e4),
	.w5(32'h394d175e),
	.w6(32'h38d1b2e5),
	.w7(32'h382d630c),
	.w8(32'h391c4701),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba305b2b),
	.w1(32'hba8da2f3),
	.w2(32'hb9bb1e45),
	.w3(32'hba507ba9),
	.w4(32'hba3f464f),
	.w5(32'hb98c60b1),
	.w6(32'hb9a5ed8d),
	.w7(32'hb8dfdc94),
	.w8(32'hb8734eaf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925f027),
	.w1(32'hb8301cd4),
	.w2(32'h38822f08),
	.w3(32'hb8076f13),
	.w4(32'h391bc52c),
	.w5(32'h38dcb4e1),
	.w6(32'hb8b89971),
	.w7(32'h39026dea),
	.w8(32'h38dfe5e4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a6cdf),
	.w1(32'hb95a28b8),
	.w2(32'hb95c4daf),
	.w3(32'hb981e814),
	.w4(32'h38fd278e),
	.w5(32'h3937de0f),
	.w6(32'hb86b7f70),
	.w7(32'h389b813a),
	.w8(32'h38ffef1a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea7ced),
	.w1(32'hb91793fa),
	.w2(32'h39862b68),
	.w3(32'hb8fd13a2),
	.w4(32'hb91d7935),
	.w5(32'h378a3823),
	.w6(32'hb8f27840),
	.w7(32'h36aa7826),
	.w8(32'h3919489e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c7b12),
	.w1(32'hba7da558),
	.w2(32'hba94426c),
	.w3(32'hba1c42ff),
	.w4(32'hba6c366e),
	.w5(32'hba8cc03b),
	.w6(32'hb9b27943),
	.w7(32'hb98c6daf),
	.w8(32'hb9577deb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70e5aaa),
	.w1(32'hb8f361db),
	.w2(32'h3811b402),
	.w3(32'h362dd32d),
	.w4(32'hb87da1e5),
	.w5(32'h38c3c9b4),
	.w6(32'hb720ecda),
	.w7(32'h37de0122),
	.w8(32'h384dae52),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37995d39),
	.w1(32'hb76b9c4f),
	.w2(32'h3896940e),
	.w3(32'h385c76af),
	.w4(32'h3731a062),
	.w5(32'h37074b3f),
	.w6(32'h3896adda),
	.w7(32'h386c7b72),
	.w8(32'h3912ee4d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ba62e),
	.w1(32'hb843c04c),
	.w2(32'h35039926),
	.w3(32'h38c0579c),
	.w4(32'h39063a9d),
	.w5(32'h38c32ead),
	.w6(32'h390315f3),
	.w7(32'h39067024),
	.w8(32'h38aa0ca7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906e07c),
	.w1(32'h38243fe3),
	.w2(32'h37dbf1fe),
	.w3(32'hb93852e5),
	.w4(32'hb78ce762),
	.w5(32'h392e0884),
	.w6(32'hb84ac674),
	.w7(32'h38fe717b),
	.w8(32'h38a3f76f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374894ac),
	.w1(32'hb790d45a),
	.w2(32'hb8898539),
	.w3(32'hb72bd1ea),
	.w4(32'hb840e812),
	.w5(32'hb881fff6),
	.w6(32'h372f07dc),
	.w7(32'h37576e8f),
	.w8(32'hb88261a9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f994d),
	.w1(32'hba20a19b),
	.w2(32'hba244988),
	.w3(32'hba109c0c),
	.w4(32'hba2074a3),
	.w5(32'hba214120),
	.w6(32'hb9685809),
	.w7(32'hb8d19f5d),
	.w8(32'hb930a520),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a844d),
	.w1(32'hb9818d61),
	.w2(32'hb89ca3bf),
	.w3(32'hb8be191a),
	.w4(32'h375e787b),
	.w5(32'h3419c568),
	.w6(32'hb91ef2ec),
	.w7(32'hb8a9ceff),
	.w8(32'hb8d6e20f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378c7841),
	.w1(32'h37c6c9f0),
	.w2(32'h37c9a547),
	.w3(32'h37e934fa),
	.w4(32'h37b7d826),
	.w5(32'h3795672d),
	.w6(32'hb708a9df),
	.w7(32'h376aa649),
	.w8(32'hb683e944),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3588b164),
	.w1(32'h36e96940),
	.w2(32'h3701aa65),
	.w3(32'hb62f377b),
	.w4(32'h37404124),
	.w5(32'h37244859),
	.w6(32'h347531ae),
	.w7(32'h3621025a),
	.w8(32'h36424dcc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7341e90),
	.w1(32'hb6dcfa93),
	.w2(32'hb7563cb2),
	.w3(32'hb611dec3),
	.w4(32'h36cf355b),
	.w5(32'hb68d50da),
	.w6(32'hb71c3d55),
	.w7(32'h35f4df37),
	.w8(32'hb6e3cd3d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d3786),
	.w1(32'h380bc888),
	.w2(32'h38e25bdb),
	.w3(32'hb6db3034),
	.w4(32'h382f938a),
	.w5(32'h38d7e3dc),
	.w6(32'h38007b62),
	.w7(32'h3846dd26),
	.w8(32'h38d45e2e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a42a1a),
	.w1(32'hb88c20ec),
	.w2(32'hb885f4be),
	.w3(32'hb875bab2),
	.w4(32'hb89c82da),
	.w5(32'hb70877f1),
	.w6(32'hb7e4ec9d),
	.w7(32'h37c627b1),
	.w8(32'h372a4a9a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964d068),
	.w1(32'hb9849501),
	.w2(32'hb997c839),
	.w3(32'hb991542c),
	.w4(32'hb96188b0),
	.w5(32'hb922174b),
	.w6(32'hb8a27cf0),
	.w7(32'hb7d2c33d),
	.w8(32'hb8f3259f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac28ab),
	.w1(32'hb9313bf0),
	.w2(32'h394d6f77),
	.w3(32'hb9d5f4cc),
	.w4(32'hb8983eba),
	.w5(32'h389d7ea4),
	.w6(32'hb9babdae),
	.w7(32'hb9071a2e),
	.w8(32'hb8832d78),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68db9c8),
	.w1(32'hb6842500),
	.w2(32'hb6ac2e1d),
	.w3(32'hb419ace9),
	.w4(32'h37246905),
	.w5(32'h361edc21),
	.w6(32'h3718ef17),
	.w7(32'h37231ed2),
	.w8(32'h37221b73),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68e6a45),
	.w1(32'hb4c2305b),
	.w2(32'hb4e52980),
	.w3(32'hb659eef0),
	.w4(32'h366fcb55),
	.w5(32'h363d87df),
	.w6(32'h36a68996),
	.w7(32'h367014fc),
	.w8(32'h36ae12b8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5aca3),
	.w1(32'h376e2c0a),
	.w2(32'h35cd69f4),
	.w3(32'h36cbec2c),
	.w4(32'h3695b5aa),
	.w5(32'hb6929ecd),
	.w6(32'hb70607d0),
	.w7(32'hb5f56447),
	.w8(32'h36298831),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb608bf20),
	.w1(32'h35e96d17),
	.w2(32'hb718a896),
	.w3(32'hb581ef27),
	.w4(32'hb6cb7b2f),
	.w5(32'hb705d0bc),
	.w6(32'hb58cdb8e),
	.w7(32'hb6f89d6c),
	.w8(32'hb7361aca),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4afb96),
	.w1(32'hb9db2c8b),
	.w2(32'hb980dccb),
	.w3(32'hba93c6f8),
	.w4(32'hba5dfed2),
	.w5(32'hba1dfee4),
	.w6(32'hb9f21984),
	.w7(32'hb9a73f41),
	.w8(32'hb917962c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fa9e2),
	.w1(32'hb9cf4076),
	.w2(32'hba01c716),
	.w3(32'hba1f84be),
	.w4(32'h38670764),
	.w5(32'h3888d609),
	.w6(32'hb93d1505),
	.w7(32'hb988fa16),
	.w8(32'hb9e568f8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb19c2),
	.w1(32'hb9e0c942),
	.w2(32'hb93204e6),
	.w3(32'hba0f4e0d),
	.w4(32'hb8c555b0),
	.w5(32'h39051c79),
	.w6(32'hb8fa4c3f),
	.w7(32'hb884f0ea),
	.w8(32'hb90bd6e0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86311cf),
	.w1(32'h39535ea2),
	.w2(32'h3962e1d5),
	.w3(32'h3988c232),
	.w4(32'h3a199637),
	.w5(32'h39f4369d),
	.w6(32'h391fb000),
	.w7(32'h39d655ca),
	.w8(32'h394f2f25),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bb13b4),
	.w1(32'hb68acf86),
	.w2(32'hb6eabce1),
	.w3(32'h372ce96b),
	.w4(32'h3618ab90),
	.w5(32'hb5dae74e),
	.w6(32'hb6929464),
	.w7(32'hb6f235a7),
	.w8(32'hb67b9ce7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3595f079),
	.w1(32'hb4e4eb45),
	.w2(32'h35d87d2c),
	.w3(32'h36b033ee),
	.w4(32'hb67b33be),
	.w5(32'hb5711267),
	.w6(32'h359aa96c),
	.w7(32'h34fc461b),
	.w8(32'hb514c7cd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e5258b),
	.w1(32'hb6d62915),
	.w2(32'hb5e4d1f0),
	.w3(32'hb7064470),
	.w4(32'hb6a85557),
	.w5(32'hb66e87a6),
	.w6(32'h35d0d81f),
	.w7(32'h368ff6e5),
	.w8(32'hb64070b1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949ea23),
	.w1(32'hb9830e00),
	.w2(32'hb96437e3),
	.w3(32'hb940e770),
	.w4(32'hb9582776),
	.w5(32'hb9618e05),
	.w6(32'hb90bd4c0),
	.w7(32'hb8dca3fa),
	.w8(32'hb8bc097a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81323cf),
	.w1(32'hb88c2049),
	.w2(32'hb7599af1),
	.w3(32'hb717b938),
	.w4(32'hb76507d1),
	.w5(32'h37987fcc),
	.w6(32'h33db0efb),
	.w7(32'h36f43195),
	.w8(32'h37b8cdf7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a0711),
	.w1(32'hb98a3c90),
	.w2(32'hb99bf129),
	.w3(32'hb90a2ba8),
	.w4(32'hb9b59814),
	.w5(32'hb9c74d89),
	.w6(32'hb896744b),
	.w7(32'h376e0990),
	.w8(32'h383397b8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9902b17),
	.w1(32'hb9a388ad),
	.w2(32'hb9ebf895),
	.w3(32'hb925cf35),
	.w4(32'hb928fa28),
	.w5(32'hba03e121),
	.w6(32'hb9574762),
	.w7(32'h383b5d04),
	.w8(32'hb92524b2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952d3e6),
	.w1(32'h398b1aac),
	.w2(32'h393672c9),
	.w3(32'hb8ab61fe),
	.w4(32'h395542d5),
	.w5(32'h38d0d1a9),
	.w6(32'hb97eccb0),
	.w7(32'h3906d9e6),
	.w8(32'h38f9e291),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952a4aa),
	.w1(32'hb95acf78),
	.w2(32'hb92d2a49),
	.w3(32'hb930f6f3),
	.w4(32'hb8b36723),
	.w5(32'hb93e2e50),
	.w6(32'hb87a2ec4),
	.w7(32'h3777a4be),
	.w8(32'hb7b405d7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98235b7),
	.w1(32'hb8eaafba),
	.w2(32'hb41c320c),
	.w3(32'hb9cdd845),
	.w4(32'hb9bb6acf),
	.w5(32'hb88f3380),
	.w6(32'hb959a9de),
	.w7(32'hb88df2e0),
	.w8(32'hb885649a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5e1d0),
	.w1(32'h3851d6ed),
	.w2(32'h394fb31c),
	.w3(32'hb834e948),
	.w4(32'h37ea484e),
	.w5(32'h38b35b70),
	.w6(32'hb901381a),
	.w7(32'h37626d7c),
	.w8(32'h38824e2a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fef18),
	.w1(32'hb99ee039),
	.w2(32'hb9aa521f),
	.w3(32'hb97380dd),
	.w4(32'hb997ac72),
	.w5(32'hb99c31c1),
	.w6(32'hb9131588),
	.w7(32'hb87e568b),
	.w8(32'hb7f4543c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fc6277),
	.w1(32'hb71a49a7),
	.w2(32'hb67f3651),
	.w3(32'h36314cb2),
	.w4(32'hb6ed02a9),
	.w5(32'hb6329871),
	.w6(32'hb75a9f90),
	.w7(32'hb710c16c),
	.w8(32'hb7656741),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f0a9c),
	.w1(32'h369bbdb9),
	.w2(32'hb508dca1),
	.w3(32'hb68745be),
	.w4(32'h36a9a06f),
	.w5(32'h357f2072),
	.w6(32'hb63e885f),
	.w7(32'hb67b5e43),
	.w8(32'h354608d9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb50c496a),
	.w1(32'hb71ea5a1),
	.w2(32'h369757d3),
	.w3(32'hb42014ef),
	.w4(32'hb786c518),
	.w5(32'h36eaf99e),
	.w6(32'hb790fcbf),
	.w7(32'hb5ee79e1),
	.w8(32'h3651adeb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ded66a),
	.w1(32'h3799b96e),
	.w2(32'h37d5f5a6),
	.w3(32'h38279ea9),
	.w4(32'h382b3150),
	.w5(32'h3829507f),
	.w6(32'hb70adebb),
	.w7(32'h3704818c),
	.w8(32'h37379718),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ea312),
	.w1(32'h39829f08),
	.w2(32'h3976f8f9),
	.w3(32'h392d1d6f),
	.w4(32'h3982abcf),
	.w5(32'h398087c1),
	.w6(32'hb7af3902),
	.w7(32'h3840a132),
	.w8(32'h38d089f1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3719b5eb),
	.w1(32'hb6e1df32),
	.w2(32'h38011ece),
	.w3(32'h36f133bc),
	.w4(32'hb7914cc6),
	.w5(32'h3817bdbc),
	.w6(32'hb7945bc1),
	.w7(32'hb7cb15d5),
	.w8(32'h37cb9284),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36eeb784),
	.w1(32'hb73056db),
	.w2(32'hb6f8e22f),
	.w3(32'hb7f10bd6),
	.w4(32'h395f10f8),
	.w5(32'h38c2ad80),
	.w6(32'h38950f8d),
	.w7(32'h39062497),
	.w8(32'hb8c77baf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05dce7),
	.w1(32'hb9baa377),
	.w2(32'hb9d10055),
	.w3(32'hb9beed56),
	.w4(32'hb9b917c7),
	.w5(32'hb9e12060),
	.w6(32'hb9825468),
	.w7(32'hb91e41ba),
	.w8(32'hb8cdedf3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91be7f7),
	.w1(32'h3894f1ab),
	.w2(32'h392a3629),
	.w3(32'h385601d2),
	.w4(32'h3920cf6a),
	.w5(32'h398f6d84),
	.w6(32'hb96f9687),
	.w7(32'hb9019213),
	.w8(32'h3866c53f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9785b77),
	.w1(32'hb99f5d59),
	.w2(32'hb936012d),
	.w3(32'hba15938c),
	.w4(32'hba0d530a),
	.w5(32'hba1a61fd),
	.w6(32'hb9ab8cda),
	.w7(32'h38939d11),
	.w8(32'h380d3243),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9265dbd),
	.w1(32'hb8922eb7),
	.w2(32'hb8a79bf3),
	.w3(32'h375779e2),
	.w4(32'h38f593f9),
	.w5(32'h38d35ec1),
	.w6(32'h38fe2ff0),
	.w7(32'h39788255),
	.w8(32'h394a12cc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3718b),
	.w1(32'hb95d43f1),
	.w2(32'hb7b91dcb),
	.w3(32'hb9ab45ad),
	.w4(32'hb91ad382),
	.w5(32'hb961eab8),
	.w6(32'hb919bbcf),
	.w7(32'h37b1535e),
	.w8(32'h37caefda),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d9532),
	.w1(32'h39953882),
	.w2(32'h39b82c12),
	.w3(32'hb5dbdcbc),
	.w4(32'h393cb04a),
	.w5(32'h3929a88b),
	.w6(32'hb834cbff),
	.w7(32'h3900660d),
	.w8(32'h391ec8f4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38735009),
	.w1(32'h3961bf46),
	.w2(32'h3905da2b),
	.w3(32'h396b9584),
	.w4(32'h399e8bab),
	.w5(32'h396b7007),
	.w6(32'hb9741ac6),
	.w7(32'h377d8603),
	.w8(32'h389f8522),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885bd20),
	.w1(32'h37eb400e),
	.w2(32'hb6c05f90),
	.w3(32'h389df3a2),
	.w4(32'h3880091c),
	.w5(32'h38448651),
	.w6(32'h388777a2),
	.w7(32'h383cf4aa),
	.w8(32'h3823eabc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f27624),
	.w1(32'hb9aac4c8),
	.w2(32'hb9647ebc),
	.w3(32'hb85d51a5),
	.w4(32'h3870950a),
	.w5(32'hb90f5d1e),
	.w6(32'h39517de8),
	.w7(32'h39b8b18f),
	.w8(32'h380bc3b9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b000c2),
	.w1(32'hb9b389c7),
	.w2(32'h37b6c0b7),
	.w3(32'hb927875f),
	.w4(32'hb92a12ba),
	.w5(32'h397c9b21),
	.w6(32'h396ac4da),
	.w7(32'h398e5ef8),
	.w8(32'h3a3cdb18),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82f9ec5),
	.w1(32'h3864276d),
	.w2(32'hba3c8695),
	.w3(32'hb9eedeb7),
	.w4(32'hb81477e6),
	.w5(32'hb8dfe0a8),
	.w6(32'hba13c1af),
	.w7(32'h3933f656),
	.w8(32'h39c6e276),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913260e),
	.w1(32'h39467353),
	.w2(32'h3a122527),
	.w3(32'h39562a44),
	.w4(32'h39985fca),
	.w5(32'h3a265c75),
	.w6(32'hb889441d),
	.w7(32'h39439a50),
	.w8(32'h39ebac58),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0971f),
	.w1(32'h39b0616c),
	.w2(32'h391f1a2e),
	.w3(32'h39393790),
	.w4(32'h39facae3),
	.w5(32'h38d6acb0),
	.w6(32'h39a7ae47),
	.w7(32'h39f83ac4),
	.w8(32'h39d4fa8b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391263f2),
	.w1(32'hb9b40f2e),
	.w2(32'hb95ebd10),
	.w3(32'hb999e34e),
	.w4(32'hb9d511e1),
	.w5(32'hb990131c),
	.w6(32'hb9bef69e),
	.w7(32'h394de891),
	.w8(32'h39969a09),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be305d),
	.w1(32'hb942ab10),
	.w2(32'h38ab584e),
	.w3(32'h3890a8e9),
	.w4(32'h38b82bbd),
	.w5(32'h39472a82),
	.w6(32'h3999b528),
	.w7(32'h399c1a76),
	.w8(32'h3964715a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb9c7e),
	.w1(32'h399d3ccd),
	.w2(32'hb9ef5d88),
	.w3(32'hb90e4679),
	.w4(32'h39303836),
	.w5(32'hb7e98e24),
	.w6(32'hb9a42198),
	.w7(32'h38fecb63),
	.w8(32'h39edec11),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93209fc),
	.w1(32'hb9673fe4),
	.w2(32'hb907cb47),
	.w3(32'hb986e3d4),
	.w4(32'hb8f1f860),
	.w5(32'h387c2546),
	.w6(32'hb951ac3f),
	.w7(32'h37411113),
	.w8(32'h384b97b8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a2abcf),
	.w1(32'h38114bbe),
	.w2(32'h37fbc63e),
	.w3(32'h37676e40),
	.w4(32'h38086879),
	.w5(32'h37c3e039),
	.w6(32'h36b748cc),
	.w7(32'h37ad9485),
	.w8(32'h37448e80),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb822942b),
	.w1(32'h3958d4f9),
	.w2(32'h3914c377),
	.w3(32'h36b056c1),
	.w4(32'h3788aca2),
	.w5(32'h38d30b2e),
	.w6(32'hb7d1bcb2),
	.w7(32'h37d21c15),
	.w8(32'hb792dbca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6e661),
	.w1(32'hb99abdfd),
	.w2(32'hb997a3f4),
	.w3(32'hb8c22329),
	.w4(32'hb950e64e),
	.w5(32'hb9a2c21f),
	.w6(32'h39232fc7),
	.w7(32'h39137cb0),
	.w8(32'h38c859f1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9369e1d),
	.w1(32'h389e5904),
	.w2(32'h37eacad7),
	.w3(32'hb8860bf6),
	.w4(32'h39531388),
	.w5(32'h392d5435),
	.w6(32'hb8879e8f),
	.w7(32'h39375563),
	.w8(32'h3900fa1c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f48f3),
	.w1(32'hb5dfdd67),
	.w2(32'h38dd6278),
	.w3(32'h38d56907),
	.w4(32'h3885eb75),
	.w5(32'h38e4837a),
	.w6(32'hb8eff351),
	.w7(32'hb79ef0d6),
	.w8(32'hb89cafa3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f7e8a6),
	.w1(32'h38c16883),
	.w2(32'h3927e6c2),
	.w3(32'h395c1670),
	.w4(32'h398cf209),
	.w5(32'h381740d4),
	.w6(32'h392183e2),
	.w7(32'h397dfcab),
	.w8(32'h392379d0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d10a48),
	.w1(32'hb9ce28bf),
	.w2(32'hb9876351),
	.w3(32'hb9c799f1),
	.w4(32'h39214e4b),
	.w5(32'h3904dbba),
	.w6(32'hb9a42b7c),
	.w7(32'hb918b85c),
	.w8(32'h38436935),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6ee9b),
	.w1(32'h39274f8b),
	.w2(32'h394b2719),
	.w3(32'hb9b3314e),
	.w4(32'hb8a11022),
	.w5(32'hb981acb1),
	.w6(32'hb9a4408c),
	.w7(32'hb88ed1a2),
	.w8(32'hb5f83143),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8151e55),
	.w1(32'hb70727c7),
	.w2(32'h3767ed5f),
	.w3(32'hb8248c2f),
	.w4(32'h385ec07c),
	.w5(32'h38818ef2),
	.w6(32'h37c1ab6b),
	.w7(32'h38c0a927),
	.w8(32'h38afbead),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3670fb64),
	.w1(32'hb5e6083a),
	.w2(32'hb6001767),
	.w3(32'h36a8c4f4),
	.w4(32'hb6b2fd45),
	.w5(32'hb651ea6f),
	.w6(32'h3664ac97),
	.w7(32'h36bad0a1),
	.w8(32'h368e8504),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a9cfef),
	.w1(32'h38c7336e),
	.w2(32'h38463f08),
	.w3(32'hb77bc22b),
	.w4(32'h381ff623),
	.w5(32'hb62d3390),
	.w6(32'hb7d677c7),
	.w7(32'h38076e84),
	.w8(32'hb703d75f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3687675f),
	.w1(32'h362b147f),
	.w2(32'hb6177362),
	.w3(32'h36c24c91),
	.w4(32'h36bafa05),
	.w5(32'h360d77c4),
	.w6(32'h36f025d0),
	.w7(32'h3716607e),
	.w8(32'h370c82cd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3720db8),
	.w1(32'h3709e16f),
	.w2(32'h36231fb0),
	.w3(32'hb6a221ee),
	.w4(32'hb5940c57),
	.w5(32'hb75f0219),
	.w6(32'hb6792692),
	.w7(32'hb67a8e47),
	.w8(32'h3780f020),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9067798),
	.w1(32'hb8381ed2),
	.w2(32'h368eacfc),
	.w3(32'hb8f674a5),
	.w4(32'h38ab9d6c),
	.w5(32'h38f55f3b),
	.w6(32'hb8b62828),
	.w7(32'h388adfcb),
	.w8(32'h38ad5334),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb745dc35),
	.w1(32'hb82d3cd6),
	.w2(32'hb8079ab0),
	.w3(32'hb7ef98f0),
	.w4(32'hb86ac530),
	.w5(32'hb7f67235),
	.w6(32'hb790109c),
	.w7(32'hb7fbca39),
	.w8(32'hb5ed824a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cd8d3),
	.w1(32'hb99c3f57),
	.w2(32'hb99e7527),
	.w3(32'hb9755aef),
	.w4(32'hb983d9c8),
	.w5(32'hb9760aa4),
	.w6(32'hb93e336a),
	.w7(32'hb89b3cdb),
	.w8(32'hb7f2cdbd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38977f76),
	.w1(32'h39c85f4e),
	.w2(32'h39bca5d2),
	.w3(32'h3991f71b),
	.w4(32'h39de66cb),
	.w5(32'h399b3ccc),
	.w6(32'hb92d3b7f),
	.w7(32'h38764ff2),
	.w8(32'h386b3954),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3577cdb6),
	.w1(32'h378ac19a),
	.w2(32'h371180ba),
	.w3(32'h36712043),
	.w4(32'h372e3644),
	.w5(32'hb67d6798),
	.w6(32'h370ccf1b),
	.w7(32'h3793f50d),
	.w8(32'h37ed4f73),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38149b0c),
	.w1(32'h35cb44bd),
	.w2(32'h35c41ba4),
	.w3(32'h36465ed6),
	.w4(32'hb527de3e),
	.w5(32'h34965dcc),
	.w6(32'h37304327),
	.w7(32'h360c0a65),
	.w8(32'h3686172a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74969d2),
	.w1(32'hb5f17d8e),
	.w2(32'h37845176),
	.w3(32'hb6afbeac),
	.w4(32'hb6533cdb),
	.w5(32'h37550e9e),
	.w6(32'hb7693a9b),
	.w7(32'h350d8c3c),
	.w8(32'h3715d6a6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3713ac7c),
	.w1(32'h397858c1),
	.w2(32'hba96b85e),
	.w3(32'hb595e27e),
	.w4(32'hba01db0d),
	.w5(32'hbababd80),
	.w6(32'h3a208f44),
	.w7(32'hbab88026),
	.w8(32'hba0de717),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d07ad),
	.w1(32'h388e7eeb),
	.w2(32'hba3b780b),
	.w3(32'hb9c37989),
	.w4(32'h39a227fa),
	.w5(32'hba1db73b),
	.w6(32'h39542057),
	.w7(32'hb98a0644),
	.w8(32'h3a18d766),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b8bb6),
	.w1(32'h3aa5f9ec),
	.w2(32'h3a846710),
	.w3(32'hb8d5d8b1),
	.w4(32'h3a1196cf),
	.w5(32'hb916a057),
	.w6(32'hbae7671e),
	.w7(32'hb9885e19),
	.w8(32'hbaa4cef4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fc6ef),
	.w1(32'h3a279e97),
	.w2(32'h390ea2de),
	.w3(32'hbaa45f2d),
	.w4(32'hb858a9e9),
	.w5(32'hb92fbf11),
	.w6(32'h3a20056f),
	.w7(32'h3a17a5fa),
	.w8(32'hb8baf5d6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9caf0ac),
	.w1(32'hba3b8dbb),
	.w2(32'hba0d04ca),
	.w3(32'hba99b5d5),
	.w4(32'hba62f0ca),
	.w5(32'hba27c3cd),
	.w6(32'hba0a0c89),
	.w7(32'hb979f1b3),
	.w8(32'hb903e58f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e0c8c),
	.w1(32'h3a999eba),
	.w2(32'h3a8920e6),
	.w3(32'hb9f18c5f),
	.w4(32'h3a735053),
	.w5(32'h39d36070),
	.w6(32'h39e3f584),
	.w7(32'hba37dc2f),
	.w8(32'hbae2d873),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba674a),
	.w1(32'h3afbabc6),
	.w2(32'h3b2b61b2),
	.w3(32'hba8b9c6f),
	.w4(32'h3b308427),
	.w5(32'h3b30ed9b),
	.w6(32'h3af7feb6),
	.w7(32'h3ac73e4e),
	.w8(32'h3ad20983),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd6372),
	.w1(32'h3a56daf5),
	.w2(32'hb94220d0),
	.w3(32'h3af97093),
	.w4(32'h398ab873),
	.w5(32'hba9431b1),
	.w6(32'hb8e09916),
	.w7(32'hbab776f1),
	.w8(32'h39b7a495),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7df4d6e),
	.w1(32'hba9dc910),
	.w2(32'hbad542b8),
	.w3(32'hb96b2554),
	.w4(32'hba9f25ba),
	.w5(32'hba7869cd),
	.w6(32'hbad01013),
	.w7(32'hbabf56bf),
	.w8(32'hba11945d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8d399),
	.w1(32'h3adb33d9),
	.w2(32'h399321dc),
	.w3(32'hba783b0d),
	.w4(32'h3a8f0122),
	.w5(32'hb85e1923),
	.w6(32'h3a5ce1f0),
	.w7(32'hb90ff126),
	.w8(32'h3a27b855),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacd510),
	.w1(32'h39a923c4),
	.w2(32'hba3e4487),
	.w3(32'h3a1e1600),
	.w4(32'h39a3c1a2),
	.w5(32'hba3f1f8a),
	.w6(32'hb9abd090),
	.w7(32'hba7f9cb4),
	.w8(32'hb73efab9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5f4f3),
	.w1(32'hb9f4bf29),
	.w2(32'hba9bef99),
	.w3(32'h39201517),
	.w4(32'hbaa5d6db),
	.w5(32'hbad18691),
	.w6(32'hba99cda5),
	.w7(32'hbaea2c19),
	.w8(32'hbb11f88b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab132ae),
	.w1(32'hbb70b845),
	.w2(32'hbb96cd62),
	.w3(32'hbab736d0),
	.w4(32'hb8def3ec),
	.w5(32'h39aaf091),
	.w6(32'hb99c3742),
	.w7(32'hb945e833),
	.w8(32'hba4bf31e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd40b6f),
	.w1(32'hb9cde126),
	.w2(32'hb7ebc775),
	.w3(32'hbaebf8bc),
	.w4(32'hba8fd96e),
	.w5(32'hbacae16b),
	.w6(32'hba385429),
	.w7(32'hbade8f25),
	.w8(32'hba80756e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a6ff8),
	.w1(32'hbab1c36a),
	.w2(32'hbabafd3f),
	.w3(32'hba8c89c2),
	.w4(32'hba772ad0),
	.w5(32'hba5bc2aa),
	.w6(32'hb9ef8a4a),
	.w7(32'hb9f119d1),
	.w8(32'hb76c47eb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47a653),
	.w1(32'h3b1814f5),
	.w2(32'hb910bf40),
	.w3(32'h398f4ebd),
	.w4(32'h3b063c73),
	.w5(32'h386ad687),
	.w6(32'h39a57115),
	.w7(32'hba90ea49),
	.w8(32'hba1692ed),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39972fea),
	.w1(32'h39ffcfc7),
	.w2(32'h3ad5ff42),
	.w3(32'h3a05350c),
	.w4(32'h3b3463ee),
	.w5(32'h3ae79e8c),
	.w6(32'h3a25adc6),
	.w7(32'hb93cefe8),
	.w8(32'h3aff4a93),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bd125),
	.w1(32'hb999fa99),
	.w2(32'hba798360),
	.w3(32'h3a83fc76),
	.w4(32'hb970598d),
	.w5(32'hba87924c),
	.w6(32'hb9f83b97),
	.w7(32'hba75f947),
	.w8(32'hb9097bc8),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa1bf8),
	.w1(32'h3a9f6a3a),
	.w2(32'hb9b241ee),
	.w3(32'hb8faa7cf),
	.w4(32'h3b55fbdc),
	.w5(32'h3ad939e3),
	.w6(32'h3b70af9a),
	.w7(32'h3a825411),
	.w8(32'hba805f08),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b7a83),
	.w1(32'hb9a7f4cf),
	.w2(32'hba5220d4),
	.w3(32'hba8fdc42),
	.w4(32'hba848a8e),
	.w5(32'hba094a94),
	.w6(32'hbaa2024e),
	.w7(32'hba565687),
	.w8(32'hba2920a5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba351e34),
	.w1(32'hb8b75d0f),
	.w2(32'h399a1124),
	.w3(32'hba934412),
	.w4(32'hb948d046),
	.w5(32'h3886b0f7),
	.w6(32'h39d83188),
	.w7(32'h3a7156dd),
	.w8(32'h3a978277),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6a930),
	.w1(32'h39901381),
	.w2(32'hba15b69f),
	.w3(32'hb9be3d4e),
	.w4(32'h39842d5d),
	.w5(32'hb9d4f1d3),
	.w6(32'hb8f80db5),
	.w7(32'hba73721b),
	.w8(32'hb958dbaf),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57f916f),
	.w1(32'h3a6f9f27),
	.w2(32'hba94fb12),
	.w3(32'h39636a22),
	.w4(32'hba9f2827),
	.w5(32'hbb29c719),
	.w6(32'h3a00780d),
	.w7(32'hbb2758a9),
	.w8(32'hba9dc93e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f62a05),
	.w1(32'h3a3058ca),
	.w2(32'h3ac43f14),
	.w3(32'hba5c4769),
	.w4(32'h38760e98),
	.w5(32'h3ab792de),
	.w6(32'hba888b11),
	.w7(32'h38e32eab),
	.w8(32'h3a3f494a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09dcf5),
	.w1(32'h3a44ae70),
	.w2(32'hbbb3638c),
	.w3(32'h3a87e5e2),
	.w4(32'h3a5b17ad),
	.w5(32'hbbd0152d),
	.w6(32'h39cda962),
	.w7(32'hbbb03df4),
	.w8(32'hbb0f1595),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050254),
	.w1(32'h3a7ce059),
	.w2(32'hb8fd7e15),
	.w3(32'hbb5501af),
	.w4(32'h3a2fcd34),
	.w5(32'hba0dfad0),
	.w6(32'h3a11bd75),
	.w7(32'hb96b5f63),
	.w8(32'h39a008e9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f53ff1),
	.w1(32'h3aa6fae4),
	.w2(32'hba5fe698),
	.w3(32'h3a40b09a),
	.w4(32'h3a8d28d1),
	.w5(32'hba8ef323),
	.w6(32'h3a8d23f2),
	.w7(32'hb9efbfac),
	.w8(32'hb9cb6054),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcf012),
	.w1(32'h3ae0368b),
	.w2(32'h3a8d35be),
	.w3(32'hba07d702),
	.w4(32'h3b7b2179),
	.w5(32'h3b4c6c61),
	.w6(32'hb9957a64),
	.w7(32'hb98b22e1),
	.w8(32'hba62bffe),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3846f8fb),
	.w1(32'h3a2c2862),
	.w2(32'hb9a61d52),
	.w3(32'h3abc9b37),
	.w4(32'h39e9d659),
	.w5(32'h397941f8),
	.w6(32'h396e882f),
	.w7(32'hba704901),
	.w8(32'hb86cb25a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d25c61),
	.w1(32'hba0f5534),
	.w2(32'hbafcf977),
	.w3(32'h39f9f1c1),
	.w4(32'hba555471),
	.w5(32'hbae3f8bc),
	.w6(32'hba6b01a2),
	.w7(32'hbae8a182),
	.w8(32'hbb16ca48),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053b7c),
	.w1(32'h3b7f6f7d),
	.w2(32'hbb454ed8),
	.w3(32'hbae1fe87),
	.w4(32'h3b9d6c13),
	.w5(32'hbb29400e),
	.w6(32'h3b89f10d),
	.w7(32'hbb72f463),
	.w8(32'h3a202a12),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904e0fe),
	.w1(32'h3b1cbadd),
	.w2(32'h3b509658),
	.w3(32'h38e8d648),
	.w4(32'h3b59ec78),
	.w5(32'h3b39e6ce),
	.w6(32'h3bb21f02),
	.w7(32'h3bfce2a0),
	.w8(32'h3bc2f4ff),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19bd03),
	.w1(32'hb937393c),
	.w2(32'hbaa02a0d),
	.w3(32'h3adaf2cf),
	.w4(32'hba102643),
	.w5(32'hbabdf963),
	.w6(32'h38ab3a15),
	.w7(32'hbaae6020),
	.w8(32'hb9a374d1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39838f73),
	.w1(32'hb99eac7b),
	.w2(32'hba366406),
	.w3(32'hb83c4fcd),
	.w4(32'hba69db14),
	.w5(32'hba8870b2),
	.w6(32'hba26e71f),
	.w7(32'hba8fab24),
	.w8(32'hb9f66fcf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db0ffc),
	.w1(32'h3a3bc473),
	.w2(32'hba3f7d12),
	.w3(32'hba45b5b6),
	.w4(32'hba5a3f62),
	.w5(32'hba2eb31c),
	.w6(32'h3a07dbf5),
	.w7(32'hbb09113a),
	.w8(32'hbaa25198),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7fe44),
	.w1(32'h3b240b4b),
	.w2(32'h3b1193eb),
	.w3(32'hba245150),
	.w4(32'h3ace3a74),
	.w5(32'h3b1ad516),
	.w6(32'h3ad06764),
	.w7(32'h3a871496),
	.w8(32'hbb13f98f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2251b4),
	.w1(32'hbaa5344d),
	.w2(32'hbab28a4f),
	.w3(32'hbac42e29),
	.w4(32'hbab97ff8),
	.w5(32'hba7fa50e),
	.w6(32'hba927981),
	.w7(32'hba62a680),
	.w8(32'hbad96cc7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1508d),
	.w1(32'hb9a0e8f3),
	.w2(32'hba7c2c89),
	.w3(32'hbad6503c),
	.w4(32'hba1d0d36),
	.w5(32'hbae3c086),
	.w6(32'hba0ba002),
	.w7(32'hbb0874d1),
	.w8(32'hba8355d4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987c7d6),
	.w1(32'hba3ec7d8),
	.w2(32'hbac13751),
	.w3(32'hba70aa01),
	.w4(32'hb9fd0b0b),
	.w5(32'hba5dc1fe),
	.w6(32'h39a87e1e),
	.w7(32'h392acd8e),
	.w8(32'h3a343032),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba441377),
	.w1(32'h3a921f18),
	.w2(32'h3a3179ed),
	.w3(32'hbaa05ffc),
	.w4(32'h3a29d3c0),
	.w5(32'h3a351449),
	.w6(32'h3a06deaa),
	.w7(32'h3a180d1c),
	.w8(32'h398295e0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e7cb0),
	.w1(32'h3a92bd3f),
	.w2(32'hb982a0f4),
	.w3(32'hb9c3ae4e),
	.w4(32'h3a60b1f5),
	.w5(32'hb9ae7731),
	.w6(32'h3a3c851c),
	.w7(32'hb9a79120),
	.w8(32'h39bc3b46),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ed638),
	.w1(32'hb99d5500),
	.w2(32'hb88c8209),
	.w3(32'h39e4ceb7),
	.w4(32'hb9934b33),
	.w5(32'h399b9fe9),
	.w6(32'h38d663ab),
	.w7(32'h3a2e3250),
	.w8(32'h3a44068b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97d2e7d),
	.w1(32'hba5433b8),
	.w2(32'h3b858ec3),
	.w3(32'hb9d66552),
	.w4(32'h3907c791),
	.w5(32'h3b17078a),
	.w6(32'h3b262ece),
	.w7(32'h3c04c29e),
	.w8(32'h3be4cd0d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb42ac0),
	.w1(32'hbae90f09),
	.w2(32'hba7fb676),
	.w3(32'h3b64e447),
	.w4(32'hbb125f31),
	.w5(32'hbab32994),
	.w6(32'hba54fd7a),
	.w7(32'hb91faeeb),
	.w8(32'hb8f57d54),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ee84),
	.w1(32'hba83b499),
	.w2(32'hbabfc54d),
	.w3(32'hbad72dc4),
	.w4(32'hba6cc4ce),
	.w5(32'hbab8d789),
	.w6(32'hbab42126),
	.w7(32'hbae73a44),
	.w8(32'hb9b91e9d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e240f),
	.w1(32'h3882ac8b),
	.w2(32'h39803bdf),
	.w3(32'hba34a5f6),
	.w4(32'h3862f404),
	.w5(32'h3a7e3061),
	.w6(32'hbaae4ff1),
	.w7(32'hba9eed4f),
	.w8(32'hbb5f3215),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb137afe),
	.w1(32'h39385d89),
	.w2(32'hb8fc71cc),
	.w3(32'hbaa1ab64),
	.w4(32'hb9a6fe5b),
	.w5(32'hb9885baa),
	.w6(32'hba530bcf),
	.w7(32'hba8843e4),
	.w8(32'hbae41960),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40dcd7),
	.w1(32'hba79b980),
	.w2(32'hba442805),
	.w3(32'hbb05d654),
	.w4(32'hba6c554e),
	.w5(32'hba26256c),
	.w6(32'hbaabd9c3),
	.w7(32'hbab3a663),
	.w8(32'hba95e0f0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe49a6),
	.w1(32'h3a241dc1),
	.w2(32'h3a3d6382),
	.w3(32'hbac54c17),
	.w4(32'h3aa6c202),
	.w5(32'h3ad19fa2),
	.w6(32'h39837aad),
	.w7(32'hba8e2f17),
	.w8(32'h3a27ab15),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af761c8),
	.w1(32'h3aa17441),
	.w2(32'hbb2c6d45),
	.w3(32'h39ba010d),
	.w4(32'h3b6d116d),
	.w5(32'hbac910c3),
	.w6(32'h3b5a1f26),
	.w7(32'hb9d0c183),
	.w8(32'h39f8a0a5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd4709),
	.w1(32'hb9feb94a),
	.w2(32'hba93b317),
	.w3(32'hb97a77ae),
	.w4(32'hba23ecf2),
	.w5(32'hba76d2a5),
	.w6(32'hba8835a7),
	.w7(32'hbae5e3fa),
	.w8(32'hba2fec44),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba411cc9),
	.w1(32'h3ac9f5b4),
	.w2(32'h39b40ca5),
	.w3(32'hb9eec8b5),
	.w4(32'h3a964f39),
	.w5(32'h3981e1a9),
	.w6(32'h3a6ac15e),
	.w7(32'h39737367),
	.w8(32'h3a322eef),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98b216),
	.w1(32'h3a854042),
	.w2(32'h3988ca04),
	.w3(32'h3a3e07ea),
	.w4(32'h3aba4070),
	.w5(32'h3a03b252),
	.w6(32'h3a0b5197),
	.w7(32'h3a05293d),
	.w8(32'hb942ea62),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c9479),
	.w1(32'h39d4d983),
	.w2(32'hba9fe94e),
	.w3(32'h3a248c40),
	.w4(32'h3ad5004e),
	.w5(32'hb997f419),
	.w6(32'hb9c5af33),
	.w7(32'h392d7765),
	.w8(32'hbae416f6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38b10b),
	.w1(32'h3aa55185),
	.w2(32'h3a204822),
	.w3(32'hbb63edf3),
	.w4(32'h3a039975),
	.w5(32'hb9e56bce),
	.w6(32'h3ad204ed),
	.w7(32'h39b5ed29),
	.w8(32'h3add8a05),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad504cd),
	.w1(32'h3a1c6657),
	.w2(32'h3a8fa80b),
	.w3(32'h3a6fe258),
	.w4(32'h3ad194b5),
	.w5(32'h3aa690e8),
	.w6(32'h3646afb4),
	.w7(32'hba2ea6bf),
	.w8(32'hb9dc3e9e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26ec4d),
	.w1(32'h3b5ff394),
	.w2(32'h3b442e23),
	.w3(32'hb9a9ed1f),
	.w4(32'h3b5d87f5),
	.w5(32'h3b4ba1c1),
	.w6(32'h3b9e8013),
	.w7(32'h3b5e198f),
	.w8(32'h3a5433db),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386847c7),
	.w1(32'h3b53b179),
	.w2(32'h3b8e6355),
	.w3(32'h3a918cac),
	.w4(32'h3b3c34bd),
	.w5(32'h3a7e4bbe),
	.w6(32'h3b19e238),
	.w7(32'h3bc80209),
	.w8(32'h3c56e96c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c510c75),
	.w1(32'h3af9cf83),
	.w2(32'h3b5df8e3),
	.w3(32'h3beccca1),
	.w4(32'h3ae5c416),
	.w5(32'h3b2d60d3),
	.w6(32'h3b075234),
	.w7(32'h3b861ae8),
	.w8(32'h3b1f368c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982c63),
	.w1(32'h3a503142),
	.w2(32'h3acbc2a1),
	.w3(32'h3ac7cfd5),
	.w4(32'h3a832052),
	.w5(32'h3a16e4a0),
	.w6(32'h39169bca),
	.w7(32'h3a58a3e3),
	.w8(32'h3ad46b75),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b4562),
	.w1(32'h39b38220),
	.w2(32'hba138f9f),
	.w3(32'h3a2042e0),
	.w4(32'h38fe1fd3),
	.w5(32'hb8ec7a6d),
	.w6(32'h3981dd6c),
	.w7(32'h388e863f),
	.w8(32'hb96f372f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bf02),
	.w1(32'h388f88de),
	.w2(32'hbab1ed99),
	.w3(32'hbb001751),
	.w4(32'hb912106e),
	.w5(32'hbaa61d6b),
	.w6(32'h39af42b8),
	.w7(32'hb9fcbed2),
	.w8(32'hb9004282),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ded897),
	.w1(32'hba01e471),
	.w2(32'h3a22c9c7),
	.w3(32'h39229598),
	.w4(32'hba77d10a),
	.w5(32'hb951205d),
	.w6(32'hb99b7724),
	.w7(32'h3a6ef275),
	.w8(32'h3a304b69),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b6b32f),
	.w1(32'h39f52109),
	.w2(32'hba30c2e2),
	.w3(32'hb9f26319),
	.w4(32'h39c65d11),
	.w5(32'hb98d5489),
	.w6(32'hb9cd6fa0),
	.w7(32'hba32a555),
	.w8(32'hb956506d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9190a78),
	.w1(32'h3b2f1887),
	.w2(32'h3b26afdc),
	.w3(32'hb907dfa8),
	.w4(32'h3ab7d3d0),
	.w5(32'h3b477a16),
	.w6(32'h38e4df6e),
	.w7(32'h3a316e04),
	.w8(32'h3ac7bfce),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c31d4e),
	.w1(32'hb9e57d6d),
	.w2(32'hb8e10832),
	.w3(32'h3a7a6c12),
	.w4(32'hb9a26b8b),
	.w5(32'h39db6aa5),
	.w6(32'hba8c1507),
	.w7(32'hba7e80a5),
	.w8(32'hbb10fdeb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac926b0),
	.w1(32'h3a593771),
	.w2(32'hb9e0695b),
	.w3(32'hba61473b),
	.w4(32'h3929d926),
	.w5(32'hba17ee98),
	.w6(32'h38ab478d),
	.w7(32'hbaa5c756),
	.w8(32'h384cb505),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9824e6b),
	.w1(32'h37b00661),
	.w2(32'hba9c39dd),
	.w3(32'hb920e6f3),
	.w4(32'h39ab296a),
	.w5(32'hb99752cf),
	.w6(32'h3a7b0b24),
	.w7(32'h397ae2a3),
	.w8(32'h398b7cea),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1449a),
	.w1(32'hba2907d3),
	.w2(32'h3b5b3fbd),
	.w3(32'hb8151f57),
	.w4(32'hba312906),
	.w5(32'h3b396c61),
	.w6(32'h3b0fcde8),
	.w7(32'h3c0f4586),
	.w8(32'h3c0febe5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9bd8b),
	.w1(32'hbaeb4b6c),
	.w2(32'hbaee77f1),
	.w3(32'h3b6f9728),
	.w4(32'hbaa942aa),
	.w5(32'hbb2cb0eb),
	.w6(32'hbadc924a),
	.w7(32'hbabef747),
	.w8(32'hbac305ec),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d8265),
	.w1(32'h38c2ab27),
	.w2(32'hb8604c74),
	.w3(32'hba8f9365),
	.w4(32'hb979671b),
	.w5(32'hb98fdff1),
	.w6(32'hb88e915d),
	.w7(32'hba179eaf),
	.w8(32'h39842d1a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a070030),
	.w1(32'hba6fc777),
	.w2(32'hbb0707ae),
	.w3(32'hb9168524),
	.w4(32'hbaac6f3b),
	.w5(32'hbb14b905),
	.w6(32'hbac672f6),
	.w7(32'hbb14dac9),
	.w8(32'hbb4349eb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb137e96),
	.w1(32'hb937e3e0),
	.w2(32'hb9bca75e),
	.w3(32'hbb17f2e0),
	.w4(32'hb9cbb7e8),
	.w5(32'h394c60bc),
	.w6(32'hb9f56dcc),
	.w7(32'h399d366d),
	.w8(32'hb957a7fb),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7530d6),
	.w1(32'h3903047b),
	.w2(32'hb9134d3f),
	.w3(32'hba973668),
	.w4(32'h38ad3683),
	.w5(32'hb770be29),
	.w6(32'h3904f3e7),
	.w7(32'hba1370ad),
	.w8(32'hb8bcaf39),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a66b48),
	.w1(32'h3a7b0968),
	.w2(32'hb9f650a9),
	.w3(32'h39be510d),
	.w4(32'h3a2398ee),
	.w5(32'hba262a99),
	.w6(32'h39b900a2),
	.w7(32'hb9d1eee5),
	.w8(32'h39a0102c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35035f),
	.w1(32'hb9cd16a2),
	.w2(32'hba585f70),
	.w3(32'h39871660),
	.w4(32'hba49aa13),
	.w5(32'hbab83af2),
	.w6(32'hba052c88),
	.w7(32'hbae1dcb9),
	.w8(32'hba125d58),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392462fe),
	.w1(32'hb7c6ea5d),
	.w2(32'hba847927),
	.w3(32'hba109694),
	.w4(32'hb9acdc3b),
	.w5(32'hba46cf72),
	.w6(32'h38006f8c),
	.w7(32'hb99276de),
	.w8(32'h38539f87),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00308b),
	.w1(32'h3a56b915),
	.w2(32'h3b3d7869),
	.w3(32'hba1fe10b),
	.w4(32'h3a2fe5c7),
	.w5(32'h3b13d933),
	.w6(32'h3a8457ea),
	.w7(32'h3af3731f),
	.w8(32'h39d95430),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0eb5d),
	.w1(32'h3b276144),
	.w2(32'hb8e7bfa5),
	.w3(32'hb99c9916),
	.w4(32'h3b0004d7),
	.w5(32'hb9b3c113),
	.w6(32'h3a6bdc03),
	.w7(32'hbac23245),
	.w8(32'hb9962771),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5642b),
	.w1(32'h3a54d1ea),
	.w2(32'h3ad1c847),
	.w3(32'h3a96c4b2),
	.w4(32'h37b9dc9d),
	.w5(32'h3a8aaa2a),
	.w6(32'h3ab7b197),
	.w7(32'h3b133d9e),
	.w8(32'h3ad8b1d3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f8a8d7),
	.w1(32'h3b7cfab7),
	.w2(32'h3aa223c5),
	.w3(32'h392cb78c),
	.w4(32'h3ba7d9b0),
	.w5(32'h3aede269),
	.w6(32'h3b995bc2),
	.w7(32'h3a799615),
	.w8(32'hbb041dca),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad793),
	.w1(32'h3a505e3d),
	.w2(32'hbacabb56),
	.w3(32'hba2d573d),
	.w4(32'h3872ebb5),
	.w5(32'hbafd96cc),
	.w6(32'h3a976cc4),
	.w7(32'hbae09d32),
	.w8(32'hb94aa900),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a054b4b),
	.w1(32'hbab21302),
	.w2(32'h39aa23ce),
	.w3(32'h38949d9b),
	.w4(32'hbadc8052),
	.w5(32'hbaecede9),
	.w6(32'h3ab39504),
	.w7(32'h3b346472),
	.w8(32'h3b93f65f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8e7e),
	.w1(32'h3a2b8c5a),
	.w2(32'h395b7f8d),
	.w3(32'h3aba048e),
	.w4(32'hba15f908),
	.w5(32'h390f8993),
	.w6(32'h3a5c1b47),
	.w7(32'h3a07a543),
	.w8(32'h39ffe158),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d33492),
	.w1(32'h3a75faa9),
	.w2(32'h3a41fcb0),
	.w3(32'hba4aea29),
	.w4(32'h3aa87d6d),
	.w5(32'h398c680b),
	.w6(32'h3b0c5880),
	.w7(32'h3af6d6f6),
	.w8(32'h3b333a61),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa96e2),
	.w1(32'h396c26cc),
	.w2(32'h39ae6b5d),
	.w3(32'h3a5a384b),
	.w4(32'hb920ddf2),
	.w5(32'h397daf47),
	.w6(32'h398a1072),
	.w7(32'h3960aa42),
	.w8(32'hb88ee1bc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c74213),
	.w1(32'hbbbadd04),
	.w2(32'hbb8641ac),
	.w3(32'hba3702d1),
	.w4(32'hba1ba9f6),
	.w5(32'hb9e987bf),
	.w6(32'hb9aa491e),
	.w7(32'hb9c4a6ef),
	.w8(32'hbac7ed31),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9faa),
	.w1(32'h3ac68bf7),
	.w2(32'h3b216478),
	.w3(32'hbad6d963),
	.w4(32'hb9b78110),
	.w5(32'h3aa9b28f),
	.w6(32'h3b11a54f),
	.w7(32'h3b86f88b),
	.w8(32'h3b6bcc47),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2dcd3),
	.w1(32'hb86c869a),
	.w2(32'h3a2e82b4),
	.w3(32'h369b4a76),
	.w4(32'hba9587fe),
	.w5(32'hb93b0e3e),
	.w6(32'hba8c9c1c),
	.w7(32'h3a77192f),
	.w8(32'h3823602d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391efe98),
	.w1(32'h38e6d70c),
	.w2(32'hba38b4b4),
	.w3(32'hba98251d),
	.w4(32'hb9f4c025),
	.w5(32'hba97f4a2),
	.w6(32'h39da1a06),
	.w7(32'hba8164f1),
	.w8(32'hb97ea4da),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09d5b7),
	.w1(32'h3b2551fe),
	.w2(32'h3b2312dd),
	.w3(32'h38b1feb2),
	.w4(32'h3b262fa2),
	.w5(32'h3b416045),
	.w6(32'h3b67e63a),
	.w7(32'h3b3fbc58),
	.w8(32'h3a80eb23),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385fa8e3),
	.w1(32'hb8968978),
	.w2(32'hbae096dc),
	.w3(32'h3aaa0943),
	.w4(32'hba87cd8b),
	.w5(32'hbaec5d64),
	.w6(32'hb9b9dff7),
	.w7(32'hbae37656),
	.w8(32'hba032818),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b67ef),
	.w1(32'hbaa25463),
	.w2(32'hbaf87276),
	.w3(32'hb9ad5b92),
	.w4(32'hbaf33a66),
	.w5(32'hbb0e5788),
	.w6(32'hba087364),
	.w7(32'hba7dc119),
	.w8(32'hb7f99da1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb34cd),
	.w1(32'hba18042b),
	.w2(32'hb8ba7081),
	.w3(32'hba8798f1),
	.w4(32'hba6cf02b),
	.w5(32'h395b2525),
	.w6(32'hba5711b0),
	.w7(32'hb99592ee),
	.w8(32'hb992244a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba257b36),
	.w1(32'h3a85f780),
	.w2(32'h3a92b43f),
	.w3(32'h398c7633),
	.w4(32'h380707e0),
	.w5(32'h3998b481),
	.w6(32'h3b009e01),
	.w7(32'h3adec637),
	.w8(32'h3aace12d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8571d),
	.w1(32'h3b5cb1a6),
	.w2(32'h39fd45d1),
	.w3(32'h39ef3979),
	.w4(32'h3b06f97c),
	.w5(32'hbb46d7d9),
	.w6(32'h3b669db6),
	.w7(32'hb9468271),
	.w8(32'h3b392f82),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c5c38),
	.w1(32'hba542bdd),
	.w2(32'hb93d6a2a),
	.w3(32'h393fcb47),
	.w4(32'hba8071c7),
	.w5(32'hba1967c6),
	.w6(32'hb970e76f),
	.w7(32'h3994176b),
	.w8(32'h3a03b7c9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899c61b),
	.w1(32'hbae83469),
	.w2(32'hbaf62118),
	.w3(32'hb9cf7493),
	.w4(32'hbac84a6a),
	.w5(32'hbafcf190),
	.w6(32'hbb0fb028),
	.w7(32'hbb4f3d43),
	.w8(32'hbadbf671),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafc55d),
	.w1(32'h3a92ec4e),
	.w2(32'hb8858a39),
	.w3(32'hbb0c73d4),
	.w4(32'hb8bb4fce),
	.w5(32'hbaa7496f),
	.w6(32'h3943f502),
	.w7(32'hbaf4f698),
	.w8(32'hbb253f86),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9efc71),
	.w1(32'h39aa85fb),
	.w2(32'h39617e5d),
	.w3(32'hbaf7c02b),
	.w4(32'hb974af42),
	.w5(32'h39c1ada0),
	.w6(32'hb9aca445),
	.w7(32'hb8fad8b6),
	.w8(32'hbad00b62),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddad33),
	.w1(32'h396044c5),
	.w2(32'h39f7cb15),
	.w3(32'hba50f5ea),
	.w4(32'hba57d7cf),
	.w5(32'h3a036f39),
	.w6(32'h3a9e6b66),
	.w7(32'h3ae041e2),
	.w8(32'h3ad8eec1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de216c),
	.w1(32'h3a82153a),
	.w2(32'hbad00712),
	.w3(32'hb9e78e16),
	.w4(32'hb899ba66),
	.w5(32'hbaf1e84c),
	.w6(32'h3ad87d84),
	.w7(32'hb922d0dd),
	.w8(32'h3a7af4ec),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219fc4),
	.w1(32'h3b2f31fa),
	.w2(32'h3b493632),
	.w3(32'hba0074e2),
	.w4(32'h3b2d921f),
	.w5(32'h3ae70973),
	.w6(32'h3a665145),
	.w7(32'h3ac2bac1),
	.w8(32'h3aec62f4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7cfa3),
	.w1(32'hb9ef5e54),
	.w2(32'h3ad0d602),
	.w3(32'h399759f2),
	.w4(32'hba8df0c6),
	.w5(32'h3a8882c8),
	.w6(32'h37e74db9),
	.w7(32'h3a7903da),
	.w8(32'h39c3d502),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab58f0f),
	.w1(32'h3b4856ad),
	.w2(32'hba69a8a6),
	.w3(32'h3ade537b),
	.w4(32'h3b1f34ac),
	.w5(32'hba920fc1),
	.w6(32'h3a692d5d),
	.w7(32'hbb190f7b),
	.w8(32'hba431d38),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5024c),
	.w1(32'h3a535866),
	.w2(32'h36e0c424),
	.w3(32'h3ad19696),
	.w4(32'h39dc6bf3),
	.w5(32'hb8be853b),
	.w6(32'h3a2d06d9),
	.w7(32'hb9fc4df5),
	.w8(32'h39bd512c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cf7ad),
	.w1(32'h3aeb147b),
	.w2(32'hb93b15a8),
	.w3(32'h3a8d0cb5),
	.w4(32'h3ab06f3e),
	.w5(32'hb9daf760),
	.w6(32'h3a34c04d),
	.w7(32'hba9fbffd),
	.w8(32'hb99f4a3c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f23e9),
	.w1(32'h35bcb6e5),
	.w2(32'hba872d2a),
	.w3(32'h3a06faa2),
	.w4(32'hb8f64869),
	.w5(32'hba7ae4f9),
	.w6(32'hb9c4c127),
	.w7(32'hbad40b42),
	.w8(32'hb9dabf50),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e13db0),
	.w1(32'hb9457360),
	.w2(32'hb9685148),
	.w3(32'h38a47c09),
	.w4(32'hba523423),
	.w5(32'hb946b25b),
	.w6(32'h39d1e5d7),
	.w7(32'h3a0e663c),
	.w8(32'h3a39c123),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03df82),
	.w1(32'h39b63164),
	.w2(32'hba8cd416),
	.w3(32'hba5513a1),
	.w4(32'hba9512ed),
	.w5(32'hbb06ac80),
	.w6(32'h39cf36ca),
	.w7(32'hbaae43b1),
	.w8(32'hb8be2d83),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09faca),
	.w1(32'h3af757ab),
	.w2(32'hb91d11d6),
	.w3(32'hba4e7ec0),
	.w4(32'h3ab28849),
	.w5(32'hb9b2f5da),
	.w6(32'h3a2d9b1a),
	.w7(32'hbaa2488a),
	.w8(32'hb9945b55),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84b331),
	.w1(32'h3aa2a2f1),
	.w2(32'h3a6e685d),
	.w3(32'h3a79c0e9),
	.w4(32'h38ccc189),
	.w5(32'h39c8f7cf),
	.w6(32'h3a380361),
	.w7(32'h38abe040),
	.w8(32'hb98050a8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e18f3c),
	.w1(32'h3a852e11),
	.w2(32'hba17e8df),
	.w3(32'hba325d1c),
	.w4(32'h3a0077cc),
	.w5(32'hba9ad93a),
	.w6(32'hb9471c27),
	.w7(32'hba7ac418),
	.w8(32'h388803f7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945682),
	.w1(32'h3b1cac75),
	.w2(32'h3aea865a),
	.w3(32'hba694e73),
	.w4(32'h3b0d6431),
	.w5(32'h3a3165e3),
	.w6(32'hba3a82f1),
	.w7(32'h3ab55db9),
	.w8(32'hba2903ce),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48928d),
	.w1(32'h396811d5),
	.w2(32'hba78503d),
	.w3(32'hbb30ccbe),
	.w4(32'h3985285c),
	.w5(32'hba9bcee5),
	.w6(32'h39297804),
	.w7(32'hba50ae89),
	.w8(32'h38d6fd4d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37315d2c),
	.w1(32'hbae405c2),
	.w2(32'hbac83091),
	.w3(32'hba46e099),
	.w4(32'hbabc2c62),
	.w5(32'hba9b9e32),
	.w6(32'hba1defcf),
	.w7(32'hb8a6a3d9),
	.w8(32'hb9426086),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f184c),
	.w1(32'h3a5ca9ca),
	.w2(32'h3a29acfc),
	.w3(32'hba7fc612),
	.w4(32'h3a5ca853),
	.w5(32'h39addda1),
	.w6(32'h393176b8),
	.w7(32'h38bf0fcf),
	.w8(32'h3a9117a8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcdee7),
	.w1(32'h3b38a724),
	.w2(32'hb92287a9),
	.w3(32'hb80d55f9),
	.w4(32'h3b069d42),
	.w5(32'hba0c987f),
	.w6(32'h3a85bcd1),
	.w7(32'hbaea3ab3),
	.w8(32'hba018fe3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4d592),
	.w1(32'h3a146c7c),
	.w2(32'hb9d65fba),
	.w3(32'h3aaa83ce),
	.w4(32'h39f58d9f),
	.w5(32'hb9f2f2c8),
	.w6(32'h39d948ed),
	.w7(32'hb9c28d23),
	.w8(32'h3a4bfd49),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a456957),
	.w1(32'h3a7b643b),
	.w2(32'hb9af8d2e),
	.w3(32'h3a20fc29),
	.w4(32'h3a1ccbe0),
	.w5(32'hba0a3f76),
	.w6(32'h3a1372a9),
	.w7(32'hba2f4a77),
	.w8(32'h3a3f9bf9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30fa20),
	.w1(32'hbacc1b7e),
	.w2(32'hbafe7733),
	.w3(32'h399dfcdd),
	.w4(32'hba8a2de6),
	.w5(32'hbae3bbe0),
	.w6(32'hbb260721),
	.w7(32'hbb2b592a),
	.w8(32'hbac77c8b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb178b26),
	.w1(32'h39b0481d),
	.w2(32'hb89495d8),
	.w3(32'hbadc5ac5),
	.w4(32'h3a267092),
	.w5(32'hb9239042),
	.w6(32'h3a132e83),
	.w7(32'h3993b16d),
	.w8(32'h3a85ccaf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32ec52),
	.w1(32'hb8964347),
	.w2(32'hbaaef9c1),
	.w3(32'hb580ba7e),
	.w4(32'hba7924d9),
	.w5(32'hbb26e659),
	.w6(32'hba1554c5),
	.w7(32'hbb18fa0a),
	.w8(32'hba01bcbd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079165),
	.w1(32'hba4711b8),
	.w2(32'hbaa96023),
	.w3(32'hba92408c),
	.w4(32'hbaa89230),
	.w5(32'hbac5283d),
	.w6(32'hba038b8f),
	.w7(32'hba280fd0),
	.w8(32'hb970cf0b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2360f9),
	.w1(32'h3a9d7534),
	.w2(32'h361dde78),
	.w3(32'hba68b96d),
	.w4(32'h3a6c9bf1),
	.w5(32'hb96405ed),
	.w6(32'h3a373d83),
	.w7(32'hb9399591),
	.w8(32'h39cc3775),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a733117),
	.w1(32'hb91e49e1),
	.w2(32'hb99a4ad8),
	.w3(32'h39d5091e),
	.w4(32'hba814954),
	.w5(32'hba58c58c),
	.w6(32'hbb131022),
	.w7(32'hbb0113ea),
	.w8(32'hbad8ca3c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba720607),
	.w1(32'h3a4737ae),
	.w2(32'hba67b514),
	.w3(32'hbac06184),
	.w4(32'h3957dd5c),
	.w5(32'hba989ae5),
	.w6(32'h3ae34d43),
	.w7(32'hb9699b70),
	.w8(32'h3add6e86),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84c86f7),
	.w1(32'hb9b5b629),
	.w2(32'hbaa91984),
	.w3(32'hb9bb300d),
	.w4(32'hba5cb5aa),
	.w5(32'hbb1afaac),
	.w6(32'h394c15ec),
	.w7(32'hbad695dc),
	.w8(32'hb9799048),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8c3eb),
	.w1(32'h3a2fcda1),
	.w2(32'hbb30c552),
	.w3(32'hb8130ded),
	.w4(32'h3a6e517e),
	.w5(32'hbae63cf2),
	.w6(32'h3ae658a4),
	.w7(32'hb9e5566b),
	.w8(32'hba282602),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b8612),
	.w1(32'hb94bded7),
	.w2(32'h39ba2f94),
	.w3(32'hbada804d),
	.w4(32'hbb01dd20),
	.w5(32'hba3a3b1c),
	.w6(32'h3a4e460c),
	.w7(32'h3a8c5cbc),
	.w8(32'h3b24d880),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule