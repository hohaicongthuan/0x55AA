module layer_10_featuremap_441(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989eb53),
	.w1(32'h3a520f4f),
	.w2(32'h3aa87280),
	.w3(32'h3c043326),
	.w4(32'hbb217a23),
	.w5(32'hbba7a51f),
	.w6(32'hbb50742c),
	.w7(32'hbb2929e8),
	.w8(32'h3b65915d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0321c3),
	.w1(32'h3c1ff276),
	.w2(32'h3c29f313),
	.w3(32'h3b0fd45a),
	.w4(32'h3ab21904),
	.w5(32'h3bf02aac),
	.w6(32'h3ac89341),
	.w7(32'h3b80cb65),
	.w8(32'h3acf8956),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb504f),
	.w1(32'hbb823da5),
	.w2(32'h3ac5b9f9),
	.w3(32'hba74a43d),
	.w4(32'hba9f9b6e),
	.w5(32'hba9838cd),
	.w6(32'h3b33c0ac),
	.w7(32'hbb5c0f76),
	.w8(32'h3b048cef),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf52a0),
	.w1(32'hbc061864),
	.w2(32'h3a1f42a5),
	.w3(32'hbb0a8f3b),
	.w4(32'hbb9b0a78),
	.w5(32'h3bc0bbaa),
	.w6(32'h3b7075fb),
	.w7(32'hbaf217f4),
	.w8(32'h3b2a7286),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c2d0),
	.w1(32'h3bc03c86),
	.w2(32'hbaf3a2a0),
	.w3(32'h3a538d5c),
	.w4(32'h3bab0ad4),
	.w5(32'hbb184c39),
	.w6(32'h3b27acc6),
	.w7(32'h3a8fe85a),
	.w8(32'hbbaa4b43),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0762f4),
	.w1(32'h3c0ca03d),
	.w2(32'hbc1e4f8f),
	.w3(32'hbaef8eb9),
	.w4(32'hbbbbc9be),
	.w5(32'hb839b952),
	.w6(32'hbbb0eeb6),
	.w7(32'h3b04ecf7),
	.w8(32'hbb1e151d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd67164),
	.w1(32'hbb2dc38a),
	.w2(32'h39c0f9e6),
	.w3(32'hbbe110a4),
	.w4(32'h3b214170),
	.w5(32'h3c18e5e2),
	.w6(32'hba8af51c),
	.w7(32'h3b877f98),
	.w8(32'hba001e76),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde87b0),
	.w1(32'h3c36c8e2),
	.w2(32'h3bc21883),
	.w3(32'h3c1fe323),
	.w4(32'h3c465df3),
	.w5(32'hbc1a7bb5),
	.w6(32'hbb6a02eb),
	.w7(32'h39b65971),
	.w8(32'hbbfe2585),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db2f3),
	.w1(32'hbafe181e),
	.w2(32'h3b5ac382),
	.w3(32'hbb89e549),
	.w4(32'h3b31dc9f),
	.w5(32'h3adbd1f3),
	.w6(32'h3a4c269e),
	.w7(32'h3b552440),
	.w8(32'hb9d4d4ad),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0192e),
	.w1(32'hbbaf27dd),
	.w2(32'h3bb40f47),
	.w3(32'h3ac34cb3),
	.w4(32'h3ac8e763),
	.w5(32'h3b3ba7c2),
	.w6(32'hba628ed0),
	.w7(32'hbbc37a18),
	.w8(32'hbc19cc9e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84e9f4),
	.w1(32'h39482436),
	.w2(32'hb9c591f3),
	.w3(32'hbb83a81c),
	.w4(32'hbb7e1e0f),
	.w5(32'hba658ca7),
	.w6(32'hbbedb2d9),
	.w7(32'hbae05c4b),
	.w8(32'h3b62c36d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50ac18),
	.w1(32'h3c42d475),
	.w2(32'h3ae411e5),
	.w3(32'h3baad5e0),
	.w4(32'h3c38db22),
	.w5(32'hbc057a55),
	.w6(32'h3bb827e1),
	.w7(32'h3b842479),
	.w8(32'hbc1ee4f0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6997),
	.w1(32'hbc08b53b),
	.w2(32'hbb5763ad),
	.w3(32'h397e2904),
	.w4(32'hbb91705d),
	.w5(32'h3c183f9a),
	.w6(32'hbb008a7a),
	.w7(32'hbb594f1a),
	.w8(32'hbb57dd82),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaceb1b),
	.w1(32'h3a1c8c6f),
	.w2(32'hbb366e48),
	.w3(32'h3ae75de0),
	.w4(32'hba01b8e1),
	.w5(32'hbb86a61d),
	.w6(32'h38c73d24),
	.w7(32'hbb7d5486),
	.w8(32'hbb9b06c0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9747633),
	.w1(32'hbb8044ac),
	.w2(32'h3a99fa62),
	.w3(32'hba747cd3),
	.w4(32'hbc0989a6),
	.w5(32'hbab90ab6),
	.w6(32'hbbe415ec),
	.w7(32'hbb57edb1),
	.w8(32'hbb9c8a00),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73cd07),
	.w1(32'hbc3c53e8),
	.w2(32'hbc0e7db3),
	.w3(32'h3912934c),
	.w4(32'hbc440a58),
	.w5(32'hbc12e388),
	.w6(32'hbaf9f7de),
	.w7(32'hbc34a768),
	.w8(32'hbc37d64c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac2c5),
	.w1(32'h38c9cea5),
	.w2(32'h3b56eeb2),
	.w3(32'h3a8193b8),
	.w4(32'h3b8a84da),
	.w5(32'h3c0061ec),
	.w6(32'h3ba612fa),
	.w7(32'hbbdf969f),
	.w8(32'hbbaf951c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294de6),
	.w1(32'hbb82115f),
	.w2(32'h3b888589),
	.w3(32'h398496d6),
	.w4(32'h3bab6395),
	.w5(32'h3aadacf7),
	.w6(32'hbba81dee),
	.w7(32'h3b3b7229),
	.w8(32'hbba1c0ce),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb9785),
	.w1(32'hbb45b4f3),
	.w2(32'hbbb0d4e1),
	.w3(32'h3aec5bed),
	.w4(32'hba5e2347),
	.w5(32'hba8f58d0),
	.w6(32'hbb813edb),
	.w7(32'hbb985515),
	.w8(32'hbbaabaa0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975808),
	.w1(32'hba97372f),
	.w2(32'h3b89ca68),
	.w3(32'h392f1a6a),
	.w4(32'hbbb9adbe),
	.w5(32'hbc165d0e),
	.w6(32'h3a31c6e1),
	.w7(32'hbc2c5eaa),
	.w8(32'hbc139757),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99743df),
	.w1(32'h3b013bb1),
	.w2(32'hbbcf4984),
	.w3(32'h3a9f68e1),
	.w4(32'h3a1ce89a),
	.w5(32'h3aa2ba19),
	.w6(32'hbb80c084),
	.w7(32'h3b975c76),
	.w8(32'h39b70054),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7274),
	.w1(32'h3a807942),
	.w2(32'h3a5ec0c3),
	.w3(32'h3af4dc37),
	.w4(32'hbb8cce44),
	.w5(32'h3b0d7c74),
	.w6(32'h3a206550),
	.w7(32'hbad4f82c),
	.w8(32'h398400a9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392debf0),
	.w1(32'h3bb51efc),
	.w2(32'hbc267aba),
	.w3(32'h3bd822c4),
	.w4(32'hbc49be0a),
	.w5(32'hbc2d7f07),
	.w6(32'hb937086c),
	.w7(32'hbc20d05e),
	.w8(32'hbc85961d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170f07),
	.w1(32'hbb02c5d0),
	.w2(32'h3b4aa1a9),
	.w3(32'hbbdf595b),
	.w4(32'hba967109),
	.w5(32'h3b567278),
	.w6(32'hbb213e5c),
	.w7(32'hbc1a72db),
	.w8(32'hbb635c43),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992d0da),
	.w1(32'hbba4eafe),
	.w2(32'hbc19b42d),
	.w3(32'hb97d59a5),
	.w4(32'hbc33aff7),
	.w5(32'hbb2ee758),
	.w6(32'hbaf68bd7),
	.w7(32'hbb8f3092),
	.w8(32'hbb43df7b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a777be),
	.w1(32'h3c135811),
	.w2(32'h3bc47d16),
	.w3(32'hbbde9161),
	.w4(32'h3c08c918),
	.w5(32'hbc0ffbe4),
	.w6(32'h3b81d732),
	.w7(32'h3bf34f4f),
	.w8(32'h3b962912),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c5396),
	.w1(32'h3bf81e59),
	.w2(32'h3ccc1a2a),
	.w3(32'h3962f784),
	.w4(32'h3cabc92c),
	.w5(32'h3cd7799d),
	.w6(32'h3bc259b0),
	.w7(32'h3c9c6895),
	.w8(32'h3c35d91b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c467fae),
	.w1(32'hb98e721e),
	.w2(32'h3a146930),
	.w3(32'h3c97d0f6),
	.w4(32'h3bfc22e4),
	.w5(32'hbb2af044),
	.w6(32'h3c2cd12e),
	.w7(32'h3ae1aeec),
	.w8(32'hbbae13f7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80dce9),
	.w1(32'h3acaefdc),
	.w2(32'h3c3464d9),
	.w3(32'hbb85b3c5),
	.w4(32'h3cb70e75),
	.w5(32'h3cc7c77e),
	.w6(32'hbc551b6c),
	.w7(32'h3bf289a6),
	.w8(32'h3b78da09),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51ca38),
	.w1(32'hb92141ba),
	.w2(32'h3873fceb),
	.w3(32'h3bb88119),
	.w4(32'h3a365ce8),
	.w5(32'hbb5e5c97),
	.w6(32'hba8b598b),
	.w7(32'hb85c372f),
	.w8(32'hbb863e2a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa76ef0),
	.w1(32'hbbee4150),
	.w2(32'h3a826f04),
	.w3(32'hbba8435b),
	.w4(32'h39067109),
	.w5(32'h3b1bb17e),
	.w6(32'hbbf2b044),
	.w7(32'hbc3ab375),
	.w8(32'hbc18753f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd51caa),
	.w1(32'h3b734efe),
	.w2(32'h3beda58d),
	.w3(32'h3bc6714a),
	.w4(32'h3b5ddc7a),
	.w5(32'h3b83125c),
	.w6(32'h3b3d9b58),
	.w7(32'hba6d6371),
	.w8(32'hbb242cd1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1f7c7),
	.w1(32'hbb887d2d),
	.w2(32'hba115216),
	.w3(32'h39b0dea4),
	.w4(32'h396f42c5),
	.w5(32'h3c00b816),
	.w6(32'h3acab1c1),
	.w7(32'hbbbbaf1b),
	.w8(32'h39f91182),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5257fd),
	.w1(32'h3c1d8cf3),
	.w2(32'h3c788a11),
	.w3(32'hbb9c8a06),
	.w4(32'h3b913aba),
	.w5(32'hbb5eb8f4),
	.w6(32'hbb3896a4),
	.w7(32'h3abee15d),
	.w8(32'hbb2c52f3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b281b26),
	.w1(32'h3c3ce65c),
	.w2(32'h3b20bf8d),
	.w3(32'hbb802380),
	.w4(32'h3c173f52),
	.w5(32'hbc0ac90a),
	.w6(32'hbbf1a24d),
	.w7(32'h3c055413),
	.w8(32'hb83495b5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad362f0),
	.w1(32'hbb45c6a0),
	.w2(32'hbb2ff390),
	.w3(32'hbba1c786),
	.w4(32'hbbbfac4c),
	.w5(32'hbb3e0e7a),
	.w6(32'h3b36e8fc),
	.w7(32'hba8e7718),
	.w8(32'h3a9fc85a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f7ec),
	.w1(32'hbbd2d850),
	.w2(32'h3a0f3ec0),
	.w3(32'h3ba4bd06),
	.w4(32'hbb66f623),
	.w5(32'h3c52de60),
	.w6(32'h3ab57e2c),
	.w7(32'h3b68eb41),
	.w8(32'hbb2c0a3f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c932055),
	.w1(32'h3bbc0e4f),
	.w2(32'hbb86c07d),
	.w3(32'h3bbb4c6a),
	.w4(32'h3beeb47a),
	.w5(32'h39826f9a),
	.w6(32'hbb406a54),
	.w7(32'h3b027994),
	.w8(32'hbbbe7b6f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04a53f),
	.w1(32'h3b988f43),
	.w2(32'hbb5476d3),
	.w3(32'h3b08bedd),
	.w4(32'h3ad2e39c),
	.w5(32'hbb05fbcf),
	.w6(32'hbba0fdcf),
	.w7(32'h39855a99),
	.w8(32'h3a0d44b5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb959564),
	.w1(32'hbbcfcdab),
	.w2(32'hbb6aa396),
	.w3(32'h3b001461),
	.w4(32'hbb8b7807),
	.w5(32'hbb3bef0e),
	.w6(32'hba7f2f07),
	.w7(32'hbbf85204),
	.w8(32'hbaaabf53),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8614),
	.w1(32'h3ba7aa1b),
	.w2(32'hbc194737),
	.w3(32'hbac22486),
	.w4(32'hbbc320b4),
	.w5(32'h3b9ce3fb),
	.w6(32'h397a0f06),
	.w7(32'h3b02650f),
	.w8(32'h3b24d0c9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96440b),
	.w1(32'hb9634594),
	.w2(32'h3b60a1b6),
	.w3(32'h3be35e90),
	.w4(32'hbafe3d0e),
	.w5(32'h3c6018e3),
	.w6(32'hbac38edd),
	.w7(32'h3b279972),
	.w8(32'hbacba9f0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac810ac),
	.w1(32'h3b254417),
	.w2(32'h3a6cd80a),
	.w3(32'h3ad2fc2d),
	.w4(32'h3beaf81f),
	.w5(32'h3bb31779),
	.w6(32'h3b0b6b8e),
	.w7(32'hbb4e811a),
	.w8(32'hbb8aaa99),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ccab),
	.w1(32'hbc1bb55b),
	.w2(32'hbb39a8b5),
	.w3(32'hbb104efe),
	.w4(32'hbc4a8355),
	.w5(32'hbae348f0),
	.w6(32'h3aa91613),
	.w7(32'hbbeef902),
	.w8(32'hbb19e583),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad25f66),
	.w1(32'hba733f0b),
	.w2(32'hbb5771c9),
	.w3(32'hbaa6c0f8),
	.w4(32'h3a26d192),
	.w5(32'hba429d12),
	.w6(32'hbb2fe33e),
	.w7(32'hba9293a6),
	.w8(32'hbbde5a10),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01cc93),
	.w1(32'hbb8d4b2d),
	.w2(32'h3b9f83fd),
	.w3(32'hba2ef156),
	.w4(32'hbc1d943c),
	.w5(32'h3b777706),
	.w6(32'hbbd2ec74),
	.w7(32'hbc029d71),
	.w8(32'hbba883e5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5569bb),
	.w1(32'hbc1afcc3),
	.w2(32'hbba9664c),
	.w3(32'h3984e3b8),
	.w4(32'h3b851f5b),
	.w5(32'h3c1a59e0),
	.w6(32'h3980e81d),
	.w7(32'hbb5a57b6),
	.w8(32'hbb93539f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a5c9),
	.w1(32'hbbd38a0b),
	.w2(32'hbb20d215),
	.w3(32'h3c354307),
	.w4(32'hbbe2884b),
	.w5(32'hbbad321d),
	.w6(32'hba354b34),
	.w7(32'hbc0cd35e),
	.w8(32'hbc2c409e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005407),
	.w1(32'h3bb02edc),
	.w2(32'hbaee98e5),
	.w3(32'hbbbf462b),
	.w4(32'h3afdac99),
	.w5(32'hbc38d489),
	.w6(32'hbbd32519),
	.w7(32'hb9166866),
	.w8(32'hbba6137a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88bc60),
	.w1(32'h3c214b5c),
	.w2(32'h39a6f439),
	.w3(32'hbbc71ed3),
	.w4(32'h3c659b8f),
	.w5(32'hbc251c11),
	.w6(32'hb9235307),
	.w7(32'h3bfa1432),
	.w8(32'hbbe82af0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addb082),
	.w1(32'h3c021d30),
	.w2(32'h3aaf7ac5),
	.w3(32'hbabea0a1),
	.w4(32'h3b8a4cdd),
	.w5(32'h39a6b634),
	.w6(32'hbb0c93e0),
	.w7(32'hba8665ee),
	.w8(32'hba147f9e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3becd9),
	.w1(32'h3aea25a1),
	.w2(32'h3cf0572c),
	.w3(32'h3b4e68c3),
	.w4(32'hbc831383),
	.w5(32'h3cbb166e),
	.w6(32'h3bf5e837),
	.w7(32'hbbaa05a5),
	.w8(32'h3b9adf51),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51c2ac),
	.w1(32'h3b9d705b),
	.w2(32'hbae31568),
	.w3(32'h3c8eba5b),
	.w4(32'hbaf22cdf),
	.w5(32'hbc5512e0),
	.w6(32'h3c825fb0),
	.w7(32'hbb5f55b8),
	.w8(32'hbbbc17c5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf55ccd),
	.w1(32'h3bf0d1db),
	.w2(32'h3ba94be5),
	.w3(32'hbc0a6ab8),
	.w4(32'h3baecbcb),
	.w5(32'hbbe9b030),
	.w6(32'hbbc7f1e6),
	.w7(32'hb9d0dc26),
	.w8(32'hbb6c2107),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc3b84),
	.w1(32'h39fca715),
	.w2(32'hba93506b),
	.w3(32'hbaa4e06a),
	.w4(32'h3b13b88b),
	.w5(32'hbba3411d),
	.w6(32'h3afe4cbe),
	.w7(32'hbbb34f6d),
	.w8(32'hbc351edc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf42ddf),
	.w1(32'hbb3032b7),
	.w2(32'h3a36a745),
	.w3(32'hbbb94c1a),
	.w4(32'hbb87f380),
	.w5(32'h3b684758),
	.w6(32'hbc2b2e03),
	.w7(32'h3b586769),
	.w8(32'h3b16c11c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c441f),
	.w1(32'h39028f54),
	.w2(32'hbb1ae76e),
	.w3(32'h3b4294e8),
	.w4(32'hbacc6b94),
	.w5(32'hb8073bb5),
	.w6(32'h3b9821fd),
	.w7(32'hbb37cb85),
	.w8(32'h3a9f126f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0833f),
	.w1(32'hbbbf91d1),
	.w2(32'hbb025039),
	.w3(32'h3bf102e8),
	.w4(32'hbc8c94d5),
	.w5(32'h3bfb8135),
	.w6(32'h3adb15dd),
	.w7(32'hbbde404e),
	.w8(32'hbbb269e3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba1c33),
	.w1(32'h3c042eb3),
	.w2(32'h3b8518bb),
	.w3(32'hbba3fc41),
	.w4(32'hb78bc130),
	.w5(32'h3bf68111),
	.w6(32'h3b19129c),
	.w7(32'hbb396cae),
	.w8(32'h3b8429aa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d57ea),
	.w1(32'hbab2f05f),
	.w2(32'hbb9246f2),
	.w3(32'h3b927aab),
	.w4(32'hbbe3b9c4),
	.w5(32'hbb5ad378),
	.w6(32'hbb0680c2),
	.w7(32'hbc2375f6),
	.w8(32'hbb27747e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc498f2b),
	.w1(32'h3b25dca1),
	.w2(32'h3ccae620),
	.w3(32'hbc0bad9d),
	.w4(32'h3ccd989b),
	.w5(32'h3d0b1ac9),
	.w6(32'h3937839c),
	.w7(32'hbba5d6a3),
	.w8(32'hbb8e7f60),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6586a),
	.w1(32'hba8bd4f4),
	.w2(32'h3b2b914f),
	.w3(32'h3b8eb450),
	.w4(32'h3b4f67a9),
	.w5(32'hb94dc11f),
	.w6(32'hbbc60a28),
	.w7(32'h3a931aff),
	.w8(32'hbc04d8b1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f0f7d),
	.w1(32'hbbef1463),
	.w2(32'hbbf9d0f9),
	.w3(32'hbb069cce),
	.w4(32'hbbd83edf),
	.w5(32'h3c2db100),
	.w6(32'hbbea1b92),
	.w7(32'hb7693402),
	.w8(32'h39fcb052),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc098f7d),
	.w1(32'h3c224b06),
	.w2(32'hba08b7c9),
	.w3(32'hbba554fc),
	.w4(32'h3b74a1ad),
	.w5(32'hbbf37aee),
	.w6(32'hbb2ae7a6),
	.w7(32'hbb8651ae),
	.w8(32'hbafdd0c3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dcc55),
	.w1(32'hbb627f6b),
	.w2(32'hbb2f13c2),
	.w3(32'h3a82015e),
	.w4(32'h3983566a),
	.w5(32'hba12e319),
	.w6(32'hba3683c8),
	.w7(32'h3b8042b9),
	.w8(32'h3b20a524),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06eecb),
	.w1(32'h3bb5e220),
	.w2(32'hb7d3b27d),
	.w3(32'h3b5d1d60),
	.w4(32'hbb0dde1e),
	.w5(32'hbb8cd889),
	.w6(32'h3aaf43f4),
	.w7(32'hba9d6478),
	.w8(32'hbbe4261e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bdc46),
	.w1(32'hbb306eb2),
	.w2(32'hbb9ed81b),
	.w3(32'hbc5df2a9),
	.w4(32'h3add42df),
	.w5(32'hbbdf7db6),
	.w6(32'hbbb79445),
	.w7(32'hbb892acc),
	.w8(32'hbb1c168b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bdf20),
	.w1(32'h3baff53e),
	.w2(32'h3cf6b022),
	.w3(32'h3aa69df0),
	.w4(32'h3c9653d4),
	.w5(32'h3cd771e7),
	.w6(32'hbbd896a4),
	.w7(32'hbbfaf29a),
	.w8(32'h3acc504b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d6553),
	.w1(32'h3b7df389),
	.w2(32'h3c1a9cf1),
	.w3(32'hbb6e0ea5),
	.w4(32'h3ae98420),
	.w5(32'h3c3d12d3),
	.w6(32'hbac23b89),
	.w7(32'hbc082f0f),
	.w8(32'h3a75e925),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b929ae0),
	.w1(32'h3c4f9df2),
	.w2(32'h3c2a420e),
	.w3(32'hbbd7d565),
	.w4(32'h3b7a1316),
	.w5(32'h3b05c1e5),
	.w6(32'hbc3132aa),
	.w7(32'hbb4a9779),
	.w8(32'hbb94537f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b843a76),
	.w1(32'h3a26c65b),
	.w2(32'hbae50426),
	.w3(32'h3b679985),
	.w4(32'h39b4cdf5),
	.w5(32'hbb17ab89),
	.w6(32'h3ba57379),
	.w7(32'h3a169f1e),
	.w8(32'h3a23e349),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e196f),
	.w1(32'hbb8713e1),
	.w2(32'hbc00c2c4),
	.w3(32'hbb206375),
	.w4(32'h3c304e1f),
	.w5(32'h3cc96523),
	.w6(32'h3b2edc16),
	.w7(32'hbac10c69),
	.w8(32'hb9fcee98),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ac835),
	.w1(32'h3a6facf3),
	.w2(32'hbba5ddbd),
	.w3(32'h3c282c2d),
	.w4(32'hba467ddd),
	.w5(32'hbbdfabf5),
	.w6(32'h3a843578),
	.w7(32'hbb640dc8),
	.w8(32'hbbeae3e7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f8895),
	.w1(32'h3adaeb06),
	.w2(32'h3b285d1a),
	.w3(32'hbba8fa90),
	.w4(32'hbabd6056),
	.w5(32'hbbac6950),
	.w6(32'hbc1efdc0),
	.w7(32'h3b823b12),
	.w8(32'h3c04278e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba229587),
	.w1(32'hbaa54d1b),
	.w2(32'hbadde4e6),
	.w3(32'h3aba0db3),
	.w4(32'h3b3220d1),
	.w5(32'h3b48914d),
	.w6(32'h3af7f201),
	.w7(32'hbb495f09),
	.w8(32'hbbc13c40),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292ee4),
	.w1(32'hbb7aeaea),
	.w2(32'hbb1bdcb4),
	.w3(32'h3b2abc31),
	.w4(32'hb9ee1b98),
	.w5(32'h3ac717d0),
	.w6(32'hbbb58609),
	.w7(32'hbb852653),
	.w8(32'hba15166c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7466),
	.w1(32'hbb960b0d),
	.w2(32'hba1e4ac7),
	.w3(32'h3b88d9fd),
	.w4(32'hbbbf0022),
	.w5(32'hbb3a8011),
	.w6(32'hbb07070e),
	.w7(32'hbbb6ae6e),
	.w8(32'h3899a4d0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac610c0),
	.w1(32'h3b8cfb89),
	.w2(32'h3b47014b),
	.w3(32'h39de7224),
	.w4(32'hb71e0afb),
	.w5(32'hba611947),
	.w6(32'h3bbb97d0),
	.w7(32'hb9872bf2),
	.w8(32'h3b3dde0d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1d41),
	.w1(32'h3af7a37d),
	.w2(32'h3780fac7),
	.w3(32'h3ba2ad2f),
	.w4(32'h3aec0535),
	.w5(32'h3b7c0002),
	.w6(32'h3bbbbf0b),
	.w7(32'hbb88a867),
	.w8(32'hbba61ca4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa63a50),
	.w1(32'hbb82f7ba),
	.w2(32'h3b86eba0),
	.w3(32'h3be0d4b5),
	.w4(32'hbbad7f76),
	.w5(32'h3b2862c4),
	.w6(32'h3a175790),
	.w7(32'hbb71a301),
	.w8(32'hbb31d20f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a732439),
	.w1(32'h3b7aa0ed),
	.w2(32'hbb55f15a),
	.w3(32'hb8bbb20b),
	.w4(32'hbb1e941e),
	.w5(32'hbbfa7008),
	.w6(32'h3a823719),
	.w7(32'h39c8059f),
	.w8(32'hbb8a1b19),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28bbe3),
	.w1(32'hbb92d962),
	.w2(32'hbb956f65),
	.w3(32'hbbc1f54d),
	.w4(32'hbb386667),
	.w5(32'hbb8f142c),
	.w6(32'hbb936696),
	.w7(32'hbb9edbe2),
	.w8(32'hbb9cc011),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12944a),
	.w1(32'h3b37d62d),
	.w2(32'hbadc99ab),
	.w3(32'hbae74709),
	.w4(32'h3b26e7e1),
	.w5(32'h3c08c1b5),
	.w6(32'hb7de1bc8),
	.w7(32'hbbb9d8b6),
	.w8(32'hbba45925),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77bb2f),
	.w1(32'hba9947fd),
	.w2(32'hbae8d1fd),
	.w3(32'h3b433bf4),
	.w4(32'hbb8220df),
	.w5(32'hbb1f2ddb),
	.w6(32'hbacd2a85),
	.w7(32'h3a602c08),
	.w8(32'hbb9d570e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4c116),
	.w1(32'h3b284a27),
	.w2(32'hba8e993a),
	.w3(32'hbbcd07f4),
	.w4(32'h3ba5ef95),
	.w5(32'h3b38ee82),
	.w6(32'hba8ef3aa),
	.w7(32'h3a50e98d),
	.w8(32'h39d2c28d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5f76),
	.w1(32'hbb4dce4a),
	.w2(32'h3b0bce0c),
	.w3(32'h3a9bc969),
	.w4(32'h39b047ab),
	.w5(32'hbb01bb86),
	.w6(32'hbb4d4ac8),
	.w7(32'hbb2442f2),
	.w8(32'hbad52b18),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c52a4),
	.w1(32'h3b049863),
	.w2(32'h3a9408be),
	.w3(32'h3a135e5e),
	.w4(32'hbb37bfdf),
	.w5(32'hbabb4337),
	.w6(32'hba5e7cfb),
	.w7(32'hbab1518f),
	.w8(32'hbb41e0f6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7623c3),
	.w1(32'hbb64d594),
	.w2(32'h3aeddc66),
	.w3(32'hba9617cc),
	.w4(32'hba0a3fcd),
	.w5(32'h39d5a8bd),
	.w6(32'h3b90e4bd),
	.w7(32'h3b8c4d4a),
	.w8(32'h3c2ab0b8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a938),
	.w1(32'h3a1fe450),
	.w2(32'hba0cd3a5),
	.w3(32'h3ab0605f),
	.w4(32'hbaf33da7),
	.w5(32'hba34df3b),
	.w6(32'h3c1354b5),
	.w7(32'h3b6d4b53),
	.w8(32'hba243395),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3839b47c),
	.w1(32'h3a5bd45f),
	.w2(32'h39bf1a73),
	.w3(32'hbb7ec8d8),
	.w4(32'hbae32e17),
	.w5(32'hbb39481c),
	.w6(32'hbb43a6b8),
	.w7(32'hbba3194d),
	.w8(32'hbc144a66),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc485a),
	.w1(32'h3be68ceb),
	.w2(32'h38965d59),
	.w3(32'h3bea4283),
	.w4(32'h3bb78fca),
	.w5(32'hb9e00cdc),
	.w6(32'h3983563a),
	.w7(32'h3b93d7dc),
	.w8(32'h3b40ab23),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d824b),
	.w1(32'hbb71afca),
	.w2(32'hbc0ba47a),
	.w3(32'h3b5ac3cd),
	.w4(32'hbabcaa6e),
	.w5(32'hbc0593b2),
	.w6(32'hb9a3de44),
	.w7(32'hbb12f5cf),
	.w8(32'hbc140ec0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76360b),
	.w1(32'h3bbbb76b),
	.w2(32'hb99383cd),
	.w3(32'h39cdc90e),
	.w4(32'h3c13c59f),
	.w5(32'h3c938765),
	.w6(32'hbaf46720),
	.w7(32'hbbb0af01),
	.w8(32'hbbe8be26),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c46ec),
	.w1(32'h3bbb81fe),
	.w2(32'h3b2d1976),
	.w3(32'h3b8a10e7),
	.w4(32'hbb04217b),
	.w5(32'hbb851f1b),
	.w6(32'hbc4938ec),
	.w7(32'h3a1e5ec9),
	.w8(32'hbb2df79d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad87011),
	.w1(32'hbb638731),
	.w2(32'hbb80e5de),
	.w3(32'h3a0c1d3c),
	.w4(32'hbbd2e52b),
	.w5(32'hbbdc4df6),
	.w6(32'h395b93a5),
	.w7(32'hbb0e62ce),
	.w8(32'hba8e6063),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21441b),
	.w1(32'h3b8d3442),
	.w2(32'h3c2a0da9),
	.w3(32'hbbaeff3e),
	.w4(32'hb96a96ab),
	.w5(32'hbb1f6b54),
	.w6(32'h3afe867a),
	.w7(32'hba4a4c09),
	.w8(32'h3bd7d01b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba912142),
	.w1(32'hbb351942),
	.w2(32'h3b5706dc),
	.w3(32'h3a9d2a29),
	.w4(32'hbb0907c7),
	.w5(32'hbbb2406d),
	.w6(32'h3b39edfc),
	.w7(32'h3a86e7b8),
	.w8(32'h3ba94539),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c21fe),
	.w1(32'hbb2e0684),
	.w2(32'h3baf1a16),
	.w3(32'hb86c8eeb),
	.w4(32'hbbe643da),
	.w5(32'hbaa7474a),
	.w6(32'h3a0117e8),
	.w7(32'hbc0560ec),
	.w8(32'hbbefcde1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c4e87),
	.w1(32'hbb241e43),
	.w2(32'hbadd74d9),
	.w3(32'hbb074a35),
	.w4(32'hbbf1872a),
	.w5(32'hbb27809e),
	.w6(32'hbbc69112),
	.w7(32'hbbecee50),
	.w8(32'hbbdf7ad4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac15f32),
	.w1(32'hbb6f4b68),
	.w2(32'hb97f589c),
	.w3(32'hba5b0e69),
	.w4(32'hbb0f5432),
	.w5(32'hbbd3de4c),
	.w6(32'hbbfff02f),
	.w7(32'hbc27a1e8),
	.w8(32'hbc546649),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c979113),
	.w1(32'h3bbacf47),
	.w2(32'hba1c7ce0),
	.w3(32'h3c714a94),
	.w4(32'h3b50b457),
	.w5(32'h3b04aaea),
	.w6(32'hbb06d8d7),
	.w7(32'h3c0645ee),
	.w8(32'h3c3216be),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d0060),
	.w1(32'h3a0ab220),
	.w2(32'h3a43670f),
	.w3(32'hb98dd247),
	.w4(32'hbb74c414),
	.w5(32'h3a9f9dc4),
	.w6(32'h3b98715b),
	.w7(32'hbbb8ddcb),
	.w8(32'hbb9a9dec),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8544b2),
	.w1(32'hbb93c069),
	.w2(32'hbb935be5),
	.w3(32'h3b60b6d2),
	.w4(32'hbb064c1d),
	.w5(32'h3a664bec),
	.w6(32'hbbca1cf8),
	.w7(32'hbbedc1f8),
	.w8(32'hbb9bf3f5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be877),
	.w1(32'h3a91a42d),
	.w2(32'hbb2cd958),
	.w3(32'h39cd9034),
	.w4(32'hbac761a0),
	.w5(32'hbb2991af),
	.w6(32'h3ac5b0dd),
	.w7(32'h3b33bc1f),
	.w8(32'hbb7f923a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd0091),
	.w1(32'hbc179505),
	.w2(32'hbbebbf37),
	.w3(32'hba28688c),
	.w4(32'hbafaf09a),
	.w5(32'h3c001048),
	.w6(32'hbc0314a4),
	.w7(32'hbc04ca22),
	.w8(32'hbc181e97),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c384935),
	.w1(32'hbb542570),
	.w2(32'hbbbb7b7a),
	.w3(32'h3c1e271a),
	.w4(32'hbab983fa),
	.w5(32'hba7eb9be),
	.w6(32'h3bc25d21),
	.w7(32'hbb5f393c),
	.w8(32'h39be7b91),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b3af),
	.w1(32'h3bee4df3),
	.w2(32'h3b805f94),
	.w3(32'hba67678e),
	.w4(32'h3b003214),
	.w5(32'hbac79926),
	.w6(32'hbaaa5d55),
	.w7(32'hbb23689d),
	.w8(32'h3a38aeca),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b363be6),
	.w1(32'h3baf0d18),
	.w2(32'hbae294ab),
	.w3(32'h39e3733b),
	.w4(32'h3bcd6981),
	.w5(32'h3a356ed8),
	.w6(32'h3b8fa637),
	.w7(32'h3b7e8eaf),
	.w8(32'hbb2258a7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14d502),
	.w1(32'hbb0eef1d),
	.w2(32'hba11cb50),
	.w3(32'h3b206895),
	.w4(32'hb9824113),
	.w5(32'h3c178713),
	.w6(32'hbb05fdd9),
	.w7(32'hb9f4e275),
	.w8(32'hbad53239),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90cfd2),
	.w1(32'hba25fcf6),
	.w2(32'hba73a585),
	.w3(32'h3bb617ce),
	.w4(32'hbb852d43),
	.w5(32'h3b294357),
	.w6(32'hba4fd914),
	.w7(32'hbb5efe1c),
	.w8(32'hbb52f88f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a505363),
	.w1(32'hb808f9ac),
	.w2(32'hbb85244d),
	.w3(32'h39ffa868),
	.w4(32'h3aad5e27),
	.w5(32'hbadb22fb),
	.w6(32'hbb84993b),
	.w7(32'hbbbe79fe),
	.w8(32'hbb701f9e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9bd9c),
	.w1(32'hbb8fa1f5),
	.w2(32'hbba4f433),
	.w3(32'h3a5fa321),
	.w4(32'hbba9b1a2),
	.w5(32'hbbb0201c),
	.w6(32'hbb6bb597),
	.w7(32'hbb8b4b67),
	.w8(32'hbbb80bb0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43ff9),
	.w1(32'h3b014fba),
	.w2(32'h3bb500e0),
	.w3(32'hbae6ceb9),
	.w4(32'h3ac4d9d2),
	.w5(32'hbb9521d5),
	.w6(32'hbba41c02),
	.w7(32'hba53319a),
	.w8(32'h3aa73773),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0398f8),
	.w1(32'h3b298146),
	.w2(32'h3b9ad47c),
	.w3(32'h3b1d3449),
	.w4(32'hbc09d16a),
	.w5(32'hb955592e),
	.w6(32'hb9276d3d),
	.w7(32'hbbc49ed0),
	.w8(32'h3b5c49c6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9452fd5),
	.w1(32'hb8974299),
	.w2(32'h3af0404a),
	.w3(32'hb9deda3f),
	.w4(32'hbb2d4bd8),
	.w5(32'h3b2be7d6),
	.w6(32'h3a8d83f3),
	.w7(32'hbb02ac5e),
	.w8(32'hbbd90723),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d3fb1),
	.w1(32'h3b693c8e),
	.w2(32'h3b2e8d4c),
	.w3(32'h3a74c089),
	.w4(32'h3b872bf0),
	.w5(32'h3a068fc9),
	.w6(32'hbb2c75c9),
	.w7(32'h3af58925),
	.w8(32'h3a26729b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34749b),
	.w1(32'h3ae9b0cb),
	.w2(32'h3b81330b),
	.w3(32'h395d6cdc),
	.w4(32'h3b2b2cce),
	.w5(32'hbb6be6f3),
	.w6(32'h3a9c23f6),
	.w7(32'h392eb3da),
	.w8(32'h3b8d7b18),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3b79),
	.w1(32'h3b28a2f0),
	.w2(32'hba15a01c),
	.w3(32'h3bb2a7f0),
	.w4(32'hbb7d0d90),
	.w5(32'h3a437f46),
	.w6(32'h3b495e19),
	.w7(32'h3add15c2),
	.w8(32'hbb713577),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f899),
	.w1(32'hb98ce94b),
	.w2(32'h3b6f39d0),
	.w3(32'hbaa6dc46),
	.w4(32'hbacfad5e),
	.w5(32'hba89133b),
	.w6(32'hbbe44498),
	.w7(32'hba5e1651),
	.w8(32'h3c0ae0d8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09935e),
	.w1(32'hbbc1ab1d),
	.w2(32'hba840f00),
	.w3(32'hba22a9ca),
	.w4(32'hba1bc355),
	.w5(32'hbb05fe4e),
	.w6(32'h3ae0d8ba),
	.w7(32'hbbb678a0),
	.w8(32'hbbdb298e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd427a4),
	.w1(32'h3ac9bf55),
	.w2(32'h3a85e3aa),
	.w3(32'hbb9b206e),
	.w4(32'h39dfab66),
	.w5(32'h3a8eb598),
	.w6(32'hbafa2857),
	.w7(32'h3b28b8ff),
	.w8(32'h3ad02f82),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5fabb),
	.w1(32'h3a195536),
	.w2(32'hb8e9fc3e),
	.w3(32'h3abed605),
	.w4(32'h3a793016),
	.w5(32'hbaeff9c2),
	.w6(32'h3ba17da7),
	.w7(32'h3a822953),
	.w8(32'hbaf4ab64),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae29f9),
	.w1(32'h39aca733),
	.w2(32'hb841d3de),
	.w3(32'hbacd1382),
	.w4(32'hbb01edce),
	.w5(32'hbbc2ec68),
	.w6(32'h3a51d6b7),
	.w7(32'hba075e62),
	.w8(32'hba1b51a5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984115a),
	.w1(32'hbb0262a0),
	.w2(32'hbb529d85),
	.w3(32'hbb5abb27),
	.w4(32'h3a18a702),
	.w5(32'hbc1bff3b),
	.w6(32'h3b2ae6f1),
	.w7(32'h3a80622f),
	.w8(32'hbac57e55),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52c871),
	.w1(32'hbadf9e3e),
	.w2(32'hbaf64dce),
	.w3(32'hbb1bfe5b),
	.w4(32'h3c3f98a1),
	.w5(32'h3c93dae7),
	.w6(32'hbb9d2c4d),
	.w7(32'h3b9da1da),
	.w8(32'h3be66f9b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeff9e0),
	.w1(32'hbb613831),
	.w2(32'hbb53c517),
	.w3(32'h3bb47f49),
	.w4(32'hbb693c2a),
	.w5(32'h3c3f69f9),
	.w6(32'h3b1d2896),
	.w7(32'hbb72ffbb),
	.w8(32'hbbb120d8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b310f4a),
	.w1(32'hbb46f1e8),
	.w2(32'hbb39550e),
	.w3(32'h3beb9c91),
	.w4(32'hbbd159d5),
	.w5(32'hbbe0d1e3),
	.w6(32'hba90383b),
	.w7(32'h3a66899b),
	.w8(32'hbb3b343c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87e677),
	.w1(32'hbbb016c8),
	.w2(32'hbb3e97ab),
	.w3(32'hbbbb841d),
	.w4(32'hbb10af2a),
	.w5(32'hbb2e7e6e),
	.w6(32'hbc0a8e39),
	.w7(32'hbb910e95),
	.w8(32'hbbbb1011),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9fefb),
	.w1(32'hbbd14c16),
	.w2(32'hbba77bb3),
	.w3(32'hbb9381ad),
	.w4(32'hbbd899f3),
	.w5(32'hb9a7f40e),
	.w6(32'hbb8535d3),
	.w7(32'hbbb2816a),
	.w8(32'hbbc3656a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe75322),
	.w1(32'hbb4fa1db),
	.w2(32'hb9ff179a),
	.w3(32'hbad64e2b),
	.w4(32'hbb692bbf),
	.w5(32'h39381117),
	.w6(32'hba7a46d7),
	.w7(32'hbbabe21f),
	.w8(32'hbbab0910),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2166d),
	.w1(32'hbb8115f8),
	.w2(32'hb8bcbb99),
	.w3(32'h3bd38b66),
	.w4(32'hbb078405),
	.w5(32'hbab3c9dc),
	.w6(32'h3a809d0a),
	.w7(32'hb9b4cfa8),
	.w8(32'h3b2fa78e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe31a3),
	.w1(32'hba66f1f1),
	.w2(32'hbb135170),
	.w3(32'h3b01916a),
	.w4(32'h3b670883),
	.w5(32'h3c8d808b),
	.w6(32'h3b67bb30),
	.w7(32'hbad8575d),
	.w8(32'h3adec6b3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5636b1),
	.w1(32'h3a3cb5e9),
	.w2(32'h3aa052c0),
	.w3(32'h3c3787f0),
	.w4(32'hba8f78c0),
	.w5(32'hbb16ef36),
	.w6(32'hba0b11ae),
	.w7(32'hbac42c24),
	.w8(32'hbb4ecc59),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f12c3),
	.w1(32'h38a67021),
	.w2(32'hbad1d3e2),
	.w3(32'hbb0359f6),
	.w4(32'hbb3098c0),
	.w5(32'hbb620ea4),
	.w6(32'hbb983eab),
	.w7(32'h3a42aa7b),
	.w8(32'hb627c07b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb141839),
	.w1(32'hbbe064b5),
	.w2(32'hbb1179b7),
	.w3(32'hbaebd29a),
	.w4(32'hbbb5c999),
	.w5(32'hbbc9c0d6),
	.w6(32'hbb96dcd0),
	.w7(32'hbbc362eb),
	.w8(32'h3a838c8a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f1c1b),
	.w1(32'hb9914504),
	.w2(32'hbb2e073a),
	.w3(32'hba8a4b0e),
	.w4(32'hbb0a0eed),
	.w5(32'hbb604aed),
	.w6(32'hbb1a1941),
	.w7(32'h3bbc1657),
	.w8(32'h3ba6b27a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf72a2a),
	.w1(32'hbb8cf68e),
	.w2(32'hbb84f11b),
	.w3(32'h39521e7e),
	.w4(32'hbbb5dad1),
	.w5(32'hbbbe26cd),
	.w6(32'hb9d40534),
	.w7(32'hbae66b16),
	.w8(32'hbb940481),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbac9c),
	.w1(32'hbb84d15a),
	.w2(32'hbb8ef0c1),
	.w3(32'hbba956bc),
	.w4(32'hbaa694d3),
	.w5(32'h3b14fb22),
	.w6(32'hbc080824),
	.w7(32'hb996d906),
	.w8(32'hbbbab4ff),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c740),
	.w1(32'h39370615),
	.w2(32'h3b2e73b2),
	.w3(32'h3a685f2c),
	.w4(32'h3b92e9fb),
	.w5(32'h3be9c4e4),
	.w6(32'hbac44056),
	.w7(32'hbb000620),
	.w8(32'h3a67ff7b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf51da),
	.w1(32'hbbd3285a),
	.w2(32'hbb81ebf8),
	.w3(32'h3c19b598),
	.w4(32'hbbb8fcea),
	.w5(32'hbb2a44a6),
	.w6(32'h3b1cb16e),
	.w7(32'hbbd4ff4d),
	.w8(32'hbaa35d2e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec6c7c),
	.w1(32'h3ad30b0b),
	.w2(32'h3a8f8f67),
	.w3(32'hbb3448c6),
	.w4(32'hbac705ad),
	.w5(32'h3ac1e7ce),
	.w6(32'h396687ff),
	.w7(32'hbbb9ecd0),
	.w8(32'hbbcba0b2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45f0ee),
	.w1(32'h3b6dd549),
	.w2(32'hbad4e2dc),
	.w3(32'h3b3dbd57),
	.w4(32'h3be53bbb),
	.w5(32'h3c40f3a4),
	.w6(32'h3c01926f),
	.w7(32'hbb0a436a),
	.w8(32'hba5381cf),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9e84d),
	.w1(32'hbb01f1b6),
	.w2(32'hbacb0726),
	.w3(32'h3b656adc),
	.w4(32'h3a92f5b5),
	.w5(32'hbb45dfc5),
	.w6(32'hbb5ca00f),
	.w7(32'hb9c7719d),
	.w8(32'hbb36f295),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a065bde),
	.w1(32'hb935b8d7),
	.w2(32'h3b1ed9cb),
	.w3(32'hbb423b87),
	.w4(32'h3b41fe63),
	.w5(32'h3a0cb4a1),
	.w6(32'hbb0b7bfb),
	.w7(32'h3b4e4119),
	.w8(32'h3bd369dd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d5b7a),
	.w1(32'hbb1d814d),
	.w2(32'hbb9cf71c),
	.w3(32'h3aba34e9),
	.w4(32'hbab1fe93),
	.w5(32'hb99e2518),
	.w6(32'h3b48d27f),
	.w7(32'h370514d5),
	.w8(32'hb8092f3c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad36c4b),
	.w1(32'h39969ded),
	.w2(32'hbb6d1e53),
	.w3(32'h39e8a260),
	.w4(32'hbb96dabd),
	.w5(32'hba86ae79),
	.w6(32'h39671248),
	.w7(32'hbb1ff1d5),
	.w8(32'hb96d3d75),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22a681),
	.w1(32'h3b07c656),
	.w2(32'h3b69df72),
	.w3(32'hbbcf2f8a),
	.w4(32'hbb91c452),
	.w5(32'hbbb0a006),
	.w6(32'hbbb1f2f2),
	.w7(32'hbafda5f3),
	.w8(32'hba53c9a5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4372),
	.w1(32'hbb6fc537),
	.w2(32'hbb0acb04),
	.w3(32'hba87180f),
	.w4(32'hbb37cacc),
	.w5(32'hbbdcb055),
	.w6(32'hba916844),
	.w7(32'hbb287552),
	.w8(32'hbb6f60d4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accaeb8),
	.w1(32'h3b8918da),
	.w2(32'h3b0a7b05),
	.w3(32'hbb1959c8),
	.w4(32'hbaf2f724),
	.w5(32'hbaff2a30),
	.w6(32'hbadc2c57),
	.w7(32'h3b044b6a),
	.w8(32'h3b353a6e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b250c31),
	.w1(32'hba9bd2c6),
	.w2(32'h3ba3746a),
	.w3(32'hbb58acb8),
	.w4(32'hbb59c86f),
	.w5(32'h3b13f79b),
	.w6(32'h3b2b859f),
	.w7(32'hba8c5123),
	.w8(32'hbb1bbcc9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01d512),
	.w1(32'h3a18485d),
	.w2(32'h3acf54ae),
	.w3(32'hba58f350),
	.w4(32'hbade686d),
	.w5(32'hbb5ebdad),
	.w6(32'h3ae30173),
	.w7(32'hba90f066),
	.w8(32'h3af8630d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38caa2),
	.w1(32'hbb3ff42d),
	.w2(32'hbbb4c5db),
	.w3(32'h3b360e32),
	.w4(32'hbc06629e),
	.w5(32'hbc5551d5),
	.w6(32'h3989858f),
	.w7(32'hbb8d46b2),
	.w8(32'hbc1ff890),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd86b64),
	.w1(32'hbb62b26f),
	.w2(32'hbb343e96),
	.w3(32'hbc5e676c),
	.w4(32'hbb73868e),
	.w5(32'hbb5e7c79),
	.w6(32'hbc296edb),
	.w7(32'hbb9d4c58),
	.w8(32'hbb19bc90),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1c01),
	.w1(32'h3c0221d3),
	.w2(32'h3be33fa9),
	.w3(32'hba060ec9),
	.w4(32'h3af00301),
	.w5(32'hbb8b7c53),
	.w6(32'hb8da6b5d),
	.w7(32'h3bb10e52),
	.w8(32'h3bbeeb8b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12bf60),
	.w1(32'hbb865eda),
	.w2(32'hba7156f7),
	.w3(32'hba25106c),
	.w4(32'hbad75501),
	.w5(32'hbb832c2f),
	.w6(32'h3b966384),
	.w7(32'hbb6fd3b0),
	.w8(32'hbb3d9fbd),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24ccac),
	.w1(32'h3b45f084),
	.w2(32'hba25f184),
	.w3(32'hbb5ee82c),
	.w4(32'h3ba49791),
	.w5(32'hbb405000),
	.w6(32'h3a8daf28),
	.w7(32'h3ae3e963),
	.w8(32'hbb5103f7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1665a3),
	.w1(32'hbb169a8a),
	.w2(32'hbb9c3879),
	.w3(32'hba8d15fc),
	.w4(32'hba8f735c),
	.w5(32'hbb71d863),
	.w6(32'hbb07363c),
	.w7(32'hbb9d74f4),
	.w8(32'hbbc0df39),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5563d),
	.w1(32'h3b83f03e),
	.w2(32'hbb3f5f03),
	.w3(32'h39d12fbf),
	.w4(32'hbaaf1cd8),
	.w5(32'h3a5e0997),
	.w6(32'hbb228a27),
	.w7(32'hbb00717c),
	.w8(32'hbb2b3655),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51be56),
	.w1(32'h3a96c1f1),
	.w2(32'hbae0e1be),
	.w3(32'hb98ae3f3),
	.w4(32'h39e3e5d7),
	.w5(32'hba49c2b5),
	.w6(32'hbb1ed827),
	.w7(32'h3b33d0ae),
	.w8(32'h3b2f1fcc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b252b61),
	.w1(32'hbb2ac14d),
	.w2(32'hba739898),
	.w3(32'h389101c7),
	.w4(32'hba0524a4),
	.w5(32'hbbc0418b),
	.w6(32'h3b80b27f),
	.w7(32'h39de542d),
	.w8(32'hba00bc80),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacb768),
	.w1(32'h3b3831e8),
	.w2(32'h3bde2bd2),
	.w3(32'hbaaf41ee),
	.w4(32'hbaa9797d),
	.w5(32'hbb93f017),
	.w6(32'h3b20cd1d),
	.w7(32'hbb78a981),
	.w8(32'h3ab7ae34),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04047d),
	.w1(32'hba39d68b),
	.w2(32'h3b2b6997),
	.w3(32'h3ab77dc3),
	.w4(32'hba6b3140),
	.w5(32'hbb81f1f1),
	.w6(32'h3ba431e2),
	.w7(32'h3a877be1),
	.w8(32'h3af08e10),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabecfd),
	.w1(32'h3bc3ee3d),
	.w2(32'h39b77d6a),
	.w3(32'h3a6ed425),
	.w4(32'h3a8b8824),
	.w5(32'h3bc75058),
	.w6(32'hbb201163),
	.w7(32'hbbb68748),
	.w8(32'hbb91443e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385423c2),
	.w1(32'hba96b40b),
	.w2(32'hbb6ded6d),
	.w3(32'h3bef3798),
	.w4(32'hbad2c18b),
	.w5(32'h3ba689e9),
	.w6(32'hbb841f23),
	.w7(32'h3b05da45),
	.w8(32'hba6b1170),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac76b),
	.w1(32'h3b763de2),
	.w2(32'h3c1100fc),
	.w3(32'hbac65673),
	.w4(32'h3af329a8),
	.w5(32'h3b8df87d),
	.w6(32'hbb302f5c),
	.w7(32'h36e19cb0),
	.w8(32'h3b36d323),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3eec7),
	.w1(32'h3accd361),
	.w2(32'hba05264c),
	.w3(32'h3b950fa3),
	.w4(32'h3b86ed45),
	.w5(32'hbb28ab1d),
	.w6(32'h3bc5ae29),
	.w7(32'h3b7e1202),
	.w8(32'hba75bd31),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fa60),
	.w1(32'hba0832bc),
	.w2(32'h3b3f7c6d),
	.w3(32'h3b958838),
	.w4(32'hbb6b2388),
	.w5(32'hbbad2efc),
	.w6(32'h3c1def14),
	.w7(32'h3a4e3b36),
	.w8(32'h3b3f8700),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e26e),
	.w1(32'h3bc19a0c),
	.w2(32'hbb09169f),
	.w3(32'hbae5b567),
	.w4(32'h3ab72fc9),
	.w5(32'hb96339e9),
	.w6(32'hba4c8df2),
	.w7(32'hb7666086),
	.w8(32'hbbc5f881),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0305be),
	.w1(32'hbaa56ab4),
	.w2(32'hbb3c52eb),
	.w3(32'hba25645b),
	.w4(32'h3bc7d0c2),
	.w5(32'h3c310550),
	.w6(32'hbba10706),
	.w7(32'hbc2ce307),
	.w8(32'hbc4b2fa7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be87fe3),
	.w1(32'h3a9786b0),
	.w2(32'hba88c1a4),
	.w3(32'h3b164811),
	.w4(32'hbb53a1c9),
	.w5(32'hbbe35cf3),
	.w6(32'hbb5355ff),
	.w7(32'h3a7581b6),
	.w8(32'hbb01d92d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76a0d0),
	.w1(32'hb7bce946),
	.w2(32'hbb3d9500),
	.w3(32'hbba09b58),
	.w4(32'hbb474c55),
	.w5(32'h3bc9e6f7),
	.w6(32'hbb7b7d1a),
	.w7(32'hbba2ca47),
	.w8(32'hbbaab9d9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fef197),
	.w1(32'hbb15d1c2),
	.w2(32'hbb07b5c4),
	.w3(32'h3aa8abd2),
	.w4(32'hbb544e7c),
	.w5(32'h394d6c8d),
	.w6(32'hbad0c98d),
	.w7(32'hbb8e6715),
	.w8(32'h3af3a2ef),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0fe26),
	.w1(32'h3c04ad00),
	.w2(32'h3ba06b61),
	.w3(32'hbac28c3a),
	.w4(32'h3b2c8e7d),
	.w5(32'hbb13b5e2),
	.w6(32'hbbdd3060),
	.w7(32'h3afc44f6),
	.w8(32'hbb786edb),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a323dad),
	.w1(32'hbb3586b5),
	.w2(32'hbb85d5e3),
	.w3(32'h3b265f49),
	.w4(32'h3b552eed),
	.w5(32'h3b2717e1),
	.w6(32'hbb89a73c),
	.w7(32'hb9a41659),
	.w8(32'h3b23ce59),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a950f),
	.w1(32'h3a8c41a3),
	.w2(32'h399afc52),
	.w3(32'h39d56f68),
	.w4(32'h3ad33980),
	.w5(32'h3c0d80cd),
	.w6(32'hbbb110ff),
	.w7(32'hbbfad8bf),
	.w8(32'hbc4242ab),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbaa3a),
	.w1(32'hbb54179e),
	.w2(32'hbac7e4e6),
	.w3(32'h3bad79cd),
	.w4(32'hba7b0a38),
	.w5(32'hbb6b6980),
	.w6(32'hbb86f715),
	.w7(32'hba642e0b),
	.w8(32'hbb7c4751),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90801),
	.w1(32'h3baa377f),
	.w2(32'h3a9c0128),
	.w3(32'hbbc846f7),
	.w4(32'h3ad0de8b),
	.w5(32'hba82a1d7),
	.w6(32'hbbbe3aae),
	.w7(32'h3bee3bd5),
	.w8(32'h3bc3c76c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb746193),
	.w1(32'h3ad653e6),
	.w2(32'h3b80d878),
	.w3(32'hbc088725),
	.w4(32'h3b982717),
	.w5(32'h3b44c932),
	.w6(32'hbb9855d7),
	.w7(32'h3ac78eaf),
	.w8(32'h3b4003e6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03eb56),
	.w1(32'h3b213307),
	.w2(32'h3bbd4303),
	.w3(32'hbbad189f),
	.w4(32'h3a5bd760),
	.w5(32'h3ac89890),
	.w6(32'h3a1975f4),
	.w7(32'h3af9a511),
	.w8(32'h391dcb1e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b207d9e),
	.w1(32'hbbda327d),
	.w2(32'h3b2270a1),
	.w3(32'h3b5c953e),
	.w4(32'hbb982001),
	.w5(32'hbaccf15f),
	.w6(32'h3b76ccda),
	.w7(32'hbbe96ba6),
	.w8(32'hbbd6ade0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9228f),
	.w1(32'hbaf25dfe),
	.w2(32'hbacfcbe4),
	.w3(32'hbb096db3),
	.w4(32'hbac2145b),
	.w5(32'hbbc78b48),
	.w6(32'hbbaa1799),
	.w7(32'h3aaf2adb),
	.w8(32'hb8f6fb8d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8ba8d),
	.w1(32'hb9d3305e),
	.w2(32'hbb79cd6d),
	.w3(32'hbb833d91),
	.w4(32'hb881bd40),
	.w5(32'hbb89e1e7),
	.w6(32'hbaff2876),
	.w7(32'hba05706a),
	.w8(32'hba50bc09),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80aa92),
	.w1(32'hbb31a2f3),
	.w2(32'hbc0d0dbd),
	.w3(32'hbb015d23),
	.w4(32'hbade6a6e),
	.w5(32'hbb8cb397),
	.w6(32'h3b063abf),
	.w7(32'hbae2e432),
	.w8(32'hbc07c079),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082d3c),
	.w1(32'h397491a1),
	.w2(32'hbb7308a8),
	.w3(32'hbb7a1038),
	.w4(32'hba3a9444),
	.w5(32'hbbeb7548),
	.w6(32'hbbb33a16),
	.w7(32'hbbe7ce8d),
	.w8(32'hbc559b17),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba098c40),
	.w1(32'hb96fef09),
	.w2(32'hbb5c7e98),
	.w3(32'h3ad1917e),
	.w4(32'hbaf354cd),
	.w5(32'hbb29d716),
	.w6(32'hbb214d52),
	.w7(32'hbb9e384f),
	.w8(32'hbbd00742),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fb1d85),
	.w1(32'h3a08faa2),
	.w2(32'h3b3a1057),
	.w3(32'h3b4a3a98),
	.w4(32'hbab97a2c),
	.w5(32'h3b1483cf),
	.w6(32'hba88d3bd),
	.w7(32'h397606a7),
	.w8(32'hbb13ed65),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe5e16),
	.w1(32'hbb69773e),
	.w2(32'hbb2cdb08),
	.w3(32'h392f36ef),
	.w4(32'hbbc37626),
	.w5(32'hbb73683d),
	.w6(32'hbaa9ae74),
	.w7(32'hbbae26c5),
	.w8(32'hbb948835),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a69b),
	.w1(32'hbb71c102),
	.w2(32'hbbae38fc),
	.w3(32'h3adf4a07),
	.w4(32'hbbb99264),
	.w5(32'hbb8bb2c6),
	.w6(32'hb8b087a7),
	.w7(32'hbb46c333),
	.w8(32'hbc2f3ff2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c3833),
	.w1(32'h3c32c25b),
	.w2(32'hba403d7d),
	.w3(32'h3add1e32),
	.w4(32'h3b53f37e),
	.w5(32'hba39e509),
	.w6(32'hbba48680),
	.w7(32'hbb32e694),
	.w8(32'hbb85ff71),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba712f3a),
	.w1(32'hbb20f3a7),
	.w2(32'hbb84d1dd),
	.w3(32'hba8e0ad0),
	.w4(32'hb9656c39),
	.w5(32'hbc0b27fd),
	.w6(32'hba897e23),
	.w7(32'hb9dd77f0),
	.w8(32'hbb845a1d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964aebd),
	.w1(32'hb9bd94fd),
	.w2(32'hba27e4e0),
	.w3(32'hbab8f4cf),
	.w4(32'hbb10b057),
	.w5(32'h3b13a444),
	.w6(32'hbb669982),
	.w7(32'hbb1eef40),
	.w8(32'hbafd6572),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b795fb9),
	.w1(32'hbb1281dd),
	.w2(32'hbaad2b16),
	.w3(32'hba8fdcce),
	.w4(32'hbb73608f),
	.w5(32'hbb803de0),
	.w6(32'hbab05531),
	.w7(32'hbb52c863),
	.w8(32'hbb0563c4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff53e3),
	.w1(32'h3bdc4bad),
	.w2(32'hba2bb0f4),
	.w3(32'hbb4e43ec),
	.w4(32'h3b134b59),
	.w5(32'hba77b7be),
	.w6(32'h39d52ed5),
	.w7(32'h3b4c5095),
	.w8(32'hba125e47),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac2ff5),
	.w1(32'hbb531173),
	.w2(32'hba9c838b),
	.w3(32'h3afc0ac0),
	.w4(32'hba914d2a),
	.w5(32'hbb93bc20),
	.w6(32'h3b249993),
	.w7(32'h3b0c34ca),
	.w8(32'h3b6930bd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a2035),
	.w1(32'hbbbc60c1),
	.w2(32'hbb37ff14),
	.w3(32'hbbf68469),
	.w4(32'hbb0be083),
	.w5(32'h3af8aa03),
	.w6(32'hbc14c0d8),
	.w7(32'h3baa3496),
	.w8(32'h3b9adc1d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf85813),
	.w1(32'hbb0859a9),
	.w2(32'hbbab7a79),
	.w3(32'h3982c975),
	.w4(32'hbbf651fd),
	.w5(32'hbb444987),
	.w6(32'h3ad4bfc4),
	.w7(32'hbb00bbef),
	.w8(32'h39fbb2e1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7bc9c),
	.w1(32'hbb80edc7),
	.w2(32'h3bb476bf),
	.w3(32'hbb8dc525),
	.w4(32'hbb58229f),
	.w5(32'h3b44ade3),
	.w6(32'hbb393a5c),
	.w7(32'hbb6cd4a1),
	.w8(32'hbaff9efb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b6928),
	.w1(32'hbbb5c65d),
	.w2(32'hbb91a58f),
	.w3(32'h3a0ea24d),
	.w4(32'hbb566932),
	.w5(32'hbb499f0a),
	.w6(32'hba008546),
	.w7(32'hbbcac96b),
	.w8(32'hbc346f85),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd560),
	.w1(32'hba81263d),
	.w2(32'hbb2ba63e),
	.w3(32'h3ae8ca4e),
	.w4(32'h3a9d1572),
	.w5(32'h3b9d8c82),
	.w6(32'h3b3a656d),
	.w7(32'h3ba55a36),
	.w8(32'h3c1e49dc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c2fbb),
	.w1(32'h3b3497b3),
	.w2(32'h3aac3607),
	.w3(32'h3b16888b),
	.w4(32'hbb0cf0bd),
	.w5(32'hbb87eb01),
	.w6(32'h3b0fb3a0),
	.w7(32'h38b9c723),
	.w8(32'hbbd4ae1b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8062c6),
	.w1(32'hba8d076e),
	.w2(32'h3c2a7530),
	.w3(32'hbb96e1b1),
	.w4(32'hba80dd71),
	.w5(32'h3be229f2),
	.w6(32'hba8087ab),
	.w7(32'hbb75b5ba),
	.w8(32'h3a4e2312),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85d94b),
	.w1(32'h3a0e326a),
	.w2(32'h3a8fce12),
	.w3(32'h3ba281cf),
	.w4(32'hbac73980),
	.w5(32'hba717796),
	.w6(32'h3b6d5849),
	.w7(32'h3ab91121),
	.w8(32'hba683c97),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae60c95),
	.w1(32'hbbe273fc),
	.w2(32'hbb5a50c4),
	.w3(32'h3b72dac7),
	.w4(32'hbc0804b0),
	.w5(32'hbbb20db2),
	.w6(32'hbabf0959),
	.w7(32'hbbf1b59d),
	.w8(32'hbbdc7f5c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe07c69),
	.w1(32'h3bad04f9),
	.w2(32'h3b7390bc),
	.w3(32'hbbd1e1a9),
	.w4(32'h3b8e37df),
	.w5(32'h3b29b8af),
	.w6(32'hbbb4464d),
	.w7(32'h3b6dac64),
	.w8(32'h3a9b871a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92fc01),
	.w1(32'h3aab4de4),
	.w2(32'h3b88a424),
	.w3(32'h3b4a6dc4),
	.w4(32'h3a77ea0d),
	.w5(32'h3a743e60),
	.w6(32'h3b8134bf),
	.w7(32'hbb72b8bb),
	.w8(32'hbbb2854f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8d2c2),
	.w1(32'hba38bc27),
	.w2(32'h3b72ac78),
	.w3(32'hbac4eb1e),
	.w4(32'hbb75db50),
	.w5(32'hbb63ff2e),
	.w6(32'hbba5a327),
	.w7(32'h39403662),
	.w8(32'h3b3dadd1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c621),
	.w1(32'h3aa754d9),
	.w2(32'hba2a70dd),
	.w3(32'h3aa60da2),
	.w4(32'h3b06ef5c),
	.w5(32'hba7e0723),
	.w6(32'h39be4f65),
	.w7(32'h3b111993),
	.w8(32'hba0b1004),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba269140),
	.w1(32'hba34883e),
	.w2(32'h3b0833b2),
	.w3(32'h3ab524b6),
	.w4(32'hbb1c2727),
	.w5(32'h3a4d6edf),
	.w6(32'h3a6b84ec),
	.w7(32'hbba6eea5),
	.w8(32'hbb65d061),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1774a),
	.w1(32'h3add8c25),
	.w2(32'h3b86ddca),
	.w3(32'hba02a8f6),
	.w4(32'hbaf92aaa),
	.w5(32'h3b5442c1),
	.w6(32'hbb15e8c3),
	.w7(32'hba0cd74f),
	.w8(32'h3ae11e10),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e2cb),
	.w1(32'hba08ed02),
	.w2(32'hba94ec00),
	.w3(32'h39f7c2d4),
	.w4(32'hbb5388ca),
	.w5(32'hbb2c7761),
	.w6(32'h3aa9995b),
	.w7(32'hbacf05dc),
	.w8(32'hbb067d97),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b412193),
	.w1(32'h3b277247),
	.w2(32'hbace92cf),
	.w3(32'hb9f29758),
	.w4(32'hbac8adb4),
	.w5(32'hbb3e6da1),
	.w6(32'hbb0a417c),
	.w7(32'h3b1ee2e3),
	.w8(32'hb950720d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb40b0b),
	.w1(32'h3bb516c5),
	.w2(32'h39d13c20),
	.w3(32'h3abaa77d),
	.w4(32'h3b884df2),
	.w5(32'h3b467718),
	.w6(32'hbba24420),
	.w7(32'h3a1d634c),
	.w8(32'h3bc1135c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9224dc),
	.w1(32'hbb43bcdb),
	.w2(32'hbae29112),
	.w3(32'h3b25391b),
	.w4(32'hbbdc5f91),
	.w5(32'hbc053552),
	.w6(32'hbb12ac6a),
	.w7(32'hbc42c6c1),
	.w8(32'hbc2da06e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1115d8),
	.w1(32'hbb4adaa1),
	.w2(32'hbb66a610),
	.w3(32'hba8e55a4),
	.w4(32'h3b5f8b4d),
	.w5(32'h3c865f3c),
	.w6(32'hbba3b916),
	.w7(32'hbbfc6b54),
	.w8(32'hbac13cef),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c8bf),
	.w1(32'hbbc70e40),
	.w2(32'hbc0ef4f4),
	.w3(32'hba4ddd9c),
	.w4(32'hbabcdcd7),
	.w5(32'hbba3e114),
	.w6(32'hbb752040),
	.w7(32'hbbd9d304),
	.w8(32'hbb713983),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6df65f),
	.w1(32'hba9ae530),
	.w2(32'hbbda0c1f),
	.w3(32'hbaff99d8),
	.w4(32'h3a6f99b8),
	.w5(32'hbac6aa8f),
	.w6(32'hbb5cd2d0),
	.w7(32'hbaa87c4b),
	.w8(32'hbbc4b66a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22abc9),
	.w1(32'h3b9012b6),
	.w2(32'h3b5484f6),
	.w3(32'hba378c72),
	.w4(32'h3b784102),
	.w5(32'h3a87cf78),
	.w6(32'hbbc1f2bf),
	.w7(32'hba4bb294),
	.w8(32'h3b377059),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b415000),
	.w1(32'hbb563d47),
	.w2(32'hbb56b43e),
	.w3(32'h3c1f1498),
	.w4(32'h39fafee0),
	.w5(32'hbb8d90f1),
	.w6(32'h3c0ad64f),
	.w7(32'h3b3b5b0b),
	.w8(32'hbb222386),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bd709),
	.w1(32'hb9b4540f),
	.w2(32'h3b601eb4),
	.w3(32'hbacf7526),
	.w4(32'h3ac19455),
	.w5(32'hb9db210c),
	.w6(32'hbb9a4023),
	.w7(32'hbaf5137c),
	.w8(32'hbbd75e0c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3ec34),
	.w1(32'hb9550f50),
	.w2(32'hbc0a21d0),
	.w3(32'h3c50a8bd),
	.w4(32'h3ac31aec),
	.w5(32'h39ca8ee8),
	.w6(32'h3b8df6f8),
	.w7(32'hbb25c677),
	.w8(32'hbb14960e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1df0),
	.w1(32'h3bdd3bb4),
	.w2(32'hbb922ea5),
	.w3(32'h399f6068),
	.w4(32'h3bafaaf2),
	.w5(32'h3a37f8bd),
	.w6(32'hbb9a6f12),
	.w7(32'h3b743d6d),
	.w8(32'h3acd3216),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c6b5),
	.w1(32'h3bbe1b22),
	.w2(32'hbb0c7f25),
	.w3(32'h3b06ba2f),
	.w4(32'h3bdcfbbf),
	.w5(32'h3acbd56c),
	.w6(32'hba281fda),
	.w7(32'hba73053b),
	.w8(32'hbaf14ad2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81470b),
	.w1(32'h3b0f6d87),
	.w2(32'hba8d4e78),
	.w3(32'h3aa32afc),
	.w4(32'hbae75696),
	.w5(32'hbb669642),
	.w6(32'hba99f338),
	.w7(32'h3b260cd3),
	.w8(32'h3ba16079),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17ecbf),
	.w1(32'hbba50d78),
	.w2(32'hb98b77c3),
	.w3(32'hba3739f7),
	.w4(32'hbaf20567),
	.w5(32'h3a4ed9ef),
	.w6(32'hbabe1f65),
	.w7(32'hbb07f069),
	.w8(32'hbb85c35c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b0881),
	.w1(32'hba78678f),
	.w2(32'h3b23131b),
	.w3(32'hbb28f191),
	.w4(32'hbb3bfccb),
	.w5(32'h3b49f55b),
	.w6(32'h3ba21ac2),
	.w7(32'h3a40a0a5),
	.w8(32'hbadbc9a1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dc788),
	.w1(32'hbb70d4a6),
	.w2(32'hbb4e5081),
	.w3(32'hbb676f23),
	.w4(32'hbabe2599),
	.w5(32'hbb9f3e11),
	.w6(32'hbb98d312),
	.w7(32'hbbd35793),
	.w8(32'hbb3d30cb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cee86),
	.w1(32'hbc1a6f7c),
	.w2(32'h3a575f19),
	.w3(32'hbb68381a),
	.w4(32'hbc19a128),
	.w5(32'hb8982ef1),
	.w6(32'hbb34512c),
	.w7(32'hbc0e297d),
	.w8(32'hbb4ff12c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab3f44),
	.w1(32'hbb7ee434),
	.w2(32'h3a16c613),
	.w3(32'hba0ef568),
	.w4(32'hbbf0a132),
	.w5(32'hbc0de50d),
	.w6(32'hbb2eb91e),
	.w7(32'hba93131e),
	.w8(32'hbaf51d8d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bab4b),
	.w1(32'h3ae5fe4c),
	.w2(32'hbac81cb9),
	.w3(32'hbbae0293),
	.w4(32'hbaa0df3d),
	.w5(32'h3971c636),
	.w6(32'hbb458f23),
	.w7(32'hbae6783d),
	.w8(32'h3a203bd7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ee6e),
	.w1(32'hbb4780af),
	.w2(32'hbadddec3),
	.w3(32'hbab7ad23),
	.w4(32'hbb0ab2b3),
	.w5(32'h3b4928fe),
	.w6(32'hbb6d829e),
	.w7(32'h3b21f94b),
	.w8(32'h3bd56f6b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab65e81),
	.w1(32'h3af45d6d),
	.w2(32'h3b3ae4c0),
	.w3(32'h3ace7994),
	.w4(32'hbb27d9c5),
	.w5(32'hbbbfe3d7),
	.w6(32'h3a957e39),
	.w7(32'hbb286c66),
	.w8(32'hbb718037),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3e7b7),
	.w1(32'hb8ebc4f7),
	.w2(32'h3b657e24),
	.w3(32'h398393c2),
	.w4(32'hbb82079a),
	.w5(32'hbac65349),
	.w6(32'h39b1262a),
	.w7(32'hba2985eb),
	.w8(32'h3b6d9290),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb781db),
	.w1(32'h3a9485e6),
	.w2(32'hbac6cc3f),
	.w3(32'h3b0978cf),
	.w4(32'hba9b2158),
	.w5(32'hbaf6fe2f),
	.w6(32'h3b7d6f20),
	.w7(32'h3b1e760c),
	.w8(32'h3b3b0bcd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b27ed),
	.w1(32'h38bdbed5),
	.w2(32'h3ae8c928),
	.w3(32'h399ebb1c),
	.w4(32'h3aa7812c),
	.w5(32'h3a787261),
	.w6(32'hbb148a1b),
	.w7(32'h3ad1136e),
	.w8(32'hbaa73718),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b311223),
	.w1(32'hbaa78d6e),
	.w2(32'hbafb2f55),
	.w3(32'h3822a0fe),
	.w4(32'hbb343618),
	.w5(32'hbacf14d5),
	.w6(32'hba55a522),
	.w7(32'h39f91856),
	.w8(32'h3af73a42),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73ebf8),
	.w1(32'h3bd4a8ac),
	.w2(32'h3a8c4047),
	.w3(32'h39fd0125),
	.w4(32'h3a3b5fe7),
	.w5(32'h3b6141d7),
	.w6(32'h3aa04e21),
	.w7(32'hba3f190f),
	.w8(32'hbae47434),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20c694),
	.w1(32'h3a8ebdad),
	.w2(32'h3b3252a9),
	.w3(32'h3b7f21e1),
	.w4(32'hbaa2b725),
	.w5(32'hbb3beebb),
	.w6(32'hbb429ed4),
	.w7(32'hbac032b6),
	.w8(32'hbb87043f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd748b),
	.w1(32'hba562bc1),
	.w2(32'hbb9a3369),
	.w3(32'hbabc6bdd),
	.w4(32'hbadac3b0),
	.w5(32'hbbe939e3),
	.w6(32'hbb02353c),
	.w7(32'hbb4629dd),
	.w8(32'hbaaf46f0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50700c),
	.w1(32'h3b95f9b1),
	.w2(32'h3bc7ee75),
	.w3(32'hbba10091),
	.w4(32'h3bd09156),
	.w5(32'h3bcbe173),
	.w6(32'hbbe06d45),
	.w7(32'hbbab2619),
	.w8(32'h3a9c751a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f55e5),
	.w1(32'hbb7c8d60),
	.w2(32'hba114e0d),
	.w3(32'hbb78a55f),
	.w4(32'hbb44d829),
	.w5(32'hbb41c977),
	.w6(32'hbb922e9d),
	.w7(32'hba47f4b8),
	.w8(32'hbb9c1fd8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12551e),
	.w1(32'h3a287461),
	.w2(32'h3a98a84f),
	.w3(32'hb913633e),
	.w4(32'hbaa1c5c3),
	.w5(32'h3b2c6219),
	.w6(32'hbb3a0f2b),
	.w7(32'hbb92f08a),
	.w8(32'h3b4d8940),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c172b),
	.w1(32'hba95717e),
	.w2(32'hba62f9aa),
	.w3(32'h3b036a5c),
	.w4(32'hbb5bd0e0),
	.w5(32'h3bb076ae),
	.w6(32'hba832326),
	.w7(32'h3b42ceaf),
	.w8(32'hbb815022),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a5a89),
	.w1(32'h3ad34f13),
	.w2(32'hbae94d89),
	.w3(32'hbada953e),
	.w4(32'h3b3c1a64),
	.w5(32'h3ba113ec),
	.w6(32'hbb8ccea9),
	.w7(32'hba2cfbc5),
	.w8(32'h3bba38d6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ff232),
	.w1(32'hbb823257),
	.w2(32'hbbbb9e0b),
	.w3(32'h3ba01dd6),
	.w4(32'hbb56b8e3),
	.w5(32'hbb9c8c93),
	.w6(32'hbb2641e0),
	.w7(32'hbaaaba49),
	.w8(32'hbbafb2ea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd57383),
	.w1(32'hb9748ae5),
	.w2(32'h39c97a09),
	.w3(32'hbba9e294),
	.w4(32'h3a8702fd),
	.w5(32'h3b8b99b1),
	.w6(32'hbc0a9fc3),
	.w7(32'h377e5ff0),
	.w8(32'h3b8c691d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269816),
	.w1(32'h3b3ff44a),
	.w2(32'hba37336e),
	.w3(32'h3b82067b),
	.w4(32'h3b87f0bc),
	.w5(32'hbab766e6),
	.w6(32'h3b963789),
	.w7(32'h3aadf3b7),
	.w8(32'h39803af8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44ee2),
	.w1(32'hbb6774f6),
	.w2(32'hb8aa79ef),
	.w3(32'h380b1a45),
	.w4(32'hbb76cba1),
	.w5(32'hbb236cdb),
	.w6(32'hbb2a1149),
	.w7(32'hbb1e973a),
	.w8(32'hbb9ec980),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb215e5c),
	.w1(32'h3ad444cb),
	.w2(32'hbb110a33),
	.w3(32'hbb5d1452),
	.w4(32'h3b142fcd),
	.w5(32'hbb401c8a),
	.w6(32'hbb611843),
	.w7(32'hb97a919c),
	.w8(32'h3abd7b0e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69bcfc),
	.w1(32'h3ada881e),
	.w2(32'h391c18f0),
	.w3(32'hba868aa6),
	.w4(32'h3b0152be),
	.w5(32'hbb1f4734),
	.w6(32'h3a63f9e2),
	.w7(32'h3a8d6f8f),
	.w8(32'hbaeae3e7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac87175),
	.w1(32'hb87e6aae),
	.w2(32'h386b094d),
	.w3(32'h3abea9e9),
	.w4(32'h3b9c4679),
	.w5(32'h3a948ff0),
	.w6(32'h3a1d9a22),
	.w7(32'h3b434eb9),
	.w8(32'hbabed63e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f4076),
	.w1(32'hbb1235b1),
	.w2(32'hbb9c54f7),
	.w3(32'hbb12a1a6),
	.w4(32'hbb917c12),
	.w5(32'hba907001),
	.w6(32'h3b6fb050),
	.w7(32'h39cf2a4f),
	.w8(32'hbb7aad8b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa43e6),
	.w1(32'hbb5b7f31),
	.w2(32'hbb97883f),
	.w3(32'hbb2f2004),
	.w4(32'hbbb7f0f5),
	.w5(32'h3b04fc72),
	.w6(32'hbb2e43a3),
	.w7(32'h3b87d6a7),
	.w8(32'h3baa13ac),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996d008),
	.w1(32'hbadc053f),
	.w2(32'hbb19b030),
	.w3(32'hba88f80f),
	.w4(32'hbb837eca),
	.w5(32'hbbbd4d81),
	.w6(32'h39d27214),
	.w7(32'hbb23e5eb),
	.w8(32'hbbb6d128),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8069),
	.w1(32'hbabd9ca4),
	.w2(32'hbb017677),
	.w3(32'hbb6f6372),
	.w4(32'hbb6405e0),
	.w5(32'hbbb854c1),
	.w6(32'hbba5ee08),
	.w7(32'hbb579625),
	.w8(32'hbc30a570),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac0d75),
	.w1(32'h3b8c1204),
	.w2(32'h3bf8d3d0),
	.w3(32'hb8a2ceaf),
	.w4(32'h3c0bf560),
	.w5(32'h3c4bac8f),
	.w6(32'hbb3efac4),
	.w7(32'h3b059724),
	.w8(32'h3bae6d0b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24c6a4),
	.w1(32'h3b220ab7),
	.w2(32'hbb8beffc),
	.w3(32'h3bdb8cfd),
	.w4(32'h3b0ad843),
	.w5(32'h3b86a533),
	.w6(32'hbbc20b0b),
	.w7(32'hbb34887b),
	.w8(32'hbb49e394),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule