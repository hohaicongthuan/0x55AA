module layer_8_featuremap_99(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccebc33),
	.w1(32'hbc52339f),
	.w2(32'hbd63464a),
	.w3(32'h3c94d272),
	.w4(32'h3b59691f),
	.w5(32'hbd1dfe98),
	.w6(32'hbc20b33e),
	.w7(32'hbca3728b),
	.w8(32'hbcd961a1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec3195),
	.w1(32'hbcb64676),
	.w2(32'hbc14ee05),
	.w3(32'h3be31406),
	.w4(32'h3c87232a),
	.w5(32'h3cdb157d),
	.w6(32'h3af5027f),
	.w7(32'h3c8fea8c),
	.w8(32'h3d142b1b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7613de),
	.w1(32'h3c0cc89d),
	.w2(32'hbb79647d),
	.w3(32'h3b9c7319),
	.w4(32'h3b9440fa),
	.w5(32'hbc281c9d),
	.w6(32'h3c8790bf),
	.w7(32'h3ce2e340),
	.w8(32'h3a8efb1a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd93fd0),
	.w1(32'h3cf76e8d),
	.w2(32'h3cec2e82),
	.w3(32'hbbb7b643),
	.w4(32'hbbb833f3),
	.w5(32'hbc4e7fc4),
	.w6(32'hbbd6cf79),
	.w7(32'hbc9ea20a),
	.w8(32'h3bf35f77),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d469d4b),
	.w1(32'h3c27c23a),
	.w2(32'h3d3a0d4b),
	.w3(32'hbc916af0),
	.w4(32'h3c773603),
	.w5(32'h3cd29935),
	.w6(32'h3bf9fda3),
	.w7(32'hbbb0e1b0),
	.w8(32'hbaeb0693),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5efb81),
	.w1(32'h3c6748ea),
	.w2(32'h3cdd307c),
	.w3(32'hbadb8158),
	.w4(32'h3c0591d0),
	.w5(32'h3d343dbc),
	.w6(32'hbc88ae7a),
	.w7(32'h3cd47086),
	.w8(32'h3d20dffe),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98e52d),
	.w1(32'hbbf0bbd4),
	.w2(32'h3b228f4d),
	.w3(32'hbc39e598),
	.w4(32'hbb43badd),
	.w5(32'h3bd22b1d),
	.w6(32'hba56d396),
	.w7(32'h3c09b57d),
	.w8(32'h3c709c3a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a771e),
	.w1(32'hbc29ce78),
	.w2(32'h3c0cc3c9),
	.w3(32'h3c46cb0c),
	.w4(32'hbc3ced22),
	.w5(32'hbc51c15d),
	.w6(32'h3cd230cd),
	.w7(32'h3ba339e7),
	.w8(32'hbc56626b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85e4c),
	.w1(32'hbc42338e),
	.w2(32'hb8f414fd),
	.w3(32'h3cac1a15),
	.w4(32'h3bdc41f9),
	.w5(32'h3c544124),
	.w6(32'h3b973e57),
	.w7(32'hbbafc266),
	.w8(32'h39ffce2f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a368acc),
	.w1(32'hbd074717),
	.w2(32'hbc028503),
	.w3(32'h3cbd92ea),
	.w4(32'hbc2f0319),
	.w5(32'hbd0a4fd1),
	.w6(32'h3bd21d38),
	.w7(32'hbbac2dc7),
	.w8(32'h3b1a0ab5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf17b94),
	.w1(32'hbcc4e7f3),
	.w2(32'hbb38a14d),
	.w3(32'h3af033b4),
	.w4(32'hbcad76cb),
	.w5(32'hbd24a696),
	.w6(32'h3c574549),
	.w7(32'hbc8ee90f),
	.w8(32'hbd079d3c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db4bd),
	.w1(32'hbb883870),
	.w2(32'hbc12aa30),
	.w3(32'hb860b95f),
	.w4(32'h3a25c8e5),
	.w5(32'hbc31f5bc),
	.w6(32'hbb76af86),
	.w7(32'h3c994478),
	.w8(32'h3aab9fbc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c344fa2),
	.w1(32'h3b3803fc),
	.w2(32'h3c58229f),
	.w3(32'h3b8f4de3),
	.w4(32'h3ba607b0),
	.w5(32'h3c952ad7),
	.w6(32'hbbb7dda0),
	.w7(32'h3c172353),
	.w8(32'h3ca7e38d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0426f),
	.w1(32'h3bbe2d02),
	.w2(32'h3b9df55b),
	.w3(32'h3b541a5c),
	.w4(32'h3b9ec268),
	.w5(32'h3b5a28a2),
	.w6(32'h3c0dcaf8),
	.w7(32'h3b7eaa08),
	.w8(32'hbb3d5ab9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68bf16),
	.w1(32'h3a0641bb),
	.w2(32'h3b8df40f),
	.w3(32'hbb954944),
	.w4(32'h3b8e9ccc),
	.w5(32'hba94edb5),
	.w6(32'hbbad26f7),
	.w7(32'h3b708b04),
	.w8(32'hbb8e73b0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf1dcc),
	.w1(32'h3a73c542),
	.w2(32'hbb749b61),
	.w3(32'hbaa81427),
	.w4(32'hbb8947d6),
	.w5(32'h3ba56b69),
	.w6(32'hbb6303ae),
	.w7(32'hbbd8de68),
	.w8(32'hbbecd1fc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb110633),
	.w1(32'hbc1433d2),
	.w2(32'hbbd76bf5),
	.w3(32'h3c808271),
	.w4(32'hbac5cc6f),
	.w5(32'hbb8512b9),
	.w6(32'h3bdfc1f4),
	.w7(32'h3bc78096),
	.w8(32'hbc92bb73),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d40cf),
	.w1(32'hbbfbcb5b),
	.w2(32'h3b365167),
	.w3(32'h3cd5d000),
	.w4(32'hbab9bc40),
	.w5(32'hbd00660b),
	.w6(32'h3c93ab9d),
	.w7(32'h3ca6445c),
	.w8(32'h3bd85472),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced31e9),
	.w1(32'h3b3e3d46),
	.w2(32'hbd587533),
	.w3(32'h3d4ef7c6),
	.w4(32'hbbedbc3b),
	.w5(32'hbdf78d20),
	.w6(32'h3d76d652),
	.w7(32'hbcc18c66),
	.w8(32'hbd98e72b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c057752),
	.w1(32'hbc72afdd),
	.w2(32'h3ca90520),
	.w3(32'h3a34327d),
	.w4(32'hbb0c7a11),
	.w5(32'h3bc85baa),
	.w6(32'hbcf459c7),
	.w7(32'h3c02fecb),
	.w8(32'h3cf3fa9c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36b8b8),
	.w1(32'hbab077a8),
	.w2(32'h3bbf5b1f),
	.w3(32'h3907a9b9),
	.w4(32'h3d086ed2),
	.w5(32'h3c726563),
	.w6(32'hbcc88e2a),
	.w7(32'h3b932cbc),
	.w8(32'h3c477fff),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea4413),
	.w1(32'h3b927597),
	.w2(32'h3c63b305),
	.w3(32'h3ba93b75),
	.w4(32'hbbd55b24),
	.w5(32'h3cc98247),
	.w6(32'h3c0a782a),
	.w7(32'hbc6f99b2),
	.w8(32'hbb1642b7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ad96a),
	.w1(32'hbcbdf00b),
	.w2(32'hbd84a921),
	.w3(32'h3d073d9d),
	.w4(32'hbc267bed),
	.w5(32'hbdf9efd1),
	.w6(32'h3d20471a),
	.w7(32'hbca30a24),
	.w8(32'hbda188e1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb95b),
	.w1(32'h3b991fb7),
	.w2(32'h3c167148),
	.w3(32'hbd1d0762),
	.w4(32'h3b956020),
	.w5(32'h3bab4047),
	.w6(32'hbcfe36a5),
	.w7(32'h3ba73d98),
	.w8(32'hbadd6793),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd93ee0),
	.w1(32'hbbecb2c7),
	.w2(32'hbb4c8ff6),
	.w3(32'hbb87fc58),
	.w4(32'hbb9139f0),
	.w5(32'h3bbeaa65),
	.w6(32'hbb8585f2),
	.w7(32'hbb4fc026),
	.w8(32'h3b71ddec),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4333d2),
	.w1(32'h39d98344),
	.w2(32'h3ba5d143),
	.w3(32'h3c74245e),
	.w4(32'h3ce1bfed),
	.w5(32'h3a8decee),
	.w6(32'h3c3fd74e),
	.w7(32'h3bfdf835),
	.w8(32'hbc34d1af),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd72db),
	.w1(32'hbbe2caa4),
	.w2(32'hbb7291fb),
	.w3(32'h3bddf0a5),
	.w4(32'hbc819408),
	.w5(32'hbc8e6825),
	.w6(32'hbc80788e),
	.w7(32'hbc29900b),
	.w8(32'hb99c9fa2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb14c08),
	.w1(32'hbd24c8a4),
	.w2(32'h3cd3ec41),
	.w3(32'h3e071621),
	.w4(32'h3d1b7b83),
	.w5(32'hbe262b99),
	.w6(32'h3e7fb6f5),
	.w7(32'h3d4dfb94),
	.w8(32'hbe3ffc77),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2df2e9),
	.w1(32'hbc92a927),
	.w2(32'hbb49ea57),
	.w3(32'h3b99ed76),
	.w4(32'hbbf27964),
	.w5(32'hbc1aee23),
	.w6(32'hb904ad56),
	.w7(32'h3b7883d6),
	.w8(32'hbc27b2c9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f5e6),
	.w1(32'hbbfd8979),
	.w2(32'h3b352e68),
	.w3(32'hbbff2fb3),
	.w4(32'h3bd45f72),
	.w5(32'h3b044ca6),
	.w6(32'h3cc00c9b),
	.w7(32'h3b52c511),
	.w8(32'h3bc30ac1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaf799),
	.w1(32'hbb3666d2),
	.w2(32'hbb39d2ca),
	.w3(32'h3c1bd806),
	.w4(32'hb9c811c0),
	.w5(32'hbbf8e527),
	.w6(32'hbc834925),
	.w7(32'hbb55b09e),
	.w8(32'hbc26f0ed),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b022f4f),
	.w1(32'h3bfc2a10),
	.w2(32'h3bc8fb01),
	.w3(32'hbc1f329a),
	.w4(32'hb944e660),
	.w5(32'h3cfe03e8),
	.w6(32'hbbf465fd),
	.w7(32'hbc12dedd),
	.w8(32'hbc22f282),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63a1b4),
	.w1(32'hbbf7a3eb),
	.w2(32'hbc76f425),
	.w3(32'h3cacbfd7),
	.w4(32'hbc441432),
	.w5(32'hbc0953ab),
	.w6(32'h3c581e32),
	.w7(32'hbc667a22),
	.w8(32'h3b3b9c49),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7df49d),
	.w1(32'h3c5c9763),
	.w2(32'hbace27fe),
	.w3(32'h3c5efae2),
	.w4(32'h3b566385),
	.w5(32'hbc35e149),
	.w6(32'h3c5cc8be),
	.w7(32'hbb85beba),
	.w8(32'hbc47aacc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66c910),
	.w1(32'hbb7da648),
	.w2(32'h3b8e6aeb),
	.w3(32'h3bb9bfa1),
	.w4(32'h3c674731),
	.w5(32'h3ceaf1f7),
	.w6(32'hbc4f9d79),
	.w7(32'hbaaee26f),
	.w8(32'h3cd646fb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bc1ba),
	.w1(32'h3bf9b576),
	.w2(32'h3bb9806b),
	.w3(32'h3cd134dc),
	.w4(32'h3c831d63),
	.w5(32'hbcd05cfb),
	.w6(32'h3d0335b8),
	.w7(32'h3cd32796),
	.w8(32'h3bcf250f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc56c7f),
	.w1(32'h3c064dd0),
	.w2(32'h3b3e700b),
	.w3(32'hbd34e098),
	.w4(32'hbca504dc),
	.w5(32'hbb39f7e0),
	.w6(32'hbc8c74bd),
	.w7(32'hbc9ff381),
	.w8(32'hbc8b0ed2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68df9a),
	.w1(32'h3b8ba2c2),
	.w2(32'hbbefe1fa),
	.w3(32'h3c95347a),
	.w4(32'hbaca0016),
	.w5(32'hbb447723),
	.w6(32'h3cd33610),
	.w7(32'hbb5c438c),
	.w8(32'hba12e51e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ae60e),
	.w1(32'hbaec7854),
	.w2(32'hbc75b22a),
	.w3(32'h3bb16e65),
	.w4(32'hbc8023d6),
	.w5(32'h3bcdbd01),
	.w6(32'hbb27936a),
	.w7(32'hbc9a4a62),
	.w8(32'hbcab968a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7be865),
	.w1(32'hbbeb5ea8),
	.w2(32'hbc84fcd4),
	.w3(32'h3cb0bd21),
	.w4(32'h3bba6c37),
	.w5(32'h3bf8c59b),
	.w6(32'h3cb4aa68),
	.w7(32'h3b9a77ec),
	.w8(32'h3b814682),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42649e),
	.w1(32'hbb82c8f4),
	.w2(32'h3ce77d4d),
	.w3(32'h3d7cdc7d),
	.w4(32'h3ca3282c),
	.w5(32'h3bfdbc79),
	.w6(32'h3cc0b543),
	.w7(32'h39e4e1a3),
	.w8(32'h3cdf2e10),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5c70),
	.w1(32'h3ae2ac3d),
	.w2(32'h3c6a3c93),
	.w3(32'h3b0a766b),
	.w4(32'h3c9ded11),
	.w5(32'hbcabf010),
	.w6(32'h3adcf9c8),
	.w7(32'h3c41b2b4),
	.w8(32'h3cb1651a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5ba22),
	.w1(32'h3c0ed717),
	.w2(32'h3c195f2e),
	.w3(32'hbd163ea2),
	.w4(32'h3ab5ca00),
	.w5(32'hbb125b67),
	.w6(32'hbcdd86f0),
	.w7(32'hbbdfad15),
	.w8(32'hbbd98ba0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab19d2),
	.w1(32'h3c309240),
	.w2(32'hbac09762),
	.w3(32'h3c42368c),
	.w4(32'h3b7a0030),
	.w5(32'hbc6fe6be),
	.w6(32'h3b261431),
	.w7(32'hbb4a210f),
	.w8(32'hbc8723ea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98af0b),
	.w1(32'hba2cfb12),
	.w2(32'hbc4fc730),
	.w3(32'h3c0490de),
	.w4(32'hbc88fea6),
	.w5(32'hbd016240),
	.w6(32'h3ca8508c),
	.w7(32'hbcef3d21),
	.w8(32'hbd6f764d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd82c8),
	.w1(32'hbb38480d),
	.w2(32'hbc040bf2),
	.w3(32'h3b8b0efc),
	.w4(32'h3a12afbb),
	.w5(32'hbcce1f8b),
	.w6(32'h3caf08e4),
	.w7(32'hbc566e44),
	.w8(32'hbbde6493),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbb27e),
	.w1(32'h3c7d2fdf),
	.w2(32'hbbe4d4aa),
	.w3(32'hbc063ab0),
	.w4(32'hbc0e5234),
	.w5(32'h3bb806e3),
	.w6(32'h3bb85934),
	.w7(32'hbc3e6e7c),
	.w8(32'hbc23ef93),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b497feb),
	.w1(32'hbcaae5e9),
	.w2(32'hbcc1e077),
	.w3(32'h3c9459e2),
	.w4(32'hbcccbb7b),
	.w5(32'hbd2bacab),
	.w6(32'h3c4105f3),
	.w7(32'hbd026dde),
	.w8(32'hbd8cd64a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9ab4e),
	.w1(32'h3b4fd46a),
	.w2(32'hbc1b81f9),
	.w3(32'h3bbf50b7),
	.w4(32'hbc12cbf8),
	.w5(32'hbb37601e),
	.w6(32'h3cb6b96e),
	.w7(32'hbc5b8083),
	.w8(32'h3bef79be),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146bb1),
	.w1(32'h3c424189),
	.w2(32'hbcf3214e),
	.w3(32'h3cd151b7),
	.w4(32'hbc977ef8),
	.w5(32'hbcadf9e1),
	.w6(32'h3c748d88),
	.w7(32'hbcbb6718),
	.w8(32'hbccc823c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdf513),
	.w1(32'h3c24ccf4),
	.w2(32'h3cdd17ca),
	.w3(32'h3c019738),
	.w4(32'h3ceee679),
	.w5(32'h3d745b42),
	.w6(32'h3b85d6a3),
	.w7(32'h3c789f1a),
	.w8(32'h3da0c24b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae78f8),
	.w1(32'hbb82056e),
	.w2(32'hbbbb8138),
	.w3(32'h3cb51486),
	.w4(32'hbb992ef7),
	.w5(32'hbd10253b),
	.w6(32'h3d3e4473),
	.w7(32'hbd4f2ec8),
	.w8(32'hbd624c0d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd58d1c),
	.w1(32'h3aeaa5f3),
	.w2(32'h3bdfbf19),
	.w3(32'h3d2140e9),
	.w4(32'h3b54663c),
	.w5(32'hbc3ae38e),
	.w6(32'h3c9f6d00),
	.w7(32'h3c3224bd),
	.w8(32'h3bd2012e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc230341),
	.w1(32'hbc2c80d1),
	.w2(32'hbc9b4401),
	.w3(32'h3caa2c3b),
	.w4(32'h3c6335a5),
	.w5(32'hbcf274ba),
	.w6(32'hbbddb46f),
	.w7(32'hbbeeef36),
	.w8(32'hbc44c416),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcc0f0),
	.w1(32'h3a2aca62),
	.w2(32'hbbd1793d),
	.w3(32'hbba59820),
	.w4(32'h3b5709d7),
	.w5(32'h3c3bf1db),
	.w6(32'hb9d7212a),
	.w7(32'hba1f1138),
	.w8(32'hbc4007a9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2daffe),
	.w1(32'h3c8725cb),
	.w2(32'hbcf907ec),
	.w3(32'h3d60e32b),
	.w4(32'h3ca5d3fa),
	.w5(32'hbd283c7e),
	.w6(32'h3cb57def),
	.w7(32'h3afbbbb4),
	.w8(32'hbd3d3c18),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca28aaf),
	.w1(32'hbb8b9390),
	.w2(32'hbc544988),
	.w3(32'h3c8075d8),
	.w4(32'h3b368d89),
	.w5(32'hbc407a1e),
	.w6(32'h3c39ca0f),
	.w7(32'h3b8e224f),
	.w8(32'hb9db71aa),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb200772),
	.w1(32'hbad4f83d),
	.w2(32'h3c19cc04),
	.w3(32'h3cc6d0dd),
	.w4(32'h3c0fa918),
	.w5(32'hbcf91068),
	.w6(32'h3d140547),
	.w7(32'h3c094a15),
	.w8(32'hbc05b4f7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bfcc6),
	.w1(32'h3b3415bb),
	.w2(32'hbc5692e5),
	.w3(32'hbcef682b),
	.w4(32'h3c01909e),
	.w5(32'hbca81d3e),
	.w6(32'hbc62b520),
	.w7(32'h3b60fb66),
	.w8(32'hbcca42c1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89e9cb),
	.w1(32'h3a257c53),
	.w2(32'hbb9655c0),
	.w3(32'hbc09d5e6),
	.w4(32'hbad796d7),
	.w5(32'hbc13eed9),
	.w6(32'hbb85dd4b),
	.w7(32'hbbd05921),
	.w8(32'hbc6b70eb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a419),
	.w1(32'h3af11a58),
	.w2(32'h3c505558),
	.w3(32'h3c6fb1b0),
	.w4(32'hbb56f7b7),
	.w5(32'hbc645bf5),
	.w6(32'h3bada9df),
	.w7(32'h3b925ee7),
	.w8(32'h3c913c54),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91510a),
	.w1(32'h3cdd42e3),
	.w2(32'h3b80e164),
	.w3(32'hbd3e3308),
	.w4(32'hbc21d74f),
	.w5(32'hbcd396a5),
	.w6(32'hbc9f373c),
	.w7(32'hba58173d),
	.w8(32'hbc998397),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b95d6),
	.w1(32'hbca7be6c),
	.w2(32'h3c647ede),
	.w3(32'h3c0432b1),
	.w4(32'h3c43798d),
	.w5(32'hbc944795),
	.w6(32'hbcb2e195),
	.w7(32'h3ca56c9f),
	.w8(32'h3b734705),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1327d),
	.w1(32'hbb2c1a85),
	.w2(32'hbbd4f878),
	.w3(32'h3c9e2272),
	.w4(32'hbba796b4),
	.w5(32'h3be9f002),
	.w6(32'hbbae12b6),
	.w7(32'hbb7e1087),
	.w8(32'hbbde76c8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4d98),
	.w1(32'h3bb59ed8),
	.w2(32'h3b1035b7),
	.w3(32'h3c77e82f),
	.w4(32'h3b035781),
	.w5(32'h3b741406),
	.w6(32'h3c4a0743),
	.w7(32'h3c4846ce),
	.w8(32'h3c6d0a1f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcb82c),
	.w1(32'hbaed00db),
	.w2(32'hbacdcfec),
	.w3(32'h3c397771),
	.w4(32'h3c09f319),
	.w5(32'hba42e6f6),
	.w6(32'h3c8f226f),
	.w7(32'h3bd25989),
	.w8(32'h3c0d628c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56626a),
	.w1(32'hbb81628c),
	.w2(32'h3ce5629f),
	.w3(32'hbc6eaa38),
	.w4(32'h3a7b4bac),
	.w5(32'h3c766af8),
	.w6(32'hbc7711de),
	.w7(32'h3c01ef9f),
	.w8(32'h3c875764),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c838b67),
	.w1(32'hbb6079d5),
	.w2(32'hbc24dc15),
	.w3(32'h3ce06bd7),
	.w4(32'h3c276b75),
	.w5(32'hbbaa8726),
	.w6(32'hbb79a247),
	.w7(32'hbb14ba1e),
	.w8(32'h3c77a158),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7c654),
	.w1(32'hbbd4bf80),
	.w2(32'hbc39f8d9),
	.w3(32'hb966d161),
	.w4(32'hbb4c83ef),
	.w5(32'h3b88a827),
	.w6(32'hbc9362e4),
	.w7(32'hbc61d604),
	.w8(32'hbc8a612f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf3eae9),
	.w1(32'h3bb4ced3),
	.w2(32'hbbb1d3ef),
	.w3(32'h3ba7672a),
	.w4(32'h3c9c5538),
	.w5(32'hbdac90ea),
	.w6(32'h3d329574),
	.w7(32'hbc878397),
	.w8(32'hbda3fe69),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32222c),
	.w1(32'h3b8e7320),
	.w2(32'h3bf13175),
	.w3(32'h3b169294),
	.w4(32'hbb8cf29c),
	.w5(32'hbc5ac33a),
	.w6(32'hbb3ed951),
	.w7(32'h3c79d9f4),
	.w8(32'h3c782282),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b699c80),
	.w1(32'h3a4584a4),
	.w2(32'hbb473e33),
	.w3(32'hbc86a44a),
	.w4(32'hbc026a78),
	.w5(32'h3c01ab86),
	.w6(32'hbc95879e),
	.w7(32'hbc10bb5c),
	.w8(32'hbc0ff66b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73f034),
	.w1(32'h3cd72355),
	.w2(32'hb9da8d34),
	.w3(32'h3ceec49a),
	.w4(32'h3bfd9d22),
	.w5(32'h3b3e6df9),
	.w6(32'h3d21f8c6),
	.w7(32'h3c0a0e2a),
	.w8(32'h3b7c5ffd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be09154),
	.w1(32'h3b2c3423),
	.w2(32'hbc108235),
	.w3(32'h3c71d844),
	.w4(32'h3c370726),
	.w5(32'h38d22c90),
	.w6(32'h3c24f5a3),
	.w7(32'h3ce4dbdc),
	.w8(32'h3cea64ec),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40f69d),
	.w1(32'hbb01fe31),
	.w2(32'hbc06d910),
	.w3(32'h3b55ce08),
	.w4(32'hbcad5c38),
	.w5(32'hbca6b75d),
	.w6(32'hbb2fdaaa),
	.w7(32'hbc5f2cb2),
	.w8(32'hbcee0e29),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29c2d),
	.w1(32'hbcba4dc9),
	.w2(32'hbc4da465),
	.w3(32'h3d1b7062),
	.w4(32'h3b1191d4),
	.w5(32'hbbadec9a),
	.w6(32'hbc14dcbb),
	.w7(32'hbb9246c9),
	.w8(32'hbca4c172),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bbd63),
	.w1(32'h3c056d9a),
	.w2(32'h3b58debd),
	.w3(32'h3bb7b85f),
	.w4(32'hba034a94),
	.w5(32'h3bffa6e8),
	.w6(32'h3c2b8d53),
	.w7(32'h3b456526),
	.w8(32'h3ca22a59),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ab2f7),
	.w1(32'hbbaab913),
	.w2(32'hbb5637a8),
	.w3(32'h3c921fdb),
	.w4(32'hba8c600a),
	.w5(32'hbc5abafc),
	.w6(32'h3ccb58a5),
	.w7(32'h3b995434),
	.w8(32'h3c530f8a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfbccf8),
	.w1(32'h3c4bc95a),
	.w2(32'hbbe41ab5),
	.w3(32'h3cb196de),
	.w4(32'h3bbf8b0b),
	.w5(32'hbb6b2be0),
	.w6(32'h3d1fa5cd),
	.w7(32'h3bdedb2d),
	.w8(32'h3c4c4a2d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c733426),
	.w1(32'h3c12d145),
	.w2(32'hbbcaed6c),
	.w3(32'h3bbe0c72),
	.w4(32'hbb88d473),
	.w5(32'h3aa3ab9b),
	.w6(32'h3c9711b7),
	.w7(32'hbb9d92e0),
	.w8(32'hbb05b505),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5f2ea),
	.w1(32'hbb536d76),
	.w2(32'hbc25413a),
	.w3(32'h3a8a6538),
	.w4(32'hbad59eb9),
	.w5(32'h3a692b7d),
	.w6(32'hba729618),
	.w7(32'hbb92429b),
	.w8(32'h3b403560),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf6988),
	.w1(32'hbc3e3871),
	.w2(32'h3a98336b),
	.w3(32'hba8196fc),
	.w4(32'h3b6f9388),
	.w5(32'hbac855ea),
	.w6(32'h3c8f5e8b),
	.w7(32'h3bcdc38a),
	.w8(32'hbc9764a7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16a93b),
	.w1(32'hbb2b7197),
	.w2(32'h3b62aaf0),
	.w3(32'h3c705e96),
	.w4(32'h3bb2b2e6),
	.w5(32'hbb5ada22),
	.w6(32'h3bf800cc),
	.w7(32'h3b6fdce1),
	.w8(32'h3bbd9758),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dbdb9),
	.w1(32'h3cc690ab),
	.w2(32'h3cf48dc9),
	.w3(32'h3d47c84e),
	.w4(32'h3c23fd86),
	.w5(32'h3d0b97c0),
	.w6(32'hbac4bca6),
	.w7(32'hbc027de1),
	.w8(32'h3d983976),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1b618),
	.w1(32'hbbe20b19),
	.w2(32'hbb4bbd3e),
	.w3(32'h3d009c46),
	.w4(32'h3c8d1e46),
	.w5(32'hbd29f088),
	.w6(32'h3d42418e),
	.w7(32'hbc59a217),
	.w8(32'hbd0b18c4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc478802),
	.w1(32'hbc9d5753),
	.w2(32'hbb80c469),
	.w3(32'h3c96ac73),
	.w4(32'h3b829931),
	.w5(32'hbb9c4ca8),
	.w6(32'h3ad30548),
	.w7(32'h3bf7327f),
	.w8(32'h3a7d736b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c711b98),
	.w1(32'h3b67a52e),
	.w2(32'hb9e2436f),
	.w3(32'h3aacc592),
	.w4(32'h3b5ab845),
	.w5(32'hbb27af4c),
	.w6(32'hba1a5d10),
	.w7(32'h3af08d31),
	.w8(32'h39e18784),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba956ffb),
	.w1(32'h3a922f02),
	.w2(32'hbb34e54e),
	.w3(32'hbad0ca09),
	.w4(32'h39b18cd9),
	.w5(32'hbbeee7c0),
	.w6(32'hb6af9f40),
	.w7(32'h3a5eb9c3),
	.w8(32'hbbb85e59),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc523a3a),
	.w1(32'hbbe2b957),
	.w2(32'hbba6f35f),
	.w3(32'hbb82c2c1),
	.w4(32'h3b045749),
	.w5(32'h3b408872),
	.w6(32'h3aa00c4d),
	.w7(32'hb9aa487b),
	.w8(32'hbb81b37d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54b29b),
	.w1(32'hba8caa67),
	.w2(32'h3b052b31),
	.w3(32'h3b8811fd),
	.w4(32'h3c5cbefc),
	.w5(32'hbbb09599),
	.w6(32'hba849bc3),
	.w7(32'h3c7bf473),
	.w8(32'h3a9f8bbf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31741e),
	.w1(32'hbc35dae4),
	.w2(32'h3c3345f0),
	.w3(32'hb89bdf7d),
	.w4(32'h3c2b7101),
	.w5(32'h3bac4c77),
	.w6(32'hbc7a2a81),
	.w7(32'h3bc03f31),
	.w8(32'hba539a0f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83cc4bf),
	.w1(32'h3a9eb62c),
	.w2(32'h3abab9c2),
	.w3(32'h3b85c1ef),
	.w4(32'hbbbb838d),
	.w5(32'hbc04e215),
	.w6(32'hbb875157),
	.w7(32'hbb5179d8),
	.w8(32'h3af7a90b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404195),
	.w1(32'hbc019ef6),
	.w2(32'h3c482511),
	.w3(32'hbc0a6034),
	.w4(32'hbb9ce7a2),
	.w5(32'h3b944ee7),
	.w6(32'hbc5a6090),
	.w7(32'hbbd43f79),
	.w8(32'hb90a912e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc83caf),
	.w1(32'hbc3bb486),
	.w2(32'h3bae1c55),
	.w3(32'h3ad4c705),
	.w4(32'h3b65f637),
	.w5(32'hbbdf04c1),
	.w6(32'hbbab8ac6),
	.w7(32'hba08610b),
	.w8(32'hbb638d3c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bbb5a),
	.w1(32'h3c4e18e8),
	.w2(32'h3c85508e),
	.w3(32'h3cb1f38a),
	.w4(32'h3c239e5f),
	.w5(32'h3d070d2f),
	.w6(32'h3c532176),
	.w7(32'h3ce54586),
	.w8(32'h3d6e88e1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdabb9e),
	.w1(32'h3beb5a58),
	.w2(32'hbc19a6c1),
	.w3(32'h3c919a3c),
	.w4(32'h3c24b41b),
	.w5(32'hbc78f012),
	.w6(32'h3d13f62d),
	.w7(32'hbc32f8aa),
	.w8(32'hbcd22657),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0116e),
	.w1(32'hbbdde2e8),
	.w2(32'h3b8f2c10),
	.w3(32'h3cc440e9),
	.w4(32'h3c319ede),
	.w5(32'h3c725334),
	.w6(32'h3bee61b1),
	.w7(32'h3c33c0fe),
	.w8(32'h3c4f254a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cc026),
	.w1(32'h3bb01500),
	.w2(32'hba203a78),
	.w3(32'h3b4f2961),
	.w4(32'hbb70eccb),
	.w5(32'hbb711332),
	.w6(32'h3b0e0d6e),
	.w7(32'hbae2ea9b),
	.w8(32'h3a22cbde),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac575fa),
	.w1(32'hbb9ffb5c),
	.w2(32'hbb8b60d0),
	.w3(32'hbb930d24),
	.w4(32'hba7bf4d6),
	.w5(32'hbbf9ef22),
	.w6(32'hbb10d163),
	.w7(32'hbb2310a7),
	.w8(32'hbc0c8b1f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f9bd),
	.w1(32'hbb90a566),
	.w2(32'h3bade342),
	.w3(32'hbbbf1aaa),
	.w4(32'h3c09f712),
	.w5(32'hba0f2c3d),
	.w6(32'hbbcec22b),
	.w7(32'h3be50f61),
	.w8(32'hb9803464),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7469fd),
	.w1(32'h3b613615),
	.w2(32'hbb39ef7c),
	.w3(32'hb8acfc70),
	.w4(32'h3b925df2),
	.w5(32'h3c46bd86),
	.w6(32'hbc06f8ab),
	.w7(32'hbbb27b5e),
	.w8(32'hba3097e2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081ea6),
	.w1(32'h3b247c62),
	.w2(32'h3c2feeb8),
	.w3(32'h3bd0d555),
	.w4(32'h3c585693),
	.w5(32'hbbe60bbd),
	.w6(32'hbac2f9c7),
	.w7(32'h3c8d9f30),
	.w8(32'hbbb9a870),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc248d6f),
	.w1(32'hbb5d12c2),
	.w2(32'h3b0d9783),
	.w3(32'hbb4c8497),
	.w4(32'h3b7cf522),
	.w5(32'hbb80188f),
	.w6(32'hbba11811),
	.w7(32'h3ba0896d),
	.w8(32'h3b4c919d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba769fa),
	.w1(32'hbc6bb60d),
	.w2(32'h3c53c532),
	.w3(32'hbc827b65),
	.w4(32'hbb7d3d9f),
	.w5(32'h3c0c367c),
	.w6(32'hbbc65826),
	.w7(32'h3a324765),
	.w8(32'hbaa41959),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3826bd),
	.w1(32'hbb9547fa),
	.w2(32'h3bbdbec3),
	.w3(32'hbb8624a8),
	.w4(32'h3ac0b7e3),
	.w5(32'h3c30b211),
	.w6(32'hbc23b032),
	.w7(32'h3bad3eac),
	.w8(32'h3c87248a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592b7e),
	.w1(32'h39b1ea52),
	.w2(32'hbbb78bcf),
	.w3(32'h3c17c7de),
	.w4(32'h3c993dfc),
	.w5(32'hbd2aa256),
	.w6(32'h3cd6afb1),
	.w7(32'h3b5b4bdd),
	.w8(32'hbd60340b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2b84),
	.w1(32'hbb2bdd94),
	.w2(32'h3b7a45d3),
	.w3(32'h3b214ad2),
	.w4(32'h3b1b04bc),
	.w5(32'hbb9e909a),
	.w6(32'hba9a0605),
	.w7(32'h3c2c9d47),
	.w8(32'h3bb0d8ff),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813f7ce),
	.w1(32'h3bfaba56),
	.w2(32'h3c5df667),
	.w3(32'hbbfcf2e7),
	.w4(32'hb86f6771),
	.w5(32'h3caf4746),
	.w6(32'hbb23c570),
	.w7(32'h3c04add2),
	.w8(32'h3d308f16),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d0de),
	.w1(32'h3baf6c4a),
	.w2(32'h3bad91dd),
	.w3(32'h3a635767),
	.w4(32'h3b65792e),
	.w5(32'hb9ef0028),
	.w6(32'h3c04fcfd),
	.w7(32'h3babdb44),
	.w8(32'hba6be9a5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc997c),
	.w1(32'hba4d8d64),
	.w2(32'h3a05fe17),
	.w3(32'h3c87b631),
	.w4(32'h3c38c304),
	.w5(32'hbb28de62),
	.w6(32'h3c367585),
	.w7(32'h3bdb1d18),
	.w8(32'h3b2b556c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc202ba),
	.w1(32'h3b989269),
	.w2(32'h3bfdf665),
	.w3(32'h3c855ddc),
	.w4(32'h3c13c4f2),
	.w5(32'h3c0ce70c),
	.w6(32'h39a3395f),
	.w7(32'h3ba68be3),
	.w8(32'h3caa5ea9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1be62f),
	.w1(32'hbb4d957a),
	.w2(32'h3c9fa5c6),
	.w3(32'h3b3b3c9e),
	.w4(32'h3ab69472),
	.w5(32'h3c613a56),
	.w6(32'h396e8bd8),
	.w7(32'h3c0e46fd),
	.w8(32'h3cb2efde),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176691),
	.w1(32'hbb0d9b96),
	.w2(32'hbac4ac4e),
	.w3(32'hbbfb97f2),
	.w4(32'hbaec8398),
	.w5(32'hb9eedf71),
	.w6(32'hbbe096b9),
	.w7(32'hbbe479ef),
	.w8(32'hbafee300),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01861c),
	.w1(32'hbbd19c18),
	.w2(32'h3b707fca),
	.w3(32'hb90f9790),
	.w4(32'h3c4061e0),
	.w5(32'h3b3c760e),
	.w6(32'hbc1752d3),
	.w7(32'h3bf381c9),
	.w8(32'hbb2f89b1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8b09),
	.w1(32'hbc271650),
	.w2(32'h3b014864),
	.w3(32'h3b960b05),
	.w4(32'h3c1c2c52),
	.w5(32'hbb43f155),
	.w6(32'hbbbdbff8),
	.w7(32'h3c182ce2),
	.w8(32'hbb387960),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130014),
	.w1(32'hbaccd331),
	.w2(32'hbb00cdc4),
	.w3(32'h3a140193),
	.w4(32'hbc29e667),
	.w5(32'h3aa18b5c),
	.w6(32'h3b1f329c),
	.w7(32'hbc39cbed),
	.w8(32'h3b13a585),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf2035),
	.w1(32'hbac02873),
	.w2(32'h3a91f9da),
	.w3(32'h3b6c44ba),
	.w4(32'h39b78cf9),
	.w5(32'hbb7027ac),
	.w6(32'h3bca795c),
	.w7(32'hba7dd65b),
	.w8(32'hbbf25708),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f089),
	.w1(32'h3ad0cd9b),
	.w2(32'h3c77c32e),
	.w3(32'h3c1d0c38),
	.w4(32'h3c02747c),
	.w5(32'h3c174f9b),
	.w6(32'h3c1b591c),
	.w7(32'h3c36091d),
	.w8(32'h3cd2675b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5da2a1),
	.w1(32'h3ba26d94),
	.w2(32'h3b5b974b),
	.w3(32'h3b2ebaf4),
	.w4(32'hbb209002),
	.w5(32'hbb816e45),
	.w6(32'h3c547f31),
	.w7(32'hbb7a6031),
	.w8(32'hbc2e08fe),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13f308),
	.w1(32'hbb17c9ef),
	.w2(32'h3adad94a),
	.w3(32'hbab50004),
	.w4(32'h3be0e333),
	.w5(32'hbc3240be),
	.w6(32'hbbe581ba),
	.w7(32'h3b9b3820),
	.w8(32'hbc3022b4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb37633),
	.w1(32'hbc98565d),
	.w2(32'hbbc6daf7),
	.w3(32'h3c4667d1),
	.w4(32'h3a17c15e),
	.w5(32'hbc45958e),
	.w6(32'hbc5a46d8),
	.w7(32'hbc09e28a),
	.w8(32'hbc27bb7f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaedbd),
	.w1(32'hbae1ec0a),
	.w2(32'h3bcfe856),
	.w3(32'h3cc33824),
	.w4(32'h3b0616a5),
	.w5(32'hbbabd4c6),
	.w6(32'h3c82b052),
	.w7(32'hb9f133f0),
	.w8(32'h3abcb5e4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c102f12),
	.w1(32'h3b01f225),
	.w2(32'h3bed2fdc),
	.w3(32'h3ba37419),
	.w4(32'hba3e9df8),
	.w5(32'h3c5c97ae),
	.w6(32'h3aa5c8ac),
	.w7(32'h3c3d9b0c),
	.w8(32'h3d1cd985),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1434ad),
	.w1(32'h3b3d8e0a),
	.w2(32'h3a773130),
	.w3(32'hb97a2eea),
	.w4(32'h39458b76),
	.w5(32'hbc81f829),
	.w6(32'h3c520a6b),
	.w7(32'hbb19373d),
	.w8(32'hbca15bdf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d86ec),
	.w1(32'hbb4844f3),
	.w2(32'h3b41b95f),
	.w3(32'hba395a56),
	.w4(32'hbbb1552d),
	.w5(32'h3c237a89),
	.w6(32'hbc29c5f4),
	.w7(32'h3b8a2de2),
	.w8(32'h3cd87b15),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ce9fa),
	.w1(32'h3c5ddc96),
	.w2(32'h3bcadbb8),
	.w3(32'h3afa83c9),
	.w4(32'h3cbbcd64),
	.w5(32'h3c24f119),
	.w6(32'h3c119750),
	.w7(32'h3bcc6b15),
	.w8(32'hbb109e00),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c503820),
	.w1(32'hbb23b0a5),
	.w2(32'h3bb6125c),
	.w3(32'h3c7cfdb8),
	.w4(32'h3bf30b36),
	.w5(32'h3c068d01),
	.w6(32'h3be4c47c),
	.w7(32'h3cb1cb89),
	.w8(32'h3c9f8eeb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40907a),
	.w1(32'h3ba186c1),
	.w2(32'h3b5ae13a),
	.w3(32'h3b82a35c),
	.w4(32'h3c0555a5),
	.w5(32'hbce20a62),
	.w6(32'h3c17ea08),
	.w7(32'h3b923737),
	.w8(32'hbc9e5e77),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule