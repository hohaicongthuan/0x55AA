module layer_10_featuremap_407(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026cbb),
	.w1(32'hba8918b3),
	.w2(32'hba04bd39),
	.w3(32'h3a3169c9),
	.w4(32'hbb2f57f1),
	.w5(32'hbabc83f0),
	.w6(32'hbb1233b2),
	.w7(32'hba9bac60),
	.w8(32'h38888cda),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb531c7d),
	.w1(32'hbb811c62),
	.w2(32'hbc57ebed),
	.w3(32'h392de5dc),
	.w4(32'h3a408d87),
	.w5(32'hbb6b106f),
	.w6(32'hbbb94adc),
	.w7(32'hbb2c0718),
	.w8(32'hbba4f308),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82907b),
	.w1(32'hbb48a932),
	.w2(32'hbc041b5c),
	.w3(32'h3b61e6e8),
	.w4(32'hba5893c3),
	.w5(32'h3b8fe99f),
	.w6(32'h3a2f38d9),
	.w7(32'hbb17c9e2),
	.w8(32'hba976326),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955584),
	.w1(32'h3aaa4fc4),
	.w2(32'h3bda3941),
	.w3(32'hbac30a34),
	.w4(32'hbb0605f3),
	.w5(32'hbbd1cc17),
	.w6(32'h3b1980f0),
	.w7(32'hbb4560e1),
	.w8(32'hbc0aa6d2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafb952),
	.w1(32'hbad8c814),
	.w2(32'hbc0505bc),
	.w3(32'h3794c3d6),
	.w4(32'h3a9da66b),
	.w5(32'hbb0be886),
	.w6(32'hb745ecac),
	.w7(32'h3b0c5aaf),
	.w8(32'h3c06df49),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9df3ba),
	.w1(32'hbb607841),
	.w2(32'hbb968fc5),
	.w3(32'hbb1735ef),
	.w4(32'h3a816ebf),
	.w5(32'h39ebcc76),
	.w6(32'h3b9b566d),
	.w7(32'h3bd5a359),
	.w8(32'h3beb4f88),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6620f0),
	.w1(32'hbbe8ef48),
	.w2(32'hbc45ccb9),
	.w3(32'h3a312c5b),
	.w4(32'hbc02a63d),
	.w5(32'h3b262788),
	.w6(32'h3b8c4b81),
	.w7(32'hbbea0e10),
	.w8(32'hbbb7d36f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc857f29),
	.w1(32'hbc20b04c),
	.w2(32'hbc473ad5),
	.w3(32'hbb9c076e),
	.w4(32'hbb6aa474),
	.w5(32'h3c1074ba),
	.w6(32'hbc369c86),
	.w7(32'hbb0613d8),
	.w8(32'h3c11d522),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d4e2b),
	.w1(32'hbb8899df),
	.w2(32'hbbb4f2eb),
	.w3(32'h3b590471),
	.w4(32'h39babb96),
	.w5(32'hbbde86bc),
	.w6(32'h3b5bda48),
	.w7(32'hbaee5317),
	.w8(32'hbb3e87bd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0ca2a),
	.w1(32'hbbb43628),
	.w2(32'hbc03447d),
	.w3(32'hbb927a5f),
	.w4(32'h3bc33686),
	.w5(32'hbbb308d2),
	.w6(32'hbbeba09c),
	.w7(32'h3a45ac47),
	.w8(32'hbbb6bd2b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc224b5a),
	.w1(32'hbb2fdeef),
	.w2(32'hbb456f5e),
	.w3(32'h369a6e38),
	.w4(32'h3a35e974),
	.w5(32'hb992ef38),
	.w6(32'h3b76dded),
	.w7(32'hb8dd5860),
	.w8(32'h3a9042cb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab34d6),
	.w1(32'h3b895801),
	.w2(32'hba2ff943),
	.w3(32'hbb7f8978),
	.w4(32'h3b534230),
	.w5(32'hba9b7a9e),
	.w6(32'h3976197a),
	.w7(32'hbb8f5711),
	.w8(32'hbb81628b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847dfc),
	.w1(32'hb8640f08),
	.w2(32'hba90a573),
	.w3(32'h3a6d6681),
	.w4(32'h36e1f208),
	.w5(32'hbbf5ede6),
	.w6(32'hbbd422a8),
	.w7(32'hbbeb2e76),
	.w8(32'hbc72b283),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e33a6),
	.w1(32'hbbe3895a),
	.w2(32'hbc047081),
	.w3(32'hb93ecf3a),
	.w4(32'hbbc5e10d),
	.w5(32'hbba785b9),
	.w6(32'hbbcf451d),
	.w7(32'hbbdf99a3),
	.w8(32'hbba06fda),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eee8e),
	.w1(32'h3814ad63),
	.w2(32'hbac5caf1),
	.w3(32'hbb833015),
	.w4(32'hba3f2a59),
	.w5(32'h3a53ee2f),
	.w6(32'hbb736e67),
	.w7(32'hbb0afe9e),
	.w8(32'hbc1cdf3f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00c601),
	.w1(32'h38f8b769),
	.w2(32'h3ba1c2f9),
	.w3(32'hbaa05220),
	.w4(32'hbae38026),
	.w5(32'h3919b105),
	.w6(32'hbc862bb2),
	.w7(32'hbc03b017),
	.w8(32'hbc38aaf4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba643b3f),
	.w1(32'h3bcf72e0),
	.w2(32'h3bd914f2),
	.w3(32'hbaae2510),
	.w4(32'h3a8d0211),
	.w5(32'h3b273919),
	.w6(32'hbbae634c),
	.w7(32'h3bc0fa23),
	.w8(32'h3bd605af),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c163),
	.w1(32'hbac26818),
	.w2(32'hbc096ad1),
	.w3(32'hbab0acab),
	.w4(32'hbb837658),
	.w5(32'hbb8c16ac),
	.w6(32'hbab3399f),
	.w7(32'h3b32781b),
	.w8(32'hba0f3c87),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3a53e),
	.w1(32'hbb90a7c0),
	.w2(32'hbb899d51),
	.w3(32'hba19456d),
	.w4(32'hbbc02533),
	.w5(32'hbbdc9be2),
	.w6(32'hb9b191ae),
	.w7(32'hbb68bf5b),
	.w8(32'hba69df8c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc5cfc),
	.w1(32'h3be554b4),
	.w2(32'hbba4b1f9),
	.w3(32'hba4f89b8),
	.w4(32'hbbab7b58),
	.w5(32'hbbb0b539),
	.w6(32'hbb583274),
	.w7(32'h3b1b9a0a),
	.w8(32'hbbc7c093),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8261c8),
	.w1(32'hbb59c831),
	.w2(32'hbc4dfae9),
	.w3(32'h3b04adc3),
	.w4(32'h39853515),
	.w5(32'hbaec57b2),
	.w6(32'hba13cdc4),
	.w7(32'h39412952),
	.w8(32'h3ba45e8a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16ed63),
	.w1(32'h3a155eda),
	.w2(32'hbba39abd),
	.w3(32'h39bc148f),
	.w4(32'h3a6e3cb0),
	.w5(32'hbb825977),
	.w6(32'hb94bbf8e),
	.w7(32'h3b4df3f6),
	.w8(32'hbb9c0a17),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8442),
	.w1(32'hbc010f59),
	.w2(32'hbafb9401),
	.w3(32'hbbe8d0bf),
	.w4(32'hbb229644),
	.w5(32'hb9d6e3c9),
	.w6(32'hbccd21c9),
	.w7(32'hbb7661fa),
	.w8(32'hbc505d9d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e0f84),
	.w1(32'hba1f11bc),
	.w2(32'hba473f49),
	.w3(32'h3c01296d),
	.w4(32'h3b0f77de),
	.w5(32'h3b2b840f),
	.w6(32'hbb648d70),
	.w7(32'h3baa55a1),
	.w8(32'h3b98275c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6639a4),
	.w1(32'h3bcb98b1),
	.w2(32'h39f0c86d),
	.w3(32'h3b28786a),
	.w4(32'h3ba83ee4),
	.w5(32'hbb85996f),
	.w6(32'h3aa2e9f5),
	.w7(32'hbbc0834d),
	.w8(32'hbc52f28f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fea41),
	.w1(32'hbb46fb3c),
	.w2(32'hbb89d8ae),
	.w3(32'hbb968bdf),
	.w4(32'h3c4525a0),
	.w5(32'h3b11233c),
	.w6(32'h3ba7399b),
	.w7(32'h3c32bb5d),
	.w8(32'h3c0b8e44),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ba0d),
	.w1(32'hba22f814),
	.w2(32'hbbfb9f8d),
	.w3(32'h3bc7c562),
	.w4(32'hbbcf5a6b),
	.w5(32'hbb024fe6),
	.w6(32'h3b482453),
	.w7(32'h3c5b1ce5),
	.w8(32'h3c9be36f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb84a6a),
	.w1(32'hbbbf6cf4),
	.w2(32'hbbe90c48),
	.w3(32'h3ca2da88),
	.w4(32'hbba57764),
	.w5(32'hbc36e457),
	.w6(32'h3cdcca6c),
	.w7(32'hbc1cbf9f),
	.w8(32'hbc30e4cc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda444),
	.w1(32'hbab92101),
	.w2(32'h3ba1e1c9),
	.w3(32'hbbd1147c),
	.w4(32'hbba6c7ce),
	.w5(32'hbbfecc26),
	.w6(32'hbb336732),
	.w7(32'hbbaaeeab),
	.w8(32'hbb5c34ca),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca69227),
	.w1(32'h3bd1296e),
	.w2(32'hbc0773a0),
	.w3(32'h3bca8894),
	.w4(32'h3b4c4ff1),
	.w5(32'hbbabee73),
	.w6(32'h3b56df65),
	.w7(32'hbba11fbd),
	.w8(32'hbc266c54),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58650d),
	.w1(32'hbbf64783),
	.w2(32'hbbde5693),
	.w3(32'hbb586aaa),
	.w4(32'hbb9b8c4a),
	.w5(32'hbbbf4954),
	.w6(32'hbb442dcf),
	.w7(32'hbbf45e57),
	.w8(32'hb931a5d5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74acd),
	.w1(32'hba09f57c),
	.w2(32'hbb620e7d),
	.w3(32'hb9835730),
	.w4(32'h3b82a07d),
	.w5(32'h3ba6ea3a),
	.w6(32'hbaa80e21),
	.w7(32'hbb7c166a),
	.w8(32'hbad34fd9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6227e),
	.w1(32'hbb3d6d1a),
	.w2(32'hbc1a0d6b),
	.w3(32'hba5097c0),
	.w4(32'h3bad2c3f),
	.w5(32'h3988e7dc),
	.w6(32'h39a83668),
	.w7(32'h3a92e01f),
	.w8(32'h3ad4b123),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9ce75),
	.w1(32'hbba29d27),
	.w2(32'hbbe6c1f9),
	.w3(32'hbbcbda97),
	.w4(32'hb9befe06),
	.w5(32'h3b38d3e1),
	.w6(32'h39c466c0),
	.w7(32'h3b58f3e4),
	.w8(32'h3b913716),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba622b5),
	.w1(32'hbacf7b09),
	.w2(32'hbbca42f2),
	.w3(32'hba7d1eb1),
	.w4(32'hb8e47841),
	.w5(32'hbc0de6e7),
	.w6(32'h3b8c34bf),
	.w7(32'h3badd6a8),
	.w8(32'h3b8dd2d1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dcc61),
	.w1(32'hbb8a1466),
	.w2(32'hbb605484),
	.w3(32'hbc16b23b),
	.w4(32'hbaf74025),
	.w5(32'hbae3a229),
	.w6(32'h3b68b789),
	.w7(32'h3a644380),
	.w8(32'hba80ed3a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac722c),
	.w1(32'hbbd43b95),
	.w2(32'hbc61f5e8),
	.w3(32'hbb3e674f),
	.w4(32'h3be958ad),
	.w5(32'h3b73cc62),
	.w6(32'hbb484147),
	.w7(32'h3b3cca89),
	.w8(32'hbbd655c1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d5f70),
	.w1(32'h3ab97f32),
	.w2(32'hbc77a803),
	.w3(32'h3bf575a0),
	.w4(32'h3bca234d),
	.w5(32'hba1fe6af),
	.w6(32'hbb58e053),
	.w7(32'hbbfb0ec0),
	.w8(32'hbc931998),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8da9c1),
	.w1(32'h3b522d22),
	.w2(32'hbbdff00a),
	.w3(32'h3c8edb70),
	.w4(32'h3aa0f122),
	.w5(32'hbc2c5258),
	.w6(32'h3c21328d),
	.w7(32'hbbe421f9),
	.w8(32'hbccb3327),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bab23),
	.w1(32'hbba55c9d),
	.w2(32'h39431200),
	.w3(32'h3bd0e965),
	.w4(32'hba659545),
	.w5(32'h3b0e2fbb),
	.w6(32'hbbcd40f4),
	.w7(32'h39dd4785),
	.w8(32'hbb6d57de),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba040938),
	.w1(32'hbaf7895a),
	.w2(32'h3c1abade),
	.w3(32'h3959b77d),
	.w4(32'hbbfc5dd2),
	.w5(32'hbbe4ab43),
	.w6(32'h3b005eec),
	.w7(32'hbbca7708),
	.w8(32'hbc00d0c3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64f667),
	.w1(32'h3b0b9a17),
	.w2(32'hbabd3982),
	.w3(32'hbb640de6),
	.w4(32'hb9ab50fd),
	.w5(32'h3a4deddb),
	.w6(32'hbae87949),
	.w7(32'hbb8ca5d7),
	.w8(32'h3ab7c0be),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d5c33),
	.w1(32'h3bc73aad),
	.w2(32'h3b6bddfc),
	.w3(32'h3be6e216),
	.w4(32'h3b85c905),
	.w5(32'h3b23ebf2),
	.w6(32'hba3f1f0c),
	.w7(32'hb9a9093c),
	.w8(32'hbb98417f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a404),
	.w1(32'h3ba13742),
	.w2(32'h3c051a1b),
	.w3(32'hbba17796),
	.w4(32'h3ba59533),
	.w5(32'h3a7de38c),
	.w6(32'hbc339e73),
	.w7(32'hbac3bd76),
	.w8(32'hbb9cd008),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97149f),
	.w1(32'hb9d3eedb),
	.w2(32'hbbe5e8f8),
	.w3(32'h3b343d58),
	.w4(32'h3bb56d19),
	.w5(32'hbb42e3f2),
	.w6(32'hbb88ec3e),
	.w7(32'hba8e378a),
	.w8(32'hbc1088ef),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009038),
	.w1(32'h3bb8fb80),
	.w2(32'h3b0366d6),
	.w3(32'hba7f576f),
	.w4(32'hb98a3a12),
	.w5(32'h3afbed93),
	.w6(32'hbc0814db),
	.w7(32'hbc39324c),
	.w8(32'hbc6e0506),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77647),
	.w1(32'hb9b751bc),
	.w2(32'h3b1980f9),
	.w3(32'hbb4d0005),
	.w4(32'hbabc399a),
	.w5(32'hbb204857),
	.w6(32'hbc3b3494),
	.w7(32'hbbc5e596),
	.w8(32'hbbb4c076),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8001a4),
	.w1(32'hba1e0f17),
	.w2(32'h38312a41),
	.w3(32'hbab714e5),
	.w4(32'hbc0b3dff),
	.w5(32'hbbb7447c),
	.w6(32'hbbbdf39c),
	.w7(32'hbbfafb8c),
	.w8(32'hbc629b8a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3b923),
	.w1(32'hbbcd7ee1),
	.w2(32'hbc54189e),
	.w3(32'h3ba5583c),
	.w4(32'hbb11dd36),
	.w5(32'hbbce6119),
	.w6(32'hbabb55c9),
	.w7(32'h3a67da70),
	.w8(32'h3ade3c93),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324842),
	.w1(32'h3b09436f),
	.w2(32'hbbb78bf3),
	.w3(32'hbbe0eb10),
	.w4(32'h3c1d8197),
	.w5(32'h3bf68ea6),
	.w6(32'hba2bb5c7),
	.w7(32'h3bd11883),
	.w8(32'h3bc0ae27),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc386290),
	.w1(32'hbb23d01d),
	.w2(32'h3a77a865),
	.w3(32'hbab61aed),
	.w4(32'hbba2554e),
	.w5(32'hbb8b88b0),
	.w6(32'h3c03cc15),
	.w7(32'hbb7e29b5),
	.w8(32'h3a6ede7c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8543dd),
	.w1(32'hbbf735cb),
	.w2(32'hbb5aa719),
	.w3(32'hbb1a97e7),
	.w4(32'hb99f79b8),
	.w5(32'h3b23bbac),
	.w6(32'hbbef7238),
	.w7(32'hbb6c99ce),
	.w8(32'h3a9ec671),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dd4eb),
	.w1(32'hbb244bd2),
	.w2(32'hbbdd3940),
	.w3(32'h3b91c6d6),
	.w4(32'h39d5584b),
	.w5(32'h3b97c18f),
	.w6(32'hbb1ad521),
	.w7(32'h3b131853),
	.w8(32'h3bb5eccb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aaf1a),
	.w1(32'hbb3ca50e),
	.w2(32'hbc8579db),
	.w3(32'hbbd844bf),
	.w4(32'h3b413984),
	.w5(32'hb9a965a3),
	.w6(32'h39d58dea),
	.w7(32'h3b98d4a2),
	.w8(32'h3b94bd82),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa639),
	.w1(32'h3a9fd9ea),
	.w2(32'hbb1f820f),
	.w3(32'hbbc43d9e),
	.w4(32'h3a070176),
	.w5(32'h3a393d51),
	.w6(32'h3acadd70),
	.w7(32'h3ba43298),
	.w8(32'hbb1a7e35),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eecfd),
	.w1(32'h395fe841),
	.w2(32'hbbd4aeed),
	.w3(32'hbb79be15),
	.w4(32'h3b70fe66),
	.w5(32'h3c10c91a),
	.w6(32'h3b317055),
	.w7(32'hbb01408a),
	.w8(32'hbabe268c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22993a),
	.w1(32'hbb075cb7),
	.w2(32'hbb87c16d),
	.w3(32'hbae1d9a2),
	.w4(32'hb8fad501),
	.w5(32'hba6668a5),
	.w6(32'hbaa87055),
	.w7(32'h3a8299fa),
	.w8(32'h3bd027e4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3fd32),
	.w1(32'hbc02c3f1),
	.w2(32'h39dcf8bc),
	.w3(32'h3bcf997f),
	.w4(32'hbb97772c),
	.w5(32'h3b1933bb),
	.w6(32'h3ab1bec3),
	.w7(32'hbafed5ac),
	.w8(32'h3a712de4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3487d),
	.w1(32'h3a92f615),
	.w2(32'h3bfa50ba),
	.w3(32'hbb056b11),
	.w4(32'h3b4e6375),
	.w5(32'h3b264127),
	.w6(32'hbaab4790),
	.w7(32'h3a46175e),
	.w8(32'h38a08dac),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c3712),
	.w1(32'h3acbb738),
	.w2(32'hbae9bce6),
	.w3(32'h3c17b227),
	.w4(32'hbb36fada),
	.w5(32'hba5d1cf3),
	.w6(32'h3b91c53a),
	.w7(32'hb9cd97c3),
	.w8(32'hbac98d53),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefc708),
	.w1(32'h3ae6f037),
	.w2(32'hb9e7dc27),
	.w3(32'h3b68bfa1),
	.w4(32'h39f488d3),
	.w5(32'hbb51abea),
	.w6(32'h3bbe931a),
	.w7(32'h3c423939),
	.w8(32'h3c5f0dca),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a865ac0),
	.w1(32'hbba3cf35),
	.w2(32'hbc1b3682),
	.w3(32'h3983367b),
	.w4(32'hba9f0613),
	.w5(32'hbc070763),
	.w6(32'h3baedc4a),
	.w7(32'h3bc09e2a),
	.w8(32'h3a6978ef),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde3875),
	.w1(32'h3ba88190),
	.w2(32'h3bf0e387),
	.w3(32'hbbd551ee),
	.w4(32'h3a5af12b),
	.w5(32'hba44b336),
	.w6(32'hbba36412),
	.w7(32'hbbcf3bcb),
	.w8(32'hbc5fb138),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae99507),
	.w1(32'h3b66feeb),
	.w2(32'h3a8e6f7f),
	.w3(32'hbb5c50a7),
	.w4(32'h3b002232),
	.w5(32'hb9134276),
	.w6(32'hbbdb8660),
	.w7(32'h3b10d454),
	.w8(32'h3bab1466),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822262),
	.w1(32'hbaf14249),
	.w2(32'hbbe1716e),
	.w3(32'h3a733f7b),
	.w4(32'h3bc3a450),
	.w5(32'h3b8cff34),
	.w6(32'h3a8caa1e),
	.w7(32'h3c041142),
	.w8(32'h3c188b97),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe66e4c),
	.w1(32'hbb31930e),
	.w2(32'hbbea970f),
	.w3(32'hbb512598),
	.w4(32'h38f6d697),
	.w5(32'h3b4b59ee),
	.w6(32'h3b19d7b1),
	.w7(32'h3a443d23),
	.w8(32'hba46aa67),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38204f),
	.w1(32'hbb1e5233),
	.w2(32'hbba136ea),
	.w3(32'h3af40f0f),
	.w4(32'h39f354f6),
	.w5(32'hbbaea06d),
	.w6(32'hbb22d261),
	.w7(32'hbb326e29),
	.w8(32'hba538019),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb150c45),
	.w1(32'h3a0a2941),
	.w2(32'hbabb7da7),
	.w3(32'hbb6222d9),
	.w4(32'h3ab8405c),
	.w5(32'h3a15c62c),
	.w6(32'hbc414a50),
	.w7(32'hbb2456a2),
	.w8(32'hbb38af96),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7cc1f),
	.w1(32'h3b97a9eb),
	.w2(32'hbadadac5),
	.w3(32'hbc047d4c),
	.w4(32'h3a98cb16),
	.w5(32'hbc2262da),
	.w6(32'hbc818114),
	.w7(32'hbbb2a9c5),
	.w8(32'hbc5f7654),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1cc21),
	.w1(32'h3bdce70b),
	.w2(32'hbbb611c0),
	.w3(32'h3b5d966a),
	.w4(32'h3c1892d8),
	.w5(32'hb9dec2fc),
	.w6(32'hbb793b48),
	.w7(32'hbb5b939e),
	.w8(32'hbc5324a8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37882551),
	.w1(32'hb83f8d65),
	.w2(32'h38b60350),
	.w3(32'h3819db2e),
	.w4(32'hb72eb57d),
	.w5(32'h38fb5c3a),
	.w6(32'h38c62a9f),
	.w7(32'h3884f576),
	.w8(32'h39442633),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddf66a),
	.w1(32'h37dc5f69),
	.w2(32'h392b29f9),
	.w3(32'h38ef4a24),
	.w4(32'h37fefdc8),
	.w5(32'h3950e5b9),
	.w6(32'h3972c4b2),
	.w7(32'h3910be69),
	.w8(32'h39a376d3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39036269),
	.w1(32'hb843c324),
	.w2(32'h391a5b6c),
	.w3(32'h391c03a0),
	.w4(32'hb8040646),
	.w5(32'h39377fa4),
	.w6(32'h3975493e),
	.w7(32'h38be0fa5),
	.w8(32'h398dbcfb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f23da6),
	.w1(32'h3a17f6f2),
	.w2(32'hb8a90b6e),
	.w3(32'hb9c628ae),
	.w4(32'h39ca1a77),
	.w5(32'hb9f76f06),
	.w6(32'hba9f6835),
	.w7(32'h39f76259),
	.w8(32'h39063b0e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac93b6),
	.w1(32'hb817a157),
	.w2(32'h391d7f1f),
	.w3(32'h3896feb7),
	.w4(32'hb8cb5f55),
	.w5(32'h3883403d),
	.w6(32'h3907f89f),
	.w7(32'hb7a8c91b),
	.w8(32'h390e6164),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49c48f),
	.w1(32'hbb2c6e8c),
	.w2(32'hbae0d526),
	.w3(32'hbb2a892c),
	.w4(32'hbb5d5eae),
	.w5(32'hba888a8a),
	.w6(32'hbb0bf278),
	.w7(32'hbae9edfc),
	.w8(32'hba9f950f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed1813),
	.w1(32'hbb4fa126),
	.w2(32'hbb4d1615),
	.w3(32'hbb7f8229),
	.w4(32'hbb90969a),
	.w5(32'hbb56c947),
	.w6(32'hbc02696d),
	.w7(32'hbafef3aa),
	.w8(32'hbb12497c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad46baa),
	.w1(32'h3a009ecc),
	.w2(32'hba9bc042),
	.w3(32'hb93df980),
	.w4(32'h3b2e04df),
	.w5(32'h3acfe1cd),
	.w6(32'hbb0ff548),
	.w7(32'hba73c5c2),
	.w8(32'hbb275f3d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc3f90),
	.w1(32'h3a66c4d9),
	.w2(32'hbaee027a),
	.w3(32'hbac20236),
	.w4(32'h3b036d9c),
	.w5(32'hba9b5cc5),
	.w6(32'hbb2a9120),
	.w7(32'h3a7cfdad),
	.w8(32'hbab62347),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270c15),
	.w1(32'hba26d4c4),
	.w2(32'hbac08290),
	.w3(32'hb9d60789),
	.w4(32'hb5323e18),
	.w5(32'h39843a8d),
	.w6(32'hb97b94d1),
	.w7(32'hb7ae5a3d),
	.w8(32'hba170b17),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8819fa),
	.w1(32'h39c412cb),
	.w2(32'hbae82fd0),
	.w3(32'hba55df78),
	.w4(32'h3aaf93a1),
	.w5(32'hba064cfb),
	.w6(32'hbaa71925),
	.w7(32'hba121ac6),
	.w8(32'hbae20194),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d5a71),
	.w1(32'hba682afc),
	.w2(32'hbb13175c),
	.w3(32'hbb05fc44),
	.w4(32'hba709863),
	.w5(32'hbb22cf86),
	.w6(32'hbb2aa710),
	.w7(32'hba046b54),
	.w8(32'hbb2b1c0f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a28799),
	.w1(32'hb75b8f1e),
	.w2(32'h35166acb),
	.w3(32'h37f3bb71),
	.w4(32'hb714e28e),
	.w5(32'h36bdc81b),
	.w6(32'h382a838c),
	.w7(32'h3731e532),
	.w8(32'h37c07354),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b08aa0),
	.w1(32'hb8773b61),
	.w2(32'hb81bcaa4),
	.w3(32'hb838bcce),
	.w4(32'h3683e7a6),
	.w5(32'h38a03238),
	.w6(32'hb89c9e02),
	.w7(32'hb79c0d82),
	.w8(32'h36b33bf4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795a356),
	.w1(32'h38b7eaf1),
	.w2(32'h394b2a2b),
	.w3(32'hb89e2432),
	.w4(32'h39178fad),
	.w5(32'h39267176),
	.w6(32'hb820dfdb),
	.w7(32'h38ace572),
	.w8(32'h3939daa4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaa0bb),
	.w1(32'h3a0505c5),
	.w2(32'hb9258c60),
	.w3(32'h3a781bfd),
	.w4(32'hb8dc3da2),
	.w5(32'hba889604),
	.w6(32'h3a97c11f),
	.w7(32'hb99fc93e),
	.w8(32'hba911fd6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11eb3a),
	.w1(32'h3a390ca3),
	.w2(32'hbb4b47ce),
	.w3(32'hbb1889b6),
	.w4(32'h3b1699bf),
	.w5(32'hb901528e),
	.w6(32'hbbac00bd),
	.w7(32'hbb107521),
	.w8(32'hbb9a5bf3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0846b2),
	.w1(32'h3a8a6d32),
	.w2(32'h39371a68),
	.w3(32'h39b141b4),
	.w4(32'h3a6b7f91),
	.w5(32'h3940bbda),
	.w6(32'hb990dc09),
	.w7(32'h39d9c764),
	.w8(32'hb926e9d7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35e6ce),
	.w1(32'h3a0eab96),
	.w2(32'hb8f86da5),
	.w3(32'hba4499f5),
	.w4(32'h3aa4ec6b),
	.w5(32'h3a93a52f),
	.w6(32'hbb9bfcee),
	.w7(32'hbaeb1e6e),
	.w8(32'hbb05a85f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbead35a),
	.w1(32'hbac043ab),
	.w2(32'hbb56706c),
	.w3(32'hbbec466b),
	.w4(32'hbb5ec9b3),
	.w5(32'hbb9a407e),
	.w6(32'hbc04eee2),
	.w7(32'hbb078169),
	.w8(32'hbbbea91e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c272209),
	.w1(32'h3b60d1f6),
	.w2(32'hbaf571cc),
	.w3(32'h3bcbc798),
	.w4(32'hb9c79f7d),
	.w5(32'hbbc15043),
	.w6(32'h3b8e7c4a),
	.w7(32'hbb43a0eb),
	.w8(32'hbc14584f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6f498),
	.w1(32'hbb81ea5b),
	.w2(32'hba96f07b),
	.w3(32'hb93ec6a8),
	.w4(32'hb91e87f1),
	.w5(32'h3a54344a),
	.w6(32'hbbe2f43a),
	.w7(32'hbb810139),
	.w8(32'hbb99e3db),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4c8c),
	.w1(32'h3a314eac),
	.w2(32'hbb892226),
	.w3(32'h3a4f955a),
	.w4(32'hbac5b77f),
	.w5(32'hbbadaf86),
	.w6(32'hbadd3e81),
	.w7(32'hbb7ef4e0),
	.w8(32'hbbefbabf),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e50a),
	.w1(32'h3a2ce103),
	.w2(32'hbae6fe56),
	.w3(32'hbb4b7bab),
	.w4(32'h3bb69512),
	.w5(32'h3b1ccaab),
	.w6(32'hbbedf449),
	.w7(32'hb988b2af),
	.w8(32'hba32471e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0df953),
	.w1(32'hba003fff),
	.w2(32'hba83a4ef),
	.w3(32'hb9272316),
	.w4(32'h3acf639a),
	.w5(32'h3a6dbfec),
	.w6(32'hbb1fb51f),
	.w7(32'hbaaf598f),
	.w8(32'hbb893664),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1754e),
	.w1(32'h3b08e596),
	.w2(32'hbb1d92d3),
	.w3(32'h3b68d777),
	.w4(32'h3aa7ac33),
	.w5(32'hbb5df10a),
	.w6(32'h3b2842a3),
	.w7(32'hbb2c4249),
	.w8(32'hbbe14093),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a58cf1),
	.w1(32'hb98e4ced),
	.w2(32'hb85816f1),
	.w3(32'hba03f4dd),
	.w4(32'hba02d61b),
	.w5(32'h396ce6a7),
	.w6(32'hb984f6fd),
	.w7(32'hb98c5fe2),
	.w8(32'h39414692),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81d463),
	.w1(32'hb92b1957),
	.w2(32'hbb5c798f),
	.w3(32'hbb86885b),
	.w4(32'h3abf59fa),
	.w5(32'hbacda5e5),
	.w6(32'hbbe4c859),
	.w7(32'hbaa54df7),
	.w8(32'hbb5c4d33),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f23b2),
	.w1(32'hbaf80d2f),
	.w2(32'hbada3e02),
	.w3(32'hbb535b93),
	.w4(32'hbb386fcd),
	.w5(32'hbb1ae50d),
	.w6(32'hbb98b49c),
	.w7(32'hbba2cd56),
	.w8(32'hbbabaf91),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc657b46),
	.w1(32'hbc011377),
	.w2(32'hbbdfe2ed),
	.w3(32'hbbc5a276),
	.w4(32'hbba50a69),
	.w5(32'h3b82902d),
	.w6(32'hbc6ed74a),
	.w7(32'h39eb7585),
	.w8(32'hb9fb5093),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9d6a),
	.w1(32'h3b79ce20),
	.w2(32'hbb904ba5),
	.w3(32'h3bbb86df),
	.w4(32'h3b4dde0d),
	.w5(32'hbb9381fa),
	.w6(32'hbb739ddb),
	.w7(32'hbbcf91ef),
	.w8(32'hbc79878a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a629a11),
	.w1(32'h3b4c10b6),
	.w2(32'hbb40fb49),
	.w3(32'hba756e3b),
	.w4(32'h3b863189),
	.w5(32'h3a295b39),
	.w6(32'hbbae6e20),
	.w7(32'hb9c780b5),
	.w8(32'hbb8a4e91),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06808e),
	.w1(32'hbba5174c),
	.w2(32'hbba27d09),
	.w3(32'hbb6bb544),
	.w4(32'hbb7389c2),
	.w5(32'h3abd105c),
	.w6(32'hbbbfe2ad),
	.w7(32'h394e7721),
	.w8(32'hba0f0eb1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d14574),
	.w1(32'hba240b69),
	.w2(32'h39afb9c8),
	.w3(32'h38949e14),
	.w4(32'hba81ca10),
	.w5(32'h39eaac17),
	.w6(32'hba102bfa),
	.w7(32'hba99f7bb),
	.w8(32'h39497139),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc716281),
	.w1(32'hbbfd52e7),
	.w2(32'hbc37cda8),
	.w3(32'hbbc902c1),
	.w4(32'hbb196af9),
	.w5(32'h3b205353),
	.w6(32'hbb69b847),
	.w7(32'h3a614330),
	.w8(32'hbb75d472),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba879ec6),
	.w1(32'hba20a547),
	.w2(32'hbb7e08cc),
	.w3(32'hbaca2b87),
	.w4(32'hbad77902),
	.w5(32'hbb5fffc5),
	.w6(32'hbb0e31a3),
	.w7(32'hbb2ac4d4),
	.w8(32'hba8daa73),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aa652),
	.w1(32'hb911ab89),
	.w2(32'hb9b8da37),
	.w3(32'h3a1bdbcd),
	.w4(32'hb8ee8b7a),
	.w5(32'hb992f06b),
	.w6(32'h3a2fcede),
	.w7(32'hb83dfa7b),
	.w8(32'hb977b53d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9d146),
	.w1(32'hba78d74c),
	.w2(32'hba0033d4),
	.w3(32'hbaa6575c),
	.w4(32'h39d3bc54),
	.w5(32'h39b58d4f),
	.w6(32'hbb31e3be),
	.w7(32'hba74f79a),
	.w8(32'hbaa34999),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb505a2d),
	.w1(32'h3787ccad),
	.w2(32'hba9e7cbf),
	.w3(32'hbaf6b2e3),
	.w4(32'h3a034fb8),
	.w5(32'hba4a23c5),
	.w6(32'hbb94fc80),
	.w7(32'hba3eabf8),
	.w8(32'hbb24e6dc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a0188),
	.w1(32'h3b3fd5e9),
	.w2(32'hba820b82),
	.w3(32'h3a4040c5),
	.w4(32'h3b0b4d55),
	.w5(32'hb9044c97),
	.w6(32'hbab1549b),
	.w7(32'hba1c93cd),
	.w8(32'hbb41dd19),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb105af),
	.w1(32'h3a028a75),
	.w2(32'hbb6db481),
	.w3(32'h3ba31a53),
	.w4(32'h3a4bd556),
	.w5(32'hbb8ccbd7),
	.w6(32'h3b912eab),
	.w7(32'hbb183387),
	.w8(32'hbc0c1830),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f96c52),
	.w1(32'h3a0072be),
	.w2(32'hba0a89ea),
	.w3(32'h3b09a6bd),
	.w4(32'h3b4a30b8),
	.w5(32'h3b0f6cad),
	.w6(32'hba35a031),
	.w7(32'hba14c6ba),
	.w8(32'hbb28510f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7a07c),
	.w1(32'h3ac5ef71),
	.w2(32'h3a82e54b),
	.w3(32'hbae18f2d),
	.w4(32'h3a2b1bde),
	.w5(32'h3aae5ad1),
	.w6(32'hbbe5b3ff),
	.w7(32'hbad64532),
	.w8(32'h38bc1503),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7be9e),
	.w1(32'hbb438145),
	.w2(32'hbb270bff),
	.w3(32'hbb317abe),
	.w4(32'h3af8e6ac),
	.w5(32'hb91c6dce),
	.w6(32'hbbe99246),
	.w7(32'hba53a72d),
	.w8(32'hbb19f735),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e2e58a),
	.w1(32'h3ab8ef41),
	.w2(32'hba8e96f7),
	.w3(32'hb9d685ae),
	.w4(32'h3ab1e5b2),
	.w5(32'hba2d8e1f),
	.w6(32'hbb2ee7cb),
	.w7(32'hba78a627),
	.w8(32'hbb229396),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9066916),
	.w1(32'hb8c6ec5f),
	.w2(32'h3769d0ad),
	.w3(32'hb8ff5963),
	.w4(32'hb811756b),
	.w5(32'h384fea83),
	.w6(32'hb91ba2ab),
	.w7(32'hb8d380fb),
	.w8(32'hb7845419),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47060b),
	.w1(32'hb9007ec8),
	.w2(32'hb8a2f9d0),
	.w3(32'hb7eee400),
	.w4(32'h3a112ead),
	.w5(32'h3a436d25),
	.w6(32'hba331259),
	.w7(32'hb964da2b),
	.w8(32'hb8b31c4f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387b8d4d),
	.w1(32'h385aae78),
	.w2(32'h3880e10f),
	.w3(32'h38613c5d),
	.w4(32'h38146ca2),
	.w5(32'h388ea028),
	.w6(32'h3891e18b),
	.w7(32'h3842e072),
	.w8(32'h3871c1d7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7829f),
	.w1(32'h39f63fa9),
	.w2(32'h39600e31),
	.w3(32'hb91e0c33),
	.w4(32'hb814f203),
	.w5(32'hb96f1b77),
	.w6(32'hb76aac69),
	.w7(32'h38c87f52),
	.w8(32'hb9a28b33),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00310d),
	.w1(32'h3acdb92d),
	.w2(32'hbaa86098),
	.w3(32'hba31856c),
	.w4(32'h3b195abd),
	.w5(32'h39f5e892),
	.w6(32'hbb5ac09a),
	.w7(32'hba15fea9),
	.w8(32'hbb30da28),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf5efe),
	.w1(32'h394a65e8),
	.w2(32'hb9505ccd),
	.w3(32'h3a035c54),
	.w4(32'h38ebbc99),
	.w5(32'hba2c9d69),
	.w6(32'h39a731b8),
	.w7(32'h38d42beb),
	.w8(32'hba6d5982),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bc549),
	.w1(32'hbb042ae3),
	.w2(32'hba93ffb7),
	.w3(32'hbb09a12d),
	.w4(32'hbb02d48b),
	.w5(32'hba82feca),
	.w6(32'hbb1493a5),
	.w7(32'hbaad4fa8),
	.w8(32'hba4831a3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19a27b),
	.w1(32'h3961ae1d),
	.w2(32'hbb56f49c),
	.w3(32'h3b201aa2),
	.w4(32'h3b0cbf5a),
	.w5(32'hba85a254),
	.w6(32'h39b9e23f),
	.w7(32'hbb395a34),
	.w8(32'hbbc3ed84),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac8136),
	.w1(32'h379bcaf4),
	.w2(32'h36eb961f),
	.w3(32'h3913a471),
	.w4(32'h38d70df5),
	.w5(32'h3848bcf0),
	.w6(32'h3951ac2f),
	.w7(32'h39045064),
	.w8(32'h38818cd3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e6944),
	.w1(32'h399b24f6),
	.w2(32'hb78b1ac3),
	.w3(32'h38417ece),
	.w4(32'h396fd2a2),
	.w5(32'h383bef4a),
	.w6(32'hb7798fe0),
	.w7(32'h38dfa697),
	.w8(32'hb9351f2a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385fa4bc),
	.w1(32'h37bfd031),
	.w2(32'h3709e830),
	.w3(32'h38404988),
	.w4(32'h380b0673),
	.w5(32'hb3b23ac6),
	.w6(32'h380c1ba7),
	.w7(32'h37e759f7),
	.w8(32'h36ab0629),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e92d4),
	.w1(32'h395c3dd0),
	.w2(32'hb90a44a6),
	.w3(32'hb9320514),
	.w4(32'h395db105),
	.w5(32'hb9400717),
	.w6(32'hba9320fc),
	.w7(32'hba1addf9),
	.w8(32'hba1320e4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b022323),
	.w1(32'hbb094667),
	.w2(32'h3a7eda5e),
	.w3(32'hba21c730),
	.w4(32'hb9b07e5a),
	.w5(32'hb96faaa5),
	.w6(32'hbb9940ee),
	.w7(32'h392cbc75),
	.w8(32'h39a227a4),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03dde7),
	.w1(32'h3a1b194a),
	.w2(32'hbb8e0da6),
	.w3(32'hbb437a95),
	.w4(32'h39192062),
	.w5(32'hbb722c3b),
	.w6(32'hbb77ac05),
	.w7(32'hb9850729),
	.w8(32'hbb528088),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8725da),
	.w1(32'hb95d9ff9),
	.w2(32'hb90bc403),
	.w3(32'hb8b6fdc4),
	.w4(32'hb8dfcfbe),
	.w5(32'h38a276a8),
	.w6(32'hba01343a),
	.w7(32'hb9c10216),
	.w8(32'hb9b9fc32),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac955ac),
	.w1(32'hba0a0c6b),
	.w2(32'hbaf3c357),
	.w3(32'hba3542d6),
	.w4(32'h37fa9d6a),
	.w5(32'hba86e86c),
	.w6(32'hbb38898c),
	.w7(32'h39c71a57),
	.w8(32'hba823b37),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bf43f),
	.w1(32'hb986b92e),
	.w2(32'hba4c4dbf),
	.w3(32'hb94de626),
	.w4(32'h394ac741),
	.w5(32'hba0340be),
	.w6(32'hba402f23),
	.w7(32'hba60f3d1),
	.w8(32'hbadea18b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0bbf),
	.w1(32'h3a69a8e8),
	.w2(32'hba90eca1),
	.w3(32'hba43d9e3),
	.w4(32'h3b21e861),
	.w5(32'h39fba6b3),
	.w6(32'hbaec3a32),
	.w7(32'h3a311670),
	.w8(32'h390f237c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dbc0e),
	.w1(32'hb8d37274),
	.w2(32'hbb637dda),
	.w3(32'hbaeed6fe),
	.w4(32'h3b0cf45c),
	.w5(32'hbaa861eb),
	.w6(32'hbb2312c8),
	.w7(32'hbab808c4),
	.w8(32'hbb5e46b8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98e72f),
	.w1(32'hbb3d16ae),
	.w2(32'hbb7b3df7),
	.w3(32'hbb8e0be0),
	.w4(32'hbaee6a0b),
	.w5(32'hbb8ff3d9),
	.w6(32'hbb97bb89),
	.w7(32'hba81e430),
	.w8(32'hbb936b79),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54c993),
	.w1(32'h3a81c6eb),
	.w2(32'hba808094),
	.w3(32'h394f3d96),
	.w4(32'h3afa1ca6),
	.w5(32'h393fc51e),
	.w6(32'hba85812e),
	.w7(32'hbad23fed),
	.w8(32'hbb3f4936),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440db0),
	.w1(32'hbaaf5fda),
	.w2(32'h38863454),
	.w3(32'hbb076e43),
	.w4(32'h39cfd865),
	.w5(32'h3a348541),
	.w6(32'hbba49449),
	.w7(32'hbab75e37),
	.w8(32'hbad5ad97),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac88ec),
	.w1(32'hbb2722e7),
	.w2(32'hbb5c124d),
	.w3(32'hbb9ffb44),
	.w4(32'hbb2dbcc4),
	.w5(32'hbb33a4a8),
	.w6(32'hbb99ae16),
	.w7(32'hb9b1c094),
	.w8(32'hbb217a3c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c2ea0),
	.w1(32'hb994b2b1),
	.w2(32'hb9a44f91),
	.w3(32'hba98f834),
	.w4(32'h3ac6c88d),
	.w5(32'h3b30b342),
	.w6(32'hbbba14c0),
	.w7(32'hba8a9fca),
	.w8(32'hba349808),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb208745),
	.w1(32'hba2f7492),
	.w2(32'hbac56d93),
	.w3(32'hba82f794),
	.w4(32'h3a199bcd),
	.w5(32'hb9ce9294),
	.w6(32'hbb7fc141),
	.w7(32'hbad65cf6),
	.w8(32'hbb355607),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f4cf25),
	.w1(32'h39c2bb61),
	.w2(32'hba1939f6),
	.w3(32'h382b9348),
	.w4(32'h3a155ac2),
	.w5(32'hb90cccc3),
	.w6(32'hba404b1b),
	.w7(32'hb9352229),
	.w8(32'hba755554),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90cac8),
	.w1(32'h3b0cc191),
	.w2(32'hb9b16eda),
	.w3(32'h3c4ef112),
	.w4(32'hbafd4502),
	.w5(32'hbbd410f3),
	.w6(32'h3c24b921),
	.w7(32'hbb9db593),
	.w8(32'hbc2c9400),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc26ca),
	.w1(32'h3818214e),
	.w2(32'hba86e509),
	.w3(32'hbadaf656),
	.w4(32'hb983e77b),
	.w5(32'hba74e3f4),
	.w6(32'hbb0f5fe5),
	.w7(32'hba1d03b7),
	.w8(32'hbad80369),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e0056),
	.w1(32'hb8fa8569),
	.w2(32'hb866c93b),
	.w3(32'hb906745a),
	.w4(32'hb903f7ba),
	.w5(32'hb88a06bb),
	.w6(32'hb941809c),
	.w7(32'hb912c902),
	.w8(32'hb7873186),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f28989),
	.w1(32'hb844fbea),
	.w2(32'h38002b38),
	.w3(32'h390421e6),
	.w4(32'h37278e16),
	.w5(32'h386a1322),
	.w6(32'h38f2d860),
	.w7(32'hb69b8a69),
	.w8(32'hb7a19898),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacddb2b),
	.w1(32'hb9be17b0),
	.w2(32'hba3fe64a),
	.w3(32'hba6d745f),
	.w4(32'hb943d6e8),
	.w5(32'hb8dbd1e4),
	.w6(32'hbaccca98),
	.w7(32'hb9928148),
	.w8(32'hb9e1fa07),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1e843),
	.w1(32'h3a6341c7),
	.w2(32'hba8a5fe7),
	.w3(32'hb96d24d2),
	.w4(32'h3b26ca01),
	.w5(32'h3b074c7e),
	.w6(32'hbb57e7de),
	.w7(32'hbb0fe895),
	.w8(32'hbb9314b4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62436a),
	.w1(32'h3a8c5030),
	.w2(32'hba961969),
	.w3(32'hbad619ad),
	.w4(32'h3adddcda),
	.w5(32'hb8a7e5c5),
	.w6(32'hbb609c56),
	.w7(32'h39cf536d),
	.w8(32'hbadcdc3a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ba4684),
	.w1(32'hb6c19ed5),
	.w2(32'h37ecb462),
	.w3(32'h363f64f8),
	.w4(32'h3659448b),
	.w5(32'h37f940a5),
	.w6(32'h37837b58),
	.w7(32'h3802e35e),
	.w8(32'h384ed0fd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506a32),
	.w1(32'h3a4ffce4),
	.w2(32'hbb590edf),
	.w3(32'hbab09e63),
	.w4(32'h3a5523a6),
	.w5(32'hbaf6920c),
	.w6(32'hbb6ff0ac),
	.w7(32'hbb042e94),
	.w8(32'hbb81a24f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf74d26),
	.w1(32'h39c9fbb7),
	.w2(32'hbac039b1),
	.w3(32'hba92649a),
	.w4(32'h3a34b248),
	.w5(32'hb99401be),
	.w6(32'hbb7d42bd),
	.w7(32'hbab7b003),
	.w8(32'hbb13c12d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd452aa),
	.w1(32'hbb16d7ab),
	.w2(32'hba9a1e97),
	.w3(32'hbb81c9f2),
	.w4(32'hbb25a773),
	.w5(32'hba290f07),
	.w6(32'hbb8bf99a),
	.w7(32'hbaeb4cf7),
	.w8(32'hbb1a21d6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28f1d6),
	.w1(32'h3a7556fa),
	.w2(32'hbb9b6393),
	.w3(32'h3c2744ce),
	.w4(32'h3b4eb39c),
	.w5(32'hbb158ea1),
	.w6(32'h3c15a860),
	.w7(32'hbaeabf13),
	.w8(32'hbc1672cf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3bff2),
	.w1(32'hb98fdbb5),
	.w2(32'hbab15cd5),
	.w3(32'hbac48776),
	.w4(32'h39e44b03),
	.w5(32'hba8c47a0),
	.w6(32'hbac729df),
	.w7(32'hb8ccf55f),
	.w8(32'hba9c18ad),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c24e8),
	.w1(32'h39baace3),
	.w2(32'h3a4a6c41),
	.w3(32'hba1cf850),
	.w4(32'hb811501b),
	.w5(32'h3a68cb6d),
	.w6(32'hba073b8d),
	.w7(32'hba41fe08),
	.w8(32'h382794af),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b674097),
	.w1(32'h3b45bcb2),
	.w2(32'h3a06d27e),
	.w3(32'h3b31e8b7),
	.w4(32'h3b416cb3),
	.w5(32'h3a8fb9ae),
	.w6(32'hb904479c),
	.w7(32'hb815b6a4),
	.w8(32'hbb096096),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8137d7),
	.w1(32'hb9568612),
	.w2(32'hbb2506a1),
	.w3(32'hbaa4d2c7),
	.w4(32'h3af27be4),
	.w5(32'hbada6a1d),
	.w6(32'hbb7180e7),
	.w7(32'hbb0869e2),
	.w8(32'hbbb9abf0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6720),
	.w1(32'h3b020515),
	.w2(32'hbaa5ab96),
	.w3(32'h3acc2095),
	.w4(32'h3ad58e71),
	.w5(32'hba9f0b9f),
	.w6(32'h39827ebb),
	.w7(32'hb9f0295e),
	.w8(32'hbb5ae9c5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa98639),
	.w1(32'hb9e319ef),
	.w2(32'hba0a5ecc),
	.w3(32'hba59a96a),
	.w4(32'hba50d3ce),
	.w5(32'hb9832dc1),
	.w6(32'hbabecdd4),
	.w7(32'hba35c29b),
	.w8(32'hba7a98b4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc4dcf),
	.w1(32'hb93f2b28),
	.w2(32'hb994abfb),
	.w3(32'hb9617eab),
	.w4(32'h387bfb9f),
	.w5(32'h394b6362),
	.w6(32'hba0364a5),
	.w7(32'hb96676b4),
	.w8(32'hb984205e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65eda8),
	.w1(32'hba400670),
	.w2(32'hbb320e1d),
	.w3(32'hbb18e823),
	.w4(32'h38bc3b57),
	.w5(32'hba37e9f6),
	.w6(32'hbb731c88),
	.w7(32'hb91cbf85),
	.w8(32'hbb09fd70),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35bf32),
	.w1(32'h3802261f),
	.w2(32'hba1022a6),
	.w3(32'h39b12968),
	.w4(32'hb9bfb831),
	.w5(32'hba8c1380),
	.w6(32'h3a1edddf),
	.w7(32'hba51abc3),
	.w8(32'hba954999),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d5d1),
	.w1(32'h3ac27a4f),
	.w2(32'h380232f0),
	.w3(32'h3ab06bd9),
	.w4(32'h39b11df7),
	.w5(32'hb94cd31b),
	.w6(32'h39be7385),
	.w7(32'hba40f7a6),
	.w8(32'hbb19ccee),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39972bd7),
	.w1(32'h393e1bb4),
	.w2(32'hb8c2e4d5),
	.w3(32'h39e18822),
	.w4(32'h39a2ee88),
	.w5(32'hb9158dd3),
	.w6(32'h39c7ab31),
	.w7(32'h39bd88b4),
	.w8(32'h38a561fe),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0658f8),
	.w1(32'h3b1579ab),
	.w2(32'hbb28556f),
	.w3(32'h3ac7e1bb),
	.w4(32'h3a4823af),
	.w5(32'hbb877b28),
	.w6(32'hb98e81a0),
	.w7(32'hb8fd51ab),
	.w8(32'hbba0d932),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38042232),
	.w1(32'hb868b8ad),
	.w2(32'h38a32a5d),
	.w3(32'h37c0f7ca),
	.w4(32'hb7d508bd),
	.w5(32'h36a1f3f1),
	.w6(32'hb78dc594),
	.w7(32'hb80713d4),
	.w8(32'h381c2df7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c86835),
	.w1(32'hb838643c),
	.w2(32'hb890e2e9),
	.w3(32'hb9e3c99f),
	.w4(32'hb887d1f3),
	.w5(32'hb94965a8),
	.w6(32'hba0f30a5),
	.w7(32'hb9259058),
	.w8(32'hb9cc1245),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a05de),
	.w1(32'h3ac40d69),
	.w2(32'hbab18eb5),
	.w3(32'h3abb39b0),
	.w4(32'h3ae6fddb),
	.w5(32'h39ce86ca),
	.w6(32'hba74cb6c),
	.w7(32'hba8dfe86),
	.w8(32'hbb1f6949),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32bb90),
	.w1(32'hba4a3e9d),
	.w2(32'hbb60e14c),
	.w3(32'hbb5d89e1),
	.w4(32'hbaa9e674),
	.w5(32'hbbb84338),
	.w6(32'hbc35f1e6),
	.w7(32'hbb6eba46),
	.w8(32'hbbc1b817),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982d584),
	.w1(32'h39a3b67b),
	.w2(32'hba9779a3),
	.w3(32'hb94827ff),
	.w4(32'h3914398c),
	.w5(32'hba9744dc),
	.w6(32'hba115a1e),
	.w7(32'hb84d102e),
	.w8(32'hba95afce),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be3e38),
	.w1(32'h3a7968ea),
	.w2(32'hbb38dad9),
	.w3(32'hba0fb191),
	.w4(32'h3a366338),
	.w5(32'hbb01ef74),
	.w6(32'hbabf3499),
	.w7(32'hbabb4890),
	.w8(32'hbb72de61),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8958c),
	.w1(32'hba0bc07b),
	.w2(32'hba3ada7c),
	.w3(32'h3aa30a20),
	.w4(32'hba3c7426),
	.w5(32'hbacce97b),
	.w6(32'h3b10d3db),
	.w7(32'hba96faa2),
	.w8(32'hba88b3b9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a11e7),
	.w1(32'hb8dcea0f),
	.w2(32'hbb64989f),
	.w3(32'hbb9ca551),
	.w4(32'h3afc6652),
	.w5(32'hbb9b5a47),
	.w6(32'hbbab0b25),
	.w7(32'hb8214839),
	.w8(32'hbbb082b8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81647f),
	.w1(32'h39e0a1cb),
	.w2(32'hbb78e321),
	.w3(32'hbb0fcf50),
	.w4(32'h3ae9737a),
	.w5(32'hbaf178fb),
	.w6(32'hbb92ec3e),
	.w7(32'hbad5d743),
	.w8(32'hbb73b125),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac53e15),
	.w1(32'h3a35e87c),
	.w2(32'hbb535b81),
	.w3(32'hbb28d1a9),
	.w4(32'h3a2c38a3),
	.w5(32'hbb3c7856),
	.w6(32'hbb8bfe37),
	.w7(32'hb932a574),
	.w8(32'hbb7c7536),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932c798),
	.w1(32'h395e17c5),
	.w2(32'h3961bc86),
	.w3(32'h39b516d2),
	.w4(32'h38b7d282),
	.w5(32'h393a181c),
	.w6(32'h399c9be7),
	.w7(32'h392589c9),
	.w8(32'h3912735f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0758d),
	.w1(32'hba28b405),
	.w2(32'hbaadbfe8),
	.w3(32'hba477aac),
	.w4(32'h3a1fd0a8),
	.w5(32'hba023bda),
	.w6(32'hba22ea69),
	.w7(32'h39a63853),
	.w8(32'hb999c24d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3858861b),
	.w1(32'h36da6a34),
	.w2(32'h381753ec),
	.w3(32'h37fd0d80),
	.w4(32'hb6d9fc6b),
	.w5(32'h37d947e0),
	.w6(32'h38df347e),
	.w7(32'h3898a874),
	.w8(32'h38dd334c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff0d57),
	.w1(32'h3a883a17),
	.w2(32'h39c7a318),
	.w3(32'h397406f8),
	.w4(32'h3a5ecea1),
	.w5(32'h3a0d8402),
	.w6(32'hba844e09),
	.w7(32'hb99f2536),
	.w8(32'hba3b5dfb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a6c05e),
	.w1(32'h390cc89d),
	.w2(32'h387a253c),
	.w3(32'hb9cbb632),
	.w4(32'h39d79c6b),
	.w5(32'h393433e2),
	.w6(32'h38080f48),
	.w7(32'h3902e330),
	.w8(32'hb99cf365),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2ea9),
	.w1(32'h3952c09a),
	.w2(32'h38005325),
	.w3(32'hbb0ccc16),
	.w4(32'h3b1d2652),
	.w5(32'h3904892b),
	.w6(32'hbb9cfa92),
	.w7(32'hba81cb41),
	.w8(32'hbafce7f2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fdc446),
	.w1(32'h373108e3),
	.w2(32'h3788f59b),
	.w3(32'h36dda21d),
	.w4(32'h370a1419),
	.w5(32'h37cfebec),
	.w6(32'h38126e4e),
	.w7(32'h382f7dcf),
	.w8(32'h3836a6b5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39272f0c),
	.w1(32'h3879711c),
	.w2(32'h387f1f67),
	.w3(32'h37d4c39b),
	.w4(32'hb80eb287),
	.w5(32'h383ee2b3),
	.w6(32'h38b072c5),
	.w7(32'hb78adaa9),
	.w8(32'h37394915),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bb9c2),
	.w1(32'hb9132241),
	.w2(32'hba2c11f9),
	.w3(32'h3adec138),
	.w4(32'h3ac3d038),
	.w5(32'h3abb2747),
	.w6(32'h3a88822b),
	.w7(32'h39705692),
	.w8(32'hb92bfb63),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3cd56),
	.w1(32'hba8a38a5),
	.w2(32'hbb4f570f),
	.w3(32'hbb97386f),
	.w4(32'h3a297b14),
	.w5(32'hbb083cb1),
	.w6(32'hbb7638c5),
	.w7(32'h3a43bc38),
	.w8(32'hba9fd67d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafcb81),
	.w1(32'hbb92a301),
	.w2(32'hbb627ecb),
	.w3(32'hbb4d0b68),
	.w4(32'hbb61b5f1),
	.w5(32'h39bac5ff),
	.w6(32'hbb05006a),
	.w7(32'hbb3d4dd7),
	.w8(32'hbb3066db),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a69c47),
	.w1(32'h39c0b709),
	.w2(32'hb93020da),
	.w3(32'hb9c457b2),
	.w4(32'h398aaf87),
	.w5(32'hba12b16b),
	.w6(32'hb9c9d4a1),
	.w7(32'hb9ea5234),
	.w8(32'hba70a4f8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1758f5),
	.w1(32'h39837b80),
	.w2(32'hbb31eaa1),
	.w3(32'hbb994706),
	.w4(32'h39fbe2a5),
	.w5(32'hbb797ef1),
	.w6(32'hbbfe82c6),
	.w7(32'h3b459647),
	.w8(32'hbb102362),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7852d6),
	.w1(32'h3a9ca5a3),
	.w2(32'hbb49b107),
	.w3(32'h3b79032f),
	.w4(32'h3b8db939),
	.w5(32'h39e7483b),
	.w6(32'h3b58fc9e),
	.w7(32'hba5b277b),
	.w8(32'hbb8deecf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69dc7ea),
	.w1(32'hb9fb683a),
	.w2(32'hba75c62c),
	.w3(32'h398fcd35),
	.w4(32'hba149528),
	.w5(32'hba5e63e3),
	.w6(32'h3a3fae6d),
	.w7(32'hba7b5b65),
	.w8(32'hba5ac82f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a651c2),
	.w1(32'hb84cbccd),
	.w2(32'hb750d3bc),
	.w3(32'hb8294734),
	.w4(32'hb8024d32),
	.w5(32'hb6288165),
	.w6(32'h37ae19bb),
	.w7(32'h381f9b67),
	.w8(32'h372aeaec),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b42004),
	.w1(32'hb7ac936e),
	.w2(32'hb7a42b59),
	.w3(32'h3949cff1),
	.w4(32'hb83e2f57),
	.w5(32'h38827b5a),
	.w6(32'h38a97cd0),
	.w7(32'hb78ad194),
	.w8(32'hb7d728a8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d9e543),
	.w1(32'h37d09c8a),
	.w2(32'h38270cfe),
	.w3(32'h3773067a),
	.w4(32'h3743e305),
	.w5(32'h37b469d4),
	.w6(32'h388f7ac9),
	.w7(32'h3861b9d4),
	.w8(32'h3886e97b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915469c),
	.w1(32'hba80ec06),
	.w2(32'hbac92e91),
	.w3(32'hba1d3d37),
	.w4(32'hbad7de46),
	.w5(32'hba60412a),
	.w6(32'hbaa9f51b),
	.w7(32'hba1acfc3),
	.w8(32'hba5fc1c4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacec960),
	.w1(32'h3a46a3f8),
	.w2(32'hba708c71),
	.w3(32'hba365516),
	.w4(32'h3af1e124),
	.w5(32'h3a0da208),
	.w6(32'hbb84aa6b),
	.w7(32'hbadfd23c),
	.w8(32'hbb7e40ed),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02599d),
	.w1(32'h3aa2e657),
	.w2(32'hbb054205),
	.w3(32'hba9ec6fd),
	.w4(32'h3b62bd1e),
	.w5(32'h3acd19f5),
	.w6(32'hbb476cad),
	.w7(32'h397555a5),
	.w8(32'hbb3eeb69),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74b0fc),
	.w1(32'h3a78f3b8),
	.w2(32'hb95c5aeb),
	.w3(32'h3a9ff04c),
	.w4(32'h3a898176),
	.w5(32'hb99acc33),
	.w6(32'hba6b6005),
	.w7(32'hb9aa7967),
	.w8(32'hbace082b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7580bf),
	.w1(32'hb96e351a),
	.w2(32'hbb474cc5),
	.w3(32'hbb07a86d),
	.w4(32'h3ab0f4d5),
	.w5(32'hbacf920e),
	.w6(32'hbbbfbfd5),
	.w7(32'hba320db0),
	.w8(32'hbb79a2b4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf52046),
	.w1(32'hbae47344),
	.w2(32'hbb271fe6),
	.w3(32'hbaa2773c),
	.w4(32'hbadbb4a2),
	.w5(32'hbabac8ef),
	.w6(32'hbb0d3f2f),
	.w7(32'hba897748),
	.w8(32'hb8fd8999),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387cddeb),
	.w1(32'h37471c89),
	.w2(32'h38c4c6e4),
	.w3(32'h3886aebb),
	.w4(32'h375de2e1),
	.w5(32'h38d0503c),
	.w6(32'h38ef3704),
	.w7(32'h388f8265),
	.w8(32'h3913d885),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6aa4),
	.w1(32'hbac9b225),
	.w2(32'hbb1c8728),
	.w3(32'hb92f3a97),
	.w4(32'hba839ceb),
	.w5(32'hba6a22b2),
	.w6(32'hb9a754ee),
	.w7(32'h39885b85),
	.w8(32'h3a857453),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390acccc),
	.w1(32'h378f3844),
	.w2(32'h393c1e12),
	.w3(32'h3915bd31),
	.w4(32'h38039296),
	.w5(32'h394130b5),
	.w6(32'h398f93fc),
	.w7(32'h392cb7b5),
	.w8(32'h399bd45e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3999e),
	.w1(32'h38a71b64),
	.w2(32'hbb02f0e9),
	.w3(32'hba928184),
	.w4(32'h3a11973b),
	.w5(32'hbaff36c6),
	.w6(32'hbb665db2),
	.w7(32'hba6376d4),
	.w8(32'hbb5835cf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90c2ce),
	.w1(32'h3af2d9c1),
	.w2(32'hbb7f582b),
	.w3(32'hba0ea62e),
	.w4(32'h3b895ecb),
	.w5(32'hba91f1e8),
	.w6(32'hbb97e323),
	.w7(32'hbaaf57b2),
	.w8(32'hbbdccdb4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba654597),
	.w1(32'h3aae7ca1),
	.w2(32'hbb0f1e6a),
	.w3(32'hb97c5a63),
	.w4(32'h3b144b20),
	.w5(32'hba75927b),
	.w6(32'hbb6b3492),
	.w7(32'hbaf20a55),
	.w8(32'hbb9a9a0d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfb47e),
	.w1(32'h38ff5664),
	.w2(32'hba5cff24),
	.w3(32'h3994e27d),
	.w4(32'h395809e3),
	.w5(32'hba5338c5),
	.w6(32'hb992b131),
	.w7(32'hb9a6371a),
	.w8(32'hba8f3586),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e8ded),
	.w1(32'h399fbd44),
	.w2(32'hbb57b008),
	.w3(32'h3b0d2208),
	.w4(32'h3b66b41e),
	.w5(32'hb9559ef2),
	.w6(32'hba9323de),
	.w7(32'hbac482cf),
	.w8(32'hbbab466b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101468),
	.w1(32'hb99583c0),
	.w2(32'hbae8cee2),
	.w3(32'hbac9b5a9),
	.w4(32'h3a457b92),
	.w5(32'hb90ea954),
	.w6(32'hbb4d5495),
	.w7(32'hba132e44),
	.w8(32'hba04bd91),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9219e2),
	.w1(32'h3a9e65a7),
	.w2(32'hbab23aca),
	.w3(32'hbb0270d3),
	.w4(32'h3ae37c57),
	.w5(32'hba5afe1a),
	.w6(32'hbba6dc91),
	.w7(32'hb97740cc),
	.w8(32'hbb4ae151),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38028f42),
	.w1(32'hb681a11f),
	.w2(32'h38ae4754),
	.w3(32'h375b9634),
	.w4(32'hb801565c),
	.w5(32'h388c73f8),
	.w6(32'h3878d17c),
	.w7(32'h37b1a5d7),
	.w8(32'h38d938d3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f97976),
	.w1(32'h390e4c2f),
	.w2(32'h38c9149f),
	.w3(32'h391b8f11),
	.w4(32'hb90d0afe),
	.w5(32'hb9cc1eec),
	.w6(32'h39a62436),
	.w7(32'hb882fc2d),
	.w8(32'hb9991b24),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4d0a),
	.w1(32'hba31d8fb),
	.w2(32'hbb717a56),
	.w3(32'hba28d2ec),
	.w4(32'h3a88fa0d),
	.w5(32'hb980d8a6),
	.w6(32'hbc12ce1e),
	.w7(32'hbb064684),
	.w8(32'hbb4c6e00),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4a74),
	.w1(32'h3755275b),
	.w2(32'hbb66901d),
	.w3(32'hbb3b3e33),
	.w4(32'hb83b3737),
	.w5(32'hbba2814b),
	.w6(32'hbc1d1c09),
	.w7(32'hbb40f0fd),
	.w8(32'hbbbe9098),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb346e47),
	.w1(32'h3a6990b4),
	.w2(32'hbaf827d2),
	.w3(32'hbababf9f),
	.w4(32'h3b8205b1),
	.w5(32'h3b0d1f2c),
	.w6(32'hbbb323b1),
	.w7(32'hb8b0f47a),
	.w8(32'hbb24d5ae),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eba3a),
	.w1(32'hb9f6dbb8),
	.w2(32'h3b51b9f4),
	.w3(32'hba9fad0c),
	.w4(32'hbb2b596b),
	.w5(32'h3a290e7b),
	.w6(32'h39a688fd),
	.w7(32'hba159ec5),
	.w8(32'h39cb71f6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36584ad7),
	.w1(32'hb978ddba),
	.w2(32'hb91a3c2a),
	.w3(32'hba207a61),
	.w4(32'hb8812705),
	.w5(32'hb9f45b2c),
	.w6(32'hba466249),
	.w7(32'hb983965c),
	.w8(32'hb95640cc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30c8da),
	.w1(32'hb9b3ec03),
	.w2(32'hb9f30154),
	.w3(32'hb8243eb0),
	.w4(32'h3994b3dd),
	.w5(32'h3a1dfa69),
	.w6(32'hb990b1b9),
	.w7(32'h3a024899),
	.w8(32'h3a2bc4b3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59ef32),
	.w1(32'hbb6678cd),
	.w2(32'hbbb64578),
	.w3(32'hbb0c2134),
	.w4(32'hbbe32d64),
	.w5(32'hbb9eab3e),
	.w6(32'hbbd101bc),
	.w7(32'hbb600ff0),
	.w8(32'hbb0d1dda),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885cfd),
	.w1(32'hbabcca27),
	.w2(32'hbb309719),
	.w3(32'hbb99c60a),
	.w4(32'hba34451e),
	.w5(32'hbb47246f),
	.w6(32'hbb9ab39e),
	.w7(32'h3ab90b76),
	.w8(32'hbb1743f4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4b930),
	.w1(32'hbb6d14d1),
	.w2(32'hbad19b7a),
	.w3(32'hbb7c9d94),
	.w4(32'hbb458120),
	.w5(32'hb9e93f07),
	.w6(32'hbbd5f49b),
	.w7(32'hb8935ed6),
	.w8(32'hbade1a7f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1f0b9),
	.w1(32'h3b37f567),
	.w2(32'hba9e7fe1),
	.w3(32'h3b4f6590),
	.w4(32'h3a37fb61),
	.w5(32'hbb2aaad9),
	.w6(32'h3a65a94d),
	.w7(32'hbb11c24c),
	.w8(32'hbbc57fa2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2db359),
	.w1(32'h39200193),
	.w2(32'hbb93c026),
	.w3(32'h3ad56bd7),
	.w4(32'h3b5c8530),
	.w5(32'hbab6280a),
	.w6(32'hba932267),
	.w7(32'hbb1f9e1d),
	.w8(32'hbbdce000),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380fcb9d),
	.w1(32'h3775a670),
	.w2(32'h381e9246),
	.w3(32'h3805646e),
	.w4(32'h3781fd36),
	.w5(32'h38092ff6),
	.w6(32'h3852a1c1),
	.w7(32'h380d1a3b),
	.w8(32'h38544bb7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a41f3),
	.w1(32'h37b17b85),
	.w2(32'h3855f2f9),
	.w3(32'h384e01db),
	.w4(32'h376feaaf),
	.w5(32'h38453318),
	.w6(32'h38a4714e),
	.w7(32'h384681bd),
	.w8(32'h38a43dd1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af58666),
	.w1(32'h3ae100cf),
	.w2(32'h3ae61aaa),
	.w3(32'h3aa5c18d),
	.w4(32'h3a113e8e),
	.w5(32'h39f97963),
	.w6(32'h3a4aa8a1),
	.w7(32'h3a0dd5d7),
	.w8(32'h39a7c68f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ea3a8),
	.w1(32'hb6537dc1),
	.w2(32'h385ff6ac),
	.w3(32'h3880a781),
	.w4(32'hb4e42369),
	.w5(32'h385bc100),
	.w6(32'h38dd2e3a),
	.w7(32'h385219e9),
	.w8(32'h38ef2fd0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38348b4a),
	.w1(32'hba8824d5),
	.w2(32'hbb0b95a3),
	.w3(32'hb8ef41dc),
	.w4(32'hba9d5e4c),
	.w5(32'hbb130e23),
	.w6(32'hb8fd4dfe),
	.w7(32'hba6cc1e7),
	.w8(32'hbaab1c54),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34a3b6),
	.w1(32'hbac8399d),
	.w2(32'hba74b53e),
	.w3(32'hbb0b7cbc),
	.w4(32'h3a1b5d8d),
	.w5(32'hb9e60581),
	.w6(32'hbbdb3ba8),
	.w7(32'hba91e4ce),
	.w8(32'hbb43f85a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8725d),
	.w1(32'h3a745d48),
	.w2(32'hba57ae7a),
	.w3(32'hba775394),
	.w4(32'h3a830bf5),
	.w5(32'hba3536e4),
	.w6(32'hbb5c5570),
	.w7(32'hbaab0aa0),
	.w8(32'hbb13bb9d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3771ba0a),
	.w1(32'h3760c14e),
	.w2(32'h38410cdf),
	.w3(32'h3807741e),
	.w4(32'h380f8a7b),
	.w5(32'h3883a577),
	.w6(32'h3890705d),
	.w7(32'h38418a11),
	.w8(32'h3883bac7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc218adf),
	.w1(32'hbb777fe8),
	.w2(32'hbb9a2aec),
	.w3(32'hbbe8292c),
	.w4(32'hbb5e57ee),
	.w5(32'hbaca93c5),
	.w6(32'hbc045886),
	.w7(32'h3a8a3d16),
	.w8(32'hb9d8bcb7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad71675),
	.w1(32'h382d62a3),
	.w2(32'hb9965142),
	.w3(32'hbac20d17),
	.w4(32'h39e7e0ad),
	.w5(32'hb9de2e9b),
	.w6(32'hbb186a93),
	.w7(32'h38c69b18),
	.w8(32'hbaa731a4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c8307),
	.w1(32'h3989ead1),
	.w2(32'hb9b627f5),
	.w3(32'h39b00af5),
	.w4(32'hb805af01),
	.w5(32'hb9dd9de8),
	.w6(32'hb8dec82e),
	.w7(32'hb90771c0),
	.w8(32'hb9d18c64),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b7ee2),
	.w1(32'hba43ecce),
	.w2(32'hba934c5d),
	.w3(32'hba92c2fa),
	.w4(32'hba0d0f3c),
	.w5(32'hbabfd9f5),
	.w6(32'hbae9f197),
	.w7(32'hba21287f),
	.w8(32'hba42c252),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38852544),
	.w1(32'hb7ea37d5),
	.w2(32'hb7b4c070),
	.w3(32'h37a5e56d),
	.w4(32'hb841d0e7),
	.w5(32'h38203819),
	.w6(32'h370912ba),
	.w7(32'hb836bfdf),
	.w8(32'h37327fa5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d6528),
	.w1(32'hb9b9d29c),
	.w2(32'hb8d06919),
	.w3(32'hb79909a7),
	.w4(32'hb7b251a1),
	.w5(32'hb81199c8),
	.w6(32'hba5cbe1f),
	.w7(32'hba311b61),
	.w8(32'hb9e5238e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907c939),
	.w1(32'h3911ba40),
	.w2(32'h3924ed07),
	.w3(32'h390f4818),
	.w4(32'h390ba80d),
	.w5(32'h3910ba26),
	.w6(32'h389cb627),
	.w7(32'h38b3d745),
	.w8(32'h38f5b270),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38839770),
	.w1(32'h3637770c),
	.w2(32'hb69181da),
	.w3(32'h3754c3d9),
	.w4(32'hb769725b),
	.w5(32'hb7514d98),
	.w6(32'h3835b441),
	.w7(32'h3710896f),
	.w8(32'h38bb6104),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39906203),
	.w1(32'h3a3c31f0),
	.w2(32'hb920bf27),
	.w3(32'hbac2c446),
	.w4(32'hba826934),
	.w5(32'hba9da4bc),
	.w6(32'hbb1bf5e3),
	.w7(32'hbb0ed8a6),
	.w8(32'hbb2c1e14),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99fc85),
	.w1(32'h39771549),
	.w2(32'hbb092957),
	.w3(32'hbb287816),
	.w4(32'h3af1809e),
	.w5(32'hbb3c18cd),
	.w6(32'hbbb0df32),
	.w7(32'hbafb51a5),
	.w8(32'hbb9c7b38),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4abec),
	.w1(32'hb9f1a376),
	.w2(32'hbb627654),
	.w3(32'hbad1fa83),
	.w4(32'h3979a22c),
	.w5(32'hbb0a28a4),
	.w6(32'hbb21ee2a),
	.w7(32'h3a1648ab),
	.w8(32'hba77e383),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a03cf),
	.w1(32'hbad6ceb7),
	.w2(32'hbb180d5a),
	.w3(32'hbb45e503),
	.w4(32'hbaaa9d39),
	.w5(32'hbb135c6b),
	.w6(32'hbb6d115e),
	.w7(32'hbaee3778),
	.w8(32'hbb506de8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a29d1),
	.w1(32'h395a8848),
	.w2(32'hb8d3a1b1),
	.w3(32'h392ac13e),
	.w4(32'h39587f57),
	.w5(32'hb856dfb9),
	.w6(32'h378f0ee6),
	.w7(32'h38b6d616),
	.w8(32'hb8a63709),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988e20d),
	.w1(32'hb9328497),
	.w2(32'hb874a5af),
	.w3(32'h3935784a),
	.w4(32'h38b2496e),
	.w5(32'h39d1b9be),
	.w6(32'hb7f1dc68),
	.w7(32'h38f636d8),
	.w8(32'h395e3b4d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38162b9b),
	.w1(32'h38a34fb1),
	.w2(32'h3892ac32),
	.w3(32'h37c3fc81),
	.w4(32'h38dcfe10),
	.w5(32'h3906c8bd),
	.w6(32'h38586cbb),
	.w7(32'h387a0297),
	.w8(32'h38979ad6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39029d5d),
	.w1(32'h38b7965d),
	.w2(32'h386d368f),
	.w3(32'h386bd198),
	.w4(32'h386bfb75),
	.w5(32'h388b8c8d),
	.w6(32'h37f8aad7),
	.w7(32'h377a7d18),
	.w8(32'h382dd109),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbaf4d),
	.w1(32'hbae6ba6e),
	.w2(32'hbb15d70e),
	.w3(32'hbb6c50d9),
	.w4(32'h3ade93ea),
	.w5(32'hba42d839),
	.w6(32'hbb859409),
	.w7(32'h3a4a814b),
	.w8(32'hb9923b5a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af95e8),
	.w1(32'h3880da10),
	.w2(32'h389ed025),
	.w3(32'h3964299d),
	.w4(32'h380f1970),
	.w5(32'h389e8b83),
	.w6(32'h39618a69),
	.w7(32'h36005366),
	.w8(32'h382c73f5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd9be0),
	.w1(32'h3a4b6da0),
	.w2(32'hbaa25bf1),
	.w3(32'h39d7b5f2),
	.w4(32'h3a3935f9),
	.w5(32'hba9ee15c),
	.w6(32'hb9d61eeb),
	.w7(32'hb90971f7),
	.w8(32'hbaebe4b0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3796b),
	.w1(32'hba4273ce),
	.w2(32'hbb1d35d6),
	.w3(32'hbb199bcc),
	.w4(32'hba91d2f1),
	.w5(32'hbae9590e),
	.w6(32'hba94cc41),
	.w7(32'hb913b9da),
	.w8(32'hba6040e5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902ab32),
	.w1(32'h383c5aa1),
	.w2(32'h369909b9),
	.w3(32'h385600ca),
	.w4(32'hb8804310),
	.w5(32'hb858df34),
	.w6(32'h38a8e434),
	.w7(32'hb8053dcd),
	.w8(32'hb870ac5e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f383),
	.w1(32'hb66e74da),
	.w2(32'h384e37fd),
	.w3(32'hb9fdbfc4),
	.w4(32'h391f926d),
	.w5(32'h38b3a80a),
	.w6(32'hbaa4a778),
	.w7(32'hb9659df4),
	.w8(32'hb9f260fa),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbcf89),
	.w1(32'hb9472cb2),
	.w2(32'hb9d0163e),
	.w3(32'h38f45dd8),
	.w4(32'h394eb27b),
	.w5(32'hb9d42733),
	.w6(32'hb92886d5),
	.w7(32'hb8bcbb0f),
	.w8(32'hba0f18e2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd55acf),
	.w1(32'h38a4c62d),
	.w2(32'hbafe491a),
	.w3(32'hbb8c8a0e),
	.w4(32'h3b7f022f),
	.w5(32'hba5f26d5),
	.w6(32'hbb9930d2),
	.w7(32'h3a260601),
	.w8(32'h3656bca0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903cf60),
	.w1(32'hb6ca081b),
	.w2(32'hb8a86f37),
	.w3(32'h38c4f546),
	.w4(32'hb714df8e),
	.w5(32'hb92e8fdc),
	.w6(32'h38a24c1b),
	.w7(32'h38348c46),
	.w8(32'hb8987d01),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b5aae),
	.w1(32'h3b23082b),
	.w2(32'h3996bf77),
	.w3(32'hba5a98f3),
	.w4(32'h3a5af308),
	.w5(32'h3a0c80fa),
	.w6(32'hbbd892f1),
	.w7(32'h382ebd88),
	.w8(32'h39ea0707),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule