module layer_8_featuremap_113(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c1b1),
	.w1(32'h3b0ea2dc),
	.w2(32'h3be4d1ba),
	.w3(32'hbae80eeb),
	.w4(32'hbb8ed05d),
	.w5(32'hbb443578),
	.w6(32'hbb0d0e21),
	.w7(32'hbb8c6546),
	.w8(32'hbb1fb8da),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afec6c2),
	.w1(32'h3aad1fc5),
	.w2(32'h3b13270d),
	.w3(32'h3b0ffbac),
	.w4(32'h3ac43081),
	.w5(32'h3afa195d),
	.w6(32'h3b2ff97d),
	.w7(32'h3b2288ac),
	.w8(32'h3b2cc46a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb472390),
	.w1(32'hbaf2548b),
	.w2(32'hbadb548c),
	.w3(32'hba62d521),
	.w4(32'h3a495c83),
	.w5(32'h3a8d2a14),
	.w6(32'h3ad4cbb5),
	.w7(32'h3add53fb),
	.w8(32'h3ad9a5ff),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be210fd),
	.w1(32'h3c7b8a1c),
	.w2(32'h3c568b2b),
	.w3(32'h3bf6ed48),
	.w4(32'h3bed4170),
	.w5(32'h3c4fe5d6),
	.w6(32'h3b9dd717),
	.w7(32'h3affcfce),
	.w8(32'h3c071c15),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4391b2),
	.w1(32'h3b351f89),
	.w2(32'h3a86c2f3),
	.w3(32'hb9bb6b2e),
	.w4(32'hba4e57c3),
	.w5(32'hba85eb15),
	.w6(32'hbad9c6eb),
	.w7(32'hbb2516b3),
	.w8(32'hbb0e5a14),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9df473),
	.w1(32'hbb15738d),
	.w2(32'hbbcc21f4),
	.w3(32'hbb38c903),
	.w4(32'hbb4517c9),
	.w5(32'h3ba54788),
	.w6(32'hbab59d9b),
	.w7(32'h3a1f1fee),
	.w8(32'h3b809435),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ca81f),
	.w1(32'h380e88d6),
	.w2(32'h37575666),
	.w3(32'hb8197253),
	.w4(32'hb8bc90f6),
	.w5(32'hb7c6d966),
	.w6(32'hb8b88c89),
	.w7(32'hb8e69d8a),
	.w8(32'hb547b850),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ba583),
	.w1(32'h3afde63d),
	.w2(32'h3bffa58a),
	.w3(32'h3bb3854e),
	.w4(32'h3bbf50b0),
	.w5(32'h3bedeb8d),
	.w6(32'h3adda671),
	.w7(32'h3afd5d94),
	.w8(32'h3b1dcf01),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a094a),
	.w1(32'h3b6d84f1),
	.w2(32'h3b6b5422),
	.w3(32'h3a1963b1),
	.w4(32'hbac099c8),
	.w5(32'hbae21e94),
	.w6(32'h3b7f6bb2),
	.w7(32'h3b259b06),
	.w8(32'h3a8114b9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f814),
	.w1(32'h3c02dc86),
	.w2(32'h3c7b7ae2),
	.w3(32'h3bb2a9bf),
	.w4(32'h3b8a93b8),
	.w5(32'h3b3ee4b4),
	.w6(32'h3a8171c7),
	.w7(32'h3b2a7c0d),
	.w8(32'h3bd826be),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430f6f),
	.w1(32'h3b810cbc),
	.w2(32'h3bb287e2),
	.w3(32'hbb557c76),
	.w4(32'hba91d17b),
	.w5(32'h3b87742d),
	.w6(32'hbab01c2d),
	.w7(32'hbbaeb4fe),
	.w8(32'hbb020a28),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa051b),
	.w1(32'h3c176e66),
	.w2(32'h3c800ee2),
	.w3(32'h3bfeec1c),
	.w4(32'h3a11b41f),
	.w5(32'h3ba057eb),
	.w6(32'h3ae28eed),
	.w7(32'h3abfeaaf),
	.w8(32'h3b243555),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcd178),
	.w1(32'h39ac9123),
	.w2(32'h3b52104e),
	.w3(32'h399fd59c),
	.w4(32'h3ab75d7f),
	.w5(32'h3b528fc7),
	.w6(32'h3b5d0f4f),
	.w7(32'h3b0a52dc),
	.w8(32'h3c20974a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01b922),
	.w1(32'h3b5416db),
	.w2(32'h3982fe99),
	.w3(32'h3adae17a),
	.w4(32'hbbbad7af),
	.w5(32'h3b3f4ea1),
	.w6(32'h3b3d2608),
	.w7(32'hbbe791ed),
	.w8(32'hba9be00a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f43a9),
	.w1(32'h3b55162b),
	.w2(32'hba739b6d),
	.w3(32'hb9f6c566),
	.w4(32'hbbd08108),
	.w5(32'h3ab81a85),
	.w6(32'h3b54f573),
	.w7(32'hbbf76924),
	.w8(32'hb6be3fc0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bc3ee),
	.w1(32'h3bb61e64),
	.w2(32'hba76e7bb),
	.w3(32'h3b865ac4),
	.w4(32'h3b73b45c),
	.w5(32'hbb08504e),
	.w6(32'h3bb89930),
	.w7(32'h3b609822),
	.w8(32'hbbfe9ae8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc184898),
	.w1(32'hbb16c4fa),
	.w2(32'hbc1836e9),
	.w3(32'h3b9cf53c),
	.w4(32'h3b386268),
	.w5(32'hbc55a751),
	.w6(32'hba66a2ea),
	.w7(32'h3b1f5755),
	.w8(32'hba1b1877),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39c820),
	.w1(32'h3c63fc75),
	.w2(32'h3c6d7bdc),
	.w3(32'h3aa67f35),
	.w4(32'hbc067a52),
	.w5(32'h3c77f156),
	.w6(32'h3bbd87c2),
	.w7(32'hbca05447),
	.w8(32'h3bce4db7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd699d0),
	.w1(32'h3c873719),
	.w2(32'h3d6dedbe),
	.w3(32'h3b48e036),
	.w4(32'hba9b8b79),
	.w5(32'h3c04e5e5),
	.w6(32'hbcb3835c),
	.w7(32'hbbf8939f),
	.w8(32'hbbf83efc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91b327),
	.w1(32'h3b622673),
	.w2(32'h3c02baa8),
	.w3(32'hbc040a89),
	.w4(32'hba98caf4),
	.w5(32'hbc1f5af3),
	.w6(32'hbce46927),
	.w7(32'hbbbb1b74),
	.w8(32'hbc3ec646),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db945e),
	.w1(32'hbbca2a9e),
	.w2(32'h3cc0acb3),
	.w3(32'h3ba9f16a),
	.w4(32'hba95e0a3),
	.w5(32'hbceacc27),
	.w6(32'h3b2a1e79),
	.w7(32'h3cde4ade),
	.w8(32'hbd65d515),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf61d27),
	.w1(32'h3bb119bc),
	.w2(32'hbc647e36),
	.w3(32'h3b02cff9),
	.w4(32'hbbe6ac61),
	.w5(32'hbc187a90),
	.w6(32'h3c0831a3),
	.w7(32'hbbe682bd),
	.w8(32'hbc8b3dfb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c0ef0),
	.w1(32'h3c3726d5),
	.w2(32'h3ce5841c),
	.w3(32'hbc2f46a4),
	.w4(32'hbc6dd761),
	.w5(32'h3c640dbf),
	.w6(32'hbb4782f7),
	.w7(32'hbc2a3f3a),
	.w8(32'h3c1c77d6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ed860),
	.w1(32'h3b5812a0),
	.w2(32'h3b6d68f8),
	.w3(32'h3c13470c),
	.w4(32'h3b613b93),
	.w5(32'hbc4685dc),
	.w6(32'h3c0444f2),
	.w7(32'hb8cf0d84),
	.w8(32'hbb499e2e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e7db),
	.w1(32'h3b953026),
	.w2(32'h3c17296b),
	.w3(32'h3b94b074),
	.w4(32'hbb4eccaa),
	.w5(32'hb5e7106a),
	.w6(32'h3c107eb4),
	.w7(32'h3a85ba19),
	.w8(32'hbbbf2acb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcc246),
	.w1(32'h3bc93809),
	.w2(32'h3ceed9a1),
	.w3(32'h3be59d0d),
	.w4(32'h3c833d15),
	.w5(32'hbd1a4e38),
	.w6(32'hbb3a8422),
	.w7(32'h3c84ead9),
	.w8(32'hbd7c9260),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c5274),
	.w1(32'h3ca3da2f),
	.w2(32'h3a3d95b7),
	.w3(32'h3c9017dc),
	.w4(32'h3a673301),
	.w5(32'hbb7ad5fe),
	.w6(32'h3c8f0e93),
	.w7(32'hbb3f852c),
	.w8(32'hbbbfa33c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf2e73f),
	.w1(32'hbd40bcb7),
	.w2(32'h3d80d7d1),
	.w3(32'h3c3b518a),
	.w4(32'hbcc3c892),
	.w5(32'hbd014cce),
	.w6(32'h3c9bd5ff),
	.w7(32'hbbdda5b1),
	.w8(32'hbd186043),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4aaa5b),
	.w1(32'h3c486f1d),
	.w2(32'h3c283c44),
	.w3(32'h3c2b2c64),
	.w4(32'hb8dd91c2),
	.w5(32'h3bb125e0),
	.w6(32'h3bd4315a),
	.w7(32'hbbaaf9f9),
	.w8(32'hbc300a38),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc698399),
	.w1(32'hbaa543b3),
	.w2(32'h3ca022b2),
	.w3(32'h3c465baf),
	.w4(32'h3a642374),
	.w5(32'h3c8d8efe),
	.w6(32'h3c476ac1),
	.w7(32'h3ae6aa8f),
	.w8(32'hbcb3c8f0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1958c5),
	.w1(32'h3ba5d9f9),
	.w2(32'h3b938de4),
	.w3(32'h391a42ac),
	.w4(32'h3a090085),
	.w5(32'h3bba8a92),
	.w6(32'h3ce5c7eb),
	.w7(32'h3b85c76f),
	.w8(32'h3c17f09d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14767f),
	.w1(32'h3be76d5a),
	.w2(32'hbb0fe1fa),
	.w3(32'h3c0d402e),
	.w4(32'hbb3fa43e),
	.w5(32'hbadc464a),
	.w6(32'h3c187880),
	.w7(32'hb920add4),
	.w8(32'hba53cf11),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d3d1),
	.w1(32'hbb5f181d),
	.w2(32'hbbc13ac0),
	.w3(32'hbbc26d34),
	.w4(32'h3bd14717),
	.w5(32'h3b8ee903),
	.w6(32'hbb558aca),
	.w7(32'hbc25da88),
	.w8(32'h3c614c77),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfbc7e),
	.w1(32'hbb95f80c),
	.w2(32'hbc05372d),
	.w3(32'hbc5cf9bb),
	.w4(32'hba9d040f),
	.w5(32'h3be37196),
	.w6(32'hbbc79665),
	.w7(32'hbc5d35aa),
	.w8(32'hba9476ee),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7cdbdf),
	.w1(32'hbbc0bb05),
	.w2(32'h39f4465e),
	.w3(32'hbb16f5e2),
	.w4(32'h3b2f1f05),
	.w5(32'hbc36efef),
	.w6(32'h3bd532fb),
	.w7(32'h3c0baf36),
	.w8(32'hbc20b5d2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82dba3),
	.w1(32'hbbb0ac56),
	.w2(32'h3c9d384d),
	.w3(32'h3a4efe83),
	.w4(32'hbc29657b),
	.w5(32'h3d11aa91),
	.w6(32'hbb637463),
	.w7(32'hbb91484d),
	.w8(32'h3c1fd946),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e8201),
	.w1(32'hbca26744),
	.w2(32'h3bfbb260),
	.w3(32'hbc34a8e5),
	.w4(32'hbbfdebf6),
	.w5(32'hbae42f14),
	.w6(32'hbca7d220),
	.w7(32'hba805dbc),
	.w8(32'hbbdad19e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009eac),
	.w1(32'h3bd1027d),
	.w2(32'hbbc39c15),
	.w3(32'hba0c20f4),
	.w4(32'hbc0883b4),
	.w5(32'h3cb28880),
	.w6(32'h3b7367b9),
	.w7(32'hbb8ec17e),
	.w8(32'h3d38d6fd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d7ccd),
	.w1(32'hbbb3a55c),
	.w2(32'hbb7f4e69),
	.w3(32'h3b41b131),
	.w4(32'hbc25983d),
	.w5(32'hbb7a4538),
	.w6(32'h3beb40f4),
	.w7(32'hbafbf5c7),
	.w8(32'hbc91b5e5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e6f5),
	.w1(32'h3b52edd5),
	.w2(32'hbbb29c63),
	.w3(32'h3afc884d),
	.w4(32'hbb66842a),
	.w5(32'hbb3394ea),
	.w6(32'h39d4ba05),
	.w7(32'hba70b183),
	.w8(32'hba33490c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad57eb),
	.w1(32'h3cd18179),
	.w2(32'h3cdccd3d),
	.w3(32'h3c769a60),
	.w4(32'h3ca84216),
	.w5(32'h3cbd0bad),
	.w6(32'h3b29af43),
	.w7(32'hbb48e965),
	.w8(32'h3c5bbbd5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03b924),
	.w1(32'h3bca23c5),
	.w2(32'h3c51d814),
	.w3(32'hbba0879b),
	.w4(32'h399755da),
	.w5(32'hbb2e2036),
	.w6(32'h3c3c1af4),
	.w7(32'h3c51244d),
	.w8(32'hbc58c442),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac23d2),
	.w1(32'hba622cf2),
	.w2(32'hbc6eb263),
	.w3(32'hba02a013),
	.w4(32'hbc22fd24),
	.w5(32'h3c7f7f85),
	.w6(32'h3b70931e),
	.w7(32'hbbff5bf1),
	.w8(32'h3d17ea08),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8f06b),
	.w1(32'hbbe5f4d0),
	.w2(32'h3be0be4e),
	.w3(32'hbca842ef),
	.w4(32'hb92b9b1d),
	.w5(32'h3be68adb),
	.w6(32'hbc6ead09),
	.w7(32'hbbbc0be6),
	.w8(32'h3b635d6b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83dd3a0),
	.w1(32'h3c489bf3),
	.w2(32'h3cd36638),
	.w3(32'h3b1573aa),
	.w4(32'h3c244677),
	.w5(32'h3ba6985e),
	.w6(32'h3b1b4157),
	.w7(32'h3baa1d48),
	.w8(32'hbccde068),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97b727),
	.w1(32'h3b897d01),
	.w2(32'hbc49ec82),
	.w3(32'h3b0075da),
	.w4(32'hbc129dfb),
	.w5(32'h3d05ee33),
	.w6(32'hba14085a),
	.w7(32'hbccfa1de),
	.w8(32'h3d86d3c2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5eb97),
	.w1(32'hbc05e515),
	.w2(32'hbaedc6a1),
	.w3(32'hbc8bc97c),
	.w4(32'h3b800cd2),
	.w5(32'hbbf534df),
	.w6(32'hbca0cd2a),
	.w7(32'h3a9af15a),
	.w8(32'hbc1be0eb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc864372),
	.w1(32'hbc44ce0b),
	.w2(32'h3cc3715b),
	.w3(32'hba95f83b),
	.w4(32'h3ae5abde),
	.w5(32'h3ba14890),
	.w6(32'hbc2118ba),
	.w7(32'hbba4d2a6),
	.w8(32'hbbf7b8cc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7c512),
	.w1(32'hbc9e35d7),
	.w2(32'h3bc95ec0),
	.w3(32'hbc4276dd),
	.w4(32'hbb8ba8b0),
	.w5(32'hbc164810),
	.w6(32'hbca05432),
	.w7(32'hbbcb257e),
	.w8(32'hbca58baa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7876cd),
	.w1(32'h3c0ed8dd),
	.w2(32'hba9988ba),
	.w3(32'h3c84b5c5),
	.w4(32'hbc80f72a),
	.w5(32'h388deb33),
	.w6(32'h3bba4ce2),
	.w7(32'hbc8680ea),
	.w8(32'hbbabc2e0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48fba),
	.w1(32'hbbb703d1),
	.w2(32'h3c758b90),
	.w3(32'hbbca7ab3),
	.w4(32'h3c205ef9),
	.w5(32'hbb26e552),
	.w6(32'hbba30058),
	.w7(32'h3bcf26df),
	.w8(32'h3d193a7e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7dda8),
	.w1(32'h3bb18824),
	.w2(32'h3cb79a08),
	.w3(32'h3c440f8c),
	.w4(32'h3d18bc70),
	.w5(32'h3c636bff),
	.w6(32'h3b71d8ea),
	.w7(32'h3be2a9d1),
	.w8(32'hba9da6f1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd12e7),
	.w1(32'h3cec3ff5),
	.w2(32'hbc0108e1),
	.w3(32'h3ac1a048),
	.w4(32'h3cae26a3),
	.w5(32'h3a6c471f),
	.w6(32'h3bb87760),
	.w7(32'h3b3ec8eb),
	.w8(32'h3b00fab7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc139dab),
	.w1(32'h3c593f31),
	.w2(32'h3c91b425),
	.w3(32'hbc71ba9d),
	.w4(32'h3ab13421),
	.w5(32'h3a87614b),
	.w6(32'h3baeedaf),
	.w7(32'h3b5dcb55),
	.w8(32'h3c1cd302),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f0356),
	.w1(32'h3aebee06),
	.w2(32'h3abe6aac),
	.w3(32'h39eeb990),
	.w4(32'h3b48cb19),
	.w5(32'hbb33d70a),
	.w6(32'h3af3b7a7),
	.w7(32'h3c3912d2),
	.w8(32'hbc425644),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b620),
	.w1(32'h3c9c03f5),
	.w2(32'h3d0eeaed),
	.w3(32'h3c3dec3d),
	.w4(32'h3b2b70aa),
	.w5(32'h3c1b5b7a),
	.w6(32'h3c28d0cf),
	.w7(32'h3c900696),
	.w8(32'h3d0cfa5c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88aeaa),
	.w1(32'hbb5ce9ca),
	.w2(32'h3adf4302),
	.w3(32'hbbf7b052),
	.w4(32'hba3be45a),
	.w5(32'h3b71ef9f),
	.w6(32'hbbafbcd3),
	.w7(32'hba80d089),
	.w8(32'h3be289e7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c3ea6),
	.w1(32'h3bc0d007),
	.w2(32'h3bd56207),
	.w3(32'h3bc26403),
	.w4(32'hbbae71d3),
	.w5(32'hbc15acc5),
	.w6(32'h3c46175d),
	.w7(32'hbaaa98d0),
	.w8(32'hbb1241b9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc214006),
	.w1(32'hbb863d42),
	.w2(32'h3b36ddaa),
	.w3(32'hbbb3ab4d),
	.w4(32'hbb8d5f46),
	.w5(32'h3b21ae79),
	.w6(32'hbc0b17f8),
	.w7(32'hbbe8face),
	.w8(32'h3aa1be14),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fc1ae),
	.w1(32'h3c7df883),
	.w2(32'h3bad8cac),
	.w3(32'h3b872d91),
	.w4(32'h3c9803a2),
	.w5(32'hbc9e8e35),
	.w6(32'h3c21ba9c),
	.w7(32'h3c92e1f5),
	.w8(32'h3be7c947),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c800b79),
	.w1(32'h39a834f8),
	.w2(32'hb9bfb520),
	.w3(32'h3c0ea730),
	.w4(32'hbc459369),
	.w5(32'h3d13bc62),
	.w6(32'hbca6f676),
	.w7(32'h3b070858),
	.w8(32'h3d1598a5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1a8f),
	.w1(32'h3c252f89),
	.w2(32'h3b8a21e3),
	.w3(32'hbc70ab79),
	.w4(32'hba1cc2cd),
	.w5(32'h3a2c3b28),
	.w6(32'hbb14c83d),
	.w7(32'h3a03010f),
	.w8(32'hbb01a542),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40e1c4),
	.w1(32'h3cf76dc6),
	.w2(32'h3cf16e52),
	.w3(32'h3cb67acc),
	.w4(32'h3ccf6dbf),
	.w5(32'h3c0161bf),
	.w6(32'h3b7927e1),
	.w7(32'h3b9e5f5d),
	.w8(32'hbb43b640),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7b565),
	.w1(32'h3bfa64ca),
	.w2(32'hbb4797e4),
	.w3(32'h3b89815d),
	.w4(32'h3b87175b),
	.w5(32'h3bf747ac),
	.w6(32'h3c55fe9f),
	.w7(32'h3ba8314b),
	.w8(32'h3c0fe0da),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff18b),
	.w1(32'h3c059633),
	.w2(32'h3c254d1d),
	.w3(32'h3ba3d8da),
	.w4(32'h3ba02336),
	.w5(32'h3aee7f38),
	.w6(32'h3c3feefc),
	.w7(32'h3c4e98ef),
	.w8(32'h3ae44c2d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0778ac),
	.w1(32'hba3bc363),
	.w2(32'hbba5fdb8),
	.w3(32'h3bb88fe7),
	.w4(32'hbc4db445),
	.w5(32'hbabd1fa9),
	.w6(32'h3bddfdcc),
	.w7(32'hbc31020f),
	.w8(32'h3bc7943c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd95fb3),
	.w1(32'h3baf9404),
	.w2(32'hbb76a124),
	.w3(32'hbb93f352),
	.w4(32'h3b181f9a),
	.w5(32'h3b9efc40),
	.w6(32'h3ac7abd3),
	.w7(32'hbbc0b168),
	.w8(32'h3ac47ba9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb3252),
	.w1(32'h3c8f1187),
	.w2(32'hb91c0ca4),
	.w3(32'h3c7a5a78),
	.w4(32'h3c5bd4f8),
	.w5(32'h3c0441e4),
	.w6(32'h3bd83ddc),
	.w7(32'hbbb5080e),
	.w8(32'hba37485e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffed2e),
	.w1(32'h3c56f30c),
	.w2(32'hbbefb88e),
	.w3(32'hbc59b435),
	.w4(32'hbab73e5c),
	.w5(32'hbc63ffbc),
	.w6(32'h3aa69dd7),
	.w7(32'hbab114f6),
	.w8(32'hbc971d38),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb1545),
	.w1(32'hbc882858),
	.w2(32'h3b920a89),
	.w3(32'h39e38444),
	.w4(32'hbc48f90f),
	.w5(32'h3b55c294),
	.w6(32'hbba2b339),
	.w7(32'hba9f84bc),
	.w8(32'h3b9a8e67),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8302c5),
	.w1(32'h3c318056),
	.w2(32'hbc0a9ec2),
	.w3(32'hbc4bb221),
	.w4(32'hbba75b71),
	.w5(32'hbbf390dc),
	.w6(32'hbc587824),
	.w7(32'hbc63027d),
	.w8(32'hbc050ce7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf34db),
	.w1(32'hbb253639),
	.w2(32'hbb9ff38b),
	.w3(32'hbc1f7a9b),
	.w4(32'hbcb215f7),
	.w5(32'h3c64718f),
	.w6(32'hbbf298a8),
	.w7(32'hbca4ace5),
	.w8(32'h3c204d23),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b6e5c),
	.w1(32'hbc84d241),
	.w2(32'h3a4d3c87),
	.w3(32'h3ab2bef3),
	.w4(32'hbbae1915),
	.w5(32'hbbe3da07),
	.w6(32'hbc5387ca),
	.w7(32'hbc072aba),
	.w8(32'hbb95f34b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53102f),
	.w1(32'h3ca88029),
	.w2(32'h3c83c17a),
	.w3(32'h3c8898ec),
	.w4(32'h3cbbd5f2),
	.w5(32'hbc4d2030),
	.w6(32'h3c3b3403),
	.w7(32'h3b6bc7ab),
	.w8(32'h3c251148),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89bfd8),
	.w1(32'hbc6ae3a6),
	.w2(32'hbb0b6819),
	.w3(32'h3c0a247d),
	.w4(32'hbba022c2),
	.w5(32'hbbe7185e),
	.w6(32'h3afa3c9d),
	.w7(32'h3ba90e59),
	.w8(32'hbbc03f15),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eeb65),
	.w1(32'hba52dd1c),
	.w2(32'h3c4ae850),
	.w3(32'hbb27267f),
	.w4(32'hbcac0d68),
	.w5(32'hb8add9ac),
	.w6(32'h3b410d87),
	.w7(32'hba7bbbed),
	.w8(32'h3c7ffc6e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01ab2a),
	.w1(32'h3c17dcfc),
	.w2(32'hb9851ce1),
	.w3(32'hbc7b86a8),
	.w4(32'h3a0c572c),
	.w5(32'hb93aa678),
	.w6(32'hbbc75eb8),
	.w7(32'h3b0fedac),
	.w8(32'h3a6977f7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801a71),
	.w1(32'h3af0df60),
	.w2(32'h3c1520cc),
	.w3(32'h3a6ca19a),
	.w4(32'hb8b462f1),
	.w5(32'h3b4124b1),
	.w6(32'hbb8c3f4e),
	.w7(32'hbc1426d0),
	.w8(32'hbbd810f7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba299ff4),
	.w1(32'h3bad73c8),
	.w2(32'h3c92587d),
	.w3(32'h3bf678f7),
	.w4(32'h3bbdaafd),
	.w5(32'h3bd7c3cb),
	.w6(32'h39efcb1f),
	.w7(32'h3b1d0e15),
	.w8(32'h3b8eff2a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f303d),
	.w1(32'hbb33d3a5),
	.w2(32'hb92e3423),
	.w3(32'hbac84df0),
	.w4(32'hbb289335),
	.w5(32'hbba59ad3),
	.w6(32'hbb5aac1a),
	.w7(32'h3b947961),
	.w8(32'h3b06047a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3c795),
	.w1(32'h3a87d881),
	.w2(32'h39adaada),
	.w3(32'hbbdba54e),
	.w4(32'hbb5a6ded),
	.w5(32'hb8a8bf4e),
	.w6(32'hbaeb3d40),
	.w7(32'hbbcbecc8),
	.w8(32'hbb6237ba),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a2b74),
	.w1(32'h3a17d039),
	.w2(32'hbb52bcc0),
	.w3(32'hbba6a3ea),
	.w4(32'hbb77b2ed),
	.w5(32'h3b23c7cf),
	.w6(32'h3b155e06),
	.w7(32'h3a634549),
	.w8(32'hbacffe01),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16c8db),
	.w1(32'h3a8d8fee),
	.w2(32'h3c782263),
	.w3(32'h3b62734b),
	.w4(32'h3b0b1969),
	.w5(32'h3b604cec),
	.w6(32'hbbfbf1cc),
	.w7(32'hbc103a4a),
	.w8(32'hbba570ad),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d56caa0),
	.w1(32'h3d65d14b),
	.w2(32'h3d4f444f),
	.w3(32'h3ce0e7bb),
	.w4(32'h3d1aa3db),
	.w5(32'h3d3ba6be),
	.w6(32'hbaef076f),
	.w7(32'hbb781471),
	.w8(32'h3cc11240),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d2dec),
	.w1(32'h3c7aec56),
	.w2(32'h3cdf206b),
	.w3(32'h3c8a3d15),
	.w4(32'h3bc68a1e),
	.w5(32'h3be363c2),
	.w6(32'h3b647b0a),
	.w7(32'h3b541e56),
	.w8(32'h3c29722d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a0802),
	.w1(32'h3c70b0db),
	.w2(32'h3c91ddf6),
	.w3(32'hbc35c3d1),
	.w4(32'h3c183792),
	.w5(32'h3c6f6aab),
	.w6(32'hb90a8a70),
	.w7(32'h3b1435b8),
	.w8(32'h3ba929ff),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea38e5),
	.w1(32'h3bb6b021),
	.w2(32'hbba8bdd9),
	.w3(32'h3b50cd9d),
	.w4(32'hb8e14fc8),
	.w5(32'h3ad10ad2),
	.w6(32'h3a9172ff),
	.w7(32'hbb9c462a),
	.w8(32'hbb25cf96),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e5606),
	.w1(32'h398c6e62),
	.w2(32'h3a9a2350),
	.w3(32'hba82ca9e),
	.w4(32'hb96a2d4b),
	.w5(32'hba5acb73),
	.w6(32'hbb4f07d4),
	.w7(32'h3a785f0c),
	.w8(32'hba83cfd6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4613af),
	.w1(32'h3a27d8d3),
	.w2(32'hba7e300d),
	.w3(32'h39986c59),
	.w4(32'hba3a59c7),
	.w5(32'hba12c8f2),
	.w6(32'hb9fdf5f9),
	.w7(32'h3acadb8b),
	.w8(32'h39dae378),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b4d6),
	.w1(32'h3b0e977f),
	.w2(32'h3b83c94f),
	.w3(32'hbb1fd2e9),
	.w4(32'h3b3f5aa1),
	.w5(32'h3a76b463),
	.w6(32'hbb6856ff),
	.w7(32'hbc03def8),
	.w8(32'hbc0afa9a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3658),
	.w1(32'h3b532026),
	.w2(32'h3b5cdd33),
	.w3(32'h3bfb831b),
	.w4(32'h3b9e046c),
	.w5(32'h3b91be3b),
	.w6(32'hbaec82cb),
	.w7(32'h3bb9bab5),
	.w8(32'h3b80198f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc3788),
	.w1(32'hbb57fd1a),
	.w2(32'h3b96cceb),
	.w3(32'hbbb0e6df),
	.w4(32'h3b632f09),
	.w5(32'h3bb896d6),
	.w6(32'hba4349b4),
	.w7(32'hbbb86f9b),
	.w8(32'hbbeda65a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb2438),
	.w1(32'h3b6e4c1c),
	.w2(32'h3a811123),
	.w3(32'h3c01e37c),
	.w4(32'h3c130713),
	.w5(32'hbb89b8fb),
	.w6(32'hbae9b07f),
	.w7(32'h3b03322c),
	.w8(32'h3b39e72b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b34e9),
	.w1(32'h3bfcc422),
	.w2(32'h3b8deaea),
	.w3(32'h3bd3a37a),
	.w4(32'h3c0c4b70),
	.w5(32'h3c4adfcd),
	.w6(32'h3b0f35bc),
	.w7(32'hbae7eff6),
	.w8(32'h3a5cdae0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eabff),
	.w1(32'hbad3536d),
	.w2(32'h3b905ef0),
	.w3(32'h3afd40ab),
	.w4(32'h38e95c49),
	.w5(32'h3af35b9e),
	.w6(32'h3c104458),
	.w7(32'h3ab63314),
	.w8(32'h3b869937),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ff680),
	.w1(32'h3a272ce4),
	.w2(32'h3c2e2d71),
	.w3(32'hbaada2e3),
	.w4(32'h3b87559f),
	.w5(32'h3b546307),
	.w6(32'hbb96b360),
	.w7(32'h3c3f3bca),
	.w8(32'h3c5e08bf),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b506095),
	.w1(32'h3c80adcd),
	.w2(32'h3b9035d0),
	.w3(32'h3b0b7939),
	.w4(32'hbbb98c5d),
	.w5(32'hbc0a0b7e),
	.w6(32'h3bd02cde),
	.w7(32'hbc317094),
	.w8(32'hbbe55bb6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba556cc9),
	.w1(32'h3accc6b8),
	.w2(32'hb989d21a),
	.w3(32'hbc0902af),
	.w4(32'hbb2fc015),
	.w5(32'hbba2a895),
	.w6(32'hbb9a5165),
	.w7(32'hbb208f7d),
	.w8(32'hbb807f2f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c021f),
	.w1(32'hbb75ed46),
	.w2(32'h3bdda00e),
	.w3(32'hbb4843c1),
	.w4(32'h3ba4abbf),
	.w5(32'h3b9f4372),
	.w6(32'hbb9ee694),
	.w7(32'h3b614803),
	.w8(32'h3a38b9b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c0778),
	.w1(32'h3b40477a),
	.w2(32'hb995306e),
	.w3(32'h3b70b039),
	.w4(32'h3ac79c1b),
	.w5(32'h3b21e643),
	.w6(32'h3abe27ab),
	.w7(32'hba9fb117),
	.w8(32'h37a01397),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb6de1),
	.w1(32'h3af8bb61),
	.w2(32'h3be658f4),
	.w3(32'h39948b51),
	.w4(32'h3c051d66),
	.w5(32'h3c0180b2),
	.w6(32'h3ab8043f),
	.w7(32'h3c647915),
	.w8(32'h3c557598),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc9106),
	.w1(32'h3c2d6af2),
	.w2(32'hba60bc20),
	.w3(32'h3bd907c9),
	.w4(32'h3a2c827b),
	.w5(32'hbb540189),
	.w6(32'h3c0f4552),
	.w7(32'hbb501805),
	.w8(32'hbbb0c502),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55539f),
	.w1(32'hbb32c425),
	.w2(32'h3b8002ba),
	.w3(32'hbb8836bb),
	.w4(32'h3b858146),
	.w5(32'hbb1ad3f7),
	.w6(32'hbc02859c),
	.w7(32'h3bd6206a),
	.w8(32'h3c415ccc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d5663),
	.w1(32'h3bd4a05d),
	.w2(32'hbb327cb5),
	.w3(32'hbbb3d29b),
	.w4(32'h39e9d87e),
	.w5(32'h39af48de),
	.w6(32'h3c2859f7),
	.w7(32'h3aa5e860),
	.w8(32'h3b613bee),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a238673),
	.w1(32'h3ab16eb1),
	.w2(32'hbba8c75b),
	.w3(32'hba99cf67),
	.w4(32'hbb0e8066),
	.w5(32'hbb6be7ed),
	.w6(32'h39d72cbc),
	.w7(32'h3c0ed29a),
	.w8(32'h3b968acc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c259),
	.w1(32'hbb425edb),
	.w2(32'h3bfcdac3),
	.w3(32'hbb0b5dd6),
	.w4(32'h3af4ebda),
	.w5(32'h3be43bed),
	.w6(32'h3b572ffa),
	.w7(32'h3b0af6c9),
	.w8(32'hba530466),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84f87a),
	.w1(32'h395797f5),
	.w2(32'h3b38add3),
	.w3(32'hbb7dfa70),
	.w4(32'hbb720f1e),
	.w5(32'hbc274e98),
	.w6(32'hbb55b518),
	.w7(32'hbc3178bc),
	.w8(32'hbc5994f6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf94f04),
	.w1(32'h3a737ae6),
	.w2(32'hbb46c25e),
	.w3(32'hbbb724b3),
	.w4(32'h3a3ccd95),
	.w5(32'hba4a1348),
	.w6(32'hbc461033),
	.w7(32'h3b7070c7),
	.w8(32'h3a9cb4de),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb130e5a),
	.w1(32'hbb48c01f),
	.w2(32'hbb7b3509),
	.w3(32'h3a410fd6),
	.w4(32'h3b446a90),
	.w5(32'hbb14ebab),
	.w6(32'h3b1712b4),
	.w7(32'h3b14e4f2),
	.w8(32'h3c0b8381),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00aefb),
	.w1(32'h3c01c4d6),
	.w2(32'h3b9da80a),
	.w3(32'hbb8fecd6),
	.w4(32'hbb00ea02),
	.w5(32'h3b65130d),
	.w6(32'hbafd3ad1),
	.w7(32'hbaef8b6c),
	.w8(32'hbbaa2050),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dbba3),
	.w1(32'h3ac2549a),
	.w2(32'h3ba31e9d),
	.w3(32'h39ee1658),
	.w4(32'h3b93cef7),
	.w5(32'hba8ce067),
	.w6(32'hbbbc3b90),
	.w7(32'hbb8df392),
	.w8(32'hbc0a602a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5879d),
	.w1(32'hbb693214),
	.w2(32'hbb5669d9),
	.w3(32'h3c555b1d),
	.w4(32'hbb9b54bd),
	.w5(32'hbb193418),
	.w6(32'h3ba37b4d),
	.w7(32'hbbb1bb24),
	.w8(32'hbbaeda28),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17068e),
	.w1(32'hbbfa5907),
	.w2(32'h39c8f466),
	.w3(32'hbb91923b),
	.w4(32'h39af5199),
	.w5(32'h3976d4fe),
	.w6(32'hbc059b16),
	.w7(32'h3be3da83),
	.w8(32'h3c1b115d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1e77a),
	.w1(32'h3b1bc5c2),
	.w2(32'h399a1a4a),
	.w3(32'hbaa40030),
	.w4(32'h3ae3d397),
	.w5(32'hbb4db20c),
	.w6(32'h3a9bbb59),
	.w7(32'h3c07e170),
	.w8(32'h3bd2e976),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb7cb1),
	.w1(32'h3c12bfb4),
	.w2(32'h3c52bc59),
	.w3(32'h3ad99f73),
	.w4(32'h3a36a83d),
	.w5(32'h3bc1dc33),
	.w6(32'h3bfa9024),
	.w7(32'hba1668c6),
	.w8(32'hbb595b96),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e2b56),
	.w1(32'h3b270d09),
	.w2(32'h3b4e6556),
	.w3(32'h3b3b3c01),
	.w4(32'hba63d8aa),
	.w5(32'h3b0a866a),
	.w6(32'hbb9df30b),
	.w7(32'h3a9ff4b6),
	.w8(32'h3b117b9d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea91c5),
	.w1(32'h397a29b3),
	.w2(32'hbbffb8f2),
	.w3(32'h3a23d1db),
	.w4(32'hbbce5480),
	.w5(32'hbbc0825e),
	.w6(32'h3b096e16),
	.w7(32'hbac94564),
	.w8(32'hbb8998e9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6a88),
	.w1(32'h3abeb481),
	.w2(32'h3bdfb7dc),
	.w3(32'h3b584293),
	.w4(32'h3b2f7efb),
	.w5(32'h3bbbb473),
	.w6(32'h3b90ec7b),
	.w7(32'h3ad2f2ec),
	.w8(32'h3af2e6c9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0451),
	.w1(32'hbaa4daab),
	.w2(32'h3bbe0aa5),
	.w3(32'hb8b469f7),
	.w4(32'h3bc1bafe),
	.w5(32'h3bc4cd7c),
	.w6(32'h39ac699b),
	.w7(32'h39fe945b),
	.w8(32'hbb45ffc0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370467),
	.w1(32'h39e0d4f0),
	.w2(32'h3bd0da70),
	.w3(32'h3bb5a3d8),
	.w4(32'hbab91520),
	.w5(32'hb95b4a31),
	.w6(32'h3b4f9df3),
	.w7(32'h3bbc1948),
	.w8(32'h3a3d502e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7343ee),
	.w1(32'h3c522b79),
	.w2(32'h3bf23648),
	.w3(32'h3bb0cfc0),
	.w4(32'h3bd88596),
	.w5(32'h3b759510),
	.w6(32'h3c013c49),
	.w7(32'h3c01e1af),
	.w8(32'h3c347d4e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3d72),
	.w1(32'hba88904f),
	.w2(32'h3b55e977),
	.w3(32'hbb52b4a6),
	.w4(32'hbb4ea093),
	.w5(32'h3a9c6341),
	.w6(32'hbbe6ed1a),
	.w7(32'hbc28fd34),
	.w8(32'hbc16921c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18da88),
	.w1(32'hbb972821),
	.w2(32'hbaacf685),
	.w3(32'h3b78d795),
	.w4(32'h3a8c5b28),
	.w5(32'h39f5290b),
	.w6(32'hbb883128),
	.w7(32'h3b58a60a),
	.w8(32'h3b23e005),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c868b),
	.w1(32'hbba544c4),
	.w2(32'h3b3779ed),
	.w3(32'hbad017a9),
	.w4(32'hbb549f4d),
	.w5(32'h3b2551f1),
	.w6(32'h39d3a2bd),
	.w7(32'h3b94d8c4),
	.w8(32'hbae9e960),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac40f),
	.w1(32'h3b92c891),
	.w2(32'hbb96bdc0),
	.w3(32'hba93c5b3),
	.w4(32'hbb628289),
	.w5(32'hbb4ae176),
	.w6(32'hbbc01ffd),
	.w7(32'hbb14065b),
	.w8(32'hbb3efaa4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991b28b),
	.w1(32'hbc04fb9c),
	.w2(32'h3a2cfabc),
	.w3(32'h3a8df5fd),
	.w4(32'h39962b73),
	.w5(32'hbb1d486c),
	.w6(32'h3bd76515),
	.w7(32'hb9ceb22c),
	.w8(32'hbb8e8d41),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cd209),
	.w1(32'hbb5ecf4a),
	.w2(32'h3c2fd903),
	.w3(32'hbb956d64),
	.w4(32'h398f0013),
	.w5(32'hba0f2ee4),
	.w6(32'hbc033012),
	.w7(32'hbb7d0f14),
	.w8(32'hbb4b8acc),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc078636),
	.w1(32'hbc14147d),
	.w2(32'hbb5fba4c),
	.w3(32'hbbb91878),
	.w4(32'hbbefac3e),
	.w5(32'hbbd019bf),
	.w6(32'h3a260d0b),
	.w7(32'hbb8e805d),
	.w8(32'hbbbf6b6f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule