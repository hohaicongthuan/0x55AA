module layer_10_featuremap_220(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb54b5b55),
	.w1(32'h350b668c),
	.w2(32'h362002cc),
	.w3(32'hb2a11220),
	.w4(32'hb647efb9),
	.w5(32'h35cd2cc5),
	.w6(32'h35d3b152),
	.w7(32'h35fd246d),
	.w8(32'h34ea5f82),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd7a2e),
	.w1(32'h38a9dcf8),
	.w2(32'h389b7c41),
	.w3(32'h3911c967),
	.w4(32'h3934306c),
	.w5(32'h38c0932e),
	.w6(32'h37f2d539),
	.w7(32'h38fb2db3),
	.w8(32'h3884d54e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351eeea9),
	.w1(32'hb5b764e3),
	.w2(32'hb5a36d01),
	.w3(32'h3534febc),
	.w4(32'hb58c21b6),
	.w5(32'hb5e939f7),
	.w6(32'hb589cfea),
	.w7(32'h34fd2c8e),
	.w8(32'h358f6a51),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b8e65d),
	.w1(32'h35deeae3),
	.w2(32'h36fdca9f),
	.w3(32'h3633ba29),
	.w4(32'h368a26e6),
	.w5(32'h36abf9ba),
	.w6(32'h367bddfc),
	.w7(32'h368749ee),
	.w8(32'h3591c08c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d993f2),
	.w1(32'h381975e5),
	.w2(32'h38235988),
	.w3(32'h369698c9),
	.w4(32'h37b1dbab),
	.w5(32'h37c7db2e),
	.w6(32'hb682890d),
	.w7(32'h3492ea4d),
	.w8(32'h37b650d1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370401c1),
	.w1(32'h371ff9b7),
	.w2(32'h3616e784),
	.w3(32'h373ad4b1),
	.w4(32'h3713ad16),
	.w5(32'h368ac095),
	.w6(32'h36efd343),
	.w7(32'h36ad2ec1),
	.w8(32'hb54ba99c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9055053),
	.w1(32'h388accba),
	.w2(32'hb83a3597),
	.w3(32'hb848ee07),
	.w4(32'h3782b088),
	.w5(32'h38110593),
	.w6(32'h38034e4c),
	.w7(32'h388544d1),
	.w8(32'h3903d2e1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d0efd1),
	.w1(32'h393d8580),
	.w2(32'h38820d5d),
	.w3(32'h39114d63),
	.w4(32'h3951e432),
	.w5(32'h39300fe2),
	.w6(32'h39974f12),
	.w7(32'h38ee58be),
	.w8(32'h3821e616),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ffd53),
	.w1(32'h37856150),
	.w2(32'h37764f37),
	.w3(32'h381e23c6),
	.w4(32'h36069e4e),
	.w5(32'hb74c0561),
	.w6(32'h3884f97f),
	.w7(32'hb6776816),
	.w8(32'hb627b77e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384f942a),
	.w1(32'h37128742),
	.w2(32'h39817d22),
	.w3(32'h37f6da63),
	.w4(32'h39877417),
	.w5(32'h398203d0),
	.w6(32'h39dfe635),
	.w7(32'h39f103be),
	.w8(32'h39d533b2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390baab1),
	.w1(32'h38fbff05),
	.w2(32'h38fb4fb6),
	.w3(32'h38d11b04),
	.w4(32'h38a9e66d),
	.w5(32'h38b319f1),
	.w6(32'h38960bb3),
	.w7(32'h38dabcaa),
	.w8(32'h38f492ea),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8444d9e),
	.w1(32'hb93b3508),
	.w2(32'hb9105396),
	.w3(32'hb95e1dad),
	.w4(32'hb9b888d9),
	.w5(32'hb9338544),
	.w6(32'hb8a91a35),
	.w7(32'hb9784803),
	.w8(32'hb91f44d9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d34852),
	.w1(32'hb901125b),
	.w2(32'h39b0072a),
	.w3(32'hb9be487d),
	.w4(32'h392bbb16),
	.w5(32'h39f7f043),
	.w6(32'h3989116a),
	.w7(32'h3a07dabb),
	.w8(32'h3a0461b9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887d0a8),
	.w1(32'h386d8700),
	.w2(32'h37b62565),
	.w3(32'h37f48916),
	.w4(32'h3864b993),
	.w5(32'h367ec646),
	.w6(32'h3713cadc),
	.w7(32'hb7a96f36),
	.w8(32'h37efa039),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c228e5),
	.w1(32'hb85113e2),
	.w2(32'h37bb842e),
	.w3(32'h39259fd2),
	.w4(32'h374ae55f),
	.w5(32'h37d653d9),
	.w6(32'h38c98e6a),
	.w7(32'h3824c436),
	.w8(32'hb6f3786e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86afbfc),
	.w1(32'hb84dc05f),
	.w2(32'h395912b5),
	.w3(32'h390e31df),
	.w4(32'h398216f1),
	.w5(32'h3992bdb9),
	.w6(32'h38e9040b),
	.w7(32'h39b424c7),
	.w8(32'h3991068b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3792ea85),
	.w1(32'hb711ce5f),
	.w2(32'hb60f3326),
	.w3(32'hb7a312ef),
	.w4(32'hb81b1354),
	.w5(32'hb7d9b02d),
	.w6(32'hb68f9603),
	.w7(32'hb7451b02),
	.w8(32'hb72f8423),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a5ef7),
	.w1(32'h3972766a),
	.w2(32'h399c4ac9),
	.w3(32'h37c6d9d9),
	.w4(32'h3988d262),
	.w5(32'h39540475),
	.w6(32'h3919d626),
	.w7(32'h3991edd1),
	.w8(32'h39a96b5d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80051dc),
	.w1(32'h3785a3e8),
	.w2(32'h3924420c),
	.w3(32'hb8fc0128),
	.w4(32'h3931c847),
	.w5(32'h3945d0b0),
	.w6(32'h390921cc),
	.w7(32'h395ae3cb),
	.w8(32'h3992ad3e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4768c63),
	.w1(32'hb55c14f1),
	.w2(32'hb5571360),
	.w3(32'h351ce750),
	.w4(32'h35d30ea3),
	.w5(32'h35af2af2),
	.w6(32'hb5944a51),
	.w7(32'h3552afc7),
	.w8(32'hb53ae891),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb695a0af),
	.w1(32'hb61da37e),
	.w2(32'hb64b95ee),
	.w3(32'hb5edd741),
	.w4(32'h34de4d77),
	.w5(32'hb4b11cbe),
	.w6(32'hb600fbe5),
	.w7(32'hb5f79ebc),
	.w8(32'hb65a54ba),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f81249),
	.w1(32'h383bd94e),
	.w2(32'h37bd1be8),
	.w3(32'hb85f7384),
	.w4(32'hb79c7b1f),
	.w5(32'hb7f0575c),
	.w6(32'hb7aab1d7),
	.w7(32'h37b9d136),
	.w8(32'h36ec0f46),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db0834),
	.w1(32'h39be694a),
	.w2(32'h3953a5f8),
	.w3(32'h3a322c81),
	.w4(32'h3a0e96be),
	.w5(32'h390ae8b4),
	.w6(32'h3a2c939f),
	.w7(32'h3a2b46d7),
	.w8(32'h39adfec5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384bd90d),
	.w1(32'h38b738a0),
	.w2(32'h399bfb80),
	.w3(32'h38fb22bc),
	.w4(32'h39661a52),
	.w5(32'h3985691f),
	.w6(32'h39bd9070),
	.w7(32'h39a09359),
	.w8(32'h39b0daa0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f5722),
	.w1(32'h38a17f36),
	.w2(32'h39a0b3a0),
	.w3(32'h38480d67),
	.w4(32'h38fcf2ca),
	.w5(32'h398f9b55),
	.w6(32'h38f2a5b8),
	.w7(32'h39817716),
	.w8(32'h39ab48ed),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61ba901),
	.w1(32'hb7bcd107),
	.w2(32'hb76fd036),
	.w3(32'h37adc635),
	.w4(32'hb7d47ff1),
	.w5(32'hb7129317),
	.w6(32'h3637661a),
	.w7(32'hb735759b),
	.w8(32'hb80e6040),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34afe142),
	.w1(32'hb635917f),
	.w2(32'hb6a34143),
	.w3(32'h369701b5),
	.w4(32'h35993ef4),
	.w5(32'hb4b20373),
	.w6(32'hb6d3aead),
	.w7(32'hb6cb0083),
	.w8(32'hb69837f0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc3c21),
	.w1(32'hb9957cb1),
	.w2(32'hb87f2119),
	.w3(32'hb8ff575e),
	.w4(32'hb932f99b),
	.w5(32'h39202b63),
	.w6(32'h38854bc0),
	.w7(32'h38b2dc6f),
	.w8(32'h38cf730e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6387d),
	.w1(32'h38275d73),
	.w2(32'h3884bf7c),
	.w3(32'h38061ea0),
	.w4(32'hb849423a),
	.w5(32'hb7dda455),
	.w6(32'h37d77897),
	.w7(32'hb7eb8ede),
	.w8(32'hb6375df9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80abf16),
	.w1(32'hb890bf89),
	.w2(32'h382c7ea9),
	.w3(32'h38a0d494),
	.w4(32'h37ff8367),
	.w5(32'h38adda0f),
	.w6(32'h3951ef99),
	.w7(32'h39184bd3),
	.w8(32'h38efc78c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb436e894),
	.w1(32'hb6489c11),
	.w2(32'hb63b26e7),
	.w3(32'hb5c32872),
	.w4(32'hb69bba47),
	.w5(32'hb69100ce),
	.w6(32'hb65ffa52),
	.w7(32'hb6b2346c),
	.w8(32'hb67a20ce),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6162d79),
	.w1(32'h368f8e7a),
	.w2(32'h35b3fa16),
	.w3(32'hb6930875),
	.w4(32'hb65773d1),
	.w5(32'hb6f9747b),
	.w6(32'hb5d2206d),
	.w7(32'hb627dd08),
	.w8(32'hb702f2e6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8427f),
	.w1(32'h388436e2),
	.w2(32'h3949f13f),
	.w3(32'hb756ddad),
	.w4(32'h38c853ac),
	.w5(32'h392654c0),
	.w6(32'h38519e24),
	.w7(32'h38f12eae),
	.w8(32'h396bee4e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df4ddc),
	.w1(32'h3898779d),
	.w2(32'h38bcaf22),
	.w3(32'h39562e5f),
	.w4(32'h38be2539),
	.w5(32'h389b537f),
	.w6(32'h38971129),
	.w7(32'h36b49c1e),
	.w8(32'hb7ab50bf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38205736),
	.w1(32'h3833aba4),
	.w2(32'h37a37e70),
	.w3(32'h3863c3df),
	.w4(32'h384c50a9),
	.w5(32'h3786324c),
	.w6(32'h37e3c289),
	.w7(32'h38204919),
	.w8(32'h37762b2a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dbce16),
	.w1(32'h37d32ddf),
	.w2(32'h3894bb3f),
	.w3(32'hb8dcf4ae),
	.w4(32'h38a08b82),
	.w5(32'h38b226c0),
	.w6(32'h38827ab9),
	.w7(32'h39202d19),
	.w8(32'h3901a07d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d9f8c),
	.w1(32'h3991f80b),
	.w2(32'h3982f961),
	.w3(32'h3a17771c),
	.w4(32'h3a2f296a),
	.w5(32'h39dbbd78),
	.w6(32'h3a177406),
	.w7(32'h3a30d12b),
	.w8(32'h39a2a041),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d686c),
	.w1(32'h388f670b),
	.w2(32'hb84cdd29),
	.w3(32'h39c4ecd4),
	.w4(32'hb8f1e104),
	.w5(32'hb80e71e1),
	.w6(32'h392003db),
	.w7(32'hb9276f67),
	.w8(32'hb700b25f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8030c),
	.w1(32'h398f271f),
	.w2(32'h38cfd75b),
	.w3(32'h39786eec),
	.w4(32'h38e4e275),
	.w5(32'h37d5d382),
	.w6(32'h39d7fc7b),
	.w7(32'h39944818),
	.w8(32'h392db53d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd8dc5),
	.w1(32'hb8e2129b),
	.w2(32'h37c06fc5),
	.w3(32'hb8d382a8),
	.w4(32'hb90458bf),
	.w5(32'h37f44354),
	.w6(32'hb8dbd202),
	.w7(32'hb8a73810),
	.w8(32'h37b35532),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36aad057),
	.w1(32'hb5313a7c),
	.w2(32'h370a949a),
	.w3(32'h36d72520),
	.w4(32'hb4bef5b3),
	.w5(32'h370155e0),
	.w6(32'hb6147b3a),
	.w7(32'h3678311b),
	.w8(32'hb69a68f6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73a3756),
	.w1(32'hb7586e22),
	.w2(32'hb76d15a8),
	.w3(32'hb6a0d144),
	.w4(32'hb66dd211),
	.w5(32'hb6d72601),
	.w6(32'hb7340a0b),
	.w7(32'hb732b50e),
	.w8(32'hb6568ba3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed153d),
	.w1(32'hb846228a),
	.w2(32'h38c4796b),
	.w3(32'h38aed98a),
	.w4(32'hb8cc279b),
	.w5(32'h39176281),
	.w6(32'h38b5f371),
	.w7(32'hb8ab02e3),
	.w8(32'h390d8a42),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385b3b04),
	.w1(32'hb8a949bf),
	.w2(32'h39c376e7),
	.w3(32'h38e55c1d),
	.w4(32'h3951b60f),
	.w5(32'h39128a44),
	.w6(32'h3987ae22),
	.w7(32'h39a58666),
	.w8(32'h396af975),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85a4121),
	.w1(32'h3714ddad),
	.w2(32'h39195ef4),
	.w3(32'h385b79af),
	.w4(32'h38f703b7),
	.w5(32'h391d753c),
	.w6(32'h3979d151),
	.w7(32'h396d1992),
	.w8(32'h396e5815),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a3fcd),
	.w1(32'h38be6d3f),
	.w2(32'h398fac28),
	.w3(32'h36dee0bc),
	.w4(32'h3985979a),
	.w5(32'h3991ad8d),
	.w6(32'h39b502c8),
	.w7(32'h39c8ccf0),
	.w8(32'h39e7dad8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83bd9b0),
	.w1(32'hb809a8da),
	.w2(32'h36a0e078),
	.w3(32'h38681659),
	.w4(32'h36cadcfe),
	.w5(32'h3869679c),
	.w6(32'h393f64de),
	.w7(32'h389fec5c),
	.w8(32'h38964860),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6b7fc),
	.w1(32'h381b8424),
	.w2(32'h39b2aa57),
	.w3(32'h37e75e16),
	.w4(32'h3952beb2),
	.w5(32'h39ec4e04),
	.w6(32'h39984c5e),
	.w7(32'h39ad6a1d),
	.w8(32'h39e08087),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5fcd85a),
	.w1(32'hb78db93c),
	.w2(32'h362f718c),
	.w3(32'h370467ab),
	.w4(32'hb77aa57d),
	.w5(32'hb69be46c),
	.w6(32'h3759cbc0),
	.w7(32'hb6c70a87),
	.w8(32'hb6bb7943),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38041763),
	.w1(32'hb87aa785),
	.w2(32'hb835a450),
	.w3(32'h38ac0f12),
	.w4(32'hb7688f43),
	.w5(32'h3635d616),
	.w6(32'h38ec7a99),
	.w7(32'h37d6a85b),
	.w8(32'h3653c726),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79c60d2),
	.w1(32'hb7831454),
	.w2(32'h375d397c),
	.w3(32'hb812c187),
	.w4(32'hb7878650),
	.w5(32'h379125b1),
	.w6(32'hb75b6edc),
	.w7(32'hb77a0710),
	.w8(32'h36fb93f1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906607a),
	.w1(32'h37cd5115),
	.w2(32'h39d1d94f),
	.w3(32'hb8a8f434),
	.w4(32'h38ba6d19),
	.w5(32'h39f4e923),
	.w6(32'h39123817),
	.w7(32'h38f60901),
	.w8(32'h3a01f489),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381fc720),
	.w1(32'h387e886a),
	.w2(32'h3867577c),
	.w3(32'hb70970a7),
	.w4(32'h36aaf69d),
	.w5(32'h37800ca5),
	.w6(32'h378eb28e),
	.w7(32'h380eacfa),
	.w8(32'h38717c79),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d8cd4),
	.w1(32'h395b2ab5),
	.w2(32'h39763c93),
	.w3(32'h382c0d5a),
	.w4(32'h398828d4),
	.w5(32'h39a65299),
	.w6(32'h39ff165e),
	.w7(32'h39fe9e69),
	.w8(32'h39e7ecc7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382345ba),
	.w1(32'h3744a83d),
	.w2(32'hb59b0f55),
	.w3(32'h38217513),
	.w4(32'hb69d118f),
	.w5(32'hb72236a5),
	.w6(32'h380bd97f),
	.w7(32'h36b0a227),
	.w8(32'hb741c66b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60e69ba),
	.w1(32'hb6454fb2),
	.w2(32'h3608da8a),
	.w3(32'hb6041e8b),
	.w4(32'hb5c666fb),
	.w5(32'h3694a39e),
	.w6(32'hb706a5cc),
	.w7(32'hb5b24f00),
	.w8(32'hb66699d7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6391858),
	.w1(32'hb62ff5ad),
	.w2(32'hb5efde47),
	.w3(32'hb599662a),
	.w4(32'hb5fd1258),
	.w5(32'h3338378b),
	.w6(32'hb5d7ec7c),
	.w7(32'hb50261c2),
	.w8(32'hb5e07f1c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34831e8c),
	.w1(32'h35e2e388),
	.w2(32'hb6ad9617),
	.w3(32'h35881285),
	.w4(32'h35aca58d),
	.w5(32'hb6f8bb0f),
	.w6(32'h35e6fa5d),
	.w7(32'hb6260465),
	.w8(32'h3525beec),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f780f),
	.w1(32'h3787f625),
	.w2(32'h382eca04),
	.w3(32'h3815ffd4),
	.w4(32'hafb127f1),
	.w5(32'h381ab8b6),
	.w6(32'h382e9d13),
	.w7(32'h36c5037c),
	.w8(32'h388516fe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e0bf90),
	.w1(32'hb7526222),
	.w2(32'h3776c33d),
	.w3(32'hb7957ef7),
	.w4(32'hb81f9ab0),
	.w5(32'h3602a1d2),
	.w6(32'h37501870),
	.w7(32'hb793acb6),
	.w8(32'h37f66794),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8acc7e7),
	.w1(32'hb891b596),
	.w2(32'h397d5d80),
	.w3(32'hb8857c43),
	.w4(32'h38341a5f),
	.w5(32'h39739453),
	.w6(32'h394ab4e0),
	.w7(32'h39ae1504),
	.w8(32'h398f14ca),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37980066),
	.w1(32'h383f6b35),
	.w2(32'h3813f189),
	.w3(32'h38ab7cd3),
	.w4(32'h38884022),
	.w5(32'h3884375b),
	.w6(32'h380be0ca),
	.w7(32'h381314f4),
	.w8(32'h38432ba1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb606db1e),
	.w1(32'hb674b601),
	.w2(32'h3669321a),
	.w3(32'hb68d2e71),
	.w4(32'hb6f2299c),
	.w5(32'hb62f732f),
	.w6(32'hb6f79ab3),
	.w7(32'hb69de6aa),
	.w8(32'hb6cbb225),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63486da),
	.w1(32'hb5faf9c6),
	.w2(32'hb593cec4),
	.w3(32'h35dd9dfb),
	.w4(32'h3541e07c),
	.w5(32'hb2902fc7),
	.w6(32'hb47f6832),
	.w7(32'h358e75e5),
	.w8(32'h346db2bd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362afe6b),
	.w1(32'hb5b385e7),
	.w2(32'hb6a71e9b),
	.w3(32'h365980f8),
	.w4(32'hb5f3f29e),
	.w5(32'hb6ce6f70),
	.w6(32'hb52f4031),
	.w7(32'hb59ad337),
	.w8(32'hb6042eea),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ac45e8),
	.w1(32'h351eeac2),
	.w2(32'hb6ff75df),
	.w3(32'h35f140dd),
	.w4(32'h35114538),
	.w5(32'hb6b9b97a),
	.w6(32'hb6853e8a),
	.w7(32'hb6ce21c2),
	.w8(32'hb5a85455),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73bc8f6),
	.w1(32'h378b0de5),
	.w2(32'h38d586b1),
	.w3(32'hb7dcdfd0),
	.w4(32'hb8694893),
	.w5(32'hb8d15c17),
	.w6(32'h390aa623),
	.w7(32'h392ac43a),
	.w8(32'h3901748f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381db1ac),
	.w1(32'h3938c489),
	.w2(32'h39b8c0b0),
	.w3(32'hb8d7d876),
	.w4(32'h391201d9),
	.w5(32'h39a225fd),
	.w6(32'h3911f431),
	.w7(32'h39984c99),
	.w8(32'h39dbbbf4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e549a6),
	.w1(32'h3988ceea),
	.w2(32'h398ffeb3),
	.w3(32'h3949dbdc),
	.w4(32'h396d1367),
	.w5(32'h3980cb33),
	.w6(32'h395788bf),
	.w7(32'h39a0bbb8),
	.w8(32'h39abfe64),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d90e4d),
	.w1(32'h371a5cbd),
	.w2(32'h39fc7c0a),
	.w3(32'h3971fb02),
	.w4(32'h39bee23a),
	.w5(32'h3a2e2070),
	.w6(32'h39f51dea),
	.w7(32'h3a462567),
	.w8(32'h3a0b3e7f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb621d3ad),
	.w1(32'hb6aaeebf),
	.w2(32'hb60e0bc0),
	.w3(32'h361531e9),
	.w4(32'h3607e811),
	.w5(32'h368bfd55),
	.w6(32'hb52bcc83),
	.w7(32'h33e80c56),
	.w8(32'h35d5466d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c379e7),
	.w1(32'hb66f791b),
	.w2(32'hb6e369a1),
	.w3(32'hb5c476f7),
	.w4(32'h35354bb4),
	.w5(32'hb4dc3dcf),
	.w6(32'hb6a40ea6),
	.w7(32'hb659a1f2),
	.w8(32'hb69c0d30),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71b8c7f),
	.w1(32'hb68a7bf5),
	.w2(32'hb6d75b20),
	.w3(32'hb6a0b674),
	.w4(32'h3614e806),
	.w5(32'h35ca1ba2),
	.w6(32'hb64effef),
	.w7(32'hb60a8d41),
	.w8(32'hb65238b9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77cc36e),
	.w1(32'h38173f1e),
	.w2(32'h38d7f375),
	.w3(32'hb8428ee7),
	.w4(32'h38572584),
	.w5(32'h38d7e9da),
	.w6(32'h3869e454),
	.w7(32'h38cccdb7),
	.w8(32'h38ea7782),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76217fa),
	.w1(32'hb699446f),
	.w2(32'hb613bef0),
	.w3(32'hb6ee5c43),
	.w4(32'hb6349def),
	.w5(32'hb517ab02),
	.w6(32'hb682574e),
	.w7(32'hb5edf68e),
	.w8(32'h35bda965),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394072bd),
	.w1(32'h398aeec5),
	.w2(32'h3943b61f),
	.w3(32'h38811c4f),
	.w4(32'h39004871),
	.w5(32'hb78d283c),
	.w6(32'h38a36ea5),
	.w7(32'h39277bdb),
	.w8(32'h39480880),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9970e),
	.w1(32'hb95d2f22),
	.w2(32'h387d2604),
	.w3(32'h38c23ab7),
	.w4(32'hb7f64ec3),
	.w5(32'hb687045c),
	.w6(32'h390df3a8),
	.w7(32'h39aa602c),
	.w8(32'hb724b9ac),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d73465),
	.w1(32'hb8e3fa00),
	.w2(32'h399ae446),
	.w3(32'hb894f475),
	.w4(32'h3884f9b9),
	.w5(32'h39b8e2a2),
	.w6(32'h392ef1be),
	.w7(32'h39a8cd73),
	.w8(32'h39c8a31a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c8534),
	.w1(32'h39013918),
	.w2(32'h396bbc32),
	.w3(32'h3910aaf0),
	.w4(32'h391484f3),
	.w5(32'h38eb77fb),
	.w6(32'h3909d97c),
	.w7(32'h3921db08),
	.w8(32'h3939dd19),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6949026),
	.w1(32'h38ce4aca),
	.w2(32'h3922a980),
	.w3(32'hb8c076c4),
	.w4(32'h38669e99),
	.w5(32'h3889b684),
	.w6(32'h389310fc),
	.w7(32'h38ee7899),
	.w8(32'h3970245d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e8711a),
	.w1(32'h3841628c),
	.w2(32'h38c1e50b),
	.w3(32'h38b7b079),
	.w4(32'h38d74f69),
	.w5(32'h38aff903),
	.w6(32'h38fc8e91),
	.w7(32'h39073271),
	.w8(32'h38ae9b8f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b79a01),
	.w1(32'h3908c2e0),
	.w2(32'h39808e09),
	.w3(32'hb9068720),
	.w4(32'h390781fa),
	.w5(32'h394007da),
	.w6(32'hb790f3a1),
	.w7(32'h3922f9f8),
	.w8(32'h3977ce22),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6499a32),
	.w1(32'hb619267f),
	.w2(32'h34b8068f),
	.w3(32'hb6400896),
	.w4(32'hb5a95da3),
	.w5(32'h34e41044),
	.w6(32'hb64cc2b8),
	.w7(32'hb4d3a92f),
	.w8(32'hb510a469),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6189f9a),
	.w1(32'hb5640b34),
	.w2(32'hb5a6c820),
	.w3(32'h351216a8),
	.w4(32'h338c70c6),
	.w5(32'hb54dcf5b),
	.w6(32'h36481bbe),
	.w7(32'h35733553),
	.w8(32'hb5ff56fb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57c0083),
	.w1(32'hb6aea24b),
	.w2(32'h332577d0),
	.w3(32'h35458afc),
	.w4(32'hb68d3ffd),
	.w5(32'h34f5326d),
	.w6(32'hb5e23ff6),
	.w7(32'h36512ffe),
	.w8(32'h366ea46f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351ad045),
	.w1(32'hb591fd70),
	.w2(32'h36086366),
	.w3(32'h3516f7ab),
	.w4(32'hb5a3c91d),
	.w5(32'h35eea805),
	.w6(32'hb5d7c4cb),
	.w7(32'hb6150980),
	.w8(32'hb5e6c4ca),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3ce46),
	.w1(32'hb9691cc3),
	.w2(32'h376f245f),
	.w3(32'hb83de6ad),
	.w4(32'hb8f78167),
	.w5(32'hb8f15434),
	.w6(32'hb825e3de),
	.w7(32'hb8af87b6),
	.w8(32'hb8eddc78),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c90e2d),
	.w1(32'h37c5a61b),
	.w2(32'h37e9abff),
	.w3(32'h3799a377),
	.w4(32'h370ceb90),
	.w5(32'h36bd8933),
	.w6(32'hb7005d0a),
	.w7(32'h37a25710),
	.w8(32'hb657097f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84f17d4),
	.w1(32'h385b4679),
	.w2(32'h390189a0),
	.w3(32'h381dc9b0),
	.w4(32'h391a924d),
	.w5(32'h390d96a6),
	.w6(32'h398a8299),
	.w7(32'h39155c02),
	.w8(32'h38fe74ab),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a016f),
	.w1(32'h3a54a6b4),
	.w2(32'h3a0068c9),
	.w3(32'h39c15433),
	.w4(32'h38c39a8e),
	.w5(32'h38571fa3),
	.w6(32'hb8235b22),
	.w7(32'h3748fdde),
	.w8(32'h39a4d9d6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972e658),
	.w1(32'h38d29b10),
	.w2(32'h38b1abad),
	.w3(32'h38a148eb),
	.w4(32'hb89e28ee),
	.w5(32'h36a0d0c9),
	.w6(32'h3941e9ee),
	.w7(32'h380f33d9),
	.w8(32'h3851a664),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398da40c),
	.w1(32'h39725a1e),
	.w2(32'h39dda6fd),
	.w3(32'h36d278cc),
	.w4(32'h355f1520),
	.w5(32'h39e36efe),
	.w6(32'h386d54bb),
	.w7(32'h391332ad),
	.w8(32'h39e26a82),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ad606),
	.w1(32'hb8f60470),
	.w2(32'h392c7d40),
	.w3(32'hb93ea9ce),
	.w4(32'h384ab6f2),
	.w5(32'h3983dce7),
	.w6(32'hb809544d),
	.w7(32'h39800ba7),
	.w8(32'h39ca3a6e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3775bc70),
	.w1(32'hb93bb2d8),
	.w2(32'hb8d73585),
	.w3(32'h39386dcb),
	.w4(32'hb8a6a444),
	.w5(32'hb7b83390),
	.w6(32'h391dffa4),
	.w7(32'hb8e0d5c2),
	.w8(32'hb84d9f61),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b2e08),
	.w1(32'hb924aa81),
	.w2(32'h37c1f386),
	.w3(32'h3813c573),
	.w4(32'hb804f02e),
	.w5(32'h3884e938),
	.w6(32'h38fdb0b5),
	.w7(32'h38a820dc),
	.w8(32'h38f22fad),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea766b),
	.w1(32'hb92b1283),
	.w2(32'h3941ea0a),
	.w3(32'hb895b78e),
	.w4(32'hb9810263),
	.w5(32'h37dab32d),
	.w6(32'h36e4b529),
	.w7(32'hb881e34f),
	.w8(32'h390ff73e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37835c20),
	.w1(32'h3732cfbb),
	.w2(32'h36b8a0c8),
	.w3(32'h36a4a8c2),
	.w4(32'hb7568175),
	.w5(32'hb7973189),
	.w6(32'h3801ad33),
	.w7(32'h374dbb9b),
	.w8(32'hb79c78b3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b6db5),
	.w1(32'hb897e531),
	.w2(32'h38ff3323),
	.w3(32'h376d3886),
	.w4(32'h38ab5f22),
	.w5(32'h38f7affd),
	.w6(32'h399c6e89),
	.w7(32'h396e12cf),
	.w8(32'h3985b931),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86d6fe8),
	.w1(32'h395d0c8d),
	.w2(32'h396544f4),
	.w3(32'h383c2118),
	.w4(32'h398a92de),
	.w5(32'h39af99c4),
	.w6(32'h39436f26),
	.w7(32'h39e739de),
	.w8(32'h39bf1858),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e2f75),
	.w1(32'h39d10ef2),
	.w2(32'h39d5aa48),
	.w3(32'hb830e4a2),
	.w4(32'h39bf560e),
	.w5(32'h39981ee7),
	.w6(32'hb888e889),
	.w7(32'h39908088),
	.w8(32'h39d59b60),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63566c0),
	.w1(32'hb9d2b390),
	.w2(32'hb821e845),
	.w3(32'h39bc1eb7),
	.w4(32'hb982e86c),
	.w5(32'h38cfe539),
	.w6(32'h3a82dc45),
	.w7(32'h38dff93d),
	.w8(32'h39b179ae),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94be296),
	.w1(32'h36b3cd0f),
	.w2(32'h398877c6),
	.w3(32'hb7f90e51),
	.w4(32'h3964028f),
	.w5(32'h39b1a232),
	.w6(32'h398e8ae3),
	.w7(32'h39c4439b),
	.w8(32'h39e86b5d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c7fd7b),
	.w1(32'h3883f804),
	.w2(32'hb61b7c53),
	.w3(32'h3919e107),
	.w4(32'h389132b8),
	.w5(32'h38f71687),
	.w6(32'h396fcbbd),
	.w7(32'h391d4990),
	.w8(32'h38d9260d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74c9f44),
	.w1(32'hb7dff4e2),
	.w2(32'hb75ec29a),
	.w3(32'hb86c220d),
	.w4(32'hb8712d9b),
	.w5(32'hb81c1970),
	.w6(32'h3819cf4b),
	.w7(32'h37a263bb),
	.w8(32'h37bc6cba),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38169cc4),
	.w1(32'h388da988),
	.w2(32'h39b18960),
	.w3(32'h379e0dc6),
	.w4(32'h39c0f693),
	.w5(32'h39c330f8),
	.w6(32'h398c0154),
	.w7(32'h398c2913),
	.w8(32'h39f08566),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a0134),
	.w1(32'hba06af6b),
	.w2(32'h3971899d),
	.w3(32'hb9296932),
	.w4(32'hb98f3a96),
	.w5(32'h39bcf5be),
	.w6(32'hb8844a69),
	.w7(32'h38b6c661),
	.w8(32'h398449d2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6110366),
	.w1(32'h37820300),
	.w2(32'h3735716b),
	.w3(32'hb78601ac),
	.w4(32'hb4d170c2),
	.w5(32'hb61dad4a),
	.w6(32'h36f6f255),
	.w7(32'h3757ff1a),
	.w8(32'h374faf03),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f79a22),
	.w1(32'h380dd8f4),
	.w2(32'h37ffd856),
	.w3(32'h3821e780),
	.w4(32'h3838b9bb),
	.w5(32'h37f20773),
	.w6(32'h3762aa3f),
	.w7(32'hb64387c9),
	.w8(32'h37fae540),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0c242),
	.w1(32'hb8dd1495),
	.w2(32'h39350182),
	.w3(32'h387fce1f),
	.w4(32'h37f0e43c),
	.w5(32'h3927b9f9),
	.w6(32'h3945db29),
	.w7(32'h39204c72),
	.w8(32'h393a666a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ca798a),
	.w1(32'h37a99346),
	.w2(32'h396c24d4),
	.w3(32'h3855653e),
	.w4(32'h39166038),
	.w5(32'h3972116d),
	.w6(32'h394c0727),
	.w7(32'h399ac368),
	.w8(32'h3999ce2f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963166d),
	.w1(32'h374b670a),
	.w2(32'hb8e8f28f),
	.w3(32'h39a37390),
	.w4(32'h396fce11),
	.w5(32'hb881ddcf),
	.w6(32'h3927c08b),
	.w7(32'h39073bd3),
	.w8(32'hb8af6a37),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b95318),
	.w1(32'h38bdda0f),
	.w2(32'h38be820c),
	.w3(32'h392f1da6),
	.w4(32'h39a4438c),
	.w5(32'h395b627a),
	.w6(32'h37c52d4d),
	.w7(32'h398a339c),
	.w8(32'h39ca6dfc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382dce51),
	.w1(32'h36f73457),
	.w2(32'h372f9048),
	.w3(32'h36a3d948),
	.w4(32'hb7d0dafe),
	.w5(32'hb763f013),
	.w6(32'h38bd5ffc),
	.w7(32'h37c02bd5),
	.w8(32'h360e0680),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885fe4b),
	.w1(32'hb71eca12),
	.w2(32'h398ead55),
	.w3(32'h374ac5a3),
	.w4(32'h38e0cc0f),
	.w5(32'h3948e9b9),
	.w6(32'h39293ff8),
	.w7(32'h3933ef0e),
	.w8(32'h39961cce),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dd24d8),
	.w1(32'h383e5640),
	.w2(32'h391a139e),
	.w3(32'hb72b81e6),
	.w4(32'h389573dd),
	.w5(32'h391ecc85),
	.w6(32'h38a4dffd),
	.w7(32'h390d8c91),
	.w8(32'h39401b15),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352b77b3),
	.w1(32'h348e11d1),
	.w2(32'hb6634627),
	.w3(32'hb55fb063),
	.w4(32'hb6162b1f),
	.w5(32'hb667ebce),
	.w6(32'hb51a2e73),
	.w7(32'hb60f14a4),
	.w8(32'hb6af959d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb58e919f),
	.w1(32'h35d934fa),
	.w2(32'h33dbbd31),
	.w3(32'hb5a8adae),
	.w4(32'h362fa485),
	.w5(32'h36233e6c),
	.w6(32'hb6067e2c),
	.w7(32'h35833d1c),
	.w8(32'hb576960d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62b8525),
	.w1(32'h34524bda),
	.w2(32'hb59cef16),
	.w3(32'h3607f501),
	.w4(32'h3602de44),
	.w5(32'h3585b7be),
	.w6(32'h3582afeb),
	.w7(32'h3611ddcb),
	.w8(32'h35acf359),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d07c5),
	.w1(32'h3813c29d),
	.w2(32'h38163768),
	.w3(32'h379454f6),
	.w4(32'h375c1dfa),
	.w5(32'h374dba28),
	.w6(32'h3715f6ce),
	.w7(32'hb706a3bd),
	.w8(32'hb6c33417),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9066f47),
	.w1(32'hb877d6d6),
	.w2(32'h38a9cd6e),
	.w3(32'h37988869),
	.w4(32'h3890a222),
	.w5(32'h39246cf7),
	.w6(32'h39502280),
	.w7(32'h390f9334),
	.w8(32'h39231c20),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee6ba6),
	.w1(32'h38a592fc),
	.w2(32'h389cf25e),
	.w3(32'h38939af3),
	.w4(32'h380ddb86),
	.w5(32'h380c8f50),
	.w6(32'h37da4010),
	.w7(32'h36c44086),
	.w8(32'h3807d192),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7f861),
	.w1(32'h3785ce22),
	.w2(32'h3845a0d3),
	.w3(32'hb782bcea),
	.w4(32'h375ea2a5),
	.w5(32'h3870dff1),
	.w6(32'h38d12a72),
	.w7(32'h38dd03f3),
	.w8(32'h3938a681),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb6ce0),
	.w1(32'h398d7ee9),
	.w2(32'h39bbec6b),
	.w3(32'h39e4ef2b),
	.w4(32'h39e8d727),
	.w5(32'h3a1bd7f4),
	.w6(32'h388f87b6),
	.w7(32'h39d32edc),
	.w8(32'h3a3600e5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36248cff),
	.w1(32'hb6d2374a),
	.w2(32'h3729da5b),
	.w3(32'hb6eb75f8),
	.w4(32'h3724972d),
	.w5(32'h379b19e8),
	.w6(32'hb7f4f534),
	.w7(32'hb63e1a44),
	.w8(32'h387ab99d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3748ea48),
	.w1(32'h37403862),
	.w2(32'h376546d4),
	.w3(32'h375fab0b),
	.w4(32'h373f200e),
	.w5(32'h370637e0),
	.w6(32'h372fba80),
	.w7(32'h373f8938),
	.w8(32'h37534930),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb45dd1bc),
	.w1(32'hb63ed8bc),
	.w2(32'hb6385d67),
	.w3(32'hb56e5f78),
	.w4(32'hb67535c2),
	.w5(32'hb5e7e42b),
	.w6(32'hb685ae65),
	.w7(32'hb69c5a33),
	.w8(32'hb5dfab3c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3821a169),
	.w1(32'hba0ecc53),
	.w2(32'hb9b46c5e),
	.w3(32'h3861e62e),
	.w4(32'hba6038ee),
	.w5(32'hb9d58ca3),
	.w6(32'hba03a373),
	.w7(32'hb9fe5da0),
	.w8(32'hb917529d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbe4e3),
	.w1(32'h37e0fb76),
	.w2(32'hb97358b4),
	.w3(32'hb9b3e07a),
	.w4(32'hb9389ec9),
	.w5(32'hb99c9b27),
	.w6(32'hb9259e8c),
	.w7(32'hb9c96617),
	.w8(32'h38558967),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bcb68f),
	.w1(32'h3a3203d0),
	.w2(32'hbb167451),
	.w3(32'hb9603ed2),
	.w4(32'h3b0598d2),
	.w5(32'h3adc9de4),
	.w6(32'h3aa030b6),
	.w7(32'h3a27b7a9),
	.w8(32'h3a493891),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d8b6e),
	.w1(32'hba22299a),
	.w2(32'hb9ae400d),
	.w3(32'h3a667f02),
	.w4(32'hb98b32c4),
	.w5(32'hba089118),
	.w6(32'hbaa8e1be),
	.w7(32'hba97e571),
	.w8(32'hba59a1ea),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c6b80),
	.w1(32'h37cc822f),
	.w2(32'h3a5f02e3),
	.w3(32'hb9e2df35),
	.w4(32'hba08d9a0),
	.w5(32'hba0c6c5b),
	.w6(32'hbaadb2cc),
	.w7(32'hbab4e623),
	.w8(32'hbabdcc5b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fd821),
	.w1(32'hb9cdfcc0),
	.w2(32'hbb438c84),
	.w3(32'hba8840fc),
	.w4(32'hb9c7f73c),
	.w5(32'hba7c34ef),
	.w6(32'h3a4e95c8),
	.w7(32'h3a6fcc2e),
	.w8(32'h3a632a5e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba854b0a),
	.w1(32'h3a725fed),
	.w2(32'h3a625f28),
	.w3(32'hbaa1a569),
	.w4(32'h3a4508a9),
	.w5(32'h39fbe7e0),
	.w6(32'h3b1617a8),
	.w7(32'h3aa307fa),
	.w8(32'h3915b3ca),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfc6fd),
	.w1(32'hba90af8e),
	.w2(32'hba6b0d47),
	.w3(32'h384d6011),
	.w4(32'hba866931),
	.w5(32'hba709b1f),
	.w6(32'hba85e559),
	.w7(32'hba825d7e),
	.w8(32'hba149f12),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb799dc68),
	.w1(32'h3a4685f1),
	.w2(32'h3a62eb0f),
	.w3(32'hb9e5639a),
	.w4(32'h3a382ba1),
	.w5(32'h39bd5c31),
	.w6(32'h393fddf4),
	.w7(32'h396d2ae7),
	.w8(32'hb965d7bf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85c725),
	.w1(32'hb8b84afd),
	.w2(32'hb9d1652e),
	.w3(32'hba325c93),
	.w4(32'hb9a32f76),
	.w5(32'hba19692d),
	.w6(32'hb96e58f9),
	.w7(32'hba326363),
	.w8(32'hba3422a0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c513b),
	.w1(32'h399e9c58),
	.w2(32'h3a46cf14),
	.w3(32'hb9e8d3f9),
	.w4(32'hba4c325f),
	.w5(32'hb8f61567),
	.w6(32'h39c1fadc),
	.w7(32'h39b0dce5),
	.w8(32'h39823ee4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa6d69),
	.w1(32'h3a656ad6),
	.w2(32'h39933f35),
	.w3(32'hb9a24341),
	.w4(32'h3ab63445),
	.w5(32'h3a942155),
	.w6(32'h3a015c30),
	.w7(32'h38ffb68e),
	.w8(32'h3a696a48),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b9521),
	.w1(32'h3ada92a0),
	.w2(32'h3a942dc7),
	.w3(32'h3ac2f4cd),
	.w4(32'h3a727a4b),
	.w5(32'h3ae1d94e),
	.w6(32'h3a6bb594),
	.w7(32'hb9bedef9),
	.w8(32'hb868f743),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaced11),
	.w1(32'h3a173b00),
	.w2(32'hb8e230de),
	.w3(32'h3a7875db),
	.w4(32'h39f10db8),
	.w5(32'h3a428554),
	.w6(32'h3aaf65c3),
	.w7(32'h3a2a4153),
	.w8(32'h3a4d5267),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5934fb),
	.w1(32'h3990922d),
	.w2(32'h3a499913),
	.w3(32'h3a260fc1),
	.w4(32'h39a0719a),
	.w5(32'h3a90e7f9),
	.w6(32'h393b4a10),
	.w7(32'hb81e74f2),
	.w8(32'hb8f54b69),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48889b),
	.w1(32'h38af54bf),
	.w2(32'hba56013a),
	.w3(32'h3aa6c603),
	.w4(32'h381b5c3f),
	.w5(32'hba87e454),
	.w6(32'hb9b87883),
	.w7(32'hbaa0197e),
	.w8(32'hba167f24),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90838bb),
	.w1(32'h3aab2f69),
	.w2(32'hbb14aca1),
	.w3(32'hba2f7fce),
	.w4(32'h3aa712d7),
	.w5(32'h3abac633),
	.w6(32'h3b590f59),
	.w7(32'h3af24749),
	.w8(32'h3abc2966),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98c6fb),
	.w1(32'hb8250eb5),
	.w2(32'h39f23ddd),
	.w3(32'h3abf8cf7),
	.w4(32'hba57bfc2),
	.w5(32'hba209e7e),
	.w6(32'hb9758766),
	.w7(32'hb8a2495f),
	.w8(32'hb914ea76),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba165e00),
	.w1(32'hb92b5080),
	.w2(32'h3a90bb89),
	.w3(32'hba5dc7b5),
	.w4(32'hb98f50cf),
	.w5(32'hb78d6cc1),
	.w6(32'hb948eaf4),
	.w7(32'h39d59ed0),
	.w8(32'h39d79425),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970b5b1),
	.w1(32'h3a1a4c0f),
	.w2(32'h3a6959a9),
	.w3(32'h3a5c614f),
	.w4(32'h3a11cc96),
	.w5(32'h3a3c3cfc),
	.w6(32'h38305951),
	.w7(32'h39aaea89),
	.w8(32'hb8d55b41),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f50fb8),
	.w1(32'hb9f28fb9),
	.w2(32'hb9133fe4),
	.w3(32'h3a043baf),
	.w4(32'hba380bbc),
	.w5(32'hba070529),
	.w6(32'hba2d4b6a),
	.w7(32'hb9d7b25a),
	.w8(32'hb9c2b72a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52c696),
	.w1(32'h3a2369fa),
	.w2(32'h3aeaed89),
	.w3(32'hba1be179),
	.w4(32'hb8a4ea1b),
	.w5(32'h3a4ae587),
	.w6(32'h3a1d1d6e),
	.w7(32'h3a9f7067),
	.w8(32'h3a896711),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1ae8c),
	.w1(32'hba2eebf0),
	.w2(32'hba092765),
	.w3(32'h39f6c609),
	.w4(32'hbab95202),
	.w5(32'hbac6a61c),
	.w6(32'hba469c06),
	.w7(32'hba2bce6c),
	.w8(32'hba7ead6b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0ea3),
	.w1(32'h3a40b412),
	.w2(32'h3a0f38a5),
	.w3(32'hba977fda),
	.w4(32'h3ad059f8),
	.w5(32'h3afa1baa),
	.w6(32'h3a431c1a),
	.w7(32'h3a59c335),
	.w8(32'h3ab41459),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38857667),
	.w1(32'h3a16dcbb),
	.w2(32'h3af1b838),
	.w3(32'h3a1cdfd2),
	.w4(32'h39687fc0),
	.w5(32'h3a947d9f),
	.w6(32'h390f07af),
	.w7(32'h3aba1c33),
	.w8(32'h3a6fa1e5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16c87e),
	.w1(32'h38a71e4d),
	.w2(32'hb8b221d3),
	.w3(32'hb99fb4bc),
	.w4(32'hb88cecb8),
	.w5(32'hb98bc816),
	.w6(32'h38af7ccd),
	.w7(32'hb9bb5c16),
	.w8(32'hb991efa1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba220aaf),
	.w1(32'hba2496f8),
	.w2(32'h39a08b91),
	.w3(32'hba3a3e59),
	.w4(32'hba18f42f),
	.w5(32'hb966eebb),
	.w6(32'hba8039f9),
	.w7(32'hb9c14559),
	.w8(32'hb8761798),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bcc10),
	.w1(32'h3a8268fa),
	.w2(32'h3a22aca6),
	.w3(32'hb650dedd),
	.w4(32'hb89ba487),
	.w5(32'hb9c1f077),
	.w6(32'h3a820729),
	.w7(32'h3a047bce),
	.w8(32'hb8936a74),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39feb8d1),
	.w1(32'h3a45cf61),
	.w2(32'h3a8d50b9),
	.w3(32'h3881fee4),
	.w4(32'h3853722d),
	.w5(32'h398d6e30),
	.w6(32'h3a4f32a2),
	.w7(32'h3a50184c),
	.w8(32'h3a24be4a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e0dcc),
	.w1(32'hb9056f85),
	.w2(32'hb9c66771),
	.w3(32'h39ec30d2),
	.w4(32'hba023062),
	.w5(32'hb969ba99),
	.w6(32'hba04e2fb),
	.w7(32'hb93d3317),
	.w8(32'hb6996da3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38908e65),
	.w1(32'hbb0cc2e1),
	.w2(32'hba2e4d6d),
	.w3(32'h39fc6a63),
	.w4(32'hbb0fa783),
	.w5(32'hbaee2e69),
	.w6(32'hbb357654),
	.w7(32'hbae3bd9c),
	.w8(32'hb95f08fe),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6409ff),
	.w1(32'hbb37b40d),
	.w2(32'hbad8ac3c),
	.w3(32'h38ed1eaf),
	.w4(32'hbb2d12c9),
	.w5(32'hbb019f32),
	.w6(32'hbb203912),
	.w7(32'hbaf78c22),
	.w8(32'hb854da6f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39ef13),
	.w1(32'hb88c3896),
	.w2(32'h38c10e75),
	.w3(32'hb933a11a),
	.w4(32'hb9d6fc74),
	.w5(32'hba012b18),
	.w6(32'h3802874f),
	.w7(32'hb9bcf42a),
	.w8(32'hba13d7cf),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a248ae),
	.w1(32'h3a17d53f),
	.w2(32'h3a65769c),
	.w3(32'hb9a5e386),
	.w4(32'h390bda2b),
	.w5(32'h39cef138),
	.w6(32'h3a088418),
	.w7(32'h3a06189c),
	.w8(32'h3969c717),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fe6b1),
	.w1(32'h39e5de89),
	.w2(32'h3a9d5139),
	.w3(32'h39ae71e9),
	.w4(32'hb908e582),
	.w5(32'h3955b110),
	.w6(32'hb7866821),
	.w7(32'h3a5128bb),
	.w8(32'h3ab8270a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a989e2e),
	.w1(32'hb9b7c2cf),
	.w2(32'h3798152d),
	.w3(32'h3a1fd34e),
	.w4(32'hb799f518),
	.w5(32'hb7185fa6),
	.w6(32'h38ada795),
	.w7(32'hb79eff3b),
	.w8(32'hba6a3b10),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39236476),
	.w1(32'hb995fe5d),
	.w2(32'hba24a499),
	.w3(32'hb9a3df62),
	.w4(32'h391de044),
	.w5(32'h3a16e5fb),
	.w6(32'hb90b22f2),
	.w7(32'hba0c546a),
	.w8(32'hb9c3423d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8807748),
	.w1(32'h39b456f0),
	.w2(32'h39f7c5bd),
	.w3(32'h3a7ab315),
	.w4(32'hb97aac69),
	.w5(32'hb91494e5),
	.w6(32'h3a15d60d),
	.w7(32'h3a2297e6),
	.w8(32'h39914771),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394685bf),
	.w1(32'h396014df),
	.w2(32'hb8c6205a),
	.w3(32'h38aa2432),
	.w4(32'h3a88c3f2),
	.w5(32'h3a40a6a9),
	.w6(32'hba0447cf),
	.w7(32'hba00de80),
	.w8(32'hba37cce9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dbe84),
	.w1(32'hb9444a23),
	.w2(32'h395a577b),
	.w3(32'h3868d935),
	.w4(32'hb9817a5c),
	.w5(32'hba13e5e4),
	.w6(32'hba586ebb),
	.w7(32'hba2fa44e),
	.w8(32'hba6a5738),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b7e31),
	.w1(32'h38a32aa0),
	.w2(32'h36f45086),
	.w3(32'hba41b47b),
	.w4(32'hb8f787e8),
	.w5(32'hb98fc269),
	.w6(32'hb99c6312),
	.w7(32'hb9d385f7),
	.w8(32'hb9cdd1a5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fc01a),
	.w1(32'h3796bd00),
	.w2(32'hba15d611),
	.w3(32'hb9681a30),
	.w4(32'h39e6662f),
	.w5(32'h38dadf9e),
	.w6(32'hb95d528b),
	.w7(32'hba4fe8a9),
	.w8(32'hba696d6e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bcfd8),
	.w1(32'hbb266427),
	.w2(32'hbb1b8af0),
	.w3(32'hb96d4500),
	.w4(32'hbafb2d98),
	.w5(32'hbb0731bd),
	.w6(32'hbaa5b8d8),
	.w7(32'hbab84f7d),
	.w8(32'hb8e1cdbb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6f104),
	.w1(32'hba02aa49),
	.w2(32'hb9411e48),
	.w3(32'hbab9b65b),
	.w4(32'hba9aa731),
	.w5(32'hba342191),
	.w6(32'hba7eea53),
	.w7(32'hba7c351d),
	.w8(32'hba9587e7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66a8a4),
	.w1(32'h3a523012),
	.w2(32'h3a95c22c),
	.w3(32'hba3cfd8b),
	.w4(32'h3a393ee0),
	.w5(32'h3ab5bd55),
	.w6(32'h3a27b695),
	.w7(32'h3a413612),
	.w8(32'h3a0e832b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a851438),
	.w1(32'h3aef8035),
	.w2(32'h39853c14),
	.w3(32'h3a35c903),
	.w4(32'h3b2f98f6),
	.w5(32'h3a79ea43),
	.w6(32'h3ad82566),
	.w7(32'h39084105),
	.w8(32'h3a9f06e2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9893e9),
	.w1(32'h3a9c2aaf),
	.w2(32'h39fe7f90),
	.w3(32'h3af87512),
	.w4(32'h3a6491ce),
	.w5(32'h38ecdcc9),
	.w6(32'h3ae823eb),
	.w7(32'h3b0ca05f),
	.w8(32'h3aed8cc1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab32688),
	.w1(32'h3a9c5a06),
	.w2(32'h3a90ff76),
	.w3(32'hb9ef0d11),
	.w4(32'h39b12934),
	.w5(32'hb9f23cb5),
	.w6(32'h3a6106d3),
	.w7(32'h3a6ca12b),
	.w8(32'h39524001),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b9eb8),
	.w1(32'h3a4de738),
	.w2(32'hbb12d0aa),
	.w3(32'hba95a7ec),
	.w4(32'h3a8c6aa6),
	.w5(32'h3ae0ddfe),
	.w6(32'h3b13a7b1),
	.w7(32'h3ac11923),
	.w8(32'h3ab144d4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5699c7),
	.w1(32'hba284046),
	.w2(32'h3aab22e7),
	.w3(32'h3a5749c0),
	.w4(32'hbaaf4876),
	.w5(32'hba1d5062),
	.w6(32'hbaffcbc0),
	.w7(32'hba05d8b1),
	.w8(32'hb95f2168),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54cd6e),
	.w1(32'h3a753bc8),
	.w2(32'h3abe8a8a),
	.w3(32'h37cc9ba8),
	.w4(32'h3a1c5ee3),
	.w5(32'h3a9d7c7a),
	.w6(32'h3a7a6c4a),
	.w7(32'h3a669f30),
	.w8(32'h3a26c995),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fa732),
	.w1(32'hb781831f),
	.w2(32'hb9b92fc0),
	.w3(32'h3a27f874),
	.w4(32'hb91de2df),
	.w5(32'hba32e79e),
	.w6(32'hb9a5e5ce),
	.w7(32'hba5d5d89),
	.w8(32'hba43fa6a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afde66),
	.w1(32'h3a7692bf),
	.w2(32'h3a6a60c7),
	.w3(32'hb9fc5b95),
	.w4(32'h3a58a6ff),
	.w5(32'h39cc5494),
	.w6(32'h394a5d8a),
	.w7(32'hb9f89232),
	.w8(32'hb9fad2dc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f8107a),
	.w1(32'h39dabf6a),
	.w2(32'h3b2a2123),
	.w3(32'h38ad1997),
	.w4(32'hba395b8c),
	.w5(32'h3a2e71d9),
	.w6(32'hba6d7479),
	.w7(32'h3a7481b7),
	.w8(32'h39e9a0e3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7465d8),
	.w1(32'hb9bb8645),
	.w2(32'h39b5404f),
	.w3(32'hba648584),
	.w4(32'hba48b576),
	.w5(32'hba8f7e4d),
	.w6(32'hba29448b),
	.w7(32'hba7e73eb),
	.w8(32'hba389b6d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6849b0),
	.w1(32'h3ad6ba57),
	.w2(32'h3ad0f9be),
	.w3(32'hba86fb2c),
	.w4(32'h3ac21262),
	.w5(32'h396a838d),
	.w6(32'h3b1535d8),
	.w7(32'h3ad28395),
	.w8(32'h3a41c619),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f77c00),
	.w1(32'h39e72ba0),
	.w2(32'h380186c1),
	.w3(32'h39cf03d5),
	.w4(32'h39ddb16d),
	.w5(32'hb94d820e),
	.w6(32'h396f4d0e),
	.w7(32'hb872bb72),
	.w8(32'h386bdd59),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f37ea),
	.w1(32'hbb1acb48),
	.w2(32'hbaf1001b),
	.w3(32'h38ba38a3),
	.w4(32'hbafa6812),
	.w5(32'hbb03ac38),
	.w6(32'hbad990c1),
	.w7(32'hbae3bd0f),
	.w8(32'hb96d7a72),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabb263),
	.w1(32'hba6aeb47),
	.w2(32'h39443b1f),
	.w3(32'hb9d15e5d),
	.w4(32'hbaafe5fc),
	.w5(32'hbac553be),
	.w6(32'hba8cc619),
	.w7(32'hbaafad15),
	.w8(32'hba8e91da),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba284aa0),
	.w1(32'h3a3edef0),
	.w2(32'h3a9d1505),
	.w3(32'hbad92495),
	.w4(32'h3a60baab),
	.w5(32'h3aafbf55),
	.w6(32'h3a881a98),
	.w7(32'h3ac305b5),
	.w8(32'hba5e4392),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae727b2),
	.w1(32'hb9b538a7),
	.w2(32'hb9dbe9e6),
	.w3(32'hba8c6184),
	.w4(32'h388d9f52),
	.w5(32'hba01e551),
	.w6(32'hba34a4ea),
	.w7(32'hba367fc7),
	.w8(32'hba15fc49),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8705dc),
	.w1(32'hb8d94321),
	.w2(32'h3a561788),
	.w3(32'hba62c5d6),
	.w4(32'h3a0a90f2),
	.w5(32'h3a4a9137),
	.w6(32'h3a72dbc6),
	.w7(32'h3ab49b2a),
	.w8(32'h3a21a407),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920e117),
	.w1(32'hba414912),
	.w2(32'hba450c45),
	.w3(32'hb8eeabc9),
	.w4(32'hb987d8f7),
	.w5(32'hba756789),
	.w6(32'hb9f34a7b),
	.w7(32'hba8b5267),
	.w8(32'hba9083b5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6be8),
	.w1(32'h37d74357),
	.w2(32'hb9bea919),
	.w3(32'hba79d2d6),
	.w4(32'hb95332ab),
	.w5(32'hba22bed8),
	.w6(32'hb8fed73e),
	.w7(32'hba21bfa1),
	.w8(32'hba304f02),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9b467),
	.w1(32'h3a3f1554),
	.w2(32'h3a630e45),
	.w3(32'hba2dd89d),
	.w4(32'hb8a1ad06),
	.w5(32'h3a6bcb11),
	.w6(32'h3a299cce),
	.w7(32'h396dc0d7),
	.w8(32'hb71a4514),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ce246),
	.w1(32'h3aa46742),
	.w2(32'h38f7846a),
	.w3(32'hb9640e6f),
	.w4(32'h3aeee382),
	.w5(32'h3a4fb43a),
	.w6(32'h3a8ddec3),
	.w7(32'h394101d9),
	.w8(32'h3a79bdf1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7356ae),
	.w1(32'hb9c729ea),
	.w2(32'h372c5334),
	.w3(32'h3ac318c6),
	.w4(32'hb9bd59b9),
	.w5(32'h39821f82),
	.w6(32'hba06d4f5),
	.w7(32'h39ed45d3),
	.w8(32'h3a1ef329),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a730c0),
	.w1(32'hba1fcdcb),
	.w2(32'h3ab2551b),
	.w3(32'h39aa641b),
	.w4(32'h37be1503),
	.w5(32'h3a24ed4d),
	.w6(32'hba0afb4f),
	.w7(32'h38bdd0ad),
	.w8(32'hba291bba),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba833558),
	.w1(32'hbb501c22),
	.w2(32'hbad32b43),
	.w3(32'hba8340b8),
	.w4(32'hbb22d2ea),
	.w5(32'hbafc640f),
	.w6(32'hbb2a9b8f),
	.w7(32'hbb149a4e),
	.w8(32'hbad200f8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21672a),
	.w1(32'hba1ce497),
	.w2(32'hba20e781),
	.w3(32'hbb001f75),
	.w4(32'hba00ddb2),
	.w5(32'hba514911),
	.w6(32'hb9dfd44a),
	.w7(32'h39546195),
	.w8(32'hb92801d4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a24a9),
	.w1(32'h3823b7fa),
	.w2(32'h39fe10a4),
	.w3(32'hbaa623ae),
	.w4(32'hb9f4ede9),
	.w5(32'hba2d2d5c),
	.w6(32'hb9b7ae02),
	.w7(32'hb9f2b1fe),
	.w8(32'hba00d12e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba399b2f),
	.w1(32'h3aa7ffe7),
	.w2(32'h3afc927b),
	.w3(32'hba494333),
	.w4(32'h3ad45aeb),
	.w5(32'h3ad62d11),
	.w6(32'h3ab3f5a4),
	.w7(32'h3ac59bd8),
	.w8(32'h3a6da294),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ee02a),
	.w1(32'hb9725150),
	.w2(32'h359b6cd6),
	.w3(32'h398db1b4),
	.w4(32'hb9abbb4b),
	.w5(32'hb9899d66),
	.w6(32'hb9a872c5),
	.w7(32'hb9f4752f),
	.w8(32'hb9c7f797),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379d8f34),
	.w1(32'h3806f6b7),
	.w2(32'h39dbe2cf),
	.w3(32'hb94f403a),
	.w4(32'h38fd258d),
	.w5(32'h38bf50b3),
	.w6(32'h383d8cb1),
	.w7(32'hb8ada7ae),
	.w8(32'hb6e97a95),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395db41b),
	.w1(32'h390d4fd5),
	.w2(32'h3943e670),
	.w3(32'h38baee1b),
	.w4(32'hb8159de6),
	.w5(32'hb90dbd93),
	.w6(32'hb936e53e),
	.w7(32'hb97b1bc8),
	.w8(32'hb9553a15),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d18472),
	.w1(32'h3a6996b6),
	.w2(32'h3a8c087a),
	.w3(32'hb9c272de),
	.w4(32'h3a009bb6),
	.w5(32'h39e8c7d5),
	.w6(32'h3a1c2d5d),
	.w7(32'h3a25fe4e),
	.w8(32'h38a41a58),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89cb59),
	.w1(32'hba40c176),
	.w2(32'h39c871d6),
	.w3(32'h39a6855a),
	.w4(32'hba13cf9d),
	.w5(32'hb8e487a1),
	.w6(32'hba89195b),
	.w7(32'hba3c8f2a),
	.w8(32'h38e23947),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00fa0e),
	.w1(32'h3a078a6a),
	.w2(32'h3a086156),
	.w3(32'hb9ba917f),
	.w4(32'hba4f20dd),
	.w5(32'h3a0100e4),
	.w6(32'hb9c5c16a),
	.w7(32'h38c74585),
	.w8(32'h390c6f76),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba570de2),
	.w1(32'h3a0572a4),
	.w2(32'h360014f3),
	.w3(32'hba0993c2),
	.w4(32'h39a6eb92),
	.w5(32'hb92dd2cf),
	.w6(32'h3a00327e),
	.w7(32'hb9bae9eb),
	.w8(32'hb828e031),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7804d),
	.w1(32'hbad82f7f),
	.w2(32'hb9a4ae7c),
	.w3(32'h394ec59d),
	.w4(32'hbb0c142c),
	.w5(32'hbac1160b),
	.w6(32'hbb056e1b),
	.w7(32'hbae28142),
	.w8(32'hba9ef959),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d134a),
	.w1(32'h3a9797e4),
	.w2(32'hb9bcc31c),
	.w3(32'hba83bb4c),
	.w4(32'h3a453948),
	.w5(32'h3a6980c1),
	.w6(32'h3a65491f),
	.w7(32'hb977c919),
	.w8(32'h3a6659f3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3148d5),
	.w1(32'hb9a5a52e),
	.w2(32'hb9c71ac7),
	.w3(32'h3aa6394b),
	.w4(32'hba740946),
	.w5(32'hba97ca8f),
	.w6(32'h382488d5),
	.w7(32'hba1f9fc1),
	.w8(32'hba39fac5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba128dc4),
	.w1(32'hbaf55d34),
	.w2(32'hba4b352a),
	.w3(32'hbaaeeb8c),
	.w4(32'hbaa3de69),
	.w5(32'hba994a1d),
	.w6(32'hba77708e),
	.w7(32'hb8d05047),
	.w8(32'hb9d69bed),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7404f),
	.w1(32'hbadf9ee2),
	.w2(32'hba0b7251),
	.w3(32'hbaebc67f),
	.w4(32'hbae05f6d),
	.w5(32'hbae60749),
	.w6(32'hbb1fa8bb),
	.w7(32'hbb0032c5),
	.w8(32'hbaf156dd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac27223),
	.w1(32'hba398bc4),
	.w2(32'hb84fbed0),
	.w3(32'hbab9bfc0),
	.w4(32'hba5b0e19),
	.w5(32'hba8286ff),
	.w6(32'hba65d01a),
	.w7(32'hb9fef80a),
	.w8(32'hb91713f3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980b0ec),
	.w1(32'hba28fc35),
	.w2(32'hba2010df),
	.w3(32'hb97c551e),
	.w4(32'hb96bd429),
	.w5(32'hba61f3b1),
	.w6(32'hb9e94af8),
	.w7(32'hb95defcd),
	.w8(32'hb91eb534),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f30a4a),
	.w1(32'h3a0b7bb7),
	.w2(32'h3ab6523a),
	.w3(32'hba2175a1),
	.w4(32'hb94d3a6b),
	.w5(32'h39f11fcc),
	.w6(32'hb9462d02),
	.w7(32'hba58b30e),
	.w8(32'hba836c3d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d4393),
	.w1(32'hbac853ee),
	.w2(32'h39948065),
	.w3(32'hbaa20bac),
	.w4(32'hbacf98ef),
	.w5(32'hbaa152d9),
	.w6(32'hbad091ed),
	.w7(32'hba88f009),
	.w8(32'hba5427f2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c278d),
	.w1(32'hba3c6a2f),
	.w2(32'hb8d69b53),
	.w3(32'hbaa386a4),
	.w4(32'hb9c42b70),
	.w5(32'hb8fa1ea6),
	.w6(32'hba9be47b),
	.w7(32'hba93f313),
	.w8(32'hb969f7ae),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0210af),
	.w1(32'hb93bd299),
	.w2(32'hb701f5a9),
	.w3(32'h39ef1190),
	.w4(32'hb9d9f6fe),
	.w5(32'hba1b4151),
	.w6(32'hb90577bc),
	.w7(32'hb9b19978),
	.w8(32'hba12e74d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919d22d),
	.w1(32'h39505a7f),
	.w2(32'h39a00a59),
	.w3(32'hb9cf33c7),
	.w4(32'h399526aa),
	.w5(32'hb9cd0f26),
	.w6(32'h3925f27e),
	.w7(32'hb8172d8e),
	.w8(32'hb8293ef2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9976510),
	.w1(32'hb6c073ab),
	.w2(32'hb7245116),
	.w3(32'hb92fffac),
	.w4(32'hba480fed),
	.w5(32'hba2d532c),
	.w6(32'h389feb41),
	.w7(32'hb8f14b7b),
	.w8(32'hb9d1890b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da4f76),
	.w1(32'h3998adba),
	.w2(32'h3a5cef96),
	.w3(32'hba92ef11),
	.w4(32'h39cddf90),
	.w5(32'h39f2d95c),
	.w6(32'h3a11a4ae),
	.w7(32'h3a11b3bc),
	.w8(32'h3882c852),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd5bb2),
	.w1(32'h3944f7d9),
	.w2(32'h3a635aac),
	.w3(32'h369b51cb),
	.w4(32'hb7ebf822),
	.w5(32'hb8ff835c),
	.w6(32'h39841c5b),
	.w7(32'h39bf958f),
	.w8(32'h3942f805),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392134a2),
	.w1(32'hbabf6200),
	.w2(32'hba8045d8),
	.w3(32'h382ca67f),
	.w4(32'hbab0a771),
	.w5(32'hbab4a4c5),
	.w6(32'hbaaecb6e),
	.w7(32'hba9a0124),
	.w8(32'hba2c7b07),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9832e88),
	.w1(32'hbab05da8),
	.w2(32'hbaa3304b),
	.w3(32'hba086928),
	.w4(32'hba97c234),
	.w5(32'hbaae3e22),
	.w6(32'hbaad5058),
	.w7(32'hba582eba),
	.w8(32'h38e0d8f7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f5b4a),
	.w1(32'hb98e6a94),
	.w2(32'h39c05895),
	.w3(32'hba6bd202),
	.w4(32'hb98c8e8a),
	.w5(32'hb966c5ee),
	.w6(32'hba52d054),
	.w7(32'hba6365e5),
	.w8(32'hba8258dd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a6fc6),
	.w1(32'h38f58f86),
	.w2(32'h3a5566f1),
	.w3(32'hb9ef991e),
	.w4(32'h3a8d5d93),
	.w5(32'h3a4a0465),
	.w6(32'hb8fc4519),
	.w7(32'hba102954),
	.w8(32'h397c4c48),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ec421),
	.w1(32'h39f39de0),
	.w2(32'h3ad7d30a),
	.w3(32'h3a00649b),
	.w4(32'h39dec518),
	.w5(32'h3a98e257),
	.w6(32'h398c41ad),
	.w7(32'h3b136a35),
	.w8(32'h391d4f26),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cd871e),
	.w1(32'hb9d84f79),
	.w2(32'hbabe5a1f),
	.w3(32'h38fdfd59),
	.w4(32'hbac261ee),
	.w5(32'hba79a8e7),
	.w6(32'hba3bbbec),
	.w7(32'hbabf052c),
	.w8(32'hb9adf2fa),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a9966),
	.w1(32'hba160223),
	.w2(32'hb971d596),
	.w3(32'hba5c6e2b),
	.w4(32'hba2575c1),
	.w5(32'hba84556d),
	.w6(32'hbaa20e94),
	.w7(32'hbac0ec92),
	.w8(32'hbacf103f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa89758),
	.w1(32'hbaa29ec4),
	.w2(32'hb956e2aa),
	.w3(32'hba9052f1),
	.w4(32'hbad6f549),
	.w5(32'hbac3da09),
	.w6(32'hbab04969),
	.w7(32'hbaa2a59a),
	.w8(32'hba0ef1e8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba173dfd),
	.w1(32'h3aa16078),
	.w2(32'h3a98fbac),
	.w3(32'hba566beb),
	.w4(32'h39e5a917),
	.w5(32'h3ab61ab9),
	.w6(32'h3aba42d1),
	.w7(32'h3a2b8500),
	.w8(32'hb9dbb482),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57deb1),
	.w1(32'h3a4f7dfd),
	.w2(32'h3b4ffe1a),
	.w3(32'hb94e6c03),
	.w4(32'h3af3b4d3),
	.w5(32'h3b39732a),
	.w6(32'h3aed8d05),
	.w7(32'h3aec00ab),
	.w8(32'h3a2335a4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcf40a),
	.w1(32'h3a52630d),
	.w2(32'hb5cbaea2),
	.w3(32'hb9238282),
	.w4(32'h3a147898),
	.w5(32'hb934ba2f),
	.w6(32'h3a32a80f),
	.w7(32'hb9edeb6a),
	.w8(32'hb76a30ba),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d2e79),
	.w1(32'h36e5cb13),
	.w2(32'h39d3cb9a),
	.w3(32'h38f1952a),
	.w4(32'hb8ba3ee7),
	.w5(32'hb965e9e9),
	.w6(32'h39921ee1),
	.w7(32'h38cf5674),
	.w8(32'h3968cc5b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390860e6),
	.w1(32'h39da7f60),
	.w2(32'hb8ec54ac),
	.w3(32'hb9462b22),
	.w4(32'h39875993),
	.w5(32'hb91b9135),
	.w6(32'h39a33f98),
	.w7(32'hb99267d7),
	.w8(32'hb7f6909a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3d360),
	.w1(32'h3a1fcb4b),
	.w2(32'h3a6f4079),
	.w3(32'h38e6f160),
	.w4(32'hb9399ece),
	.w5(32'h39247e14),
	.w6(32'h3a15ea4b),
	.w7(32'h3a3b5a7d),
	.w8(32'h3a389d5a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e12180),
	.w1(32'hb9b02f77),
	.w2(32'h39f22ac9),
	.w3(32'h39ad84dd),
	.w4(32'hba792cf9),
	.w5(32'hba2c834f),
	.w6(32'hba6cea73),
	.w7(32'hba1845f6),
	.w8(32'hba870be7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bdeb6),
	.w1(32'hb9951693),
	.w2(32'h3766768a),
	.w3(32'hba7e4174),
	.w4(32'hb9d8b3a3),
	.w5(32'hba258780),
	.w6(32'hba07c8c4),
	.w7(32'hba389c7d),
	.w8(32'hba881e35),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5277a),
	.w1(32'h39c7099d),
	.w2(32'hb8737c29),
	.w3(32'hba17140c),
	.w4(32'h396f2e33),
	.w5(32'hb978ae33),
	.w6(32'h3997455f),
	.w7(32'hb9a02b94),
	.w8(32'hb92e5fc1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946411e),
	.w1(32'h37cf8c34),
	.w2(32'h3909c8d1),
	.w3(32'h3883cee7),
	.w4(32'h382c9a26),
	.w5(32'h395d572b),
	.w6(32'hba3b65c8),
	.w7(32'h39300473),
	.w8(32'h3a873fb8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbd63c),
	.w1(32'h39bc8e92),
	.w2(32'h3a33b19a),
	.w3(32'h39ea05dd),
	.w4(32'hb9b910b2),
	.w5(32'hba11b71f),
	.w6(32'hb937d677),
	.w7(32'hb8f30a3e),
	.w8(32'hba120013),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9e045),
	.w1(32'hba09eb99),
	.w2(32'hba6281e9),
	.w3(32'hba83de31),
	.w4(32'h3a428d5d),
	.w5(32'h3af5cffd),
	.w6(32'hba7d44d4),
	.w7(32'h3a024a91),
	.w8(32'h3b2169c8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f690f),
	.w1(32'h388e5eff),
	.w2(32'h39a56720),
	.w3(32'h3a81cec1),
	.w4(32'hba5fa61e),
	.w5(32'hba86c3e3),
	.w6(32'hb98afdd8),
	.w7(32'hb9dce302),
	.w8(32'hb99f2727),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0663f0),
	.w1(32'hba973ef2),
	.w2(32'hb9989b14),
	.w3(32'hba988d1c),
	.w4(32'hba6f41b2),
	.w5(32'hba036c5a),
	.w6(32'hbab094ea),
	.w7(32'hba91281c),
	.w8(32'hba97f5e5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f07056),
	.w1(32'h3a2418ce),
	.w2(32'h3a2c4d7f),
	.w3(32'hba516207),
	.w4(32'hb91feff5),
	.w5(32'hba13773d),
	.w6(32'h3a2352bb),
	.w7(32'h393223aa),
	.w8(32'hb9cacc72),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ce105),
	.w1(32'h3a185717),
	.w2(32'hb8f837a1),
	.w3(32'hb984dd75),
	.w4(32'h39be2536),
	.w5(32'hb9909160),
	.w6(32'h39e951f8),
	.w7(32'hb9ddbc25),
	.w8(32'hb90c8161),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bee0ce),
	.w1(32'hb9860bbd),
	.w2(32'hb9941670),
	.w3(32'h39557623),
	.w4(32'hb99c4a70),
	.w5(32'hb9945ec8),
	.w6(32'hb968a8ba),
	.w7(32'hb9e103e2),
	.w8(32'hb9f7b0aa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9281864),
	.w1(32'hb98802ec),
	.w2(32'hb9e23761),
	.w3(32'hb999b55b),
	.w4(32'hb9d46d7a),
	.w5(32'hb9c31fec),
	.w6(32'hb9b22ba6),
	.w7(32'hba262bac),
	.w8(32'hb9eea4f4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9582900),
	.w1(32'h3a9bf3eb),
	.w2(32'hb97d793e),
	.w3(32'hb9110b6c),
	.w4(32'h3ae073d7),
	.w5(32'h3a87d037),
	.w6(32'h39c4426a),
	.w7(32'h38f1ccdf),
	.w8(32'h3ab93ba2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac40505),
	.w1(32'h3a0193a9),
	.w2(32'h39bd2036),
	.w3(32'h3a0eff75),
	.w4(32'h3974df5e),
	.w5(32'hba1285f8),
	.w6(32'hb94651b4),
	.w7(32'hba503738),
	.w8(32'hba845077),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46d6f),
	.w1(32'h3a484fa2),
	.w2(32'h3abac537),
	.w3(32'hba9b3978),
	.w4(32'hb6f427a5),
	.w5(32'h38f6777e),
	.w6(32'h3a6f4de0),
	.w7(32'h3a297641),
	.w8(32'h39e77839),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867466),
	.w1(32'h39011e2c),
	.w2(32'h3a85f6f2),
	.w3(32'h3994abe8),
	.w4(32'hb8053719),
	.w5(32'h393a6061),
	.w6(32'h38ef8f4c),
	.w7(32'h391f2080),
	.w8(32'h3a143358),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6da25),
	.w1(32'h3947c3f5),
	.w2(32'hb8f8b349),
	.w3(32'h3a265764),
	.w4(32'hb80029dc),
	.w5(32'hb99b1d2e),
	.w6(32'hb840e3b3),
	.w7(32'hb9fc7d06),
	.w8(32'hb9e6dfca),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9591407),
	.w1(32'h3a9f2c2a),
	.w2(32'h3a045c75),
	.w3(32'hb9eaac27),
	.w4(32'h3b720be8),
	.w5(32'h3b129862),
	.w6(32'h3aa98ceb),
	.w7(32'h3b1fb429),
	.w8(32'h3ae70fe5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f81249),
	.w1(32'hba9b695d),
	.w2(32'hb980ef41),
	.w3(32'h3a095259),
	.w4(32'hba85fe4e),
	.w5(32'hbab62ef6),
	.w6(32'hba7d6d5d),
	.w7(32'hbabc7f96),
	.w8(32'hba7407f4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba110dbf),
	.w1(32'hb882d6bd),
	.w2(32'hb88676ee),
	.w3(32'hba792802),
	.w4(32'hb9ed3987),
	.w5(32'hba2b9b02),
	.w6(32'hb92dbe29),
	.w7(32'hba29573d),
	.w8(32'hb9c32067),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3713ba57),
	.w1(32'hbe72bafc),
	.w2(32'hbf114bae),
	.w3(32'hb8fa66e1),
	.w4(32'hbe88af6b),
	.w5(32'h3f21f0e8),
	.w6(32'hbed3ce6f),
	.w7(32'hbf20d78f),
	.w8(32'hbf111b4c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeb909e2),
	.w1(32'hbefeb932),
	.w2(32'hbf1a81cc),
	.w3(32'hbeb6e9b9),
	.w4(32'hbecbeb38),
	.w5(32'h3e4fe621),
	.w6(32'hbeb150bb),
	.w7(32'hbeadbff2),
	.w8(32'hbefe903d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule