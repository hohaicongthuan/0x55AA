module layer_8_featuremap_163(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbc899),
	.w1(32'h3cb8a8c3),
	.w2(32'hbb577e1c),
	.w3(32'hbbc55f9f),
	.w4(32'h3b06685d),
	.w5(32'h3ca1f687),
	.w6(32'hbbe89a85),
	.w7(32'h3bc86195),
	.w8(32'h3c1ff8d6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61f887),
	.w1(32'hbb0f0c3e),
	.w2(32'hba241bab),
	.w3(32'h3cce7550),
	.w4(32'hbb0b28cc),
	.w5(32'hbaa7fa76),
	.w6(32'hba59d647),
	.w7(32'h3a9e3fd0),
	.w8(32'h39fa7944),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba229445),
	.w1(32'hbbac99b7),
	.w2(32'hbc8530b4),
	.w3(32'hbb2c9e73),
	.w4(32'hbc21246c),
	.w5(32'h39c9dceb),
	.w6(32'hbc379b81),
	.w7(32'hb8312cbf),
	.w8(32'hbb635af6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb83199),
	.w1(32'hbbc8fcde),
	.w2(32'hbd15ebc8),
	.w3(32'hbb9d360e),
	.w4(32'h3ca48f8f),
	.w5(32'h3cdf79b6),
	.w6(32'hbc7ae08a),
	.w7(32'h3c0760b2),
	.w8(32'hbb38dcc2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a759a),
	.w1(32'hba8d3c46),
	.w2(32'h3aa16c64),
	.w3(32'hbc1397d8),
	.w4(32'hbb600aa3),
	.w5(32'hbb9409ed),
	.w6(32'hba2a4a8d),
	.w7(32'hbb563a5f),
	.w8(32'hbb0d481e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ecbf),
	.w1(32'hbc161073),
	.w2(32'h3c43858e),
	.w3(32'hbc039cb3),
	.w4(32'h3b8dfb57),
	.w5(32'hbc2637d3),
	.w6(32'hbacdc88f),
	.w7(32'hbb2094e9),
	.w8(32'hbb0e732f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ff4b0),
	.w1(32'hb99be2f9),
	.w2(32'h3a7b19a9),
	.w3(32'h3aec91d8),
	.w4(32'hb9aba33e),
	.w5(32'hbb389ee2),
	.w6(32'h3afca273),
	.w7(32'hba8909ed),
	.w8(32'hbb29000f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b33a1),
	.w1(32'h3c482972),
	.w2(32'hbc72ed4a),
	.w3(32'hbb46f333),
	.w4(32'hbb85320e),
	.w5(32'h3c6e9693),
	.w6(32'hbc980816),
	.w7(32'hbba5c7c9),
	.w8(32'h3c0f3ff7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d5fcb),
	.w1(32'hb87f1a09),
	.w2(32'h3beff132),
	.w3(32'h3cc2f2c0),
	.w4(32'hbada5c59),
	.w5(32'hb88268e0),
	.w6(32'h3b9643c4),
	.w7(32'h3bae62ee),
	.w8(32'h3b879ad1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb11600),
	.w1(32'hbc9c58eb),
	.w2(32'h3d2c68d8),
	.w3(32'hbbcef06c),
	.w4(32'h3b022133),
	.w5(32'hbd3db6f2),
	.w6(32'h3cb324a5),
	.w7(32'h3b6a92e7),
	.w8(32'hbc97ebde),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d66dbd1),
	.w1(32'hbc4a9fbd),
	.w2(32'hbd270afc),
	.w3(32'hbcdd20a3),
	.w4(32'h3c3aa2b3),
	.w5(32'h3ce2421b),
	.w6(32'hbc69ea97),
	.w7(32'h3c1a22bb),
	.w8(32'h3c628d74),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc954631),
	.w1(32'h3a76656a),
	.w2(32'hbb369a0b),
	.w3(32'hbb4f751e),
	.w4(32'hbb89c6eb),
	.w5(32'hbadcf591),
	.w6(32'hba6790b6),
	.w7(32'h3b70e91b),
	.w8(32'h3a1d1b2b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd838d),
	.w1(32'hbc04b59e),
	.w2(32'h3c87026b),
	.w3(32'h3b198cb4),
	.w4(32'h391869c4),
	.w5(32'hbc9fabbe),
	.w6(32'h3b84f626),
	.w7(32'h3c0d702b),
	.w8(32'h3a9c225b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03de15),
	.w1(32'h3ce7416c),
	.w2(32'h3cec1554),
	.w3(32'hbb81c981),
	.w4(32'hbca7fbe2),
	.w5(32'hbb2d7a25),
	.w6(32'hbc8e5be7),
	.w7(32'hbcd5e3e6),
	.w8(32'hbb315bd3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6ed85),
	.w1(32'h39e9d6bf),
	.w2(32'h3b6da2dc),
	.w3(32'h3cda17cd),
	.w4(32'hbb1650d2),
	.w5(32'hbad423b0),
	.w6(32'h3b280790),
	.w7(32'hba6dcdf3),
	.w8(32'hbb19c81f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56bb7),
	.w1(32'hbbb1ba0a),
	.w2(32'hbbdbc03d),
	.w3(32'hb94ad86c),
	.w4(32'hbc4f1718),
	.w5(32'h3c0b569a),
	.w6(32'hbbc237a3),
	.w7(32'h3b556216),
	.w8(32'h3bce26e1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab90c3),
	.w1(32'hbab3dc30),
	.w2(32'hb9c64710),
	.w3(32'hbb5b4dac),
	.w4(32'h3d082962),
	.w5(32'h3ca2d560),
	.w6(32'h3caea189),
	.w7(32'h3c7c8f48),
	.w8(32'h3ad31f55),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d67f5),
	.w1(32'hbbd511f6),
	.w2(32'hbc632c5c),
	.w3(32'hbbde47a5),
	.w4(32'hbc14a097),
	.w5(32'hbc22a558),
	.w6(32'h3bd82d41),
	.w7(32'h3b80e6a1),
	.w8(32'h3b67d2c7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba511374),
	.w1(32'h3b1fe27f),
	.w2(32'h3c21e524),
	.w3(32'hbb863c00),
	.w4(32'hbba91c6d),
	.w5(32'hbba73b45),
	.w6(32'h3c008f4d),
	.w7(32'hbc08dbbb),
	.w8(32'hbb910351),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34447c),
	.w1(32'hbab864bd),
	.w2(32'hb899dee5),
	.w3(32'h3c031549),
	.w4(32'h3a8962de),
	.w5(32'hbb1da1dc),
	.w6(32'h3b1fe619),
	.w7(32'hbafe7828),
	.w8(32'hbb661f94),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c16dfa),
	.w1(32'h3c35fe57),
	.w2(32'h3c00d752),
	.w3(32'hbb6b7d79),
	.w4(32'hbc9a83a8),
	.w5(32'hbb793266),
	.w6(32'hbb695e66),
	.w7(32'hbbfee658),
	.w8(32'hbbb9e27e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820844),
	.w1(32'hbc9b61f7),
	.w2(32'hbc6af25e),
	.w3(32'h3b4df556),
	.w4(32'h3b8ff4cf),
	.w5(32'h3ab8517a),
	.w6(32'hbb6359bd),
	.w7(32'h3b0eb09d),
	.w8(32'hbb62b992),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f15bd),
	.w1(32'hbc86fd20),
	.w2(32'hbbddebad),
	.w3(32'hbbed8098),
	.w4(32'hbaf53739),
	.w5(32'h3b4f445b),
	.w6(32'h3b532fa9),
	.w7(32'h3aaa4f89),
	.w8(32'hba7aaf04),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab9229),
	.w1(32'hbc039828),
	.w2(32'hbbb47b02),
	.w3(32'h3bf77e5b),
	.w4(32'h3ba1a92c),
	.w5(32'hbc28684a),
	.w6(32'hbc2cd17a),
	.w7(32'hbbc9618e),
	.w8(32'hbc1184cd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a0a3),
	.w1(32'h39f1f2de),
	.w2(32'hbb30c5b9),
	.w3(32'hbc0fe187),
	.w4(32'hbc60ff37),
	.w5(32'hbbb260ea),
	.w6(32'h3b0c260b),
	.w7(32'h3b00c342),
	.w8(32'h3b4a9c1d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec25b7),
	.w1(32'h3b8994ce),
	.w2(32'h3b2f961e),
	.w3(32'h3b66dae1),
	.w4(32'hbba04e0c),
	.w5(32'hbc52fc0e),
	.w6(32'hbbf02f5d),
	.w7(32'hbc7423fa),
	.w8(32'hbbadd29b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a887590),
	.w1(32'h3acefd2d),
	.w2(32'hbc50c6ae),
	.w3(32'hbc0a7f06),
	.w4(32'h3cac1790),
	.w5(32'h3d09657e),
	.w6(32'hba4608f9),
	.w7(32'h3caa12d7),
	.w8(32'h3cdcdc36),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cba87),
	.w1(32'hbae8b94f),
	.w2(32'hbc9f47a3),
	.w3(32'h3c4ab3d6),
	.w4(32'h3b9d52aa),
	.w5(32'h3c1b0650),
	.w6(32'hbb84f266),
	.w7(32'h3ad8fd91),
	.w8(32'h3c5ae404),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075bd3),
	.w1(32'h3b9f2b7d),
	.w2(32'h3bc6b535),
	.w3(32'hbc20003c),
	.w4(32'h3acf6bec),
	.w5(32'h3bcbc407),
	.w6(32'h39874e60),
	.w7(32'h3b265e9b),
	.w8(32'h3b344407),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a893b0d),
	.w1(32'hbacbe62c),
	.w2(32'hba3d1218),
	.w3(32'h3b424e3c),
	.w4(32'hbbf3c3cd),
	.w5(32'hbba94559),
	.w6(32'h388cb944),
	.w7(32'hbb026c70),
	.w8(32'hba3680a9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a182753),
	.w1(32'h3be43c3e),
	.w2(32'h3a401224),
	.w3(32'hbb86157c),
	.w4(32'hbb8ed4f6),
	.w5(32'h3b2bc149),
	.w6(32'hb9c912ca),
	.w7(32'hbb3b6840),
	.w8(32'h3b724ef9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012fe0),
	.w1(32'h39e16f33),
	.w2(32'h3ba353c4),
	.w3(32'h3bdee30c),
	.w4(32'hba7f5655),
	.w5(32'hbbe31cb3),
	.w6(32'h3b93f2d9),
	.w7(32'h3b079a70),
	.w8(32'hbb683588),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47e18d),
	.w1(32'h3b980373),
	.w2(32'h3caef5f1),
	.w3(32'hbc1a8fca),
	.w4(32'hbc284626),
	.w5(32'h3c878b72),
	.w6(32'h3c15a16f),
	.w7(32'h3b02e20c),
	.w8(32'hb98def29),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348790),
	.w1(32'h3beb9aff),
	.w2(32'h3bc08870),
	.w3(32'h3c0260bf),
	.w4(32'hbc301d0b),
	.w5(32'hbba56d79),
	.w6(32'h3a566d77),
	.w7(32'hbc788d38),
	.w8(32'hbad26b45),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9c185),
	.w1(32'h3b540b42),
	.w2(32'h39766354),
	.w3(32'h3c0c8f64),
	.w4(32'hbb0f15cc),
	.w5(32'hbb1b751e),
	.w6(32'h3abba178),
	.w7(32'hb917ab6c),
	.w8(32'hbad0c1cc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b682faa),
	.w1(32'hbbfcd3c5),
	.w2(32'hbbeb73ff),
	.w3(32'hba841c83),
	.w4(32'h3b78a5e9),
	.w5(32'hbc0a0761),
	.w6(32'h3bf9e98e),
	.w7(32'h3ba489d6),
	.w8(32'h3c4aed1e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c41f3),
	.w1(32'hbb468d94),
	.w2(32'hbb263c57),
	.w3(32'h3b7c7393),
	.w4(32'h3b892d10),
	.w5(32'hba8682ad),
	.w6(32'h3a9a6221),
	.w7(32'h3b90246a),
	.w8(32'h3bc3e2c0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9878),
	.w1(32'hbb323a3a),
	.w2(32'h3ad6524e),
	.w3(32'hbb213e5e),
	.w4(32'hbae2aa8f),
	.w5(32'hb68b28bb),
	.w6(32'h3b0115a5),
	.w7(32'hbae51327),
	.w8(32'hbaf4635e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b6ee),
	.w1(32'hbb6aaa13),
	.w2(32'hbb7932d6),
	.w3(32'hbb92d9f0),
	.w4(32'h3b0b914e),
	.w5(32'hbb284a6a),
	.w6(32'h3af4cd30),
	.w7(32'h3ba2f8c2),
	.w8(32'hbb99149f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c016a12),
	.w1(32'hbc111a0f),
	.w2(32'hbb90c798),
	.w3(32'hbac75c11),
	.w4(32'h3b305ba4),
	.w5(32'hbbf60188),
	.w6(32'hbba2689a),
	.w7(32'h391369aa),
	.w8(32'hbc57f463),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd03bc),
	.w1(32'h39bc9bde),
	.w2(32'hbb7e415d),
	.w3(32'hbc18bcf0),
	.w4(32'h3b460ab9),
	.w5(32'hba95f63e),
	.w6(32'h3b9a7d1b),
	.w7(32'hb8a65c52),
	.w8(32'h3aac95d6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8b7b5),
	.w1(32'h3ba9c219),
	.w2(32'h3a85f696),
	.w3(32'hba860541),
	.w4(32'h3afc20b8),
	.w5(32'hbb5f64b8),
	.w6(32'h3bbb1013),
	.w7(32'hbb389e23),
	.w8(32'hbb1d0747),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad7ac0),
	.w1(32'h3b964a17),
	.w2(32'hbc1d42a5),
	.w3(32'h3c23eb63),
	.w4(32'h3b717984),
	.w5(32'h3b3dc14a),
	.w6(32'h3a6e9185),
	.w7(32'h3aea7ceb),
	.w8(32'h3bca246a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb01f7),
	.w1(32'hbc8770f4),
	.w2(32'hbba96e4d),
	.w3(32'h3b2f76a4),
	.w4(32'h3b3e7a8c),
	.w5(32'hbc7703ec),
	.w6(32'h3c4d7dcd),
	.w7(32'h3c818487),
	.w8(32'h3c3ecf01),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71b8a2),
	.w1(32'h3c281fd7),
	.w2(32'h3be5b28a),
	.w3(32'hbbd7ffea),
	.w4(32'hbc5dbb50),
	.w5(32'h3bd5345d),
	.w6(32'hbc3f95a8),
	.w7(32'hbc03ab67),
	.w8(32'hbbe08dcf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc433bcf),
	.w1(32'hbb3c4d88),
	.w2(32'hba8fd23e),
	.w3(32'h3c70a4f5),
	.w4(32'hbafed93e),
	.w5(32'hbbc1e03d),
	.w6(32'h38c3dc97),
	.w7(32'hbab2cba8),
	.w8(32'hbb4f515e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48fab),
	.w1(32'hbb0aa82b),
	.w2(32'hbaa73595),
	.w3(32'hbbc9b46d),
	.w4(32'h3aad4f66),
	.w5(32'hbbb647b6),
	.w6(32'hbbc10e29),
	.w7(32'hbc0b6302),
	.w8(32'hbc140c99),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2b2a),
	.w1(32'hbbb4039c),
	.w2(32'hbc03f6a8),
	.w3(32'hbbe7c977),
	.w4(32'h3b9038f6),
	.w5(32'hbc6b2d46),
	.w6(32'h3b976284),
	.w7(32'h3c94da83),
	.w8(32'h3c73e6ff),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a554f),
	.w1(32'hbc41e04e),
	.w2(32'hbc8a2264),
	.w3(32'hbba5f671),
	.w4(32'hbb63fdc4),
	.w5(32'hbbf1eab5),
	.w6(32'h3c2dd025),
	.w7(32'h3c4c2cd4),
	.w8(32'h3c2c305a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f166),
	.w1(32'hbb260a88),
	.w2(32'hbbb88cb4),
	.w3(32'hbc2a85f7),
	.w4(32'h3b5e84a0),
	.w5(32'hbadb67fb),
	.w6(32'hba8f08bf),
	.w7(32'hbc057513),
	.w8(32'hbb637be1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bba2a),
	.w1(32'hb9beaf6f),
	.w2(32'h3b9bfc69),
	.w3(32'hbc40a3b7),
	.w4(32'h3acc9d49),
	.w5(32'h3bab6876),
	.w6(32'h3b1db880),
	.w7(32'h3bc32b25),
	.w8(32'h3b6726d7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36c91b),
	.w1(32'hba9c6849),
	.w2(32'hbb84a934),
	.w3(32'h3a128e01),
	.w4(32'hba7d7481),
	.w5(32'hbb9ccaee),
	.w6(32'h3b9278dd),
	.w7(32'h3a02e0c4),
	.w8(32'hbb1495a6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a7d3),
	.w1(32'hb983787f),
	.w2(32'h3b06759b),
	.w3(32'hbb9b98ca),
	.w4(32'hbaf0edfb),
	.w5(32'hba42df7d),
	.w6(32'h3af50d9e),
	.w7(32'h3b22af96),
	.w8(32'h39d3921f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192986),
	.w1(32'hbb2e36db),
	.w2(32'hbc79c52a),
	.w3(32'h3924ea28),
	.w4(32'hbbbba505),
	.w5(32'hbc65b873),
	.w6(32'h3af339a8),
	.w7(32'h3aad9cbe),
	.w8(32'hbb66497f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd661a),
	.w1(32'hbba2f2fe),
	.w2(32'h3bf2e1f0),
	.w3(32'hbc336f07),
	.w4(32'hbade2809),
	.w5(32'hbc4cde47),
	.w6(32'h3c1ba1b7),
	.w7(32'hbb8fd788),
	.w8(32'hbbadd74c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab71195),
	.w1(32'hbc62b8f3),
	.w2(32'hbc8387de),
	.w3(32'hbb401aac),
	.w4(32'hbc2a69a7),
	.w5(32'hbc8665fc),
	.w6(32'h3c0e40eb),
	.w7(32'h3bca34eb),
	.w8(32'h3ad805d7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c8a7e),
	.w1(32'hbbfad37d),
	.w2(32'h3c1d7c77),
	.w3(32'hbb52eea5),
	.w4(32'hbb671a6a),
	.w5(32'hbb3f1458),
	.w6(32'h3bc0cd11),
	.w7(32'hba955e85),
	.w8(32'hbbb235c3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6829e3),
	.w1(32'hbb562f18),
	.w2(32'hbb745bf3),
	.w3(32'h3b850ea4),
	.w4(32'h3b20b5f5),
	.w5(32'hbb9e218b),
	.w6(32'h3a71f70d),
	.w7(32'h3b1790c1),
	.w8(32'h3be46efd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0739a),
	.w1(32'h3b519f05),
	.w2(32'hba094f53),
	.w3(32'h3b6b9b9a),
	.w4(32'h3aa9fb2b),
	.w5(32'h3a5eaea2),
	.w6(32'h3aa43d79),
	.w7(32'hb808b022),
	.w8(32'h3874eb88),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad30c5a),
	.w1(32'hbca63bbb),
	.w2(32'hbc1849e0),
	.w3(32'h3972542f),
	.w4(32'hbc770075),
	.w5(32'hbc465b35),
	.w6(32'hbba4202c),
	.w7(32'hbc567860),
	.w8(32'hbc060531),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bee3d),
	.w1(32'hbb96c71c),
	.w2(32'hba98690c),
	.w3(32'hbc3a0bc7),
	.w4(32'h3a5eeb19),
	.w5(32'hbb63cd5e),
	.w6(32'h3b34de56),
	.w7(32'h3b790b1e),
	.w8(32'hbb1022e4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5d1e2),
	.w1(32'hba9e1bc7),
	.w2(32'hbb1e8e42),
	.w3(32'h3bedf9ee),
	.w4(32'h3c0c1000),
	.w5(32'h3be7b434),
	.w6(32'h3b3fe164),
	.w7(32'h3b274a2e),
	.w8(32'h3c0bc6d0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8482e8),
	.w1(32'hbad7075c),
	.w2(32'h3a2a0ffe),
	.w3(32'hbc1da286),
	.w4(32'h3b465bdc),
	.w5(32'h39283ed0),
	.w6(32'h3b15d9e7),
	.w7(32'h3b09b510),
	.w8(32'h3a22b7d7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcdffb),
	.w1(32'h3c023d55),
	.w2(32'h3b8ccc63),
	.w3(32'hbbb008d2),
	.w4(32'h3b27dfac),
	.w5(32'h3a450242),
	.w6(32'h3bcf0f66),
	.w7(32'h3aea8f7e),
	.w8(32'h39cd3867),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a5a44),
	.w1(32'h3b361cc7),
	.w2(32'h3b7f52cd),
	.w3(32'h3b18d403),
	.w4(32'h3b3410f1),
	.w5(32'h3b2647bc),
	.w6(32'h3b89a721),
	.w7(32'h3b8d8e9b),
	.w8(32'h3b3a8327),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27bff7),
	.w1(32'h3a166a69),
	.w2(32'h3aa4c84c),
	.w3(32'h3b7f3d3b),
	.w4(32'h3b6fead9),
	.w5(32'h398b39dd),
	.w6(32'hbad733d3),
	.w7(32'hbb8a56ae),
	.w8(32'hbb114b8b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821d37),
	.w1(32'h3b97b6ee),
	.w2(32'hbbf7b3a9),
	.w3(32'hbb91a2ca),
	.w4(32'hbc6aabc7),
	.w5(32'hbcbdc8c3),
	.w6(32'hbc6c235e),
	.w7(32'hbc78359b),
	.w8(32'hbbac6aca),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3ef52),
	.w1(32'hbc0072db),
	.w2(32'hbbc4bb33),
	.w3(32'hbc434a5d),
	.w4(32'hbad4a4e4),
	.w5(32'hb914f8ea),
	.w6(32'hbbc71528),
	.w7(32'hbbba93af),
	.w8(32'hbb2c8c8c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb703c7c),
	.w1(32'h3be2e9fa),
	.w2(32'h3b99dd41),
	.w3(32'hbb06046e),
	.w4(32'hbc998da4),
	.w5(32'hbbaff3f4),
	.w6(32'h3b3bb69b),
	.w7(32'hbc869acb),
	.w8(32'h3731ec52),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd064c74),
	.w1(32'hbbd28db7),
	.w2(32'hbbcb59df),
	.w3(32'h3befe5dc),
	.w4(32'hbc245810),
	.w5(32'hbc7a0148),
	.w6(32'h3b10939a),
	.w7(32'hbb437029),
	.w8(32'hbc1fbb66),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfecba6),
	.w1(32'hbaaac007),
	.w2(32'h3bcf4025),
	.w3(32'hbc1db446),
	.w4(32'h3bf0d93d),
	.w5(32'h3a3c5d4a),
	.w6(32'h3c580484),
	.w7(32'h3b58e3f0),
	.w8(32'hba191a76),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4406bc),
	.w1(32'h3c16c4dd),
	.w2(32'h3b8beee8),
	.w3(32'hbbabfefe),
	.w4(32'hbcdd97a5),
	.w5(32'hbc1a2ce6),
	.w6(32'hbc290e36),
	.w7(32'hbbe11af2),
	.w8(32'h3b844ec2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc612e08),
	.w1(32'hbb874496),
	.w2(32'hbc3c82fa),
	.w3(32'h3c4812e4),
	.w4(32'hbcc8aa26),
	.w5(32'hbc9c7a6d),
	.w6(32'hbb7ae406),
	.w7(32'h3bfae246),
	.w8(32'h3cbd1dab),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2659b9),
	.w1(32'hbc4b7e7f),
	.w2(32'h3b6b0964),
	.w3(32'hbb09630a),
	.w4(32'hbbc8c867),
	.w5(32'hbbbb014d),
	.w6(32'hbab671d8),
	.w7(32'h3bbb376c),
	.w8(32'h3b60047a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90819f),
	.w1(32'hbb8c12f0),
	.w2(32'hbbb39943),
	.w3(32'h3b13c16c),
	.w4(32'hbb816543),
	.w5(32'hbb075633),
	.w6(32'h3ba09cce),
	.w7(32'h3a8a8a28),
	.w8(32'h3bb0a793),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85964d),
	.w1(32'hbc7e4d5a),
	.w2(32'hbbb8b38f),
	.w3(32'h3b3429be),
	.w4(32'hbae822d9),
	.w5(32'hbc65ef3d),
	.w6(32'h3bac1358),
	.w7(32'h3ba510e5),
	.w8(32'h3a177f41),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf268e),
	.w1(32'hbb95eafe),
	.w2(32'hb9faa26b),
	.w3(32'hbc23de09),
	.w4(32'h3acf99d3),
	.w5(32'h3b508389),
	.w6(32'h3b4d1c5b),
	.w7(32'h39f1522c),
	.w8(32'hbb69b001),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372bd21d),
	.w1(32'h3a5b3c65),
	.w2(32'hbb528c0b),
	.w3(32'hb9ed8a81),
	.w4(32'h3ac483e3),
	.w5(32'hbab6902d),
	.w6(32'hbb313d82),
	.w7(32'hbb3253cc),
	.w8(32'hbb0d836d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c5a7),
	.w1(32'h3b9ffeae),
	.w2(32'h3b40ab2a),
	.w3(32'hbb499123),
	.w4(32'hbbe1b5ab),
	.w5(32'h3a25777d),
	.w6(32'hbbdc3f87),
	.w7(32'hbb22a939),
	.w8(32'h3baa8598),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad36eb),
	.w1(32'hba5fe60f),
	.w2(32'hbc632796),
	.w3(32'h3c3c590e),
	.w4(32'hbc4651ed),
	.w5(32'hbb6840f0),
	.w6(32'h3bbab8c2),
	.w7(32'hbbb794f0),
	.w8(32'h3b2f69fe),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3dab6),
	.w1(32'h3c9c2b21),
	.w2(32'h3c674d68),
	.w3(32'hbc0b0b47),
	.w4(32'hbb61bb76),
	.w5(32'h3cbbc9e8),
	.w6(32'hbbd6a3b8),
	.w7(32'hbbfb4183),
	.w8(32'h3bc500a0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc578a7e),
	.w1(32'h3cf8ead6),
	.w2(32'h3d0cbce7),
	.w3(32'h3cc69001),
	.w4(32'hbca8e907),
	.w5(32'h3b9035b2),
	.w6(32'h39c980de),
	.w7(32'hbc8d4b79),
	.w8(32'hbc3c2178),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f4597),
	.w1(32'hbc25edd4),
	.w2(32'h3bed8625),
	.w3(32'h3cc58062),
	.w4(32'h3bcf0d94),
	.w5(32'hbb9e32ed),
	.w6(32'h3c0dcfbf),
	.w7(32'h3b7d8d3a),
	.w8(32'h391f3b8b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca506c2),
	.w1(32'h3bed0263),
	.w2(32'h3c510f67),
	.w3(32'hbbe64469),
	.w4(32'hbb71dc27),
	.w5(32'hbbe895af),
	.w6(32'h3ba497ca),
	.w7(32'hbae3e822),
	.w8(32'hbbd3d6aa),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53f2fb),
	.w1(32'h3ceb902f),
	.w2(32'hb8477180),
	.w3(32'hbbaad170),
	.w4(32'hbc57251d),
	.w5(32'h3c81cd5c),
	.w6(32'hbcb86045),
	.w7(32'hbc9b4f4d),
	.w8(32'hbb27822b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf67098),
	.w1(32'h3c1d3f94),
	.w2(32'hbbdf0e84),
	.w3(32'h3ca06da2),
	.w4(32'hbc0d3635),
	.w5(32'hbb9878c0),
	.w6(32'hbc0de2e6),
	.w7(32'hbbfe16de),
	.w8(32'h3be22327),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc627a70),
	.w1(32'hba65c250),
	.w2(32'hbaba48e5),
	.w3(32'h3b775a92),
	.w4(32'hb9d002cd),
	.w5(32'hbbd50a48),
	.w6(32'h3ba0c62a),
	.w7(32'h3be3aa89),
	.w8(32'h3bcd9da5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c2dc),
	.w1(32'hba8b6f05),
	.w2(32'hbc04c3ac),
	.w3(32'hbb680409),
	.w4(32'h3b8f7a4e),
	.w5(32'h3b31976a),
	.w6(32'hbabbe6b4),
	.w7(32'h3b141aea),
	.w8(32'h3bb653c1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52b99),
	.w1(32'hbab6e0bd),
	.w2(32'h3b05d39d),
	.w3(32'hba168caf),
	.w4(32'hbbf7265a),
	.w5(32'hbbe7c7c7),
	.w6(32'hbaec6c89),
	.w7(32'h3b00c64d),
	.w8(32'hb90d7328),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d96dba),
	.w1(32'hbbe9049f),
	.w2(32'hbc903b97),
	.w3(32'hb9a80d00),
	.w4(32'hbc3f7d02),
	.w5(32'hbcad2573),
	.w6(32'hbc1c0a8e),
	.w7(32'hbb21558f),
	.w8(32'hbbc9eb54),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9695d7),
	.w1(32'hbba1af91),
	.w2(32'hbc8fa6e4),
	.w3(32'hbb5c489e),
	.w4(32'hbca01582),
	.w5(32'hbc3dfe4d),
	.w6(32'hbb03c1ff),
	.w7(32'h3c0f72ab),
	.w8(32'h3c32a649),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f8664),
	.w1(32'h3c94a08a),
	.w2(32'h3c0dc2d2),
	.w3(32'h3bf3c4d8),
	.w4(32'hbc45c70c),
	.w5(32'h3c4b5a92),
	.w6(32'hba4c028f),
	.w7(32'hbb9ee23d),
	.w8(32'hba90ebd7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7de495),
	.w1(32'hbada8c15),
	.w2(32'h3a41cf06),
	.w3(32'h3c7529e7),
	.w4(32'hbaad0cd4),
	.w5(32'hbaf771d1),
	.w6(32'h3884a96d),
	.w7(32'h3a1b959e),
	.w8(32'hbb5d761e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2a26),
	.w1(32'hbaeb7ca0),
	.w2(32'hbb12592b),
	.w3(32'hbb20cf46),
	.w4(32'hbab5cb3d),
	.w5(32'hba0c1b5a),
	.w6(32'hbb2ef6a7),
	.w7(32'hbaf700bc),
	.w8(32'hba88b619),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc15f),
	.w1(32'hbafafad9),
	.w2(32'hbc9340f0),
	.w3(32'hba234ece),
	.w4(32'h3c46c0bc),
	.w5(32'hbbd0a49f),
	.w6(32'h3bd6d7cd),
	.w7(32'h3a502ea8),
	.w8(32'h3b3c4399),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d52b0),
	.w1(32'h3a079ff0),
	.w2(32'h3ba3b4ea),
	.w3(32'hbbb079b5),
	.w4(32'h39c69c8c),
	.w5(32'h3b488d72),
	.w6(32'h3bafa0c3),
	.w7(32'h3b8a5f6e),
	.w8(32'h3b1845cd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990111),
	.w1(32'hbcbc0c4d),
	.w2(32'hbab59e58),
	.w3(32'h3acd63f9),
	.w4(32'h3b7edce8),
	.w5(32'hbc41a953),
	.w6(32'hbaf0fb13),
	.w7(32'h3aaf9b15),
	.w8(32'hbb528246),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf47836),
	.w1(32'hbc130b09),
	.w2(32'hbb0011a2),
	.w3(32'hbbf9c243),
	.w4(32'h3c57d476),
	.w5(32'h3bad16f5),
	.w6(32'h3acdd9cd),
	.w7(32'h3c6b43e7),
	.w8(32'h3bb7e10b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a2d36),
	.w1(32'hbb10ccb6),
	.w2(32'h3c0c0e36),
	.w3(32'h3c0ce015),
	.w4(32'h3bc1ec6d),
	.w5(32'h3ad5c979),
	.w6(32'h3c6f32a8),
	.w7(32'h3c727a75),
	.w8(32'hb9fde7d0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90b35d),
	.w1(32'h3bac851c),
	.w2(32'hbc9d321d),
	.w3(32'hba3161d2),
	.w4(32'h3cb64dfd),
	.w5(32'h3ca71608),
	.w6(32'hbc0e01ea),
	.w7(32'h3c4a93b0),
	.w8(32'h3c60bc7e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3345d4),
	.w1(32'h3c46e8f6),
	.w2(32'h3c39cc2f),
	.w3(32'hbb7ef733),
	.w4(32'hbcb6aa70),
	.w5(32'hbb407034),
	.w6(32'hbaa96924),
	.w7(32'hbb98e8d9),
	.w8(32'hbb3641c8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8470d4),
	.w1(32'hbb980748),
	.w2(32'h3bc73e75),
	.w3(32'h3cc04891),
	.w4(32'h3b1cb01e),
	.w5(32'h3c40882d),
	.w6(32'hb9adf268),
	.w7(32'h3bb7dce8),
	.w8(32'hb8eea0bb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84552b),
	.w1(32'h3d1c326f),
	.w2(32'h3ceb5613),
	.w3(32'hbb30d7ab),
	.w4(32'hbc40623a),
	.w5(32'h3d10e85b),
	.w6(32'hbc3038b7),
	.w7(32'hbc50c41b),
	.w8(32'h3b68fe81),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd3006),
	.w1(32'h3bd43e04),
	.w2(32'hba72da38),
	.w3(32'h3d3eebf9),
	.w4(32'hbc381dca),
	.w5(32'hbcb279d8),
	.w6(32'hbae30b4f),
	.w7(32'hbbe9359d),
	.w8(32'hbc1c435f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa72ff),
	.w1(32'hbc137437),
	.w2(32'h3b33813b),
	.w3(32'hbc0ae24f),
	.w4(32'h3a946ee0),
	.w5(32'h3aaae806),
	.w6(32'h3aa03b8f),
	.w7(32'hbc043025),
	.w8(32'hbb02dcc7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38d9ca),
	.w1(32'hbb99da9c),
	.w2(32'hb98b8003),
	.w3(32'hbaf235ea),
	.w4(32'hbc129b20),
	.w5(32'hbc1717b5),
	.w6(32'hbb2ae0de),
	.w7(32'hbb8502bb),
	.w8(32'hbb6a1eba),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23d122),
	.w1(32'h3bc51d30),
	.w2(32'h3ba2377d),
	.w3(32'hbabe7b0a),
	.w4(32'hbc44177a),
	.w5(32'hbc0f2375),
	.w6(32'h3bc623e9),
	.w7(32'h3a95438d),
	.w8(32'h3b68eda5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31ba63),
	.w1(32'h3c163005),
	.w2(32'hbb04c987),
	.w3(32'h3af0cd83),
	.w4(32'h3a7bb44a),
	.w5(32'hbb4fe806),
	.w6(32'hbbd4ab51),
	.w7(32'hbbd7ed61),
	.w8(32'hbb7253a6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4289d),
	.w1(32'h3c0758a2),
	.w2(32'h3a8522d0),
	.w3(32'h3c04a773),
	.w4(32'h3b811b7a),
	.w5(32'h3bce225f),
	.w6(32'h3b7652a5),
	.w7(32'h3b2883c8),
	.w8(32'h3b883d8d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c313d4),
	.w1(32'hbb04c43a),
	.w2(32'hbadec397),
	.w3(32'h3c3a9afe),
	.w4(32'hba971eda),
	.w5(32'h3a62dcd2),
	.w6(32'hbb30550a),
	.w7(32'hba33e1dc),
	.w8(32'h39d736e5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48a08),
	.w1(32'h3c4bd1ce),
	.w2(32'hbba70cfb),
	.w3(32'h38d29f7a),
	.w4(32'hbad84cb1),
	.w5(32'h3d1f3aee),
	.w6(32'hbc8fd56e),
	.w7(32'hbb4de640),
	.w8(32'hba3c87a5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb681da),
	.w1(32'hb99bd461),
	.w2(32'h3a1cb99f),
	.w3(32'h3d2eec99),
	.w4(32'h3ae01ead),
	.w5(32'hb7bb0d54),
	.w6(32'h3aed19cc),
	.w7(32'h3a57c6ad),
	.w8(32'h3aadd013),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c15eb),
	.w1(32'hbac52a74),
	.w2(32'h3c0854a5),
	.w3(32'hbaae0173),
	.w4(32'hb92121c7),
	.w5(32'h3b906cad),
	.w6(32'h3b90aabd),
	.w7(32'h3b014de6),
	.w8(32'h3ab1e633),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d9c2e),
	.w1(32'h3bcbb100),
	.w2(32'h3ca87beb),
	.w3(32'h3a93376a),
	.w4(32'hbbf8b781),
	.w5(32'hbcb3ea17),
	.w6(32'h3acc9304),
	.w7(32'hbbcae39a),
	.w8(32'hbb601b34),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8545e5),
	.w1(32'hbb907230),
	.w2(32'hbb8bd9a2),
	.w3(32'h3897924f),
	.w4(32'hbc14f261),
	.w5(32'hbc6f5bd2),
	.w6(32'hbb0abf30),
	.w7(32'h39486838),
	.w8(32'hbb1afb33),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fd2b3),
	.w1(32'hbb97c7de),
	.w2(32'hbb448375),
	.w3(32'hbbba9524),
	.w4(32'hbb79afd2),
	.w5(32'hbb534271),
	.w6(32'hbb5b5621),
	.w7(32'hbb513383),
	.w8(32'hbb3762b8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad630a3),
	.w1(32'hbb279f2e),
	.w2(32'h3b063969),
	.w3(32'hbaa25f0f),
	.w4(32'hba2cae2c),
	.w5(32'h3b8c3082),
	.w6(32'h3b9e40fc),
	.w7(32'h3ac697e5),
	.w8(32'h3b4563a2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6cb90),
	.w1(32'h3b2c9b2c),
	.w2(32'h3b4222bc),
	.w3(32'hbae63ad6),
	.w4(32'h3b5988b2),
	.w5(32'h3be1fce6),
	.w6(32'h3bf5fe0a),
	.w7(32'hb8b04d5c),
	.w8(32'h3ac9ee0e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7e012),
	.w1(32'h3cd1de34),
	.w2(32'h3cd6d4b4),
	.w3(32'hbaacac69),
	.w4(32'hbc884ab9),
	.w5(32'h3c3e432e),
	.w6(32'h3bc92a0b),
	.w7(32'hbc03f52a),
	.w8(32'hbb94d081),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcda0e1),
	.w1(32'hbbc333c7),
	.w2(32'hbb89d70a),
	.w3(32'h3ce90471),
	.w4(32'hbb2b1f3a),
	.w5(32'hbb20d78f),
	.w6(32'h3bae610a),
	.w7(32'h3af47aa5),
	.w8(32'h3b3123e5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c2d04),
	.w1(32'h3b1e1206),
	.w2(32'h3b989eb0),
	.w3(32'hbb728bde),
	.w4(32'hbbbfb5f2),
	.w5(32'h3a859157),
	.w6(32'h3bd02093),
	.w7(32'hbc01385e),
	.w8(32'h3b9d5744),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d2449),
	.w1(32'h3c250d4d),
	.w2(32'h3bb30ada),
	.w3(32'h3b8f6294),
	.w4(32'hbb907fe6),
	.w5(32'h3c3094ce),
	.w6(32'hbbc1fb29),
	.w7(32'hbbb93eb5),
	.w8(32'hbb38bd3e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7e0d),
	.w1(32'h3b4ba407),
	.w2(32'h3b1100e8),
	.w3(32'h3c1e71d0),
	.w4(32'h3a00d4b6),
	.w5(32'h3abbcd1d),
	.w6(32'h3a4aeae2),
	.w7(32'h3b1d3896),
	.w8(32'h3a18b30e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bf6e3),
	.w1(32'h3ad940c5),
	.w2(32'h3c3edcfe),
	.w3(32'h39cf238c),
	.w4(32'h3be1bbc4),
	.w5(32'h3b9531a8),
	.w6(32'h39ec2dfa),
	.w7(32'h3b96ece7),
	.w8(32'h3b7635ac),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba21eb2),
	.w1(32'hbc25ff35),
	.w2(32'h3d1b2ab3),
	.w3(32'h3b6c0b05),
	.w4(32'hbc8601e2),
	.w5(32'hbd37e269),
	.w6(32'h3cd02163),
	.w7(32'hbc0bcf82),
	.w8(32'hbcec3ad5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4ad55),
	.w1(32'hbac683de),
	.w2(32'h3b4503b2),
	.w3(32'hbc41670f),
	.w4(32'h3ba4eb7a),
	.w5(32'h3ba40d7a),
	.w6(32'h3c660e21),
	.w7(32'h3c897be7),
	.w8(32'h3b938172),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7b4d7),
	.w1(32'hbaa82bf6),
	.w2(32'hbb031e2f),
	.w3(32'h3a46f0a1),
	.w4(32'hbaae592b),
	.w5(32'hbaa5e1e3),
	.w6(32'hba8a256e),
	.w7(32'hb92f3f19),
	.w8(32'hba922fa8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb6295),
	.w1(32'h3ca8b0e9),
	.w2(32'h3c92c62a),
	.w3(32'hba7bbc6d),
	.w4(32'h3c3f399a),
	.w5(32'h3c38750a),
	.w6(32'h3c553109),
	.w7(32'h3c8cc1d5),
	.w8(32'h3c3f9620),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule