module layer_8_featuremap_171(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04660f),
	.w1(32'h3a90f248),
	.w2(32'hbaed2414),
	.w3(32'hbbc854cc),
	.w4(32'h3ba394ce),
	.w5(32'h3b7518ab),
	.w6(32'hbabda718),
	.w7(32'hba7ccfa8),
	.w8(32'hbb279741),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39857650),
	.w1(32'h3ada9c87),
	.w2(32'h3aa7d285),
	.w3(32'h3c0a1751),
	.w4(32'h3af73bf7),
	.w5(32'h3b04b973),
	.w6(32'h3996ef69),
	.w7(32'h3891ca80),
	.w8(32'h3a198545),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b423f84),
	.w1(32'h377517b9),
	.w2(32'hbb2b9f11),
	.w3(32'h3b40c079),
	.w4(32'hbaf7c03a),
	.w5(32'hbba71e15),
	.w6(32'h3baa14df),
	.w7(32'h3b14463f),
	.w8(32'h3b695cab),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1effe6),
	.w1(32'hbb11cdfb),
	.w2(32'hbc0e230a),
	.w3(32'hbb908ca9),
	.w4(32'hbb562b8e),
	.w5(32'hbbcc72b6),
	.w6(32'hbadb0104),
	.w7(32'hbb973fe4),
	.w8(32'hbb85ba09),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407cc6),
	.w1(32'hbb341870),
	.w2(32'hbacc550b),
	.w3(32'hbb2ae9d7),
	.w4(32'hbb1a579a),
	.w5(32'hba101bda),
	.w6(32'hbbb892f6),
	.w7(32'hbb67446c),
	.w8(32'hbb2a5b74),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbf122),
	.w1(32'h3b6e7d69),
	.w2(32'h3ba56d9f),
	.w3(32'hba1721a0),
	.w4(32'h3bf4abf3),
	.w5(32'h3beb4839),
	.w6(32'hbb6eb2c5),
	.w7(32'hbb449c3b),
	.w8(32'hbb0bf15e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0788d),
	.w1(32'hbb106f10),
	.w2(32'hbb0ad16e),
	.w3(32'hb963d3eb),
	.w4(32'hbb17944d),
	.w5(32'hbb10dea4),
	.w6(32'hbb04a45a),
	.w7(32'hbb051481),
	.w8(32'hbaf4d4ec),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d6246),
	.w1(32'h3a459f43),
	.w2(32'hb8a65c04),
	.w3(32'h3a2ba990),
	.w4(32'h3ac533c3),
	.w5(32'h3b134df6),
	.w6(32'hbafc809d),
	.w7(32'hba37db90),
	.w8(32'h3ab5c4b1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e178),
	.w1(32'hbad7f3b4),
	.w2(32'h3b03cf6a),
	.w3(32'h3bb4380c),
	.w4(32'hbb3f6f53),
	.w5(32'h3aa4aac0),
	.w6(32'hbb3154b1),
	.w7(32'h3a83e58a),
	.w8(32'hb91ecf54),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2bf34),
	.w1(32'h3aa409a4),
	.w2(32'hbb8919cf),
	.w3(32'h3b44ed44),
	.w4(32'h3b495c43),
	.w5(32'hbb2e9707),
	.w6(32'h3aab6612),
	.w7(32'h3b86aad4),
	.w8(32'h3b6970e7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf216ec),
	.w1(32'hbba40962),
	.w2(32'hbb69919d),
	.w3(32'hbbbe17c6),
	.w4(32'hbbf5fc49),
	.w5(32'hbaf4e23d),
	.w6(32'hbc647994),
	.w7(32'hbc24d537),
	.w8(32'hbc1ed0cb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeef09),
	.w1(32'h3ba60e9e),
	.w2(32'h3c0e0d17),
	.w3(32'hb709f1ad),
	.w4(32'h3baf3ccf),
	.w5(32'h3bddee22),
	.w6(32'hbad70be8),
	.w7(32'h3bb5bb2c),
	.w8(32'h3b842399),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12c99f),
	.w1(32'h3b0839cf),
	.w2(32'h3aecfa46),
	.w3(32'h3c102baa),
	.w4(32'h3b1f5ad2),
	.w5(32'h3a2b7ece),
	.w6(32'h3ad11d91),
	.w7(32'h3b41d34d),
	.w8(32'h3bbbd630),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6b418),
	.w1(32'hbc14123c),
	.w2(32'hbc39933b),
	.w3(32'hba61104c),
	.w4(32'hbba3ea20),
	.w5(32'hbc4743f9),
	.w6(32'hbb8a84ad),
	.w7(32'hbad263f3),
	.w8(32'h3a8a792c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c09ea),
	.w1(32'hb95d4f55),
	.w2(32'h39e71eca),
	.w3(32'hbbb64e7c),
	.w4(32'hb9ea621d),
	.w5(32'h38c35f17),
	.w6(32'hba62aaa4),
	.w7(32'h39459f1f),
	.w8(32'hba2391e0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980c1a0),
	.w1(32'hbb2b9e79),
	.w2(32'h3b722218),
	.w3(32'hb9c78304),
	.w4(32'h3b93f9f3),
	.w5(32'h3be490a0),
	.w6(32'hbb680e3f),
	.w7(32'hb941a4ca),
	.w8(32'hba5069fc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df0b2f),
	.w1(32'h3a316a52),
	.w2(32'h3b681351),
	.w3(32'hbb16dd01),
	.w4(32'h3ab9db9c),
	.w5(32'h3b8f89ed),
	.w6(32'hbb512af6),
	.w7(32'hbb440d6a),
	.w8(32'hbbc9a711),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2267d),
	.w1(32'hbb26d66f),
	.w2(32'hbc0912c0),
	.w3(32'hbbe1bad8),
	.w4(32'hbb724939),
	.w5(32'hbc134544),
	.w6(32'hbc1612d9),
	.w7(32'hbc0cfb28),
	.w8(32'hbb8cb389),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc86b6),
	.w1(32'h3c97e8c8),
	.w2(32'h3c124710),
	.w3(32'hbc0d3968),
	.w4(32'h3c516ec5),
	.w5(32'h3c45ae9f),
	.w6(32'hbc014e4b),
	.w7(32'hbb982bbe),
	.w8(32'hbc0ba32e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1713d9),
	.w1(32'hbae1888b),
	.w2(32'h3aa8aa35),
	.w3(32'hbbbccc39),
	.w4(32'hbb156782),
	.w5(32'h3a0ec69b),
	.w6(32'hbc4ad7a6),
	.w7(32'hbb62f844),
	.w8(32'hbaaa974d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb179f2b),
	.w1(32'hbbad640c),
	.w2(32'hbac0ffa1),
	.w3(32'hbb3906a9),
	.w4(32'hbb07101f),
	.w5(32'hbad8dee9),
	.w6(32'hbbe51b32),
	.w7(32'hbb59d7dc),
	.w8(32'hb9afe65b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d74b),
	.w1(32'hbb87ab8a),
	.w2(32'hbbcfa6bb),
	.w3(32'h385cb5f2),
	.w4(32'hbaa0f113),
	.w5(32'hbbbf0d9a),
	.w6(32'hbb883206),
	.w7(32'hbc10659c),
	.w8(32'hbb826ef5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16c64e),
	.w1(32'h3c03bf9f),
	.w2(32'h3b964ced),
	.w3(32'hbb2b1464),
	.w4(32'h3b5aaa9b),
	.w5(32'h3b6dd15a),
	.w6(32'hbbb28cdb),
	.w7(32'hbafe5926),
	.w8(32'hbbfc5738),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c557c),
	.w1(32'hbc3436a1),
	.w2(32'hbc501fe8),
	.w3(32'h3b83b49d),
	.w4(32'hbbf47886),
	.w5(32'hbc27462f),
	.w6(32'hbc20b03a),
	.w7(32'hbc3a016a),
	.w8(32'hbbb94487),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fe290),
	.w1(32'hbb43f097),
	.w2(32'hbb2d2c98),
	.w3(32'hbbcd7319),
	.w4(32'hbb15468c),
	.w5(32'hbb2b2251),
	.w6(32'hbb0d9399),
	.w7(32'hbb5611ba),
	.w8(32'hbadded33),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b42a7),
	.w1(32'h3bc5eb57),
	.w2(32'h3b7f81ed),
	.w3(32'hbb94ca08),
	.w4(32'h3bde4f13),
	.w5(32'h3addde49),
	.w6(32'hbbd04bbc),
	.w7(32'hbb31cf0e),
	.w8(32'hbb21c565),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c6280),
	.w1(32'h3be6dbda),
	.w2(32'h3bf84eb8),
	.w3(32'h3b5cd4f7),
	.w4(32'h3b98dd45),
	.w5(32'h3bfbe70e),
	.w6(32'h3c2226de),
	.w7(32'h3bf5b186),
	.w8(32'h3b8bed01),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989d6ea),
	.w1(32'h3cf18265),
	.w2(32'h3d209d68),
	.w3(32'hbcb67f2f),
	.w4(32'h3c45d78c),
	.w5(32'h3bfb85e2),
	.w6(32'hbce791e8),
	.w7(32'h3b2bdce5),
	.w8(32'h3c065bf3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c07ff),
	.w1(32'h3b0bf198),
	.w2(32'h3b156b83),
	.w3(32'h3b48580e),
	.w4(32'hbb3c700c),
	.w5(32'h3aed59f3),
	.w6(32'hbb592869),
	.w7(32'h39a20de9),
	.w8(32'hba71403d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc5193),
	.w1(32'hb9ee8ee5),
	.w2(32'hb9aaab81),
	.w3(32'h3a1b15fc),
	.w4(32'h3984d93b),
	.w5(32'hba0ee9c4),
	.w6(32'h3a09d913),
	.w7(32'h39c6a81a),
	.w8(32'hbb6aacd3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976821),
	.w1(32'hba3744db),
	.w2(32'h3a327f05),
	.w3(32'hbba2de5f),
	.w4(32'hba9c7709),
	.w5(32'h3a538571),
	.w6(32'hba70841c),
	.w7(32'h3afa1348),
	.w8(32'h3b5e250d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae66722),
	.w1(32'hbb8b3026),
	.w2(32'hbad97ad7),
	.w3(32'hba6305dd),
	.w4(32'hbbe906b8),
	.w5(32'hbbc31452),
	.w6(32'hbadf8a12),
	.w7(32'h3b9f211a),
	.w8(32'h3b938501),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ab20),
	.w1(32'h3bb721ed),
	.w2(32'h3ae90a75),
	.w3(32'hbba896da),
	.w4(32'h3ba6404e),
	.w5(32'h3bb3379e),
	.w6(32'h3b5ed5a4),
	.w7(32'hb9e72020),
	.w8(32'h3b2033b9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e71c),
	.w1(32'hbadf9313),
	.w2(32'hbafccab1),
	.w3(32'h3bebf8f5),
	.w4(32'hbac97625),
	.w5(32'hba75fea8),
	.w6(32'hbad2cbf1),
	.w7(32'h38d66b27),
	.w8(32'h3a8db1fd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8317c4),
	.w1(32'hb90b065e),
	.w2(32'hb9f404b1),
	.w3(32'hbb8978ca),
	.w4(32'h3acf6bce),
	.w5(32'h3a9b6649),
	.w6(32'hba8fdefd),
	.w7(32'hba167b4c),
	.w8(32'h3b5957f0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b503877),
	.w1(32'h3b9906d8),
	.w2(32'h3b956072),
	.w3(32'h3afd41ea),
	.w4(32'hbb21b412),
	.w5(32'hbae046b0),
	.w6(32'hbb067724),
	.w7(32'h3b370496),
	.w8(32'h3b317b8e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14485d),
	.w1(32'hb9de4bdd),
	.w2(32'h3a2feb53),
	.w3(32'hbb9a1a1e),
	.w4(32'hb9ca80cd),
	.w5(32'h3b001bc5),
	.w6(32'h3a0432a6),
	.w7(32'h3a8937aa),
	.w8(32'hba96b3d8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1743fe),
	.w1(32'hbb2db5bf),
	.w2(32'hbaf25e84),
	.w3(32'hba8c6aff),
	.w4(32'hbb4e671e),
	.w5(32'hbb27593e),
	.w6(32'hbacc330c),
	.w7(32'hb9b4ee1d),
	.w8(32'hbada69c7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20cc46),
	.w1(32'hbc1470e1),
	.w2(32'hbba9102d),
	.w3(32'hbb2c7e49),
	.w4(32'hbba4d406),
	.w5(32'hbb7e6079),
	.w6(32'hbbe98b45),
	.w7(32'hbb47a61b),
	.w8(32'hbb8a1c60),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72cdf0),
	.w1(32'hba0dcfe4),
	.w2(32'hba122fc8),
	.w3(32'hba6f4351),
	.w4(32'hbb0fd4cc),
	.w5(32'h396eb4ab),
	.w6(32'hbb0783e7),
	.w7(32'hbaedd2c9),
	.w8(32'hba6ce2d4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e2fa),
	.w1(32'h3c9113db),
	.w2(32'h3c34f1f0),
	.w3(32'hbc064a87),
	.w4(32'h3bb99684),
	.w5(32'h3b6788ae),
	.w6(32'hbc080ca6),
	.w7(32'h3afd5103),
	.w8(32'hba9ada36),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7a5ef),
	.w1(32'hbaec5de4),
	.w2(32'h3a325ece),
	.w3(32'h3b28ebb4),
	.w4(32'h3ab30fde),
	.w5(32'h3b682fa8),
	.w6(32'hbbe8143a),
	.w7(32'hbb525486),
	.w8(32'h399d5dbc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6ea02),
	.w1(32'hbb454c33),
	.w2(32'hbab7ab14),
	.w3(32'h3a896d5d),
	.w4(32'hbb35d5be),
	.w5(32'hb8ca16ed),
	.w6(32'hbb7e6749),
	.w7(32'hbb878bb0),
	.w8(32'hbbaf106f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78a223),
	.w1(32'hbb3cab05),
	.w2(32'hbb215774),
	.w3(32'hbb9446e6),
	.w4(32'hbbb2eff9),
	.w5(32'hbbacac04),
	.w6(32'hbc2f5af1),
	.w7(32'hbba37fec),
	.w8(32'hbbf7a590),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d558e),
	.w1(32'h3bf6ca4b),
	.w2(32'h3bd5e942),
	.w3(32'hbb72a276),
	.w4(32'h3b7588db),
	.w5(32'h3ba0e65e),
	.w6(32'hba870091),
	.w7(32'hb9f5412a),
	.w8(32'hbb968fba),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6875f),
	.w1(32'h3bb9f34a),
	.w2(32'h3b6f19f0),
	.w3(32'h3b3481c9),
	.w4(32'h3b514ddb),
	.w5(32'h3b333d22),
	.w6(32'h39e68ff0),
	.w7(32'h3af58798),
	.w8(32'h3b1184f5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb8b12),
	.w1(32'hbbabd8eb),
	.w2(32'hbba021d6),
	.w3(32'hb726db76),
	.w4(32'hbb7002d4),
	.w5(32'hbaa4ae15),
	.w6(32'hbbd04285),
	.w7(32'hbbaa0129),
	.w8(32'hbbe04c67),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55305a),
	.w1(32'hbb662711),
	.w2(32'hbc1a49fd),
	.w3(32'hbb793fa8),
	.w4(32'hbba05b30),
	.w5(32'hbc25090a),
	.w6(32'hbb85590a),
	.w7(32'hbc08d987),
	.w8(32'hbb97e980),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc325584),
	.w1(32'hbc0f84f5),
	.w2(32'hbc1f03b2),
	.w3(32'hbc1919d6),
	.w4(32'hbbddc51c),
	.w5(32'hbc19f39b),
	.w6(32'hbbc9c0e5),
	.w7(32'hbbb16ba6),
	.w8(32'hbb98f885),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2106b6),
	.w1(32'h3a0926de),
	.w2(32'h3a8ad9b5),
	.w3(32'hbc37396d),
	.w4(32'h3a4d64cc),
	.w5(32'h3b2078a0),
	.w6(32'hbbb053d3),
	.w7(32'hbc05d8e5),
	.w8(32'hbbfe9de9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb105444),
	.w1(32'h3a9191e5),
	.w2(32'h3ae5a2d3),
	.w3(32'h3c147349),
	.w4(32'h3bb364b3),
	.w5(32'h3bc99b88),
	.w6(32'h3ba94897),
	.w7(32'h3c2a2da6),
	.w8(32'h3bd38558),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c43523),
	.w1(32'h3c84ef6e),
	.w2(32'h3c3d1c72),
	.w3(32'hbbb53a2c),
	.w4(32'h3bf06860),
	.w5(32'h3c316bc4),
	.w6(32'hbc6464fd),
	.w7(32'hbbb42f9a),
	.w8(32'hbbfb39eb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbace833),
	.w1(32'h39f78f20),
	.w2(32'hba27f13f),
	.w3(32'hbb59a363),
	.w4(32'hbb167f73),
	.w5(32'hbaa79dd1),
	.w6(32'hbb894141),
	.w7(32'hbb2fa9ee),
	.w8(32'hbb2cfbc3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1babf),
	.w1(32'h3b2003f9),
	.w2(32'hbbdaebbb),
	.w3(32'hbb7e90dc),
	.w4(32'h3accc27d),
	.w5(32'hbbbf62be),
	.w6(32'hbb1d424d),
	.w7(32'hbb070ffe),
	.w8(32'hbba676eb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1483b),
	.w1(32'hbae194a7),
	.w2(32'hbbd08286),
	.w3(32'hbb759d2c),
	.w4(32'h3b07cb0c),
	.w5(32'hbad5e7b7),
	.w6(32'hbb91aad0),
	.w7(32'hbbdefed1),
	.w8(32'hbb9fc4fe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbae13),
	.w1(32'hbb6e3241),
	.w2(32'hbbbe4604),
	.w3(32'h3b1b78af),
	.w4(32'h3b15190c),
	.w5(32'hbbd2fa22),
	.w6(32'hbb0c5d96),
	.w7(32'h3ae82fb2),
	.w8(32'hb9933f40),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5da78),
	.w1(32'hbbc0b0d1),
	.w2(32'hbba33027),
	.w3(32'hbb7eeb95),
	.w4(32'h3a888c01),
	.w5(32'h3ba8d631),
	.w6(32'hbc158f92),
	.w7(32'hbbb2e4a7),
	.w8(32'hbb819b25),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90a73a),
	.w1(32'h3baea065),
	.w2(32'h3c19dbd0),
	.w3(32'h3c04b68e),
	.w4(32'h3aa6b355),
	.w5(32'h3becbefd),
	.w6(32'hbbc77e75),
	.w7(32'hbae6a970),
	.w8(32'h3a432cd1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef2fe2),
	.w1(32'hbb35afe9),
	.w2(32'hba022984),
	.w3(32'h3b0477d3),
	.w4(32'hbb8e19a9),
	.w5(32'hbb0302de),
	.w6(32'hbbc36927),
	.w7(32'hbb7d0661),
	.w8(32'hbb89856a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0da54),
	.w1(32'hbb99f436),
	.w2(32'hbc5c3075),
	.w3(32'hbbd0ecc2),
	.w4(32'hbbd2160c),
	.w5(32'hbc0dc4f7),
	.w6(32'hbc0531a5),
	.w7(32'hbc356531),
	.w8(32'hbbc8a4f0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29aad),
	.w1(32'hbaf03ee7),
	.w2(32'h3b2d47ad),
	.w3(32'hbb9975dc),
	.w4(32'hbaf02794),
	.w5(32'h3b7fec5e),
	.w6(32'hbb8d5f80),
	.w7(32'h3988fb4e),
	.w8(32'hba5cfab0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ba6ad),
	.w1(32'hba1bf9e9),
	.w2(32'hbaea8efa),
	.w3(32'h3ac94326),
	.w4(32'hb8314f52),
	.w5(32'hbae4c969),
	.w6(32'h3b89e4f0),
	.w7(32'h3b309775),
	.w8(32'h3aa88639),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba698856),
	.w1(32'hbb2c7d56),
	.w2(32'hbb147502),
	.w3(32'hbbfe0904),
	.w4(32'hbc1b73c9),
	.w5(32'hbc204cd8),
	.w6(32'hbc6b86aa),
	.w7(32'hbb00e868),
	.w8(32'hbb8c8ec7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed66ea),
	.w1(32'h3b11c75c),
	.w2(32'h3b7f6ef6),
	.w3(32'hbc5ac7c2),
	.w4(32'h3aec9ca4),
	.w5(32'h3bb01e84),
	.w6(32'h3b45b36f),
	.w7(32'h3ba6cc57),
	.w8(32'h3bca799f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd57fb),
	.w1(32'h3b5129b8),
	.w2(32'h3b4bf2eb),
	.w3(32'h3bd578fb),
	.w4(32'h3b3a86bb),
	.w5(32'h3b82be8e),
	.w6(32'h3b8c90be),
	.w7(32'h3b9be2c1),
	.w8(32'h3ba9da60),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1f386),
	.w1(32'hb94dc283),
	.w2(32'h3a07a190),
	.w3(32'h3b6c2b73),
	.w4(32'hbac8d276),
	.w5(32'hbac21fcf),
	.w6(32'hbb1744f1),
	.w7(32'hba717fa8),
	.w8(32'hba99c7d7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b3b38),
	.w1(32'h3b6886d4),
	.w2(32'h3b5bbaf3),
	.w3(32'hbac1763b),
	.w4(32'h3a89b0c4),
	.w5(32'h3ad7bab3),
	.w6(32'hbb1f604e),
	.w7(32'hbaee9659),
	.w8(32'hba678d13),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383afd66),
	.w1(32'h3be4f764),
	.w2(32'h3c065d43),
	.w3(32'hbbca2b80),
	.w4(32'h3c0f98c6),
	.w5(32'h3bde0252),
	.w6(32'h3a9768bf),
	.w7(32'h3be48a90),
	.w8(32'h3b033753),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30fae3),
	.w1(32'hbc00ced6),
	.w2(32'hbc2488e2),
	.w3(32'h3bcec59f),
	.w4(32'hbbf1d26d),
	.w5(32'hbc50046f),
	.w6(32'hbbc14b8b),
	.w7(32'hbbffd1a6),
	.w8(32'hbb9ad92f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8605ef),
	.w1(32'h3b79a836),
	.w2(32'hba65ec06),
	.w3(32'hbc98fb93),
	.w4(32'hbc16fab9),
	.w5(32'hbc348eac),
	.w6(32'hbc5c6922),
	.w7(32'hbc3555c9),
	.w8(32'hbbc0c30c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edd170),
	.w1(32'h3aafe308),
	.w2(32'hb8ff050c),
	.w3(32'hb9cb618d),
	.w4(32'hbaf8bacb),
	.w5(32'hbb3bb2ab),
	.w6(32'h3acafbdd),
	.w7(32'h3ac25d0d),
	.w8(32'h3b55abad),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e2314),
	.w1(32'hbb8f2a26),
	.w2(32'hbbf43e46),
	.w3(32'hba457696),
	.w4(32'hbc018e91),
	.w5(32'hbbfd87e7),
	.w6(32'hbb5fc705),
	.w7(32'hbb539520),
	.w8(32'hb9a2e212),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6fade),
	.w1(32'hbbe33d48),
	.w2(32'hbbf6f9c0),
	.w3(32'hbc0300ae),
	.w4(32'hbb144dd0),
	.w5(32'hbbc34ab2),
	.w6(32'h3ad9d935),
	.w7(32'h3a58914e),
	.w8(32'h3acaba6b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7648),
	.w1(32'hba556f5c),
	.w2(32'hb9ba556e),
	.w3(32'hbc267888),
	.w4(32'h3abd24dc),
	.w5(32'hb95e5b71),
	.w6(32'hbb0d6a72),
	.w7(32'h3b19b207),
	.w8(32'hba61d19d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c272),
	.w1(32'hbac50cac),
	.w2(32'hbae8a229),
	.w3(32'h3a658a23),
	.w4(32'h3a80d397),
	.w5(32'h3ab8e47f),
	.w6(32'h364a06bd),
	.w7(32'h3aba0795),
	.w8(32'h3b952fab),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a177c0d),
	.w1(32'h39f50507),
	.w2(32'hbb9ae8f4),
	.w3(32'h39d7cec3),
	.w4(32'h3bb45cb1),
	.w5(32'h39512910),
	.w6(32'hba5f9e45),
	.w7(32'hbb843bd3),
	.w8(32'hbb8beb8b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9cfd),
	.w1(32'hbb73d419),
	.w2(32'hbb5d701c),
	.w3(32'hb8ce88ea),
	.w4(32'hbabd0e4b),
	.w5(32'hb926f70e),
	.w6(32'hbb933ae9),
	.w7(32'hbb9db638),
	.w8(32'hbb83b084),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813683),
	.w1(32'h3be1e147),
	.w2(32'h3c5531d7),
	.w3(32'hbbdd9a4d),
	.w4(32'h3bd5784d),
	.w5(32'h3c512de3),
	.w6(32'hbbb02cd4),
	.w7(32'h3b98971e),
	.w8(32'h3b094151),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c142d5c),
	.w1(32'h3be86120),
	.w2(32'h3bb57af3),
	.w3(32'h3c15dcaa),
	.w4(32'h3bd2c821),
	.w5(32'h3b8b1c88),
	.w6(32'h3bbd43d1),
	.w7(32'h3b970bcc),
	.w8(32'h3b853ba6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804d70),
	.w1(32'hbb94e4f3),
	.w2(32'hba8ba9b5),
	.w3(32'h3b779eb0),
	.w4(32'hbbc00cc7),
	.w5(32'hbb6c2059),
	.w6(32'hbb71cc27),
	.w7(32'h394f0215),
	.w8(32'hbaa33e65),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a695db2),
	.w1(32'h3a91d562),
	.w2(32'hbaf8910d),
	.w3(32'h3aef9320),
	.w4(32'hb9ca5042),
	.w5(32'hbb874a19),
	.w6(32'h3b81ac03),
	.w7(32'h3b2d42c1),
	.w8(32'h3b8a6bd9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03bde2),
	.w1(32'hbc0d9eea),
	.w2(32'hbc848f4d),
	.w3(32'hbbaa4297),
	.w4(32'hbc4eb70d),
	.w5(32'hbc866103),
	.w6(32'hbc424965),
	.w7(32'hbc8d37f4),
	.w8(32'hbc09115e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cc69e),
	.w1(32'h3b933be8),
	.w2(32'h3b8af2e0),
	.w3(32'hbc6aedd9),
	.w4(32'h3b926c47),
	.w5(32'h3bae0fb5),
	.w6(32'hbc0ee39a),
	.w7(32'hbb0ce63f),
	.w8(32'hbb84eb80),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaefbcb),
	.w1(32'h3c80299b),
	.w2(32'hbb5e46e0),
	.w3(32'hbc11f8d0),
	.w4(32'h3b593075),
	.w5(32'h3b5820d8),
	.w6(32'hbc4e84e7),
	.w7(32'hbbb3a64e),
	.w8(32'hba579825),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d4bea),
	.w1(32'h3c405461),
	.w2(32'h3c1211d9),
	.w3(32'hbb5a501c),
	.w4(32'h3aa6652e),
	.w5(32'hb99c3778),
	.w6(32'hbbddae41),
	.w7(32'h3b8575d6),
	.w8(32'h3af6e8c6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d11834),
	.w1(32'h3b155833),
	.w2(32'hb9d27c68),
	.w3(32'hbc1b0b9f),
	.w4(32'hbc0c2eaf),
	.w5(32'hbc0474fe),
	.w6(32'hbc0bcae5),
	.w7(32'hbc07dbc9),
	.w8(32'hbbd311f0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab03837),
	.w1(32'hb91535e8),
	.w2(32'h3abf764f),
	.w3(32'hbbdf8770),
	.w4(32'h3abf6a73),
	.w5(32'h3b1ef94a),
	.w6(32'h393c25ba),
	.w7(32'h3aa0df50),
	.w8(32'h3b8ba3e7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba14f7a),
	.w1(32'h374784cf),
	.w2(32'h3bc1d0dc),
	.w3(32'h3bbf1d86),
	.w4(32'hba3fcc56),
	.w5(32'h3b88d7c4),
	.w6(32'hbb917ce3),
	.w7(32'hba12a525),
	.w8(32'hba5c31d1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be87450),
	.w1(32'hbaac17ee),
	.w2(32'hb8c3a8eb),
	.w3(32'h3b6ff3bb),
	.w4(32'hbb3f037d),
	.w5(32'hba9000ca),
	.w6(32'h3af4aae7),
	.w7(32'h3b7e782c),
	.w8(32'h3b5fe1c6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080630),
	.w1(32'hbc21f932),
	.w2(32'hbc47460e),
	.w3(32'hbb768f9b),
	.w4(32'hbb75e877),
	.w5(32'hbb8d6853),
	.w6(32'hbabe75e2),
	.w7(32'hbb0ecb16),
	.w8(32'h3a95453a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16d7cf),
	.w1(32'hbadbd45a),
	.w2(32'hbab42974),
	.w3(32'hbacf700a),
	.w4(32'hbb893c0c),
	.w5(32'hbb9889f0),
	.w6(32'hbb7e033b),
	.w7(32'hb9f9d792),
	.w8(32'hba8f9368),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb861ff6d),
	.w1(32'hbab4aaaf),
	.w2(32'hbb7c5cbf),
	.w3(32'hbb763b6d),
	.w4(32'hbb431a7d),
	.w5(32'hbb9cc8cc),
	.w6(32'hbb2ad784),
	.w7(32'hba6b5dec),
	.w8(32'hbb936548),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8087e),
	.w1(32'h3b951d57),
	.w2(32'h3b97b131),
	.w3(32'hbc160243),
	.w4(32'h3a295ae4),
	.w5(32'h3b369274),
	.w6(32'hbb71167f),
	.w7(32'hbad677dc),
	.w8(32'h3b1b9c69),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816f52),
	.w1(32'h3b8e895e),
	.w2(32'h3b701443),
	.w3(32'h3aa32583),
	.w4(32'h3b3c2d0c),
	.w5(32'h3b4fcc95),
	.w6(32'hbb1bb019),
	.w7(32'h386c97f7),
	.w8(32'h39aba114),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd25f1),
	.w1(32'hbb878c6b),
	.w2(32'hbac59b75),
	.w3(32'h3b86efbb),
	.w4(32'h3c007dfc),
	.w5(32'h3c17132b),
	.w6(32'hba4ac3de),
	.w7(32'hbab0437e),
	.w8(32'hbb0a5d13),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ab2fb),
	.w1(32'h3bcb4dc8),
	.w2(32'h3bc59483),
	.w3(32'h3ae78d98),
	.w4(32'h3b3a90fa),
	.w5(32'h3bf593df),
	.w6(32'hbae0a31a),
	.w7(32'h3bd08ee5),
	.w8(32'h3b9e654f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b31970),
	.w1(32'h392c877d),
	.w2(32'hbb5d1e05),
	.w3(32'hbb60005d),
	.w4(32'h3ba37d3b),
	.w5(32'h3a343418),
	.w6(32'hbbe2a44a),
	.w7(32'hbbaa3a3b),
	.w8(32'hbb8bd912),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d564e),
	.w1(32'hba904563),
	.w2(32'hbbd75bef),
	.w3(32'hb9c78d15),
	.w4(32'h3ae8e3e0),
	.w5(32'hbba91f49),
	.w6(32'hbb28d7d7),
	.w7(32'hbbd90f06),
	.w8(32'h3b366bc4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d388ca),
	.w1(32'hbbe08513),
	.w2(32'hbc08c03b),
	.w3(32'h3b9c1c18),
	.w4(32'hbba9939c),
	.w5(32'hbbfa6b93),
	.w6(32'hbbdc0f6a),
	.w7(32'hbc022c7e),
	.w8(32'hbbdbff8d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a8a3),
	.w1(32'h39c17510),
	.w2(32'h3a019f11),
	.w3(32'hbb73b848),
	.w4(32'hbbcb1a85),
	.w5(32'hb961581d),
	.w6(32'hbafa1ed0),
	.w7(32'h3b337309),
	.w8(32'h3bbee1d0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16c779),
	.w1(32'hb9792f12),
	.w2(32'h3b3abee6),
	.w3(32'h3b1e6334),
	.w4(32'hbb268b56),
	.w5(32'hbb14a837),
	.w6(32'hb957eefb),
	.w7(32'h3aec5941),
	.w8(32'hbb63b9f1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57f5dc),
	.w1(32'hbb10ea22),
	.w2(32'h3bb52256),
	.w3(32'hbb5fd9fa),
	.w4(32'hb9ea4061),
	.w5(32'h3bc8a0fe),
	.w6(32'hbbd01d67),
	.w7(32'hbb6bfdfd),
	.w8(32'hbaaac1c4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef053a),
	.w1(32'hbc0559d8),
	.w2(32'hbc222de9),
	.w3(32'h3bafd51e),
	.w4(32'hbbc8967d),
	.w5(32'hbc00536b),
	.w6(32'hbba3d83f),
	.w7(32'hbbd5bbb8),
	.w8(32'hbc0bde46),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc355d7a),
	.w1(32'hbb8696d3),
	.w2(32'hbb71d3a3),
	.w3(32'hbc78b17f),
	.w4(32'hbb93d844),
	.w5(32'h3aa394f8),
	.w6(32'hbc234f87),
	.w7(32'hbc36057d),
	.w8(32'hbc1f4046),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2341cc),
	.w1(32'hbc11b84d),
	.w2(32'hbb0d6892),
	.w3(32'h39981f66),
	.w4(32'hbbd5376b),
	.w5(32'h3b97244a),
	.w6(32'hbc14b6cf),
	.w7(32'hbbbd1ca2),
	.w8(32'hbb03a934),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8d428),
	.w1(32'h398106a0),
	.w2(32'h3aec6943),
	.w3(32'hbb90100c),
	.w4(32'hbbc7f2a0),
	.w5(32'hbbba72b6),
	.w6(32'hbc03ae2c),
	.w7(32'hbbafb45a),
	.w8(32'hbbc6b0f1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e08e),
	.w1(32'h3b127cb3),
	.w2(32'h3b91b2a4),
	.w3(32'hbb97d3af),
	.w4(32'h3b035c2d),
	.w5(32'h3ba05af0),
	.w6(32'hb9c16ebb),
	.w7(32'h3b535bf0),
	.w8(32'h3b2098ce),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5eb30),
	.w1(32'h3ac7e337),
	.w2(32'h3b75598a),
	.w3(32'hba006fd7),
	.w4(32'h3b67b5d7),
	.w5(32'h3bcfd8f3),
	.w6(32'hbb119c26),
	.w7(32'hbabc5ac4),
	.w8(32'hbb9c3ec9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ef6bf),
	.w1(32'h39b20f36),
	.w2(32'h3aab8b54),
	.w3(32'hb84d8268),
	.w4(32'hba89100a),
	.w5(32'hb9c0a00b),
	.w6(32'h3b3e6013),
	.w7(32'h3b972142),
	.w8(32'h3b8649c3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0a1e),
	.w1(32'h3a52a3de),
	.w2(32'h3a3fc3b5),
	.w3(32'h3b360b29),
	.w4(32'hb9b00662),
	.w5(32'h398c40e4),
	.w6(32'h3abce236),
	.w7(32'h3afce294),
	.w8(32'h3aaf4aee),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbfe2a),
	.w1(32'hbb0e107f),
	.w2(32'hbac2c588),
	.w3(32'hbb2d6e04),
	.w4(32'hb7ac5982),
	.w5(32'hba160bec),
	.w6(32'hbb5c7aea),
	.w7(32'hba8d3ac4),
	.w8(32'h3ab92c31),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe18614),
	.w1(32'h3b6d500e),
	.w2(32'h3bad4f32),
	.w3(32'hbc1566ee),
	.w4(32'h3b23687a),
	.w5(32'h3b93d15f),
	.w6(32'hbb61b26a),
	.w7(32'h3a6334c1),
	.w8(32'h3b6726f0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148188),
	.w1(32'hbc6f7cf2),
	.w2(32'hbc7c878f),
	.w3(32'h3b53f993),
	.w4(32'hbc571633),
	.w5(32'hbc5cb2c7),
	.w6(32'hbc2d9151),
	.w7(32'hbc21b542),
	.w8(32'hbc6794a9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d71da),
	.w1(32'hba6143d0),
	.w2(32'hbbbca45f),
	.w3(32'hbbfe8d72),
	.w4(32'hbb4e399a),
	.w5(32'hbb81c5ee),
	.w6(32'hbb6f91e0),
	.w7(32'hbbeff84a),
	.w8(32'hbb440bbd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2085f2),
	.w1(32'hbb44d18c),
	.w2(32'hbb20267c),
	.w3(32'h39145fb0),
	.w4(32'hbb5648c1),
	.w5(32'hbb281eab),
	.w6(32'hba112c20),
	.w7(32'hba17be82),
	.w8(32'hbb088773),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67a71),
	.w1(32'hba8ceac8),
	.w2(32'hbacb9173),
	.w3(32'hbb907d5b),
	.w4(32'hbac5aaca),
	.w5(32'hba7a8457),
	.w6(32'hba6bffa7),
	.w7(32'hba2ce6bb),
	.w8(32'hba967226),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e6958),
	.w1(32'h3b4b6854),
	.w2(32'h3b248594),
	.w3(32'hbb85a182),
	.w4(32'h3b1c39e4),
	.w5(32'h3a13b6dd),
	.w6(32'h3989a115),
	.w7(32'h3ad325c0),
	.w8(32'h3a53cc7d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e09ac7),
	.w1(32'hbb1dbe18),
	.w2(32'hbb5ac632),
	.w3(32'hbb51bbce),
	.w4(32'hbb0a26d9),
	.w5(32'hbb8cf05f),
	.w6(32'hbc043636),
	.w7(32'hbbabae55),
	.w8(32'hbb83fcd0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba68f66),
	.w1(32'h3af7e3b3),
	.w2(32'hbaf92604),
	.w3(32'hbba3e9c1),
	.w4(32'h3b3149e8),
	.w5(32'h3bb7f238),
	.w6(32'h3a4051d8),
	.w7(32'hbb9e0caf),
	.w8(32'hb9c9418d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a280f75),
	.w1(32'h395ea363),
	.w2(32'hba8a9445),
	.w3(32'h3b1d063f),
	.w4(32'h3b257880),
	.w5(32'hb9b55f84),
	.w6(32'hba687163),
	.w7(32'hbaa4e790),
	.w8(32'hba3e590f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb6566),
	.w1(32'hbbc7cca3),
	.w2(32'hbc46b479),
	.w3(32'hbb054c17),
	.w4(32'hbc2872ef),
	.w5(32'hbc2dda43),
	.w6(32'hbc121ec5),
	.w7(32'hbbc62d0e),
	.w8(32'hbbb9b0ad),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ef017),
	.w1(32'hba53cc40),
	.w2(32'h39e3b7db),
	.w3(32'hbc06a59b),
	.w4(32'h3b58eebe),
	.w5(32'h3b6bc239),
	.w6(32'hbacf75d7),
	.w7(32'hbb22949b),
	.w8(32'hbae9429f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10ec7a),
	.w1(32'h3ad5be94),
	.w2(32'h3ad7c0de),
	.w3(32'h3b966b3b),
	.w4(32'h3b2e5a25),
	.w5(32'h3b44de85),
	.w6(32'h3b03d47f),
	.w7(32'h3ad82fc9),
	.w8(32'h3b5c890a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8146d5),
	.w1(32'hbc62746a),
	.w2(32'hbc218079),
	.w3(32'h3bab3ba2),
	.w4(32'hbc2c95a8),
	.w5(32'hbc0ef794),
	.w6(32'hbc55714c),
	.w7(32'hbc41a322),
	.w8(32'hbbf7c0ee),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f4f72),
	.w1(32'h3aebfde0),
	.w2(32'hbb69c1a8),
	.w3(32'hbc0f1b78),
	.w4(32'h39a7b813),
	.w5(32'hbbaa215b),
	.w6(32'h39d3c09a),
	.w7(32'hbb0ee87a),
	.w8(32'hbb4c561a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff7a6),
	.w1(32'hbc0c79d0),
	.w2(32'hbc3296f7),
	.w3(32'hbb8b8a5d),
	.w4(32'hbbff8f44),
	.w5(32'hbc34ba97),
	.w6(32'hbc21d2b2),
	.w7(32'hbbf5d794),
	.w8(32'hbbb30c4f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13484c),
	.w1(32'h39953d0d),
	.w2(32'hbb7a1d2e),
	.w3(32'hbc0527aa),
	.w4(32'h3a4cfd3f),
	.w5(32'hbb57b6d3),
	.w6(32'h3821f139),
	.w7(32'hbb12a307),
	.w8(32'h3b1986a1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932b38),
	.w1(32'h3c240159),
	.w2(32'h3c6035fc),
	.w3(32'h3ae6b431),
	.w4(32'h3c7b31a8),
	.w5(32'h3c38d0b7),
	.w6(32'h3b15c8a2),
	.w7(32'h3c60ec88),
	.w8(32'h3a6d5e87),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule