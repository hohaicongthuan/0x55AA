module layer_8_featuremap_187(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03b22),
	.w1(32'h3c8eb9b9),
	.w2(32'h3ce85178),
	.w3(32'hbbd8a514),
	.w4(32'h3c8a0c5d),
	.w5(32'h3d12b3cc),
	.w6(32'hbbc98cf2),
	.w7(32'h3af9d218),
	.w8(32'h3ca21d45),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e750c),
	.w1(32'hbbb5e76d),
	.w2(32'hbc48a16b),
	.w3(32'h39558968),
	.w4(32'hbbb891be),
	.w5(32'hbc2026ec),
	.w6(32'hbc2ca313),
	.w7(32'hbc0ac0cd),
	.w8(32'hbc325db3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6c9b5),
	.w1(32'hbc9dc1c8),
	.w2(32'hbcd49ab5),
	.w3(32'hbc27c75c),
	.w4(32'hbc8780b7),
	.w5(32'hbc75931e),
	.w6(32'hbc594650),
	.w7(32'hbcb400c1),
	.w8(32'hbc883652),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56fea1),
	.w1(32'h3bb6174e),
	.w2(32'hbb098e76),
	.w3(32'h3bb04d06),
	.w4(32'hb9066b4e),
	.w5(32'h3c3e37a2),
	.w6(32'h3b6cb720),
	.w7(32'h3a442f59),
	.w8(32'hbb464169),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d8d8),
	.w1(32'hbb32e8e9),
	.w2(32'hbc01a255),
	.w3(32'h3b319169),
	.w4(32'hbb344d92),
	.w5(32'hbb92b458),
	.w6(32'hbb32ce8e),
	.w7(32'hbb886101),
	.w8(32'hb824c432),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a43b),
	.w1(32'hbc16815f),
	.w2(32'hbc07a2e8),
	.w3(32'hb9b2dc59),
	.w4(32'hbc22abf8),
	.w5(32'hbc2c49be),
	.w6(32'hbb07a5d4),
	.w7(32'hbc587a0e),
	.w8(32'hbb4b4d2e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5b006),
	.w1(32'hbc1571fb),
	.w2(32'hbc3d9560),
	.w3(32'hbb1c1b82),
	.w4(32'hbbf28359),
	.w5(32'hbc0734af),
	.w6(32'hbbc624cb),
	.w7(32'hbbf293af),
	.w8(32'hbc0660c1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7f97e),
	.w1(32'h3c007406),
	.w2(32'hbb9646ba),
	.w3(32'hbc6333fd),
	.w4(32'h3d0659d6),
	.w5(32'h3bdfb79f),
	.w6(32'hbc322da4),
	.w7(32'hbc58a56d),
	.w8(32'hbcb0cc83),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2595eb),
	.w1(32'hba6c9ba4),
	.w2(32'hbc43adae),
	.w3(32'hbc40db49),
	.w4(32'hbc30c292),
	.w5(32'hbc819af2),
	.w6(32'hbc047079),
	.w7(32'hbb099054),
	.w8(32'hbbc09b37),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f37fb),
	.w1(32'hbc5918ab),
	.w2(32'hbc9c13eb),
	.w3(32'hbc94fbfa),
	.w4(32'hbc057a52),
	.w5(32'hbcd0ae0c),
	.w6(32'hbbbed3a7),
	.w7(32'hbb8d4a0c),
	.w8(32'h3ac7d5c8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc656829),
	.w1(32'h3c22af33),
	.w2(32'h3cc1ddb0),
	.w3(32'hbc83ef97),
	.w4(32'h3cbf181c),
	.w5(32'h3d157400),
	.w6(32'h3b88de90),
	.w7(32'h3c1f8f98),
	.w8(32'h3cacae1d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf787ee),
	.w1(32'hbbada747),
	.w2(32'hbb963fa4),
	.w3(32'h3c69bdc9),
	.w4(32'hbbf8228b),
	.w5(32'hbb599154),
	.w6(32'hbbca0837),
	.w7(32'hbbed76e9),
	.w8(32'hbb36c57c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cc67f),
	.w1(32'hbbd03462),
	.w2(32'hbd036bd4),
	.w3(32'hbc2e842d),
	.w4(32'hbc81f93a),
	.w5(32'hbcb9cfe4),
	.w6(32'hb9d8cc81),
	.w7(32'hbc349ce8),
	.w8(32'hbc109679),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb3a37),
	.w1(32'hb9939e58),
	.w2(32'h3c275e46),
	.w3(32'hbb9dfe79),
	.w4(32'h3be0e077),
	.w5(32'h3c2357e7),
	.w6(32'h3bab39e3),
	.w7(32'h3b6e23cb),
	.w8(32'h3be6098a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9808cc),
	.w1(32'hb98fe929),
	.w2(32'h3ade71c8),
	.w3(32'h3c80d34d),
	.w4(32'h3a845619),
	.w5(32'h3b700516),
	.w6(32'hbb668a86),
	.w7(32'hbad8509b),
	.w8(32'hbb922728),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a245f13),
	.w1(32'h3b26c4f9),
	.w2(32'h3c421af5),
	.w3(32'h381776a9),
	.w4(32'hbb19ee95),
	.w5(32'h3cad7c35),
	.w6(32'hba802d4d),
	.w7(32'h3ba4b261),
	.w8(32'h3bdf4f45),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0c077),
	.w1(32'hbc05b62f),
	.w2(32'h3bba4807),
	.w3(32'h3cc92c48),
	.w4(32'hbbc5e3a0),
	.w5(32'h3beb41d3),
	.w6(32'hbbe99681),
	.w7(32'hbba818a4),
	.w8(32'hbc5adf57),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f04f8),
	.w1(32'hbb8e292a),
	.w2(32'hbc69abe5),
	.w3(32'hb98a0386),
	.w4(32'h3baef4d3),
	.w5(32'h3af519a3),
	.w6(32'h3ac51077),
	.w7(32'hbbf2ccee),
	.w8(32'hbaaa22a9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39a9a3),
	.w1(32'h3d4198c2),
	.w2(32'h3d03d2dd),
	.w3(32'h3be6e615),
	.w4(32'h3d910bec),
	.w5(32'h3d6dc266),
	.w6(32'hbc44bcc0),
	.w7(32'h3c020b05),
	.w8(32'h3b1ff735),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fabfe),
	.w1(32'h3cd2811f),
	.w2(32'h3cfb3b01),
	.w3(32'h3c4bd7c7),
	.w4(32'h3cb62c36),
	.w5(32'h3d23d446),
	.w6(32'hba1ba32b),
	.w7(32'h3c0ccb1c),
	.w8(32'h3c968713),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93ecf3),
	.w1(32'hbaab83d5),
	.w2(32'h3a68d1d1),
	.w3(32'hbc1b8a06),
	.w4(32'hbc5dbf7f),
	.w5(32'hbb473731),
	.w6(32'h3a075cb5),
	.w7(32'hbb5fc1f2),
	.w8(32'hb9b31459),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38c084),
	.w1(32'hbce4dbb3),
	.w2(32'hbd41a7b2),
	.w3(32'hbc763047),
	.w4(32'hbca6345c),
	.w5(32'hbcf1e3f7),
	.w6(32'hbc952b85),
	.w7(32'hbcf295dc),
	.w8(32'hbcf94132),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6d98c2),
	.w1(32'h3c4de2cf),
	.w2(32'h3cf45bcb),
	.w3(32'hbd0fa9dd),
	.w4(32'h3d01a3b2),
	.w5(32'h3d3cbf0a),
	.w6(32'hbc407b23),
	.w7(32'h3cd8824d),
	.w8(32'h3cc33f9a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4ee6e),
	.w1(32'hbca6ff3c),
	.w2(32'hbcf313ab),
	.w3(32'h3ca8da8d),
	.w4(32'hbc836516),
	.w5(32'h38b52d26),
	.w6(32'hbc3c6430),
	.w7(32'hbc0fac05),
	.w8(32'hbb8279c5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca74d91),
	.w1(32'h3ac5233c),
	.w2(32'hbbcde51c),
	.w3(32'hbc35f1ab),
	.w4(32'hbc1ca4ec),
	.w5(32'hbc6aca21),
	.w6(32'h3bdd0e8c),
	.w7(32'h3a70b467),
	.w8(32'hbace389a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb8f50),
	.w1(32'h3be9517d),
	.w2(32'h3cd7f33d),
	.w3(32'hbc9f9a1c),
	.w4(32'h3c86eb51),
	.w5(32'h3d304e95),
	.w6(32'hbc96f497),
	.w7(32'hb8ed0b5b),
	.w8(32'h3cfe93ed),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab92309),
	.w1(32'h3b4acc8e),
	.w2(32'h3aefccc4),
	.w3(32'hbbae71f1),
	.w4(32'hbbb8aaa7),
	.w5(32'h3b7b7a5e),
	.w6(32'h3bb3043b),
	.w7(32'hbbfa458e),
	.w8(32'hbae75e72),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f5978),
	.w1(32'hbbbbc3b1),
	.w2(32'h3d8cd837),
	.w3(32'h3cc58650),
	.w4(32'h3c2bdd90),
	.w5(32'h3e18bb40),
	.w6(32'h3e42b788),
	.w7(32'h3e0cf1c5),
	.w8(32'h3d7cca8f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4290),
	.w1(32'hbb7a6055),
	.w2(32'h392ee1ff),
	.w3(32'h3c606d54),
	.w4(32'h3ba6ae12),
	.w5(32'h3c43047a),
	.w6(32'hbc77caee),
	.w7(32'hbbf3d55e),
	.w8(32'hbadcace8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56385b),
	.w1(32'hbbdd6638),
	.w2(32'hbc346c49),
	.w3(32'h3b5575fb),
	.w4(32'hbccefe0b),
	.w5(32'hbcdc9c6f),
	.w6(32'hbbe8bcc0),
	.w7(32'hbbfbc141),
	.w8(32'hbbc062a0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcadaf9),
	.w1(32'h3991354d),
	.w2(32'hbad77c13),
	.w3(32'hbccc55cd),
	.w4(32'h3b8b694b),
	.w5(32'h3a4d8dfa),
	.w6(32'hbb637686),
	.w7(32'hbaeff931),
	.w8(32'hbbea4257),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc238ec4),
	.w1(32'h3bae38c7),
	.w2(32'hbbaacf76),
	.w3(32'hbc31c78b),
	.w4(32'h3b22d097),
	.w5(32'hbc162ab4),
	.w6(32'hbc17b68c),
	.w7(32'hbbca7208),
	.w8(32'hba26a19b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc49ee1),
	.w1(32'h3c0bd87c),
	.w2(32'h3c9436b9),
	.w3(32'hbbe38cb3),
	.w4(32'h3bd87061),
	.w5(32'h3cc449aa),
	.w6(32'h3bc51a82),
	.w7(32'h3c0a9515),
	.w8(32'h3b4a503b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5e1c1),
	.w1(32'hbbe7f5dc),
	.w2(32'hbbab5ec2),
	.w3(32'h3c5868dc),
	.w4(32'h3a247da7),
	.w5(32'h3bc24e24),
	.w6(32'h3bb03750),
	.w7(32'h3ae25cec),
	.w8(32'h384a0eca),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c0eed),
	.w1(32'h3bca51a7),
	.w2(32'h3c11f8aa),
	.w3(32'h3ba5c26f),
	.w4(32'hbc06e46f),
	.w5(32'hbba1aa4a),
	.w6(32'h3a1c1c7a),
	.w7(32'hbc49bbb6),
	.w8(32'hbb78bb07),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7978a7),
	.w1(32'h3c309ab7),
	.w2(32'h3cd7bb00),
	.w3(32'h3c8a0a95),
	.w4(32'h3c532a4e),
	.w5(32'h3c436e1e),
	.w6(32'h3bc31582),
	.w7(32'h3b7957a9),
	.w8(32'h3b997d28),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993c29),
	.w1(32'hb97220b1),
	.w2(32'h3aebc301),
	.w3(32'hbc53cab6),
	.w4(32'hb9b08368),
	.w5(32'hba605411),
	.w6(32'h3a5dba92),
	.w7(32'h3acd6901),
	.w8(32'h3a85a34f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bac01),
	.w1(32'hbbae46ca),
	.w2(32'hbbb6abf0),
	.w3(32'hbc2293ac),
	.w4(32'hbb59339a),
	.w5(32'hbb358682),
	.w6(32'hbc07bb4a),
	.w7(32'hbbf1a4cc),
	.w8(32'hbc426154),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be295a5),
	.w1(32'hbd0f38c7),
	.w2(32'hbd59b6f4),
	.w3(32'h3bd972df),
	.w4(32'hbcabb2e5),
	.w5(32'hbcea9b89),
	.w6(32'hbc5d6ee1),
	.w7(32'hbcff9a69),
	.w8(32'hbc97ab25),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf7f152),
	.w1(32'h3b56120d),
	.w2(32'hbb70caff),
	.w3(32'hba91172d),
	.w4(32'h3ac5b01c),
	.w5(32'h3994621d),
	.w6(32'hbb869dcd),
	.w7(32'h3b121d49),
	.w8(32'h39b45d33),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1f40a),
	.w1(32'h3cc29d66),
	.w2(32'h3d0385d5),
	.w3(32'hbb2493e5),
	.w4(32'h3ce0e654),
	.w5(32'h3d041a11),
	.w6(32'h3c8dc99c),
	.w7(32'h3c9cb102),
	.w8(32'h3cbe72fa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b34e9),
	.w1(32'h3c1a180f),
	.w2(32'hba96deea),
	.w3(32'h3ad2bc96),
	.w4(32'h3c1a625b),
	.w5(32'hb81169e8),
	.w6(32'h3a1d0ffd),
	.w7(32'hbc265148),
	.w8(32'hbc040c47),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1344d2),
	.w1(32'hbbc172f8),
	.w2(32'hbb82481d),
	.w3(32'h3bfbbf7a),
	.w4(32'hbb97668a),
	.w5(32'h3afb7af7),
	.w6(32'hbbb7ea62),
	.w7(32'hbbe99adf),
	.w8(32'hbb1a1a78),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce9fdf),
	.w1(32'hbcc3260c),
	.w2(32'hbd428484),
	.w3(32'h39ff9e19),
	.w4(32'hb9b00e05),
	.w5(32'hbc02b4d2),
	.w6(32'hbcaef730),
	.w7(32'hbcc7bb14),
	.w8(32'h3bde0c71),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3fe917),
	.w1(32'h3d306f5b),
	.w2(32'h3dd574f8),
	.w3(32'hbd069abd),
	.w4(32'h3d0acbe7),
	.w5(32'h3d8283b1),
	.w6(32'h3c57de5f),
	.w7(32'h3d1f9162),
	.w8(32'h3c975b21),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d777fd6),
	.w1(32'h3c795d8b),
	.w2(32'h3c26d569),
	.w3(32'h3d0ee8b6),
	.w4(32'h3c538658),
	.w5(32'h3bf93fa8),
	.w6(32'h3bff8437),
	.w7(32'h3b49ddbd),
	.w8(32'hba7a821c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a1c5b),
	.w1(32'hbca004d9),
	.w2(32'hbcd88585),
	.w3(32'hba95830e),
	.w4(32'hbc0b9ebb),
	.w5(32'hbc8f76d5),
	.w6(32'hbc52e54b),
	.w7(32'hbc9f567f),
	.w8(32'hbbe6b0ae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf22fa),
	.w1(32'h3cd17a0d),
	.w2(32'h3cff56b5),
	.w3(32'hbc923f96),
	.w4(32'h3cd07960),
	.w5(32'h3d051fac),
	.w6(32'h3aa807b7),
	.w7(32'h3cbeec1c),
	.w8(32'h3cb8ed3f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f0d61),
	.w1(32'h3c604b4b),
	.w2(32'h3cbc74ea),
	.w3(32'h3b7bc1e6),
	.w4(32'h3c26a56d),
	.w5(32'h3c9cc88f),
	.w6(32'h3b9c46d0),
	.w7(32'h3c116269),
	.w8(32'h3c46cba4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53321f),
	.w1(32'h3c18ef93),
	.w2(32'h3c0b57f8),
	.w3(32'h3c1d080e),
	.w4(32'h3c7536c1),
	.w5(32'h3ca54d76),
	.w6(32'hbb531e5e),
	.w7(32'hbbb05a22),
	.w8(32'h3c497ef4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f2810),
	.w1(32'hbce6c75a),
	.w2(32'hbcf077e7),
	.w3(32'hbad894f3),
	.w4(32'hbcd8beb3),
	.w5(32'hbce1ed44),
	.w6(32'hbce50571),
	.w7(32'hbce94f73),
	.w8(32'hbcf08cd7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd031830),
	.w1(32'h3be52bae),
	.w2(32'h3b899645),
	.w3(32'hbbea5f27),
	.w4(32'h3d533e2a),
	.w5(32'h3cc7fa4d),
	.w6(32'hbc962fbc),
	.w7(32'h3c46e94f),
	.w8(32'h3c5cda04),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976138),
	.w1(32'h3acb1a8c),
	.w2(32'h39d82d39),
	.w3(32'h3a6f9dac),
	.w4(32'h3cc16208),
	.w5(32'h3c92a746),
	.w6(32'hbb24c5c2),
	.w7(32'h3c41ad4d),
	.w8(32'h3c56c623),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aefd7),
	.w1(32'h3c5cb40d),
	.w2(32'h3c36c7e5),
	.w3(32'hbb56386c),
	.w4(32'h3bf7e031),
	.w5(32'h3b1e3ca6),
	.w6(32'hbbaf53b0),
	.w7(32'hbc1c1997),
	.w8(32'hbc6f034c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084907),
	.w1(32'h3b053e22),
	.w2(32'hbbabf8f1),
	.w3(32'hba8f1927),
	.w4(32'h3c2b5232),
	.w5(32'h3c910fea),
	.w6(32'h3a352331),
	.w7(32'hbb872acc),
	.w8(32'h3bbc5374),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20968e),
	.w1(32'hbcef0783),
	.w2(32'hbd07a56c),
	.w3(32'hba87997d),
	.w4(32'hbbec9b30),
	.w5(32'hbb54a827),
	.w6(32'hbd07f238),
	.w7(32'hbca1e1ee),
	.w8(32'hbc4cb2c5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc843c92),
	.w1(32'h3ac56140),
	.w2(32'h3b403eb9),
	.w3(32'hbc6e7403),
	.w4(32'h3c052eea),
	.w5(32'h3b0d1755),
	.w6(32'h3b94a5f9),
	.w7(32'h3c4436e9),
	.w8(32'h3c3d7004),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9935d4),
	.w1(32'hbc0f3cbd),
	.w2(32'hbc8cae91),
	.w3(32'h3cb157d4),
	.w4(32'h3c2fbcf5),
	.w5(32'hbbb4298b),
	.w6(32'h3b893f5e),
	.w7(32'h3b8e196c),
	.w8(32'hbab9ab2c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9e92),
	.w1(32'hb8bac151),
	.w2(32'h3be89cd4),
	.w3(32'hbc00637f),
	.w4(32'h3bc7effb),
	.w5(32'h3c161666),
	.w6(32'h3b03b0ab),
	.w7(32'h3c13d7e7),
	.w8(32'h3c52e806),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849257),
	.w1(32'hbc21db8e),
	.w2(32'hbca27c56),
	.w3(32'hbaa3b212),
	.w4(32'hbc3be647),
	.w5(32'hbbf2a30a),
	.w6(32'hbb7cb29a),
	.w7(32'hbbf07973),
	.w8(32'hbbca735f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc911b34),
	.w1(32'hbc8a1217),
	.w2(32'hbcd6a327),
	.w3(32'hbbc1780f),
	.w4(32'hbc2d873e),
	.w5(32'hbc940c4a),
	.w6(32'hbb79edb5),
	.w7(32'hbbaff6b9),
	.w8(32'h3b272aa8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfce93d),
	.w1(32'hbbc02406),
	.w2(32'hbb6a40be),
	.w3(32'hbc173c57),
	.w4(32'h3b951838),
	.w5(32'h3bc3ac42),
	.w6(32'hbc0beff7),
	.w7(32'hbc3ae6f3),
	.w8(32'hbbb74263),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc839f3b),
	.w1(32'h3caffcea),
	.w2(32'h3ccd507e),
	.w3(32'hb9216668),
	.w4(32'h3caf225b),
	.w5(32'h3cd3bed8),
	.w6(32'h3bc8b7e9),
	.w7(32'h3c462309),
	.w8(32'h3bc7fc5a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc1c28),
	.w1(32'hb7e8a447),
	.w2(32'hbaeb4b5a),
	.w3(32'hbc6383e3),
	.w4(32'hba8be5f7),
	.w5(32'hbb15218c),
	.w6(32'hbbb2ccf0),
	.w7(32'hbb790ebc),
	.w8(32'h38844509),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2ef1),
	.w1(32'h3b858912),
	.w2(32'h3c0cf48b),
	.w3(32'hbb2a52e6),
	.w4(32'h3bbab980),
	.w5(32'h3c401691),
	.w6(32'h3a3b6b97),
	.w7(32'h3b2e61f8),
	.w8(32'h3bbd0553),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56fba7),
	.w1(32'hbb400e0c),
	.w2(32'hbc52e0d7),
	.w3(32'hba6b6c69),
	.w4(32'h3922e1e2),
	.w5(32'hb90075b2),
	.w6(32'h3b825be1),
	.w7(32'h3b808736),
	.w8(32'h3b22c149),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c263c),
	.w1(32'h3b69bb89),
	.w2(32'hbc1c8071),
	.w3(32'hbc8ad86e),
	.w4(32'hbc9f22aa),
	.w5(32'hbc930c75),
	.w6(32'h3ae0bad4),
	.w7(32'h3c1caf00),
	.w8(32'hbbbb037b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24a1a),
	.w1(32'h3c66a70e),
	.w2(32'h3c191d6f),
	.w3(32'hbba6aa8c),
	.w4(32'h3bdfcdb4),
	.w5(32'h3c977c58),
	.w6(32'h3b0b9fdf),
	.w7(32'hba0edf5f),
	.w8(32'h3c41f357),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c385553),
	.w1(32'hbc3a02b5),
	.w2(32'hbcce3cb8),
	.w3(32'h3b6a43a2),
	.w4(32'hbaf97af4),
	.w5(32'hbb510f96),
	.w6(32'hbba57242),
	.w7(32'hbba061a2),
	.w8(32'hbbef32ad),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb0879),
	.w1(32'h3c46ae30),
	.w2(32'h3d054f78),
	.w3(32'hbcbf5299),
	.w4(32'h3c5c0cee),
	.w5(32'h3d4e8ce1),
	.w6(32'h3ca9bbe7),
	.w7(32'h3cc0ffb3),
	.w8(32'h3cc8b69c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b6d70),
	.w1(32'hbb2e38d6),
	.w2(32'hba80ccd8),
	.w3(32'h3af89581),
	.w4(32'hbb0936c0),
	.w5(32'h3b3db51e),
	.w6(32'h3a2293b4),
	.w7(32'hba255764),
	.w8(32'hba89a964),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab24d19),
	.w1(32'hbc05f900),
	.w2(32'hbbfade3e),
	.w3(32'hbb528a9f),
	.w4(32'hbbbda6b2),
	.w5(32'h3b48213a),
	.w6(32'hbc09846b),
	.w7(32'hbb9ac62e),
	.w8(32'h3b99c7f3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc902327),
	.w1(32'hbcdb8217),
	.w2(32'hbcbdd42a),
	.w3(32'hbb6282a5),
	.w4(32'hbba6f856),
	.w5(32'hbc79d941),
	.w6(32'hbc7fdcd2),
	.w7(32'hbc8af0e2),
	.w8(32'hbc34303a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf252e),
	.w1(32'hbbe028b9),
	.w2(32'hbc815896),
	.w3(32'hbc8ea21f),
	.w4(32'hbbb872ab),
	.w5(32'hbc19bb08),
	.w6(32'h3b6eb57b),
	.w7(32'hba615992),
	.w8(32'hbb4a57be),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba260ff),
	.w1(32'h3a8d4a77),
	.w2(32'hbc0d20f4),
	.w3(32'h3be7bd5f),
	.w4(32'h3b24b61c),
	.w5(32'h3b811c85),
	.w6(32'h3c296b21),
	.w7(32'hbba7054f),
	.w8(32'h3a764d89),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4dc33),
	.w1(32'h3894dfed),
	.w2(32'h3c2861c7),
	.w3(32'h3aaa68ad),
	.w4(32'h3bcf768e),
	.w5(32'h3ccd3c31),
	.w6(32'h3c5df35f),
	.w7(32'h3ca1bd59),
	.w8(32'h3cf72f02),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16abe0),
	.w1(32'h3bb1706f),
	.w2(32'h3b91f83c),
	.w3(32'h3cbae645),
	.w4(32'h3b1dd458),
	.w5(32'hba0898ad),
	.w6(32'h3b51348a),
	.w7(32'h3b41a886),
	.w8(32'h3bd60114),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6c11),
	.w1(32'h3c505578),
	.w2(32'h3cd1a56b),
	.w3(32'h3bce7f71),
	.w4(32'h3ce1c41c),
	.w5(32'h3d2612de),
	.w6(32'h3c25f5ba),
	.w7(32'h3ca6e4d6),
	.w8(32'h3ce3f198),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caafc07),
	.w1(32'h3c151058),
	.w2(32'h3a598eff),
	.w3(32'h3cac06a4),
	.w4(32'h3c294006),
	.w5(32'h3bc3ff7a),
	.w6(32'hbb9310c4),
	.w7(32'hbae259ab),
	.w8(32'hbbdcb0c0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4c154),
	.w1(32'hbcb808dd),
	.w2(32'hbc9c6c63),
	.w3(32'hbba91e5f),
	.w4(32'hbc0aaaa1),
	.w5(32'hbbfa8502),
	.w6(32'hbbc86987),
	.w7(32'hbbb129cd),
	.w8(32'h3bcac735),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32d962),
	.w1(32'hbc0c8dc3),
	.w2(32'hbc7a078c),
	.w3(32'h3c270cb2),
	.w4(32'h3a91bd00),
	.w5(32'hbc0fd633),
	.w6(32'h3b8c668a),
	.w7(32'hbc91c145),
	.w8(32'hbc0fc37d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08bfba),
	.w1(32'h3ae654a1),
	.w2(32'h3bfdb885),
	.w3(32'hbc1fc31e),
	.w4(32'h37937c98),
	.w5(32'h3c02e678),
	.w6(32'hba00e966),
	.w7(32'hbb163d2a),
	.w8(32'h3b8a3e22),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a03e3),
	.w1(32'h3c8c55e0),
	.w2(32'h3d0bd54c),
	.w3(32'h3bc5e631),
	.w4(32'h3cbbb76e),
	.w5(32'h3d342deb),
	.w6(32'h3b9ebb4e),
	.w7(32'h3c9ce4b7),
	.w8(32'h3cbc654e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b833431),
	.w1(32'h3be0aad2),
	.w2(32'h3c124c9c),
	.w3(32'h3cc817ea),
	.w4(32'h3cac8710),
	.w5(32'h3c86196d),
	.w6(32'h3c292095),
	.w7(32'hbb063423),
	.w8(32'hbb48fa4b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3f988),
	.w1(32'h3c73b96f),
	.w2(32'h3c9749c0),
	.w3(32'hba1663fe),
	.w4(32'h3d0c3893),
	.w5(32'h3d34e44a),
	.w6(32'h3c2fa4ad),
	.w7(32'h3ca6fe7d),
	.w8(32'h3d04dcb5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f8c1a),
	.w1(32'h3c61d0e2),
	.w2(32'h3cb97d68),
	.w3(32'hbb7493b7),
	.w4(32'h39052a05),
	.w5(32'h3cf0ec0a),
	.w6(32'h3c035b78),
	.w7(32'h3c8fc0fd),
	.w8(32'h3cf9fac1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a3e9),
	.w1(32'h3a936e1d),
	.w2(32'hbb26e0bf),
	.w3(32'h3b945b6a),
	.w4(32'h3b1d4a5e),
	.w5(32'hbb9d0346),
	.w6(32'h39b89587),
	.w7(32'h3adf0563),
	.w8(32'hbbbca166),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd52fc5),
	.w1(32'h3aec484c),
	.w2(32'h3a7d4362),
	.w3(32'hbbf05990),
	.w4(32'hbaa5ae15),
	.w5(32'hba8ceea9),
	.w6(32'h3bb20932),
	.w7(32'h3bfd1530),
	.w8(32'h3c271fc4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad3e23),
	.w1(32'hbb968723),
	.w2(32'hbbed2c8e),
	.w3(32'hbb962509),
	.w4(32'hbbc07626),
	.w5(32'hbc410349),
	.w6(32'hbaa40054),
	.w7(32'hba47036f),
	.w8(32'h3a2874af),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232ed4),
	.w1(32'hba958cc0),
	.w2(32'h3beb51e8),
	.w3(32'hbc676536),
	.w4(32'h3b24612b),
	.w5(32'hba5cfaa1),
	.w6(32'hba39a95b),
	.w7(32'hba66c7dd),
	.w8(32'h3bcbfd40),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a40e2),
	.w1(32'hbc81fcab),
	.w2(32'hbc685ce6),
	.w3(32'hbc0dcc6e),
	.w4(32'hbc7d451b),
	.w5(32'hbc63c743),
	.w6(32'hbc8f0798),
	.w7(32'hbc6c4ab5),
	.w8(32'hbc171e9c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9172b3),
	.w1(32'h3b6b360d),
	.w2(32'h3a9f1d63),
	.w3(32'hbc173fe5),
	.w4(32'h3b7a906f),
	.w5(32'h3c637b12),
	.w6(32'h3c258442),
	.w7(32'h3c5f7fc7),
	.w8(32'h3c4238f8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078eac),
	.w1(32'hbb763d3b),
	.w2(32'hbb38cdbf),
	.w3(32'h3bd0af83),
	.w4(32'hbb587c3b),
	.w5(32'hbb96862f),
	.w6(32'hbb020ce6),
	.w7(32'hbb5d14ab),
	.w8(32'hbb026efd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dda19),
	.w1(32'hbc002920),
	.w2(32'hbc286bf0),
	.w3(32'hbb9e9065),
	.w4(32'h3a58eef2),
	.w5(32'h3946b0db),
	.w6(32'hbc2bceed),
	.w7(32'hbbd9f820),
	.w8(32'hbaa9fbe2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08d79c),
	.w1(32'h3c992f50),
	.w2(32'hbac94e23),
	.w3(32'hbbb8652e),
	.w4(32'h3bb93255),
	.w5(32'h3c1dc503),
	.w6(32'h3aa43a5c),
	.w7(32'hbb934bac),
	.w8(32'hbc22ec28),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143eba),
	.w1(32'h3c046348),
	.w2(32'h3c8cf945),
	.w3(32'h3aa7180f),
	.w4(32'h3c24aee6),
	.w5(32'h3c94e251),
	.w6(32'h39823a24),
	.w7(32'h3c7d75ca),
	.w8(32'h3ca1daba),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0320b7),
	.w1(32'h3ca81c2a),
	.w2(32'h3c94ff1f),
	.w3(32'hbb398e3c),
	.w4(32'h3d0cd1de),
	.w5(32'h3ccd4f80),
	.w6(32'h3b92a7c6),
	.w7(32'h3ce09721),
	.w8(32'h3cede656),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33a3d9),
	.w1(32'hbcc2b69b),
	.w2(32'hbd0a884c),
	.w3(32'h3c3254ee),
	.w4(32'hbc32e3f8),
	.w5(32'hbca1087a),
	.w6(32'h3b4394a3),
	.w7(32'hbc89b633),
	.w8(32'hba9a4260),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dadee),
	.w1(32'hbd2173fc),
	.w2(32'hbd647d72),
	.w3(32'h3c1af877),
	.w4(32'hbcf78164),
	.w5(32'hbd11b99f),
	.w6(32'hbc902d46),
	.w7(32'hbd074812),
	.w8(32'hbc3bfc85),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe6b79),
	.w1(32'hbbcc233c),
	.w2(32'h3a23a244),
	.w3(32'hbbb5c8c7),
	.w4(32'hbc2219c4),
	.w5(32'hbb8cfec2),
	.w6(32'h3b96e494),
	.w7(32'h390803f0),
	.w8(32'h3b817133),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a73c6),
	.w1(32'h3aa606cf),
	.w2(32'h3c81320d),
	.w3(32'h3c3ec69c),
	.w4(32'hbc4a455d),
	.w5(32'hbc02beb0),
	.w6(32'h3c102556),
	.w7(32'h3bb2cc37),
	.w8(32'hbb84b845),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47ec70),
	.w1(32'h3be08217),
	.w2(32'h3b0f7508),
	.w3(32'hbc885f29),
	.w4(32'h3b26ba49),
	.w5(32'h3bcadb4b),
	.w6(32'h3bee8d2a),
	.w7(32'h3b24c345),
	.w8(32'hbc572ea6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8daa33),
	.w1(32'h3bfaa336),
	.w2(32'h3c81fb26),
	.w3(32'hbb3f1a63),
	.w4(32'h3c816be2),
	.w5(32'h3cbb7d9e),
	.w6(32'h3c234be8),
	.w7(32'h3cb7f2e2),
	.w8(32'h3b9f0f88),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c9df9),
	.w1(32'h3b57c62b),
	.w2(32'h3c0dd092),
	.w3(32'h3c65e264),
	.w4(32'h3af49599),
	.w5(32'hbb7f43b8),
	.w6(32'hb9315bb1),
	.w7(32'hba2f22ca),
	.w8(32'hbb9e89f5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3015ac),
	.w1(32'hbcc0f098),
	.w2(32'hbb695563),
	.w3(32'hbb53d451),
	.w4(32'hbc054bb7),
	.w5(32'h3bc32f36),
	.w6(32'hbb103132),
	.w7(32'hbbc77116),
	.w8(32'h3a4785ad),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f9ba9),
	.w1(32'h3a2889f2),
	.w2(32'h3bfe7585),
	.w3(32'h3c86a3ac),
	.w4(32'h3c9c26e4),
	.w5(32'h3cfaa70b),
	.w6(32'h3bcef05b),
	.w7(32'h3c255b6b),
	.w8(32'h3c96b898),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf75428),
	.w1(32'h3cb66131),
	.w2(32'h3c5502d4),
	.w3(32'h3b02520d),
	.w4(32'h3be0a6bf),
	.w5(32'h3b9935e1),
	.w6(32'h3c173c41),
	.w7(32'h3c9cd49a),
	.w8(32'h3ce0fd89),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed93bd),
	.w1(32'hbb401c2b),
	.w2(32'h3bc0792d),
	.w3(32'hbc8155be),
	.w4(32'h3b216d55),
	.w5(32'h3c290d5d),
	.w6(32'hbbb895bc),
	.w7(32'hbb5e082d),
	.w8(32'h3beb97c7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e46d),
	.w1(32'h3b636ed2),
	.w2(32'hbc0b0c58),
	.w3(32'h37afa784),
	.w4(32'hbbbd50db),
	.w5(32'hbcaa3d27),
	.w6(32'h3b1b2b2f),
	.w7(32'hbb66f852),
	.w8(32'hbbd60763),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9345f9),
	.w1(32'hbc09498f),
	.w2(32'hbc950f1f),
	.w3(32'hbcd2c2f2),
	.w4(32'hbbebc0fe),
	.w5(32'hbc84c8d3),
	.w6(32'hbc7bae48),
	.w7(32'hbc16bab7),
	.w8(32'hbc5c2ef2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98af35),
	.w1(32'h3af2ae9d),
	.w2(32'h3bc4dfce),
	.w3(32'hb9a27c7e),
	.w4(32'h3bcdcd08),
	.w5(32'h3c178dd1),
	.w6(32'hbb842e89),
	.w7(32'hbc2e7c8e),
	.w8(32'hbc57e90f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137846),
	.w1(32'h3b232152),
	.w2(32'h3b703935),
	.w3(32'h3c805cb1),
	.w4(32'h3b9ab59f),
	.w5(32'h3b18d303),
	.w6(32'h3c30d66e),
	.w7(32'hba7c8912),
	.w8(32'h39426618),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f13ba),
	.w1(32'hbc428827),
	.w2(32'hbcf81e6f),
	.w3(32'hbc1731b6),
	.w4(32'hbc38e282),
	.w5(32'hbcbe4ae7),
	.w6(32'hbc316ede),
	.w7(32'hbc996f28),
	.w8(32'hbc18b3df),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee37ec),
	.w1(32'h3aaf4ef6),
	.w2(32'h39fd9505),
	.w3(32'hbc04ce6f),
	.w4(32'h3b1d352e),
	.w5(32'h3a5e018e),
	.w6(32'hb9275380),
	.w7(32'h3b6afb8d),
	.w8(32'hbb3f93d8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b2a27),
	.w1(32'h3b0845bf),
	.w2(32'hbb5415f0),
	.w3(32'hbb9f15d5),
	.w4(32'h3b9bb6bb),
	.w5(32'hba862c2b),
	.w6(32'h3b27561f),
	.w7(32'h3b102e36),
	.w8(32'hb9af364e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f0c06),
	.w1(32'hbbea0b78),
	.w2(32'hbb89c85e),
	.w3(32'hbc6af443),
	.w4(32'hbba95142),
	.w5(32'hbb8fafba),
	.w6(32'hbb1762a7),
	.w7(32'hbb8d1ce3),
	.w8(32'hbb150956),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6c3a),
	.w1(32'h3c1d7603),
	.w2(32'h3c03c926),
	.w3(32'h3b739e27),
	.w4(32'hbb0824e6),
	.w5(32'hbb8e51fc),
	.w6(32'h3c4b6ca6),
	.w7(32'h3b3a26d3),
	.w8(32'h3bd7d92f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55a712),
	.w1(32'hbbdecb90),
	.w2(32'hbc0d4cdb),
	.w3(32'hbbdabb93),
	.w4(32'hbab7eccf),
	.w5(32'h3a464c3f),
	.w6(32'h3a8cb68d),
	.w7(32'hb9c2153c),
	.w8(32'h3a9d661f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e9e6),
	.w1(32'h3c47d739),
	.w2(32'h3bfc32a7),
	.w3(32'hbb93f2e5),
	.w4(32'h3c7567bd),
	.w5(32'h3c47403f),
	.w6(32'h3bf3c151),
	.w7(32'h3b9b63a7),
	.w8(32'h3c153e1f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8987a3),
	.w1(32'h3b8b442a),
	.w2(32'h3adbfe7b),
	.w3(32'h3c2c41cf),
	.w4(32'h3680235c),
	.w5(32'h39af4ce5),
	.w6(32'h3abd3d3a),
	.w7(32'hbb34afd2),
	.w8(32'hbb182d9b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6af9d9),
	.w1(32'hbcb2a9e3),
	.w2(32'hbd01b277),
	.w3(32'hbc0e4efb),
	.w4(32'hbca1a10f),
	.w5(32'hbc9901eb),
	.w6(32'hbcd68f19),
	.w7(32'hbbc9ebc8),
	.w8(32'hbb0f6c4a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38e864),
	.w1(32'h3bd23df7),
	.w2(32'h3ccc10e0),
	.w3(32'hbb9de073),
	.w4(32'h3c4f457d),
	.w5(32'h3c2a24be),
	.w6(32'h3bbfea76),
	.w7(32'h3c6e4856),
	.w8(32'h3bd5d803),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd89df3),
	.w1(32'h3ba08cab),
	.w2(32'h3a38f092),
	.w3(32'h3c8e0eb3),
	.w4(32'h3a8dfe8c),
	.w5(32'hba92402e),
	.w6(32'h39d1efcd),
	.w7(32'hbaaedc96),
	.w8(32'hba37e52c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837fe89),
	.w1(32'hbbbeae55),
	.w2(32'hbcaa4bc7),
	.w3(32'hba61f85c),
	.w4(32'hbc5feca4),
	.w5(32'hbca4bfdf),
	.w6(32'h3bac6569),
	.w7(32'hbbdc4b23),
	.w8(32'hbbe1f0a3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc810fe1),
	.w1(32'hbbbc5f0b),
	.w2(32'hbc127bda),
	.w3(32'hbc702c00),
	.w4(32'hbc1acf3c),
	.w5(32'hbc5ad573),
	.w6(32'hbbcc617c),
	.w7(32'hbc038b9c),
	.w8(32'h3ac4b70e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1e380),
	.w1(32'h3c748499),
	.w2(32'h3ca01153),
	.w3(32'hbc2285aa),
	.w4(32'h3c3f223d),
	.w5(32'h3c99aa2a),
	.w6(32'hba8c6468),
	.w7(32'h3c888436),
	.w8(32'h3c1b0fcf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c213fa6),
	.w1(32'h3b1f503f),
	.w2(32'hbb9ca029),
	.w3(32'hb9f6e01a),
	.w4(32'hbb31a850),
	.w5(32'hbc0b43f0),
	.w6(32'hbbe3cc09),
	.w7(32'hbbab5753),
	.w8(32'hbb9832ce),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f82ae2),
	.w1(32'h3b5b8600),
	.w2(32'h3c3eed03),
	.w3(32'hbb9181d3),
	.w4(32'h3b94d760),
	.w5(32'h3bb81eff),
	.w6(32'h3a9b2c16),
	.w7(32'h3bc527bb),
	.w8(32'h3bd77bff),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule