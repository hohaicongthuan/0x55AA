module layer_8_featuremap_36(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa01b9),
	.w1(32'h3ae16e1f),
	.w2(32'hbd2a3c32),
	.w3(32'h3baaf858),
	.w4(32'hbc153e01),
	.w5(32'hbd3e46ca),
	.w6(32'hbb0acd32),
	.w7(32'hbca56665),
	.w8(32'hbca0dfe8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb434a93),
	.w1(32'hbbdd01bb),
	.w2(32'hbbd1abfb),
	.w3(32'hbc0b0b49),
	.w4(32'hbc082003),
	.w5(32'hbb415a35),
	.w6(32'hbbacd29c),
	.w7(32'hbbacbf3e),
	.w8(32'hb6a0b169),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5ceda),
	.w1(32'hbc1c9b5f),
	.w2(32'hbbd1fbe4),
	.w3(32'hbbb803e6),
	.w4(32'hbc1e0303),
	.w5(32'hbaa1c8cc),
	.w6(32'hbb068ba0),
	.w7(32'hbba4c2c0),
	.w8(32'hbadaabd2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb874fce),
	.w1(32'hbc92467e),
	.w2(32'hbc048aad),
	.w3(32'h3c2127c4),
	.w4(32'hbc8b0882),
	.w5(32'hbc4cbf66),
	.w6(32'hbb19b23a),
	.w7(32'hbba09fe6),
	.w8(32'hbbd86273),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e740d),
	.w1(32'h3a5066ed),
	.w2(32'h3b9b11fb),
	.w3(32'hbc0dd19a),
	.w4(32'h3ae7632a),
	.w5(32'h3bc3862e),
	.w6(32'hbc01f380),
	.w7(32'h39ade7a9),
	.w8(32'h3b35a79d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ccd21),
	.w1(32'h3c0b251b),
	.w2(32'h3d3c54ce),
	.w3(32'hbc7eeac0),
	.w4(32'h3d15f0f6),
	.w5(32'h3d6382ae),
	.w6(32'hbc0393bd),
	.w7(32'h3d17e673),
	.w8(32'h3d0d849b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f46d2),
	.w1(32'hb965e2ea),
	.w2(32'hb9570c56),
	.w3(32'hba27aa0d),
	.w4(32'hb915ad0a),
	.w5(32'hb9857528),
	.w6(32'hb957ba51),
	.w7(32'h3785c8e7),
	.w8(32'hba101d35),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd93f01),
	.w1(32'hbbba3591),
	.w2(32'hbc928472),
	.w3(32'h3a5db99c),
	.w4(32'hbc4b02bb),
	.w5(32'hbccdb349),
	.w6(32'hbbe3e134),
	.w7(32'hbc81c0ef),
	.w8(32'hbc7ace72),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8286da),
	.w1(32'hbbc9f5c8),
	.w2(32'hbbd993f7),
	.w3(32'hbbcfc8b0),
	.w4(32'hbb8ff33e),
	.w5(32'hbbb1ee1b),
	.w6(32'hbba4bf2b),
	.w7(32'hbb89fc49),
	.w8(32'hbc0c3795),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d7c39),
	.w1(32'hbca40b11),
	.w2(32'hbd225b42),
	.w3(32'hba5c5479),
	.w4(32'hbd195cbf),
	.w5(32'hbd386a6f),
	.w6(32'h3b3e48e8),
	.w7(32'hbcca79a1),
	.w8(32'hbcaa88bf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c309560),
	.w1(32'hbc199e6f),
	.w2(32'hbcf3eac7),
	.w3(32'h3c18a6da),
	.w4(32'hbc136ef6),
	.w5(32'hbd312982),
	.w6(32'hbae1e20a),
	.w7(32'hbc9fb2ec),
	.w8(32'hbcd95603),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c429a11),
	.w1(32'h3c3cfe72),
	.w2(32'hbbfb8879),
	.w3(32'hba39a8f8),
	.w4(32'hbb85f5fd),
	.w5(32'h3b3d4a15),
	.w6(32'hbbc6b818),
	.w7(32'h3b99a43d),
	.w8(32'h3c7e54a1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7396e6),
	.w1(32'hbba04fb1),
	.w2(32'h3acaccb1),
	.w3(32'hbb196c82),
	.w4(32'hbb1510ed),
	.w5(32'h3c08d004),
	.w6(32'hbb5b68d3),
	.w7(32'h3b189e10),
	.w8(32'h3c33e263),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb7d2c),
	.w1(32'h398b9291),
	.w2(32'h3abb6e28),
	.w3(32'hba70ff74),
	.w4(32'h3ab9e0df),
	.w5(32'h3b4aa13d),
	.w6(32'hba927a77),
	.w7(32'h3b568a21),
	.w8(32'h39e36b2b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbcd67),
	.w1(32'h35834c92),
	.w2(32'h3a832941),
	.w3(32'hba0b199f),
	.w4(32'h3a8bf862),
	.w5(32'h3adb226d),
	.w6(32'h370c0da5),
	.w7(32'h3ae514f7),
	.w8(32'h38a28b77),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06c404),
	.w1(32'h3af7e6a0),
	.w2(32'hba5b6b8f),
	.w3(32'h3a3392f8),
	.w4(32'h3ab0eb66),
	.w5(32'hba21ce35),
	.w6(32'h3b093f1a),
	.w7(32'h3a846c18),
	.w8(32'hbb06183f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce8fde),
	.w1(32'h3b25725e),
	.w2(32'hbb718cd5),
	.w3(32'h3c516b7f),
	.w4(32'h3b90ae8e),
	.w5(32'hbc5022c6),
	.w6(32'h3c15992b),
	.w7(32'h3bf18460),
	.w8(32'hbaa5ed06),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae93b86),
	.w1(32'hbae23218),
	.w2(32'hbc5c48da),
	.w3(32'hbbe22f00),
	.w4(32'hbbf37039),
	.w5(32'hbc23fa23),
	.w6(32'hbc262b88),
	.w7(32'hbb970044),
	.w8(32'h3a588a47),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db48d62),
	.w1(32'h3c9ccece),
	.w2(32'hbd817007),
	.w3(32'h3d1959a0),
	.w4(32'hbc9dc683),
	.w5(32'hbdb17196),
	.w6(32'h3c0318b8),
	.w7(32'hbd771f6f),
	.w8(32'hbbc47a2d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a8eed),
	.w1(32'hbba84d6a),
	.w2(32'h3b82ede6),
	.w3(32'hbb781971),
	.w4(32'hbbd1b5d4),
	.w5(32'h3c3fbd2c),
	.w6(32'hbc45832c),
	.w7(32'hbbbf18c3),
	.w8(32'h3d00e206),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881a993),
	.w1(32'h3c9d6bd1),
	.w2(32'h3acb37c8),
	.w3(32'hbb0aa47c),
	.w4(32'h3d1dccdd),
	.w5(32'h3ca92231),
	.w6(32'h3a3f7399),
	.w7(32'h3c21fe57),
	.w8(32'h3bc64364),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4246c3),
	.w1(32'hbc82a27f),
	.w2(32'h3b52f5d3),
	.w3(32'hbc98c968),
	.w4(32'hbc7b4f6e),
	.w5(32'h3bea569e),
	.w6(32'hbc8720a9),
	.w7(32'hbc67ee92),
	.w8(32'h3b9f2c22),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d18e960),
	.w1(32'h3c6f1087),
	.w2(32'hbdd4ab9a),
	.w3(32'h3d2e9703),
	.w4(32'hbc4e1af2),
	.w5(32'hbe06ba26),
	.w6(32'h3c910748),
	.w7(32'hbd4c386f),
	.w8(32'hbda62dc8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb0af),
	.w1(32'hbc6868a2),
	.w2(32'hbb909b9a),
	.w3(32'hbc39736a),
	.w4(32'hbb9ca4e9),
	.w5(32'h3af6036d),
	.w6(32'hbc004c2c),
	.w7(32'h3a8fee11),
	.w8(32'hb97c0e02),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b306ab2),
	.w1(32'h3bdda272),
	.w2(32'h3bf75c4e),
	.w3(32'h3ba5fa9c),
	.w4(32'h3bfa46d9),
	.w5(32'h3bea04bd),
	.w6(32'h3bb51675),
	.w7(32'h3b5b294a),
	.w8(32'h3c227e4f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c415dfa),
	.w1(32'h3caa613a),
	.w2(32'hbb72b5c1),
	.w3(32'h3a78a90d),
	.w4(32'h3b851ff6),
	.w5(32'hbc6a7971),
	.w6(32'hb92a5fb6),
	.w7(32'hbc159a68),
	.w8(32'hbb21ee4d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9971e7a),
	.w1(32'hbad26d52),
	.w2(32'hbacc5369),
	.w3(32'h39e4977b),
	.w4(32'hba8aabc5),
	.w5(32'hbac6d8b8),
	.w6(32'hba990e45),
	.w7(32'hbb3bdd08),
	.w8(32'h3a4f8757),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e01913d),
	.w1(32'h3d47127b),
	.w2(32'hbdc7426e),
	.w3(32'h3d88896d),
	.w4(32'h3dffab39),
	.w5(32'hbda37f9a),
	.w6(32'h3de62d8f),
	.w7(32'h3b7db6c0),
	.w8(32'hbdafcdf5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb1955),
	.w1(32'h3a97b57d),
	.w2(32'hbc3b81e8),
	.w3(32'h3c013a21),
	.w4(32'hbb642672),
	.w5(32'hbc88dc87),
	.w6(32'hbb2df892),
	.w7(32'hbbe1d665),
	.w8(32'h39ff1eaa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0eab7),
	.w1(32'hbb15059f),
	.w2(32'hba4518e6),
	.w3(32'h37653aa9),
	.w4(32'hba6e2352),
	.w5(32'hba1d49bd),
	.w6(32'h39dd801e),
	.w7(32'hba56ad89),
	.w8(32'h3ac8a911),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf76103),
	.w1(32'hbc39868d),
	.w2(32'hbc3bae7d),
	.w3(32'hbc0b84fd),
	.w4(32'hbc0304a6),
	.w5(32'hbc2611f2),
	.w6(32'hbc078da9),
	.w7(32'hbc3013f0),
	.w8(32'hbb904488),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb1dfc),
	.w1(32'h3c42fd70),
	.w2(32'h3c74f21a),
	.w3(32'hbb1e74c4),
	.w4(32'h3c760657),
	.w5(32'h3ca94b4f),
	.w6(32'hbacb3cf7),
	.w7(32'h3ae4f726),
	.w8(32'h3b019fad),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901961),
	.w1(32'hbbdffac4),
	.w2(32'hbbeb2388),
	.w3(32'hbb7039fc),
	.w4(32'hbb6ca051),
	.w5(32'hbb9fbdde),
	.w6(32'hbb68a4f0),
	.w7(32'hbaccd1a5),
	.w8(32'h39f1a88c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231711),
	.w1(32'h3b2c38ad),
	.w2(32'hbb2cbd29),
	.w3(32'hbb28923f),
	.w4(32'hbbddd00c),
	.w5(32'hbba5b5af),
	.w6(32'h3afae13e),
	.w7(32'hbb54592d),
	.w8(32'hba55ef1f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc691a50),
	.w1(32'hbc025e44),
	.w2(32'h3c104743),
	.w3(32'hbc387b5d),
	.w4(32'hbafc5053),
	.w5(32'h3cc813fc),
	.w6(32'hba65a27f),
	.w7(32'h3c0d9bfe),
	.w8(32'h3ca2614b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c603e76),
	.w1(32'h3cb50802),
	.w2(32'hbcd65d9a),
	.w3(32'h3c44f22e),
	.w4(32'h3bd814db),
	.w5(32'hbcb7cd76),
	.w6(32'h3c29e8bc),
	.w7(32'hbc25c438),
	.w8(32'hbbd737f5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39127fe4),
	.w1(32'h38fc4923),
	.w2(32'hbae632fd),
	.w3(32'hb9a12b50),
	.w4(32'hba82280e),
	.w5(32'hbafcdce2),
	.w6(32'hb9d00dc6),
	.w7(32'hbafb4018),
	.w8(32'h3abefca8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176c9e),
	.w1(32'hbba2af96),
	.w2(32'hbb98cadb),
	.w3(32'hbb9a2f59),
	.w4(32'hbbbeebf5),
	.w5(32'hbb7ec242),
	.w6(32'hbb9f0eb1),
	.w7(32'hbbc98b04),
	.w8(32'hbb9760f7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee9e0),
	.w1(32'h37e3fb40),
	.w2(32'h3b276156),
	.w3(32'hba0b886f),
	.w4(32'h3b37c19b),
	.w5(32'h3b5f9051),
	.w6(32'h3a370ead),
	.w7(32'h3b6b56d2),
	.w8(32'h3a78347b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52afbe),
	.w1(32'h3ab06ecc),
	.w2(32'hbaaf8a19),
	.w3(32'h3b63ee08),
	.w4(32'h3ac86363),
	.w5(32'hbafec305),
	.w6(32'h3aa94f2a),
	.w7(32'hbb061c2e),
	.w8(32'hba5c1375),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1557f2),
	.w1(32'h3c7c16d5),
	.w2(32'h3d0b3e51),
	.w3(32'h3d0554fd),
	.w4(32'hbc253429),
	.w5(32'h3cca5daa),
	.w6(32'hbbbe2aa1),
	.w7(32'hbbbf7449),
	.w8(32'h3d84b6e0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d12ffaa),
	.w1(32'h3c059c55),
	.w2(32'hbc543048),
	.w3(32'h3cc984e6),
	.w4(32'h39c1e726),
	.w5(32'hbcad13cf),
	.w6(32'h3c9449ba),
	.w7(32'hbc286822),
	.w8(32'h3b0b56b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc58e5a),
	.w1(32'hbcbb27ab),
	.w2(32'hbc575cf9),
	.w3(32'h3bdf9530),
	.w4(32'hbca30ccc),
	.w5(32'hbccd6fe8),
	.w6(32'hbc890c16),
	.w7(32'hbbfa1941),
	.w8(32'h3c81e366),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf85983),
	.w1(32'h3c60a02a),
	.w2(32'hbcb681b5),
	.w3(32'h3c90882f),
	.w4(32'h3ab7994f),
	.w5(32'hbcd48303),
	.w6(32'h3c33d33e),
	.w7(32'hbc324c47),
	.w8(32'h3c2aeeea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d514771),
	.w1(32'h3c5864ab),
	.w2(32'hbd547811),
	.w3(32'h3cd7a6b8),
	.w4(32'hbc807b5b),
	.w5(32'hbd9ff9f3),
	.w6(32'h3c55025a),
	.w7(32'hbd20afbd),
	.w8(32'hbcc850ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d115503),
	.w1(32'hbae9cee3),
	.w2(32'hbcf6fd36),
	.w3(32'h3caa3b65),
	.w4(32'hbc8fd7a4),
	.w5(32'hbd0b0efb),
	.w6(32'h3b75aad7),
	.w7(32'hbcbd7df9),
	.w8(32'hb9892de5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f67a3),
	.w1(32'hbbe78e61),
	.w2(32'hba656f66),
	.w3(32'h3ca2cb1a),
	.w4(32'h3afeb527),
	.w5(32'hbc4e42f9),
	.w6(32'hbc085f08),
	.w7(32'h3abc36f2),
	.w8(32'h394483a2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3f349),
	.w1(32'h3cb79af7),
	.w2(32'hbd30266b),
	.w3(32'h3c6a37a5),
	.w4(32'hbc0b5409),
	.w5(32'hbd6279d9),
	.w6(32'h3c959a8c),
	.w7(32'hbcb5750b),
	.w8(32'hbd9d2c8a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a964e),
	.w1(32'hbc47d4be),
	.w2(32'h3d201089),
	.w3(32'hbcc3c917),
	.w4(32'h3b639ea5),
	.w5(32'h3d3107b3),
	.w6(32'hbcafa21e),
	.w7(32'h3c4de522),
	.w8(32'h3cc68ef2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc86a0),
	.w1(32'hbb01619f),
	.w2(32'hbd362169),
	.w3(32'h3c2a08b8),
	.w4(32'hbcd5408a),
	.w5(32'hbd59908a),
	.w6(32'h3b6b6499),
	.w7(32'hbc9f133f),
	.w8(32'h3a67236c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c646e99),
	.w1(32'h3c23b3a4),
	.w2(32'h3b1834ca),
	.w3(32'hbc26ed4b),
	.w4(32'h3bbd29fc),
	.w5(32'h3ca0b902),
	.w6(32'hbc81485c),
	.w7(32'h3c069634),
	.w8(32'h3d4304fb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d95762f),
	.w1(32'h3cfa9cf7),
	.w2(32'hba3772ff),
	.w3(32'h3d52e89d),
	.w4(32'hbb16447a),
	.w5(32'hbd3b4fbe),
	.w6(32'h3d0bc64e),
	.w7(32'hbca97bfc),
	.w8(32'h3cbfb39f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdaded0),
	.w1(32'h3c666de5),
	.w2(32'hbbef9f4f),
	.w3(32'h3c4019e5),
	.w4(32'hbb79d158),
	.w5(32'hbc859b8d),
	.w6(32'h3c825ce6),
	.w7(32'hbbced111),
	.w8(32'h3c484e3c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0638ca),
	.w1(32'h3cb15e6f),
	.w2(32'hbc8a81dd),
	.w3(32'h3c631fc7),
	.w4(32'hbc507a8a),
	.w5(32'hbcf1e327),
	.w6(32'h3c866672),
	.w7(32'hbbe42e6b),
	.w8(32'hbbdd3ebb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79772e),
	.w1(32'hbc13c270),
	.w2(32'h3b1d77da),
	.w3(32'h3b81504f),
	.w4(32'hbaf6fa73),
	.w5(32'hbc09f2a9),
	.w6(32'h3c1f10d6),
	.w7(32'hbb1e3092),
	.w8(32'hbb86ffc8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d411336),
	.w1(32'h3d1535b7),
	.w2(32'hbd8d09f6),
	.w3(32'hbb0433a1),
	.w4(32'hbca61a69),
	.w5(32'hbd2cfc5f),
	.w6(32'h3b807350),
	.w7(32'hbcf220aa),
	.w8(32'hbca72cea),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb122d3),
	.w1(32'hbb32a505),
	.w2(32'hbc936a89),
	.w3(32'h3b6a6160),
	.w4(32'hba54b23c),
	.w5(32'hbc12c0bd),
	.w6(32'h3afd45f1),
	.w7(32'h3babbe25),
	.w8(32'h3c8bc5df),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced4563),
	.w1(32'hbbf2756a),
	.w2(32'hbc5738dd),
	.w3(32'h3c1f2ea4),
	.w4(32'hbc4e45c7),
	.w5(32'hbd137de6),
	.w6(32'h3c798dfa),
	.w7(32'hbcb4d42d),
	.w8(32'hbc48cf94),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1fad9),
	.w1(32'h3c878e6f),
	.w2(32'hbc4905b1),
	.w3(32'h3cbdead1),
	.w4(32'h3c899f34),
	.w5(32'hbca11db9),
	.w6(32'h3c8d4adf),
	.w7(32'h3ba960e5),
	.w8(32'h3bc23f67),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8dcfe),
	.w1(32'h3aafc3ea),
	.w2(32'hbc7fe85e),
	.w3(32'h3c9e37c9),
	.w4(32'hbaba928e),
	.w5(32'hbce78fb4),
	.w6(32'h3ca1420a),
	.w7(32'hbc804566),
	.w8(32'hbc8b8fc0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c436d),
	.w1(32'hbc6ca259),
	.w2(32'hbc559ba2),
	.w3(32'h3c69ce33),
	.w4(32'hbb538e36),
	.w5(32'hbc4d31a3),
	.w6(32'h3b23a9de),
	.w7(32'h3b011754),
	.w8(32'h3c45a914),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bdab6),
	.w1(32'h3b8a4b54),
	.w2(32'hbcbc020d),
	.w3(32'h3c1de811),
	.w4(32'hbbcfe42a),
	.w5(32'hbcbdf9bc),
	.w6(32'h3aa498ce),
	.w7(32'hbc73da5e),
	.w8(32'h3ce38c86),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3a004f),
	.w1(32'h3cad0019),
	.w2(32'hbc1eabdd),
	.w3(32'h3c9fbb14),
	.w4(32'hbc880757),
	.w5(32'hbc8ec324),
	.w6(32'h3c5e0ed8),
	.w7(32'hbc849e7b),
	.w8(32'h3d38f994),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b23e7),
	.w1(32'hbc61403a),
	.w2(32'hbc5f5d41),
	.w3(32'h3b982220),
	.w4(32'hbc2eb0e1),
	.w5(32'hbbbd78cd),
	.w6(32'hba1e999c),
	.w7(32'hbc36ea00),
	.w8(32'h3c3d1049),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f4286),
	.w1(32'h3b54d27d),
	.w2(32'hbc503f2e),
	.w3(32'h3bae4013),
	.w4(32'hba8f6ee6),
	.w5(32'hbc6262f0),
	.w6(32'h3bb27a25),
	.w7(32'hbc024bba),
	.w8(32'h3bafeaf7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cc192),
	.w1(32'h3be86529),
	.w2(32'hbc87b424),
	.w3(32'h3c3019b2),
	.w4(32'h38f17be6),
	.w5(32'hbc8cabdc),
	.w6(32'h3bc3decb),
	.w7(32'hbbb4a45c),
	.w8(32'h3b318bc5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f5451),
	.w1(32'h3bd772a9),
	.w2(32'h3c246bd4),
	.w3(32'h3c047022),
	.w4(32'h3b923130),
	.w5(32'h3bdb082b),
	.w6(32'h3c04f027),
	.w7(32'h3ad117c7),
	.w8(32'h3c67b323),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d009605),
	.w1(32'h3cb71e22),
	.w2(32'hbc85d3b0),
	.w3(32'h3c1835d5),
	.w4(32'h3b504abc),
	.w5(32'hbb0678d8),
	.w6(32'hbc0176a6),
	.w7(32'hbb2ba3bc),
	.w8(32'h3d198eeb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6f382),
	.w1(32'h3bcb0f77),
	.w2(32'hbc87a808),
	.w3(32'h3c283d50),
	.w4(32'hbaf2ca2a),
	.w5(32'hbcb9ab21),
	.w6(32'h3c201ead),
	.w7(32'hbc004003),
	.w8(32'h3d3f218e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9a72f9),
	.w1(32'h3d97148f),
	.w2(32'hbd783b68),
	.w3(32'h3d6d8c1e),
	.w4(32'h3d19d59f),
	.w5(32'hbdcb0b0f),
	.w6(32'h3d8c3f08),
	.w7(32'hbd0f168f),
	.w8(32'hbd7e9203),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52354a),
	.w1(32'h3bcb9b24),
	.w2(32'hbbf743ea),
	.w3(32'h3c0827fe),
	.w4(32'h3ae28b3b),
	.w5(32'hbc0f17ec),
	.w6(32'h3bedf412),
	.w7(32'hbb554782),
	.w8(32'h3c9ecfc7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9050e),
	.w1(32'hbab9e116),
	.w2(32'hbc9e2514),
	.w3(32'h3c856834),
	.w4(32'hbc05bfe2),
	.w5(32'hbcf5eb9f),
	.w6(32'h3c63e455),
	.w7(32'hbc70e0e0),
	.w8(32'h3c6ec575),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91f37e),
	.w1(32'h3ba2f54c),
	.w2(32'hbc3fb25a),
	.w3(32'h3c35491f),
	.w4(32'hbac05e8e),
	.w5(32'hbc6a7d3e),
	.w6(32'h3c2aa60b),
	.w7(32'hbb464ac8),
	.w8(32'h3bc717fc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa7af6),
	.w1(32'hb96dc2ae),
	.w2(32'hbcff3483),
	.w3(32'hbc3dfc01),
	.w4(32'hbcd47bae),
	.w5(32'hbcd2d1b8),
	.w6(32'hbb4d5594),
	.w7(32'h3be3f82d),
	.w8(32'h3ca0295e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9aaca),
	.w1(32'h3b63b0b4),
	.w2(32'hbc9d99af),
	.w3(32'h3c07abbf),
	.w4(32'hbbe80b71),
	.w5(32'hbccffdf4),
	.w6(32'h3c09ac61),
	.w7(32'hbc2b6df7),
	.w8(32'h3c0fd5da),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5df9e5),
	.w1(32'h3c1ab8f4),
	.w2(32'hbbafeab2),
	.w3(32'h3c5d3f22),
	.w4(32'h3be7a58e),
	.w5(32'hbbeb7934),
	.w6(32'h3c1b6d62),
	.w7(32'h3b4b1ff2),
	.w8(32'h3c76a7d0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75d852),
	.w1(32'h3b7a92b0),
	.w2(32'hbc62bae6),
	.w3(32'h3c03de80),
	.w4(32'hbb5de45e),
	.w5(32'hbc7de0e8),
	.w6(32'h3bbb9410),
	.w7(32'hbbfd3a19),
	.w8(32'h3d526a5f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dacacfb),
	.w1(32'h3cf4622f),
	.w2(32'hbd65e886),
	.w3(32'h3d37ab2e),
	.w4(32'hbb11875d),
	.w5(32'hbd841d43),
	.w6(32'h3cfec80d),
	.w7(32'hbcef4f49),
	.w8(32'h3c6f8553),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d599514),
	.w1(32'h3c41a749),
	.w2(32'hbd544ba5),
	.w3(32'h3d02921a),
	.w4(32'hbc48c771),
	.w5(32'hbd45e997),
	.w6(32'h3d07ef68),
	.w7(32'hbcce462f),
	.w8(32'hbb788e2c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f9df0),
	.w1(32'h3b193353),
	.w2(32'hbb9124ca),
	.w3(32'h3bdd8415),
	.w4(32'hba8b609f),
	.w5(32'hbb3f1189),
	.w6(32'h3b8ff99c),
	.w7(32'h3a3ccc64),
	.w8(32'h3c50b2cf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb228e31),
	.w1(32'hbc813051),
	.w2(32'hbc8f4665),
	.w3(32'h3b691c0e),
	.w4(32'hbbe48a13),
	.w5(32'hbcac6e82),
	.w6(32'h3bf14dd4),
	.w7(32'h3b8c0933),
	.w8(32'h3bbe044b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12f1fe),
	.w1(32'hbbe4db62),
	.w2(32'hbb8c9531),
	.w3(32'h3bbeb123),
	.w4(32'h3c24be57),
	.w5(32'hbc98213b),
	.w6(32'h3c95ce65),
	.w7(32'h3b945649),
	.w8(32'hb9dcd6a2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3e650f),
	.w1(32'h3c53036d),
	.w2(32'hbcc810ac),
	.w3(32'h3cb21ba3),
	.w4(32'hbc6056cf),
	.w5(32'hbd15a909),
	.w6(32'h3c00508c),
	.w7(32'hbcdd6865),
	.w8(32'h3c4a9deb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfc618c),
	.w1(32'h3d190cf2),
	.w2(32'h3d49dbe6),
	.w3(32'h3ce1e4f3),
	.w4(32'hbcd01229),
	.w5(32'h3cd13d6f),
	.w6(32'h3bd4418b),
	.w7(32'hbcc50fb3),
	.w8(32'h3da737de),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d47545f),
	.w1(32'h3c9574a2),
	.w2(32'hbd6b9927),
	.w3(32'h3cd533b0),
	.w4(32'hbc856fcb),
	.w5(32'hbd957227),
	.w6(32'h3bbf7a8d),
	.w7(32'hbd12a9fb),
	.w8(32'h3bf007f4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf1b1e),
	.w1(32'hbb910a29),
	.w2(32'hbcb255e7),
	.w3(32'h3cc5a07e),
	.w4(32'h3b3d6c53),
	.w5(32'hbd486e9c),
	.w6(32'h3cd25a9c),
	.w7(32'hbab7aea0),
	.w8(32'hbda26bc3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd700fdd),
	.w1(32'hbbf68e36),
	.w2(32'h3d56077a),
	.w3(32'hbcee7bb6),
	.w4(32'h3c355413),
	.w5(32'h3d63b52d),
	.w6(32'hbcadbee9),
	.w7(32'h3ccee4cc),
	.w8(32'h3bb79720),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8db63c),
	.w1(32'h3b5adec1),
	.w2(32'hbbba2c1f),
	.w3(32'hba3d185e),
	.w4(32'hbaf8f217),
	.w5(32'hbc2c9d98),
	.w6(32'h3c1ca66f),
	.w7(32'hbaee8b2b),
	.w8(32'h3d14a9fc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d040312),
	.w1(32'hbc13a83b),
	.w2(32'hbce79e0d),
	.w3(32'h3ce592bf),
	.w4(32'hbc111097),
	.w5(32'hbd0623c4),
	.w6(32'h3c4804d5),
	.w7(32'hbbd18326),
	.w8(32'hbd647d84),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd671199),
	.w1(32'hbbd403c0),
	.w2(32'h3d47894f),
	.w3(32'hbcdef0ed),
	.w4(32'h3c368c50),
	.w5(32'h3d5173ba),
	.w6(32'hbca9e08e),
	.w7(32'h3cbe4c5e),
	.w8(32'hbd4847b9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd358ce0),
	.w1(32'hbbb53184),
	.w2(32'h3d34900d),
	.w3(32'hbce3e84d),
	.w4(32'h3c5ec55a),
	.w5(32'h3d36bc85),
	.w6(32'hbc9fa82e),
	.w7(32'h3d01b898),
	.w8(32'h3c5a5611),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d4784),
	.w1(32'hbb958136),
	.w2(32'hbb6b29c7),
	.w3(32'h3bd4c7eb),
	.w4(32'hbba59849),
	.w5(32'hbc03e354),
	.w6(32'hb96792bf),
	.w7(32'hbb21fd20),
	.w8(32'h3c8d3db2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156fec),
	.w1(32'h3c320220),
	.w2(32'h3ca706b6),
	.w3(32'hbb6e9a08),
	.w4(32'hbaafc615),
	.w5(32'h3b75090a),
	.w6(32'h3c52fb85),
	.w7(32'hbb531b04),
	.w8(32'h3c42c0b3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb365f),
	.w1(32'hbc0dd40e),
	.w2(32'hbc89d4b3),
	.w3(32'h3bdfbce6),
	.w4(32'hbc65b72b),
	.w5(32'hbc94d9b2),
	.w6(32'hbaaab9fa),
	.w7(32'hbc8a7962),
	.w8(32'h3ccb89f7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1cd84d),
	.w1(32'h3c62a9c0),
	.w2(32'hbc80175d),
	.w3(32'hbcc9967c),
	.w4(32'hbc9df2cc),
	.w5(32'h3ba1c63c),
	.w6(32'h3bb7b2c6),
	.w7(32'hbc4045f0),
	.w8(32'h3d1f12ab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28ca6c),
	.w1(32'h3c4b1aa6),
	.w2(32'hbd0cb2cc),
	.w3(32'h3d47c803),
	.w4(32'h3ba0d0cf),
	.w5(32'hbd3cda15),
	.w6(32'h3cc4a7f3),
	.w7(32'hbcdaeaba),
	.w8(32'hbba557d8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cade6fc),
	.w1(32'h3c3aa4dc),
	.w2(32'h3c39ac95),
	.w3(32'h3c816e46),
	.w4(32'h3939d2b7),
	.w5(32'h3c0c0ca3),
	.w6(32'h3c3364bf),
	.w7(32'h3c29c090),
	.w8(32'h3cb641a7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ffc39),
	.w1(32'hbb906c16),
	.w2(32'hbb39b17d),
	.w3(32'hbbc568ae),
	.w4(32'hbb76eb29),
	.w5(32'hbbef5f92),
	.w6(32'h3aa8f7c7),
	.w7(32'hbab02c51),
	.w8(32'h3d37c8cb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d497c58),
	.w1(32'h3c2f5549),
	.w2(32'hbd0ac391),
	.w3(32'h3cb74e01),
	.w4(32'hbc1e6d75),
	.w5(32'hbd196ab2),
	.w6(32'h3ca50b81),
	.w7(32'hbc29712a),
	.w8(32'h3c08e525),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23cbf4),
	.w1(32'h3b4082ab),
	.w2(32'hbc292853),
	.w3(32'h3b8483a9),
	.w4(32'hbb0b491e),
	.w5(32'hbc6213d5),
	.w6(32'h3c0fc715),
	.w7(32'hbb37abc7),
	.w8(32'h3d02d98d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc854b9),
	.w1(32'hbc1ba5f4),
	.w2(32'hbcd0acb5),
	.w3(32'h3ca777cc),
	.w4(32'hbc3fe20c),
	.w5(32'hbd0a65e4),
	.w6(32'h3c0a2e0b),
	.w7(32'hbc7f99f6),
	.w8(32'h3c31b8a2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc01b8),
	.w1(32'hbb1bfc6f),
	.w2(32'hbc6ffb8b),
	.w3(32'hba66823a),
	.w4(32'hbbe69fbc),
	.w5(32'hbc51ebfc),
	.w6(32'hba510544),
	.w7(32'hbc34c6a0),
	.w8(32'h3d314629),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ccd3e),
	.w1(32'h3cb67728),
	.w2(32'hbd023daa),
	.w3(32'h3d0c15ac),
	.w4(32'h3b165a79),
	.w5(32'hbcf1f482),
	.w6(32'h3cf0252f),
	.w7(32'hbbc49446),
	.w8(32'h3ca0d347),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d521f),
	.w1(32'hbc9d1492),
	.w2(32'h39e48fd0),
	.w3(32'hba338c5a),
	.w4(32'hbc4ee2e5),
	.w5(32'hbc0706f7),
	.w6(32'h3bf4f1eb),
	.w7(32'hbbe84457),
	.w8(32'hbcc674f0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceec307),
	.w1(32'hbc225689),
	.w2(32'h3cb35e37),
	.w3(32'hbc904de9),
	.w4(32'hba6da902),
	.w5(32'h3cd31235),
	.w6(32'hbc3976c0),
	.w7(32'h3bd3d19b),
	.w8(32'h3a85b17c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf2e83),
	.w1(32'h3cf9049b),
	.w2(32'hbcad9a72),
	.w3(32'h3c703893),
	.w4(32'h3c6b6ea3),
	.w5(32'hbd1dbdbe),
	.w6(32'h3ce63145),
	.w7(32'hbb7af0e3),
	.w8(32'hbcb94f35),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80c4c7),
	.w1(32'h3b257eb0),
	.w2(32'hba2362c9),
	.w3(32'hbc9132dd),
	.w4(32'hbcdde6b2),
	.w5(32'hbbe6e6fc),
	.w6(32'hbc7e8b08),
	.w7(32'hbbf861e1),
	.w8(32'h3801f514),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfac599),
	.w1(32'hbbcfb12f),
	.w2(32'h3c2d09d9),
	.w3(32'hbc3ce814),
	.w4(32'hbb5deec0),
	.w5(32'h3c12dd73),
	.w6(32'hbb0f7c62),
	.w7(32'hbbc4ce9d),
	.w8(32'h3b901a8d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8de143),
	.w1(32'hbb1635cd),
	.w2(32'h3af61a57),
	.w3(32'hbc2b31c5),
	.w4(32'hbbed3352),
	.w5(32'hbb8ca3b0),
	.w6(32'hbb3d055b),
	.w7(32'hbbc69e72),
	.w8(32'h3b107094),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0df0ba),
	.w1(32'h3ae6a364),
	.w2(32'hbc182fad),
	.w3(32'h3b045582),
	.w4(32'hbbd12d7e),
	.w5(32'hbc2dbbb3),
	.w6(32'h3bc2d16c),
	.w7(32'hbb61010e),
	.w8(32'h3c890f11),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c101942),
	.w1(32'h3d339ca7),
	.w2(32'h3badb8bc),
	.w3(32'hbc273247),
	.w4(32'h3c148c4e),
	.w5(32'h3cf3e306),
	.w6(32'h3bf35387),
	.w7(32'hbc50b5cc),
	.w8(32'h3cd6059b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e03d8),
	.w1(32'h3b9a9ffd),
	.w2(32'h3cad773e),
	.w3(32'h3b46aca0),
	.w4(32'hbb4ee866),
	.w5(32'h3c380b41),
	.w6(32'hbb8f0000),
	.w7(32'hbbd097ff),
	.w8(32'h3c7cfffc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cee16),
	.w1(32'hbc9c7616),
	.w2(32'hbd1a0ee8),
	.w3(32'hbcee7ecb),
	.w4(32'hbd33a31a),
	.w5(32'hbcd9270c),
	.w6(32'hbc182dda),
	.w7(32'hbcd1e414),
	.w8(32'hbb515add),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add5d7b),
	.w1(32'h3b8178bd),
	.w2(32'hbacd7246),
	.w3(32'hbb524fd4),
	.w4(32'hbb1fafd8),
	.w5(32'hbbe07436),
	.w6(32'h3b2b1e92),
	.w7(32'hbb54429a),
	.w8(32'hbab9ebad),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c3d76),
	.w1(32'hb8d80c6a),
	.w2(32'h3ba6ec48),
	.w3(32'h3c0970eb),
	.w4(32'h3a8032af),
	.w5(32'hb9cf94cd),
	.w6(32'h3b1004d4),
	.w7(32'hba7d3222),
	.w8(32'hbb05903b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9bc50),
	.w1(32'hbb677aad),
	.w2(32'h3c2a35c3),
	.w3(32'h3bd18c67),
	.w4(32'h3bd85c0b),
	.w5(32'h3bc55cd3),
	.w6(32'h3b8eadac),
	.w7(32'h3bb7a2de),
	.w8(32'h3c03dacb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1515f4),
	.w1(32'h3b8ced04),
	.w2(32'h3c83ca9f),
	.w3(32'h3bbec0f5),
	.w4(32'hbc2deef8),
	.w5(32'hbb5b73f0),
	.w6(32'h3b414cb1),
	.w7(32'h3b8679fc),
	.w8(32'h3b879d07),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4210c0),
	.w1(32'h3c5dd5c1),
	.w2(32'hbb72cc55),
	.w3(32'h3bdcf074),
	.w4(32'hbbd9ea7d),
	.w5(32'hbc27835b),
	.w6(32'h3ba5526f),
	.w7(32'hbc3ace67),
	.w8(32'hbaee7d97),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a389297),
	.w1(32'h3ba8255b),
	.w2(32'h3c10e840),
	.w3(32'hbbe30aa1),
	.w4(32'hbba58aac),
	.w5(32'h3bf24eed),
	.w6(32'hbca60cca),
	.w7(32'hb99493c2),
	.w8(32'h3a15a9bd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31e94e),
	.w1(32'h3c9148ae),
	.w2(32'hbc85d383),
	.w3(32'hbb9895fc),
	.w4(32'h39ffc39a),
	.w5(32'hbba9f491),
	.w6(32'h3c04d966),
	.w7(32'hbc6c4f2c),
	.w8(32'h3c40b198),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f8364),
	.w1(32'hbc82ca58),
	.w2(32'hbc4e79cf),
	.w3(32'hbb623364),
	.w4(32'hbca7e27d),
	.w5(32'hbccaea30),
	.w6(32'h3c1a0504),
	.w7(32'hbc3bcfb6),
	.w8(32'hbc98b716),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93324a),
	.w1(32'h3c660371),
	.w2(32'h3c3dd5ad),
	.w3(32'h3c554df9),
	.w4(32'h3b936dfb),
	.w5(32'hbc3304ec),
	.w6(32'hbb80a089),
	.w7(32'h3ca234dc),
	.w8(32'h3c2ed918),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba631f1e),
	.w1(32'hbb87780e),
	.w2(32'hbd23e04f),
	.w3(32'hbcb67753),
	.w4(32'hbd1ae4ff),
	.w5(32'hbcf39b2d),
	.w6(32'hbb595389),
	.w7(32'hbcb1aa3b),
	.w8(32'h3a6d56c3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e6d18),
	.w1(32'h3c9351fb),
	.w2(32'h3c6b4e67),
	.w3(32'hbafdb9d8),
	.w4(32'h3ae717d7),
	.w5(32'h3c0e6746),
	.w6(32'h3b2f7c4f),
	.w7(32'h3b943fd5),
	.w8(32'h3b88d414),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2377f),
	.w1(32'h3bb942a6),
	.w2(32'hbc716577),
	.w3(32'hbc670c72),
	.w4(32'hbc59ec7c),
	.w5(32'h3c0cb141),
	.w6(32'h3b340c5c),
	.w7(32'hbc8f1f4d),
	.w8(32'h3b15328f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c218692),
	.w1(32'h3cdbd178),
	.w2(32'h3b75606f),
	.w3(32'h3c269550),
	.w4(32'h3c3b2030),
	.w5(32'hbb55392d),
	.w6(32'h3c8d1bbf),
	.w7(32'hbc857f90),
	.w8(32'hbbd5c2fa),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81d780),
	.w1(32'h395450af),
	.w2(32'hbb4e3183),
	.w3(32'h3b898a1c),
	.w4(32'hbae540d9),
	.w5(32'hba5d61bf),
	.w6(32'h3bc8e27b),
	.w7(32'h3ab2bccf),
	.w8(32'h3b668fe9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd2063),
	.w1(32'h3cf6a4d8),
	.w2(32'h39d07a0f),
	.w3(32'h3d02801a),
	.w4(32'h3cacaf9f),
	.w5(32'hbcd1674f),
	.w6(32'h3cd1b9f3),
	.w7(32'h3c0bbf16),
	.w8(32'hbc4b53ad),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule