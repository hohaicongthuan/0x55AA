module layer_10_featuremap_22(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de1a6),
	.w1(32'hbc3dc025),
	.w2(32'h3b7bf407),
	.w3(32'hbcd04ae4),
	.w4(32'hbc4971a6),
	.w5(32'h3c0871d4),
	.w6(32'hbcf103bb),
	.w7(32'h3c8193e8),
	.w8(32'hbb64b374),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc722e5b),
	.w1(32'h3ae8a279),
	.w2(32'hbbae476a),
	.w3(32'hbc4c1cca),
	.w4(32'h3afe19e8),
	.w5(32'hbc3e8980),
	.w6(32'hbc0ba63d),
	.w7(32'hb8f5fa83),
	.w8(32'hba0611fd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61aad6),
	.w1(32'h384d6569),
	.w2(32'hbc0b703c),
	.w3(32'hbbb3ff1a),
	.w4(32'h3afdb3bd),
	.w5(32'hbafdfc2a),
	.w6(32'hbb0f5b86),
	.w7(32'hbc0f1c8c),
	.w8(32'h3a4a3574),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4268a0),
	.w1(32'hbb2bcbbe),
	.w2(32'h3bc5b4b0),
	.w3(32'hba9055db),
	.w4(32'hba1df537),
	.w5(32'hbc8dff22),
	.w6(32'hbb96a0ed),
	.w7(32'h3bbe52b6),
	.w8(32'hbbd30e6a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f333),
	.w1(32'h3a76ddfa),
	.w2(32'hbbbc0e2c),
	.w3(32'hbab9e3c9),
	.w4(32'h3c4aa797),
	.w5(32'h3b6236a0),
	.w6(32'h3c8a285c),
	.w7(32'hbb98c93d),
	.w8(32'hbc87a359),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f04b),
	.w1(32'hbc809b4d),
	.w2(32'h3afba134),
	.w3(32'hbc9940b3),
	.w4(32'hbc62b5ed),
	.w5(32'hb94f7f1f),
	.w6(32'hbcb55cf5),
	.w7(32'hbc0e7585),
	.w8(32'hbb24cfd0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1884a),
	.w1(32'hbbb98875),
	.w2(32'hbc0a8964),
	.w3(32'h3b1af2e0),
	.w4(32'hbc0c89e0),
	.w5(32'hbc09ee75),
	.w6(32'h39707928),
	.w7(32'hbc055870),
	.w8(32'hbbceca1f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ef51),
	.w1(32'h3c2d32ee),
	.w2(32'h3badbbd6),
	.w3(32'hbb430ece),
	.w4(32'h3cb1cc52),
	.w5(32'hbb2379c3),
	.w6(32'h3a19e05a),
	.w7(32'hb98d434b),
	.w8(32'hbc2f0cd5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77df66),
	.w1(32'hbc4dfced),
	.w2(32'h3badaba9),
	.w3(32'hbc4dcac3),
	.w4(32'hbbb61e40),
	.w5(32'h3b4bc4f9),
	.w6(32'hbbd9da8d),
	.w7(32'h3b6bcf17),
	.w8(32'h3bf25e16),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02b387),
	.w1(32'h3b23c9d2),
	.w2(32'hbc276043),
	.w3(32'h3c397116),
	.w4(32'h3c40eb81),
	.w5(32'hbbcf6ef0),
	.w6(32'h3c5cd0b9),
	.w7(32'h3bfa4e10),
	.w8(32'hbbad07ef),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90a313),
	.w1(32'h3b8078a2),
	.w2(32'hba2a33e8),
	.w3(32'h3a8b7603),
	.w4(32'h3b1f8cc9),
	.w5(32'h3c37f3ca),
	.w6(32'h3b4ea26c),
	.w7(32'h3afceadf),
	.w8(32'h3c5934a8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd58538),
	.w1(32'h3c3bc663),
	.w2(32'hbb8a2513),
	.w3(32'h3ca7daea),
	.w4(32'hba133a8f),
	.w5(32'hbaff6842),
	.w6(32'hba7372ae),
	.w7(32'hba19775b),
	.w8(32'hbadb7228),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1f99d),
	.w1(32'hbb9912f3),
	.w2(32'hbc0c605c),
	.w3(32'h3b12e246),
	.w4(32'hbba7b78d),
	.w5(32'hbae45583),
	.w6(32'hba769b4f),
	.w7(32'hbb64eee0),
	.w8(32'hbae9a990),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3d8eb),
	.w1(32'h3c0d6811),
	.w2(32'hbc40ff5e),
	.w3(32'h3b94469d),
	.w4(32'h39d502a0),
	.w5(32'hbc277e7a),
	.w6(32'h3c27539a),
	.w7(32'h3ba739a2),
	.w8(32'hbc3f6e3a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc530dd5),
	.w1(32'hbc41fd38),
	.w2(32'h3bfb57f9),
	.w3(32'hbce2fde4),
	.w4(32'hbc399c39),
	.w5(32'h3bed41d4),
	.w6(32'hbb0e6a50),
	.w7(32'h3b8e48ee),
	.w8(32'h3c2c53f5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b5564),
	.w1(32'hbbcdfe94),
	.w2(32'hbc90f14e),
	.w3(32'h3b0358a8),
	.w4(32'h3b5e0284),
	.w5(32'hbc231a13),
	.w6(32'hba814fd0),
	.w7(32'h3bbb0c0b),
	.w8(32'hbc246a81),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9b789),
	.w1(32'h3b76d81c),
	.w2(32'hbc495410),
	.w3(32'h3b3ade59),
	.w4(32'h3b85236a),
	.w5(32'hbc10aedc),
	.w6(32'h3bca61da),
	.w7(32'h3bbe428a),
	.w8(32'h3b8fae93),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3614e1),
	.w1(32'h3b8917f3),
	.w2(32'hbbdab69c),
	.w3(32'h3c011754),
	.w4(32'h38932399),
	.w5(32'hbc008272),
	.w6(32'hb910a482),
	.w7(32'hbc491bb7),
	.w8(32'hbc68dcfa),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35f4d4),
	.w1(32'h3b99cf72),
	.w2(32'h3bb51a6e),
	.w3(32'h3c0f1134),
	.w4(32'h3bccb339),
	.w5(32'hbb764777),
	.w6(32'h3bd4f840),
	.w7(32'h3a514fad),
	.w8(32'hbc51a87a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba653ec),
	.w1(32'h3bedfb1d),
	.w2(32'hbbc8827a),
	.w3(32'hbaf4c011),
	.w4(32'hbbbafe4d),
	.w5(32'h3aa597dc),
	.w6(32'hba82ea16),
	.w7(32'h3b3723b3),
	.w8(32'h3be84ea2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125225),
	.w1(32'h3bbb73db),
	.w2(32'hbbf7b73c),
	.w3(32'h3c41d968),
	.w4(32'h3afaf5c2),
	.w5(32'hba89d85a),
	.w6(32'h3b1c0062),
	.w7(32'hbbffccc5),
	.w8(32'h3a5192f6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea7c2),
	.w1(32'h3a898286),
	.w2(32'h3bce2913),
	.w3(32'h39b4e876),
	.w4(32'hbc0967f7),
	.w5(32'h3baa40bc),
	.w6(32'hbaee8843),
	.w7(32'h3b8e9346),
	.w8(32'h3b232b0d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86aa9d),
	.w1(32'hbbfdc551),
	.w2(32'hbcbd2d42),
	.w3(32'h3b4f5043),
	.w4(32'hbbc3eb88),
	.w5(32'hbc86d172),
	.w6(32'hbaa6675b),
	.w7(32'hbb091d36),
	.w8(32'hbc989169),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc187),
	.w1(32'hbb8c8246),
	.w2(32'hba6003e2),
	.w3(32'hbc0bd9d9),
	.w4(32'hbb9846b3),
	.w5(32'hb92f2e23),
	.w6(32'hbb5f327c),
	.w7(32'h3b8b1b71),
	.w8(32'h3af3f879),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b15e6),
	.w1(32'h3c0f9f84),
	.w2(32'h3ca7f955),
	.w3(32'hbb4c7411),
	.w4(32'h3c12b79b),
	.w5(32'h3d001ca2),
	.w6(32'h3b0b109d),
	.w7(32'h3c3f2585),
	.w8(32'h3c230f95),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c828559),
	.w1(32'hbb933895),
	.w2(32'hbb266c83),
	.w3(32'hbc39668b),
	.w4(32'hbc427a4e),
	.w5(32'h3ba74beb),
	.w6(32'hbc163bef),
	.w7(32'h3bc12ebe),
	.w8(32'hbb8e6bde),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a21c),
	.w1(32'h3bb00e7e),
	.w2(32'h3959cdb0),
	.w3(32'h3b1a7d10),
	.w4(32'hbb82b1c6),
	.w5(32'h3b481017),
	.w6(32'hba957c28),
	.w7(32'hbbc5809e),
	.w8(32'h3a58bfe8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dfb99),
	.w1(32'hb99678e8),
	.w2(32'h3c1e34db),
	.w3(32'h3bc91c28),
	.w4(32'h3b48fe3c),
	.w5(32'h3c1b167c),
	.w6(32'h3b28dd04),
	.w7(32'hb87a721a),
	.w8(32'h3b56a8a6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dcb41),
	.w1(32'hbbe57cd9),
	.w2(32'h3b4d5f07),
	.w3(32'hbcad6132),
	.w4(32'hbcde4bae),
	.w5(32'hbc23cb1f),
	.w6(32'hbcb75902),
	.w7(32'hbc83a0ba),
	.w8(32'hbb87eb41),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819a81),
	.w1(32'h3c9dc47f),
	.w2(32'h3b6f5260),
	.w3(32'hbbce6332),
	.w4(32'h3a6b0b98),
	.w5(32'hb9d1c7ae),
	.w6(32'hbc96b562),
	.w7(32'h3b529e3c),
	.w8(32'h3b4054f5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5073),
	.w1(32'hba2c4753),
	.w2(32'hbbdcf082),
	.w3(32'hba8c266e),
	.w4(32'h3aa1eead),
	.w5(32'hbb70dd5f),
	.w6(32'hb9b6f073),
	.w7(32'h3ad60013),
	.w8(32'hbbc6d158),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf39dfe),
	.w1(32'hbb371849),
	.w2(32'hbc028168),
	.w3(32'hb9f291a7),
	.w4(32'hbb2663f1),
	.w5(32'hbc33cdf7),
	.w6(32'hbbfa4a5d),
	.w7(32'hbc3da928),
	.w8(32'hbb2fad89),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc541256),
	.w1(32'hbbc70ce4),
	.w2(32'hbaabb8e9),
	.w3(32'hbb9ac099),
	.w4(32'hbaf65120),
	.w5(32'hbb4d9b49),
	.w6(32'h39673401),
	.w7(32'hbaf1065c),
	.w8(32'hbb17ae4b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac816),
	.w1(32'hbb178387),
	.w2(32'hbb4142c6),
	.w3(32'hbc2fe7ec),
	.w4(32'hbbfc8337),
	.w5(32'hbc8529d4),
	.w6(32'hbbaa21e0),
	.w7(32'hbb85bab5),
	.w8(32'hbc0f88b2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109298),
	.w1(32'h3c08db25),
	.w2(32'h3a3a8c68),
	.w3(32'h3bfb0e17),
	.w4(32'h3c917dc2),
	.w5(32'h3b71b0c9),
	.w6(32'h3c1159df),
	.w7(32'h3c1cd43b),
	.w8(32'h3b37e256),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbbf4f),
	.w1(32'h3add47cb),
	.w2(32'h3bf753c1),
	.w3(32'h3bebdcd6),
	.w4(32'h38ae9e7c),
	.w5(32'hbb1dd14b),
	.w6(32'h3bea04c1),
	.w7(32'hbb454a35),
	.w8(32'hbc0331f3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5c414),
	.w1(32'h3bd21e9a),
	.w2(32'hbca91dd9),
	.w3(32'h3b9a6431),
	.w4(32'h3bab5308),
	.w5(32'hbcaed875),
	.w6(32'hbc8a41aa),
	.w7(32'hbc3d93cd),
	.w8(32'hbca05073),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a5e2f),
	.w1(32'h3c37b3dd),
	.w2(32'h3c9e6bcb),
	.w3(32'hbd057579),
	.w4(32'hbaba4c48),
	.w5(32'h3bdce3c2),
	.w6(32'hbc981129),
	.w7(32'h3c6195a2),
	.w8(32'h3c80c181),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65f3e3),
	.w1(32'h3c90b59c),
	.w2(32'h3cd10484),
	.w3(32'hbc18e0b2),
	.w4(32'h3ba4740c),
	.w5(32'h3d02b3df),
	.w6(32'hbc9cab64),
	.w7(32'h3c260f4b),
	.w8(32'h3d100bdc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68e56c),
	.w1(32'hbc8ae049),
	.w2(32'h3adcca34),
	.w3(32'hbc21e29e),
	.w4(32'hbc89b167),
	.w5(32'h39d3c4b0),
	.w6(32'h3ba8d2d0),
	.w7(32'hbbcc5cc3),
	.w8(32'h3996f2f0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1578),
	.w1(32'h3bdf47f0),
	.w2(32'h3b5a5ccf),
	.w3(32'h3c531bd8),
	.w4(32'h3c0bfe48),
	.w5(32'h3b95f1e4),
	.w6(32'h3b830614),
	.w7(32'h3c17e23b),
	.w8(32'hbc1d9cf3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a9625),
	.w1(32'h3c576532),
	.w2(32'hba661af5),
	.w3(32'h3c1db8e3),
	.w4(32'h3c2ab016),
	.w5(32'h3bc5500c),
	.w6(32'hbc297c27),
	.w7(32'hbb0fb39e),
	.w8(32'hba368df4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd81414),
	.w1(32'h3b1150ff),
	.w2(32'hbb60daf0),
	.w3(32'h3be6787d),
	.w4(32'h3c8b053e),
	.w5(32'hbb61131e),
	.w6(32'h3a1380f3),
	.w7(32'h3ae047e3),
	.w8(32'hbbd1aedc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c231324),
	.w1(32'hb9d7a138),
	.w2(32'hbca9ade9),
	.w3(32'h3b7d0c34),
	.w4(32'h3baca3c8),
	.w5(32'hbcc41659),
	.w6(32'h3a87acd1),
	.w7(32'hba521a64),
	.w8(32'hbcdc40dd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0326f),
	.w1(32'h3a896178),
	.w2(32'hbc780cc9),
	.w3(32'hbbf6dd4c),
	.w4(32'h3bc7f4f7),
	.w5(32'hbc9a2908),
	.w6(32'hbac9757e),
	.w7(32'h3bbd965d),
	.w8(32'hbc94d7df),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b97c7),
	.w1(32'hbaa88960),
	.w2(32'hbbe14334),
	.w3(32'hbc62cd99),
	.w4(32'hbc9eb7ef),
	.w5(32'hbaaa0438),
	.w6(32'hbcd5cd46),
	.w7(32'hbca6f433),
	.w8(32'hbbe2c24d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f9954),
	.w1(32'hbc37bc05),
	.w2(32'hbc6cf4c2),
	.w3(32'hb91a46d1),
	.w4(32'hbb966413),
	.w5(32'hbc7c2f47),
	.w6(32'hbbb822e0),
	.w7(32'hba1b6502),
	.w8(32'hbc7ed3b0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91d514),
	.w1(32'hbba2c952),
	.w2(32'hbc9ed218),
	.w3(32'h3cfa5499),
	.w4(32'h3c305f19),
	.w5(32'hbc3b6f9c),
	.w6(32'h3c221ba9),
	.w7(32'hbb9e9c55),
	.w8(32'hbcaccc07),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40d27a),
	.w1(32'hbbd1f263),
	.w2(32'h3c2368f4),
	.w3(32'h37a5f0b2),
	.w4(32'hbb332d85),
	.w5(32'h3c028fd1),
	.w6(32'hbb26d9b3),
	.w7(32'hbb878989),
	.w8(32'h3c31768c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bd374),
	.w1(32'h3b8ffea4),
	.w2(32'h3a71508a),
	.w3(32'h3b015ad1),
	.w4(32'h3af0ba1b),
	.w5(32'h3be48a33),
	.w6(32'h3b1e0869),
	.w7(32'hbb415548),
	.w8(32'h3b7151b6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3260b8),
	.w1(32'h3be262fa),
	.w2(32'hbaf08d84),
	.w3(32'h3c9bc121),
	.w4(32'h3c6a3f97),
	.w5(32'h3c8bed83),
	.w6(32'h3c62831d),
	.w7(32'h3c1f99fc),
	.w8(32'h3c502c39),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c376d89),
	.w1(32'h3c4a800c),
	.w2(32'hbbc3c321),
	.w3(32'h3cf28fd0),
	.w4(32'h3bb9d044),
	.w5(32'hbbcfb0ef),
	.w6(32'h3bd6465f),
	.w7(32'hbbbe8254),
	.w8(32'hbab00e47),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9e032),
	.w1(32'h3b694922),
	.w2(32'hbc7ea5e9),
	.w3(32'h3b786b72),
	.w4(32'h3b827bca),
	.w5(32'hbc8d4e14),
	.w6(32'h3addd1a4),
	.w7(32'h3c02031b),
	.w8(32'hbc71a502),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1ff65),
	.w1(32'hbaa8438d),
	.w2(32'hb9f35bd4),
	.w3(32'hbbcc4fae),
	.w4(32'hbbdd46bc),
	.w5(32'hbc8ed5e5),
	.w6(32'hbc6e55a5),
	.w7(32'hbcb14a3b),
	.w8(32'hbcee3242),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cdbef),
	.w1(32'h3b8c76b3),
	.w2(32'hbbf14d48),
	.w3(32'hbc2858b4),
	.w4(32'hbc2c24f5),
	.w5(32'hbc4c61f6),
	.w6(32'hbc323640),
	.w7(32'hbab500a6),
	.w8(32'hbc5758b5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2085f8),
	.w1(32'hbbf787e5),
	.w2(32'h3a110e01),
	.w3(32'hbc0fe170),
	.w4(32'hbb3d27b6),
	.w5(32'h3be5b625),
	.w6(32'hbb853fe7),
	.w7(32'h3b35d7b6),
	.w8(32'hba57dc25),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba993601),
	.w1(32'hbb1b3d88),
	.w2(32'hbb9aca99),
	.w3(32'hbbe10a99),
	.w4(32'hbb7867f5),
	.w5(32'hbb4b3ae6),
	.w6(32'hbb6500e5),
	.w7(32'hbb4fb59b),
	.w8(32'hbb0b4853),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828713),
	.w1(32'h3a2b325d),
	.w2(32'h3b05614b),
	.w3(32'hba87ab0a),
	.w4(32'h3b6d8f3b),
	.w5(32'h3b88e3d1),
	.w6(32'hbb8e9ad9),
	.w7(32'h3c098910),
	.w8(32'h3bb5ac7e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ce228),
	.w1(32'h3c838ea4),
	.w2(32'h3b52b86f),
	.w3(32'hba0752c9),
	.w4(32'h3c6aeb42),
	.w5(32'h3bda2e55),
	.w6(32'h3b210787),
	.w7(32'h3c73a4a5),
	.w8(32'h398e6b23),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ece04),
	.w1(32'hbc0a8923),
	.w2(32'h3a86f6ab),
	.w3(32'hbbcba6df),
	.w4(32'hbc0c3106),
	.w5(32'h39ffd331),
	.w6(32'hbc6bc3ae),
	.w7(32'hbc16008d),
	.w8(32'h3b50e1ad),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46bf07),
	.w1(32'h3b196501),
	.w2(32'hbc3a8053),
	.w3(32'h3c347127),
	.w4(32'h3c519bda),
	.w5(32'hba8342a9),
	.w6(32'h3b27dab9),
	.w7(32'h3b91507d),
	.w8(32'h39b4cb15),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4714e8),
	.w1(32'hbba8fdfb),
	.w2(32'hbcaafd40),
	.w3(32'h3c098261),
	.w4(32'h3b54bd47),
	.w5(32'hbc71c4ad),
	.w6(32'h3ba14eeb),
	.w7(32'hbb6b2239),
	.w8(32'hbc88e487),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5049),
	.w1(32'hbb2b2ddf),
	.w2(32'hbc0a2835),
	.w3(32'hbbe5db52),
	.w4(32'hbbbfbec3),
	.w5(32'hbbc49164),
	.w6(32'hbbdec431),
	.w7(32'hbbd15f26),
	.w8(32'hbc613a77),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d782a),
	.w1(32'hbc2e4fcd),
	.w2(32'hbb2b8d5e),
	.w3(32'hbc94d725),
	.w4(32'hbc595015),
	.w5(32'h3a87f8c5),
	.w6(32'hbce99fe2),
	.w7(32'hbcaa4fbd),
	.w8(32'h3b160f3a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491c6c),
	.w1(32'hbbbc06ff),
	.w2(32'hbc08d19b),
	.w3(32'hbaa9ace5),
	.w4(32'h3bc8a8ae),
	.w5(32'hbb7e261e),
	.w6(32'h3ac5454f),
	.w7(32'h3be9c396),
	.w8(32'hb9472689),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c254f),
	.w1(32'hbc5f267f),
	.w2(32'hbc2538b2),
	.w3(32'hbc6dc84a),
	.w4(32'hbc8730dc),
	.w5(32'hbc9ba6bc),
	.w6(32'hbc0cd1bd),
	.w7(32'hbc3019c9),
	.w8(32'hbc63cf8c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb4a9),
	.w1(32'hbc57c7b5),
	.w2(32'hbcb8a304),
	.w3(32'hbc676cf9),
	.w4(32'hbb842572),
	.w5(32'h3b130fbf),
	.w6(32'hbcd95981),
	.w7(32'hbc5b6008),
	.w8(32'hbaf59168),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0f49a),
	.w1(32'h3bebcf89),
	.w2(32'hbc7aa5b2),
	.w3(32'h3c67a6a2),
	.w4(32'h3b9a1202),
	.w5(32'hbc951bf4),
	.w6(32'h3c1f40c2),
	.w7(32'hbbd3d31d),
	.w8(32'hbcc6d032),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02cf34),
	.w1(32'hbbe32554),
	.w2(32'hbcc63fe9),
	.w3(32'hbc32bd73),
	.w4(32'hbc6fc82b),
	.w5(32'hbd095085),
	.w6(32'hbbbcfdbf),
	.w7(32'hbc8ffca2),
	.w8(32'hbd0c8ee4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf20c55),
	.w1(32'hbbd6de19),
	.w2(32'hbc14f927),
	.w3(32'hbd27b511),
	.w4(32'hbc60045e),
	.w5(32'h3a3017ed),
	.w6(32'hbd082703),
	.w7(32'hbbe66362),
	.w8(32'h3bb9cc50),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f3f8d),
	.w1(32'hbc439809),
	.w2(32'hbc161ce9),
	.w3(32'hbc39c4a7),
	.w4(32'hbba485ed),
	.w5(32'hbb254786),
	.w6(32'hbbcec176),
	.w7(32'hbc1011c5),
	.w8(32'hbb309768),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcd6e8),
	.w1(32'hbb686237),
	.w2(32'hbc1863c9),
	.w3(32'hbc29731a),
	.w4(32'hbc4a86ba),
	.w5(32'hba434bf9),
	.w6(32'hbbc3caac),
	.w7(32'hbc4db6b5),
	.w8(32'hbb94b302),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cad9a),
	.w1(32'h3b965b1d),
	.w2(32'h3a91d070),
	.w3(32'h3ca7f358),
	.w4(32'h3bbdb529),
	.w5(32'hba028476),
	.w6(32'h3bf452d7),
	.w7(32'h3c1f52f8),
	.w8(32'hbb5c6e30),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c408356),
	.w1(32'h3b7a1223),
	.w2(32'hbc0cf3a0),
	.w3(32'h3c08df8c),
	.w4(32'h3bec58f3),
	.w5(32'hbbd4a13b),
	.w6(32'h3c041d94),
	.w7(32'h3a2d9f3d),
	.w8(32'hbc0f965d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499085),
	.w1(32'hbbb066d1),
	.w2(32'h3b2e6867),
	.w3(32'hbb0d40b2),
	.w4(32'hbb911425),
	.w5(32'h3ce6a425),
	.w6(32'hbbbe229f),
	.w7(32'hbb9e17a2),
	.w8(32'h3c210d7e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0272fc),
	.w1(32'h3ba98968),
	.w2(32'hbc2f81c2),
	.w3(32'h3d8bdb33),
	.w4(32'h3d2464e0),
	.w5(32'hb9d9cc73),
	.w6(32'h3d34d49c),
	.w7(32'h3ca3c747),
	.w8(32'hbb3e7b38),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22adfd),
	.w1(32'h3c073d2e),
	.w2(32'hbb412446),
	.w3(32'h3cb9038a),
	.w4(32'h3caf9c35),
	.w5(32'h3b731479),
	.w6(32'h3c1478c3),
	.w7(32'h3c55f0b0),
	.w8(32'hbc1099db),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991f9dd),
	.w1(32'h3c47a42e),
	.w2(32'hbb932e30),
	.w3(32'h3c77cd7b),
	.w4(32'h3ccaa01b),
	.w5(32'hbbebaaef),
	.w6(32'h3c6b036d),
	.w7(32'h3ca33128),
	.w8(32'hba3da1cb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad65227),
	.w1(32'h3bb50e48),
	.w2(32'hbbb64513),
	.w3(32'h3bd9037c),
	.w4(32'h3be9d474),
	.w5(32'hbba33a5d),
	.w6(32'hbc186f7c),
	.w7(32'hbafb3a3d),
	.w8(32'hbbc173a5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecb22d),
	.w1(32'h3b493b10),
	.w2(32'hbc80e4e3),
	.w3(32'h3b01737e),
	.w4(32'h3bcb9760),
	.w5(32'hbc28261f),
	.w6(32'hba2159e0),
	.w7(32'h3a2a849f),
	.w8(32'hbbcdd513),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064043),
	.w1(32'hbb85d352),
	.w2(32'hbba64e30),
	.w3(32'hbb19f010),
	.w4(32'hb9f743d7),
	.w5(32'hbb1a2ba6),
	.w6(32'hbb3792c7),
	.w7(32'hbb521e18),
	.w8(32'h39ca0989),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ace5),
	.w1(32'h3c104bba),
	.w2(32'hbb8d92c8),
	.w3(32'h3a9ec9ac),
	.w4(32'h3bfcda37),
	.w5(32'h3c120cf6),
	.w6(32'h3b87535e),
	.w7(32'h3be1d74e),
	.w8(32'h3ab005d9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd08b),
	.w1(32'hbb9b17dc),
	.w2(32'hbc1debab),
	.w3(32'hba7276d5),
	.w4(32'hbc607409),
	.w5(32'hbc7dcda9),
	.w6(32'h3ab0551e),
	.w7(32'hbb3138b4),
	.w8(32'hbc2a6f69),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb352626),
	.w1(32'h3ad78949),
	.w2(32'h3afb83b6),
	.w3(32'hba4a1414),
	.w4(32'h3b89b7da),
	.w5(32'h3bd1f951),
	.w6(32'hbc32c89e),
	.w7(32'hbbbd0960),
	.w8(32'h3b9466f7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d0241),
	.w1(32'hbbd1cbb8),
	.w2(32'hba7d880f),
	.w3(32'h3b9583a3),
	.w4(32'h3aa19474),
	.w5(32'h3c1ce8e8),
	.w6(32'h3c1d5cb8),
	.w7(32'h3b53c730),
	.w8(32'hbc036844),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd31bb8),
	.w1(32'h3acb7476),
	.w2(32'hbab47d47),
	.w3(32'h3c6b944f),
	.w4(32'hbb47aa73),
	.w5(32'hbb812d06),
	.w6(32'h3b27c7a3),
	.w7(32'hbb069238),
	.w8(32'hbb518e21),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24dec8),
	.w1(32'hba7866df),
	.w2(32'h3ac415b1),
	.w3(32'hbc923394),
	.w4(32'hbc07a5d1),
	.w5(32'h3bbdc051),
	.w6(32'hbc55643a),
	.w7(32'hbb7b4117),
	.w8(32'h3b9bd003),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7ba5),
	.w1(32'h3c3b652f),
	.w2(32'h3b4713c5),
	.w3(32'h3c59d94c),
	.w4(32'h3c4f12c5),
	.w5(32'h3b1f29e5),
	.w6(32'h3bef50b4),
	.w7(32'h3c438150),
	.w8(32'h3bd6f051),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f1042),
	.w1(32'h3bf93a46),
	.w2(32'hbbb564ed),
	.w3(32'h3c0d33f4),
	.w4(32'h3aece6fe),
	.w5(32'hbb577c9b),
	.w6(32'h3b57d82e),
	.w7(32'hba183d10),
	.w8(32'hbc465bdd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda5b14),
	.w1(32'h3860823b),
	.w2(32'hbc93e763),
	.w3(32'h3bbfda9e),
	.w4(32'h3aeb1451),
	.w5(32'hbc39c3d9),
	.w6(32'h3bb74aa9),
	.w7(32'hbb27fdb7),
	.w8(32'h39d524f7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd08ab92),
	.w1(32'hbbf1bf15),
	.w2(32'hba161957),
	.w3(32'hbc9b4229),
	.w4(32'hbb9b3f56),
	.w5(32'hbc9d5c88),
	.w6(32'h3c5c54b9),
	.w7(32'h3c4e27d2),
	.w8(32'h3b9349ff),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce69819),
	.w1(32'hbc74c702),
	.w2(32'hbb6a8709),
	.w3(32'hbd66c934),
	.w4(32'hbd12131e),
	.w5(32'h3c213d19),
	.w6(32'hbd221a2e),
	.w7(32'hbc7c4d07),
	.w8(32'h3bc06457),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c304c0b),
	.w1(32'h3ca14568),
	.w2(32'h3be5d302),
	.w3(32'h3c6f7876),
	.w4(32'h3ccb7b95),
	.w5(32'h3ba09752),
	.w6(32'h3c422200),
	.w7(32'h3ca8061c),
	.w8(32'h3be9e4a3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c031ba6),
	.w1(32'h3b49a8ec),
	.w2(32'hbca5c031),
	.w3(32'h3b958a00),
	.w4(32'h3c0694dd),
	.w5(32'hbc38ade8),
	.w6(32'hba1d8d08),
	.w7(32'h3bb0f9f4),
	.w8(32'hbc5cfdc5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3313b8),
	.w1(32'hbbcd2751),
	.w2(32'hbbaa3c00),
	.w3(32'hba5b7f47),
	.w4(32'hba4c0167),
	.w5(32'hbb12d349),
	.w6(32'hbb6d1f0a),
	.w7(32'hbbe6e2c3),
	.w8(32'h3b97f767),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0018a),
	.w1(32'h3c28831b),
	.w2(32'h3c8db3c8),
	.w3(32'hbb834596),
	.w4(32'h3c447f00),
	.w5(32'h3cbc96d7),
	.w6(32'h3b670b2f),
	.w7(32'h3c05832f),
	.w8(32'h3ca61cce),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17e374),
	.w1(32'h3c0fa669),
	.w2(32'hb850bb5c),
	.w3(32'h3d0045be),
	.w4(32'h3c24eef5),
	.w5(32'h3bb977bd),
	.w6(32'h3bf81868),
	.w7(32'hbb96ccf6),
	.w8(32'h3c1643bc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69e19f),
	.w1(32'h3b0a8d83),
	.w2(32'hbc4b75f3),
	.w3(32'h3cb42c9f),
	.w4(32'h3c8aade3),
	.w5(32'hbca11555),
	.w6(32'h3c9e8302),
	.w7(32'h3bb2880a),
	.w8(32'hbcb9ef53),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed1ad),
	.w1(32'hbc4f4547),
	.w2(32'hbd09854d),
	.w3(32'hbb3aebb0),
	.w4(32'hbc19d369),
	.w5(32'hbd1bdbfe),
	.w6(32'hbc259355),
	.w7(32'hba5cf3db),
	.w8(32'hbcf0742e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bd9ce),
	.w1(32'h3ca03edb),
	.w2(32'hbb445d07),
	.w3(32'hbce686ac),
	.w4(32'h3bfe170b),
	.w5(32'h3a2b63ed),
	.w6(32'hbc68686c),
	.w7(32'hba7c5daf),
	.w8(32'hbc7a6b07),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a58d),
	.w1(32'h3c6495ed),
	.w2(32'h3ce29894),
	.w3(32'h3b9ce76b),
	.w4(32'h3c8e6957),
	.w5(32'h3d07bb3c),
	.w6(32'h3c053638),
	.w7(32'h3cd3ed0f),
	.w8(32'h3d18cb67),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d6add),
	.w1(32'h3c31225e),
	.w2(32'h3ad933f6),
	.w3(32'h3c3357e2),
	.w4(32'h3c596ba3),
	.w5(32'hbc2f5675),
	.w6(32'h3c4e7661),
	.w7(32'h3c71351d),
	.w8(32'hbc2dbed9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80003a),
	.w1(32'hbc3ac168),
	.w2(32'hbd0a7a1b),
	.w3(32'hbae21787),
	.w4(32'hbb8e96ea),
	.w5(32'hbcc8a717),
	.w6(32'hbc1d2931),
	.w7(32'hbc077e3e),
	.w8(32'hbcfad54f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f0a39),
	.w1(32'hbc6a5d97),
	.w2(32'hbc3c2a56),
	.w3(32'hbc469815),
	.w4(32'hbbde90ef),
	.w5(32'hbbcea371),
	.w6(32'hbc340aa9),
	.w7(32'hbb538f3e),
	.w8(32'hbc763184),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb308db),
	.w1(32'hbba10fba),
	.w2(32'hbc7c532e),
	.w3(32'hbcad9862),
	.w4(32'hbb9c2c40),
	.w5(32'hbc0a005f),
	.w6(32'hbc89ba40),
	.w7(32'h38d2286a),
	.w8(32'hbc84b7ad),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f315),
	.w1(32'hb9c9bbb3),
	.w2(32'hbb53b68f),
	.w3(32'hbb6d1c7a),
	.w4(32'hbbbae5be),
	.w5(32'h3bb01997),
	.w6(32'h3b061e92),
	.w7(32'hba9d5e18),
	.w8(32'h3b868d85),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47a632),
	.w1(32'hbbc76bb2),
	.w2(32'hbc4a7287),
	.w3(32'h3b5cce03),
	.w4(32'hbbe8fe00),
	.w5(32'hbbd9ee49),
	.w6(32'h3b8cc65a),
	.w7(32'hbb85a985),
	.w8(32'hbb0392f7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f741),
	.w1(32'h3bfb5a2c),
	.w2(32'hbbbc266d),
	.w3(32'hbc3080d3),
	.w4(32'hbb4917e1),
	.w5(32'hbac69f2c),
	.w6(32'hbc003a77),
	.w7(32'hbc16e519),
	.w8(32'hba749438),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b931942),
	.w1(32'hbb8581e1),
	.w2(32'hbba413b8),
	.w3(32'h3bffece4),
	.w4(32'hba98ae63),
	.w5(32'hbc09fbc2),
	.w6(32'h3baac68c),
	.w7(32'hbb7b354a),
	.w8(32'hbbacf4eb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfeab),
	.w1(32'h3ab13e84),
	.w2(32'h3b7e1360),
	.w3(32'hbc0263d2),
	.w4(32'hba0eab86),
	.w5(32'h3bb472c3),
	.w6(32'hbb122c6e),
	.w7(32'hba8a1dfb),
	.w8(32'h3c2c0168),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b959),
	.w1(32'h3c1e0164),
	.w2(32'h3a9cc70b),
	.w3(32'h3c4ee0ba),
	.w4(32'h3ca55db6),
	.w5(32'h3b1dc033),
	.w6(32'h3bb1c7e4),
	.w7(32'h3ca41cfb),
	.w8(32'h3c408624),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc880195),
	.w1(32'h39d74431),
	.w2(32'hbb9a5059),
	.w3(32'hbb8d7cb5),
	.w4(32'h3c381819),
	.w5(32'hbaa3c101),
	.w6(32'hbb911d82),
	.w7(32'h3c3a530f),
	.w8(32'h3ac4c21f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26fdce),
	.w1(32'h3c53a1b7),
	.w2(32'hbb295ecb),
	.w3(32'h3ba9e9f5),
	.w4(32'h3b243a21),
	.w5(32'hbbb89f55),
	.w6(32'hbbf30dfd),
	.w7(32'hbc31d3e3),
	.w8(32'hbc34d416),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473678),
	.w1(32'hbc219105),
	.w2(32'hbc7cfffd),
	.w3(32'hbbca4d7d),
	.w4(32'hbb571015),
	.w5(32'hbc681f83),
	.w6(32'hbc862805),
	.w7(32'hbb7eaba5),
	.w8(32'hbc4d5192),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a20a8),
	.w1(32'hbc16338c),
	.w2(32'hbb189387),
	.w3(32'hbca0b8f3),
	.w4(32'hbc3f6b78),
	.w5(32'hbbe7ccfb),
	.w6(32'hbc2bdd99),
	.w7(32'h3aae1596),
	.w8(32'hbc49c420),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e9e9d),
	.w1(32'h3bdcf2c2),
	.w2(32'hbbe05a7f),
	.w3(32'hbc053cad),
	.w4(32'hbb09b800),
	.w5(32'hbb86ea75),
	.w6(32'hbc72b4cd),
	.w7(32'hbbc92dee),
	.w8(32'hbbd2f899),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe83d5),
	.w1(32'hba9d55bc),
	.w2(32'h39ca5dfb),
	.w3(32'hbbbd9b61),
	.w4(32'hbc5101a5),
	.w5(32'hbb324c4c),
	.w6(32'hbc3afb7c),
	.w7(32'hbc856c34),
	.w8(32'hbc28efe6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2d74f),
	.w1(32'h3a0d1ebb),
	.w2(32'hbb8160b1),
	.w3(32'hbb139539),
	.w4(32'hbb36d130),
	.w5(32'hbc190fd6),
	.w6(32'hbc644b8f),
	.w7(32'hbc1cc84a),
	.w8(32'hbbe39fe1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5a599),
	.w1(32'hbb4c9b2c),
	.w2(32'h3bde605d),
	.w3(32'hbb7b8488),
	.w4(32'hbba1fe1c),
	.w5(32'h3c05b6b8),
	.w6(32'hbbf1cc00),
	.w7(32'hbca0d5af),
	.w8(32'h3ab78b34),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd883e0),
	.w1(32'h3bb96889),
	.w2(32'h3b92ec8b),
	.w3(32'h3bec3348),
	.w4(32'h3c2e5159),
	.w5(32'hbafd8913),
	.w6(32'h3c1a2edf),
	.w7(32'h3bb9f2ae),
	.w8(32'hbb88a5b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddc646),
	.w1(32'hbb7bce48),
	.w2(32'h39644814),
	.w3(32'hbbcdb377),
	.w4(32'hba2353f6),
	.w5(32'hbb2952d2),
	.w6(32'hbb25528d),
	.w7(32'hbb7be304),
	.w8(32'hba81f958),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9149fd),
	.w1(32'h3b03518e),
	.w2(32'h3805cbb8),
	.w3(32'h3b23b909),
	.w4(32'hba35752f),
	.w5(32'h3c0c74d1),
	.w6(32'h3a515248),
	.w7(32'hba818b3e),
	.w8(32'h3bc18445),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d6fd7),
	.w1(32'h3c5de149),
	.w2(32'h3c3a8a16),
	.w3(32'h3c8f56f4),
	.w4(32'h3cb99bb2),
	.w5(32'h3c0671b5),
	.w6(32'h3c75d02a),
	.w7(32'h3ca7197e),
	.w8(32'h3b89576b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b609d16),
	.w1(32'h3bd44b20),
	.w2(32'h3c009a46),
	.w3(32'h3bb4098b),
	.w4(32'h3c1bf2ee),
	.w5(32'h3a75ac3a),
	.w6(32'hbb620ed6),
	.w7(32'hbb29f2c8),
	.w8(32'hbbd77dbe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f6c57),
	.w1(32'hbc2a63da),
	.w2(32'h3a92b889),
	.w3(32'hbc0a9490),
	.w4(32'hbc866cbc),
	.w5(32'h3bc1b16f),
	.w6(32'hbc6bd500),
	.w7(32'hbc9765d1),
	.w8(32'h3ba7923d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef6406),
	.w1(32'hbc39cf83),
	.w2(32'hb9d705b0),
	.w3(32'h3aba3acc),
	.w4(32'hbc0f60b2),
	.w5(32'h3c0e8e66),
	.w6(32'hbbebbba4),
	.w7(32'hbc901b1e),
	.w8(32'hba26024a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828bca),
	.w1(32'hbc4d0967),
	.w2(32'h3bb93a08),
	.w3(32'h3c2b2f2d),
	.w4(32'hbb2a35a0),
	.w5(32'h3c54abc0),
	.w6(32'h3bf8ad69),
	.w7(32'h3a2e8323),
	.w8(32'h3be2d7c5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfdb9bc),
	.w1(32'h3bd48ccc),
	.w2(32'hbc19facc),
	.w3(32'h3cec7354),
	.w4(32'h3bafb34b),
	.w5(32'hbc354d6e),
	.w6(32'h3c7d53a0),
	.w7(32'hbbf422ed),
	.w8(32'hbc7fd826),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3e3f0),
	.w1(32'hbc19fef6),
	.w2(32'hbc32d05a),
	.w3(32'h3cd6fde0),
	.w4(32'h3b9ba8f8),
	.w5(32'hbb265510),
	.w6(32'h3b459cb3),
	.w7(32'hbc0d1ae0),
	.w8(32'hbc317de3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50e6fa),
	.w1(32'hbb73af2e),
	.w2(32'hbab82331),
	.w3(32'hbc48c83f),
	.w4(32'hbc22e123),
	.w5(32'hbca0c1b1),
	.w6(32'hbc3b96f4),
	.w7(32'hbc308f64),
	.w8(32'hbc3fa149),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d3210),
	.w1(32'h3b946b17),
	.w2(32'hbaea22d8),
	.w3(32'hbce71981),
	.w4(32'hbacbba27),
	.w5(32'hbb50b89b),
	.w6(32'hbc3b4dc1),
	.w7(32'hbba684ce),
	.w8(32'hb9c62598),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39885f1b),
	.w1(32'h3b0817e4),
	.w2(32'h39ec0732),
	.w3(32'h3bb730ce),
	.w4(32'h3ba4b18e),
	.w5(32'hbc2e84d3),
	.w6(32'h3be5ed46),
	.w7(32'h3b9580ab),
	.w8(32'hbc1d09fe),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba800fb6),
	.w1(32'hbaf06666),
	.w2(32'hbc400dec),
	.w3(32'hbc07c3fb),
	.w4(32'hbc3d067e),
	.w5(32'hbc04ef72),
	.w6(32'h3a2d4a06),
	.w7(32'hbb5194e3),
	.w8(32'hbc2b3b48),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc748e6b),
	.w1(32'hbb9be691),
	.w2(32'hbc77f55b),
	.w3(32'hbc8eab11),
	.w4(32'hbb8d483a),
	.w5(32'hbc56ef0c),
	.w6(32'hbc8b8205),
	.w7(32'hbc180fb3),
	.w8(32'hbc2ea308),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a5d0),
	.w1(32'hbbf68054),
	.w2(32'hbbf69403),
	.w3(32'h3b5871a2),
	.w4(32'hbbdb8112),
	.w5(32'hbc75f980),
	.w6(32'hbc14a3c7),
	.w7(32'hbc6155fe),
	.w8(32'hbc83038c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0d41),
	.w1(32'h3b98ffc8),
	.w2(32'hbc4c6d7a),
	.w3(32'hbc192839),
	.w4(32'hbbcdf998),
	.w5(32'hbb333827),
	.w6(32'hbc3fd047),
	.w7(32'hbbadd57c),
	.w8(32'h3b9f6f67),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02e8d6),
	.w1(32'hbb33d465),
	.w2(32'hbc88445f),
	.w3(32'hbc4c3a85),
	.w4(32'hbbfa94b0),
	.w5(32'hbcccf821),
	.w6(32'hbc10e182),
	.w7(32'hbc3f03fa),
	.w8(32'hbcb39755),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5327c7),
	.w1(32'hbc8a3d69),
	.w2(32'hbc3d411f),
	.w3(32'hbd20ba0a),
	.w4(32'hbd2e8281),
	.w5(32'hbc5155db),
	.w6(32'hbd079aa4),
	.w7(32'hbd0982a8),
	.w8(32'hbc1e6a32),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c23a9),
	.w1(32'h3aa3aa0d),
	.w2(32'h3ba16b44),
	.w3(32'hbc489847),
	.w4(32'hbb3cf1d9),
	.w5(32'h3baa6fc0),
	.w6(32'hbbbc8418),
	.w7(32'hbaad1425),
	.w8(32'h3c06fec1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac72554),
	.w1(32'hbbad92b5),
	.w2(32'hb9806002),
	.w3(32'h3ca9b8c2),
	.w4(32'h3b4c60a7),
	.w5(32'h3b9ab445),
	.w6(32'h3c08581a),
	.w7(32'h3b3e30b4),
	.w8(32'h3b8d2264),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4719a7),
	.w1(32'h3bf236c1),
	.w2(32'h3bd0136a),
	.w3(32'h3c72d650),
	.w4(32'h3c162f1d),
	.w5(32'h3c02d394),
	.w6(32'h3c33ccde),
	.w7(32'h3c19162b),
	.w8(32'h3c0a1670),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2222c7),
	.w1(32'h3ca47403),
	.w2(32'h3ca61e60),
	.w3(32'hbc3b21a8),
	.w4(32'h3bd3af9f),
	.w5(32'h3ca8c7a3),
	.w6(32'h3a899874),
	.w7(32'h3c015622),
	.w8(32'h3c975d33),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8395cd),
	.w1(32'h3c10cca7),
	.w2(32'hbc233808),
	.w3(32'h3bf9dc55),
	.w4(32'h3b89a638),
	.w5(32'hbc5d5c45),
	.w6(32'hbbefb8e1),
	.w7(32'hbc25a4f7),
	.w8(32'hbc60ffcc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dbbbb),
	.w1(32'hba12dc35),
	.w2(32'hba6795b8),
	.w3(32'hbc8ef953),
	.w4(32'hbb9c8a1c),
	.w5(32'hbadbca70),
	.w6(32'hbc79f272),
	.w7(32'hbc38dc30),
	.w8(32'h3a0a1b5a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849d22),
	.w1(32'h3abf416b),
	.w2(32'hbc6793e3),
	.w3(32'hbb492a59),
	.w4(32'hb936e9d3),
	.w5(32'hbc900cfa),
	.w6(32'h3a955227),
	.w7(32'h3b0744f8),
	.w8(32'hbc028fb3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb0286),
	.w1(32'hbc5bff66),
	.w2(32'h3b6c5e35),
	.w3(32'hbccb98e5),
	.w4(32'hbc913468),
	.w5(32'h3bff77d8),
	.w6(32'hbc4ebb83),
	.w7(32'hbb4687f9),
	.w8(32'h3bad66c4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a028f05),
	.w1(32'hbacf8129),
	.w2(32'h3bc2a91d),
	.w3(32'h3b033a81),
	.w4(32'h3a7035c3),
	.w5(32'h3baf99d4),
	.w6(32'h3be64913),
	.w7(32'h3c21348d),
	.w8(32'hb9a07a74),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11282d),
	.w1(32'h3a76d743),
	.w2(32'hbc1b2552),
	.w3(32'h3c841af6),
	.w4(32'h3c9763ab),
	.w5(32'hbc1b4694),
	.w6(32'h3aea8058),
	.w7(32'h3bf029e8),
	.w8(32'hbc58ebf3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd26f),
	.w1(32'hbbc2655a),
	.w2(32'h3c1ce394),
	.w3(32'hbb6b1b4a),
	.w4(32'hbb3b4c50),
	.w5(32'h3c9f100b),
	.w6(32'hbc02c5f1),
	.w7(32'hbba87907),
	.w8(32'h3be8b36d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c623f6f),
	.w1(32'h3b96b3bd),
	.w2(32'hbbca1605),
	.w3(32'h3cb26cdc),
	.w4(32'h3c676bb7),
	.w5(32'h3c3e52c2),
	.w6(32'h3c801aed),
	.w7(32'h3c03be68),
	.w8(32'hbaa136c7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c843271),
	.w1(32'h3b8d74eb),
	.w2(32'hb99d44d4),
	.w3(32'h3d35b8d0),
	.w4(32'h3cf2b046),
	.w5(32'hbadfe2ae),
	.w6(32'h3ce0d6b0),
	.w7(32'h3c87330c),
	.w8(32'hbb22c2da),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedcae8),
	.w1(32'hbb0f7b1d),
	.w2(32'hbbad6486),
	.w3(32'h3bd97745),
	.w4(32'hbb43ca66),
	.w5(32'hb98840bb),
	.w6(32'h3a1036eb),
	.w7(32'hbc07713d),
	.w8(32'hba8e8fbf),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3a1f5),
	.w1(32'h3b103c69),
	.w2(32'hbc7640e7),
	.w3(32'h3a31018d),
	.w4(32'h3b22f3bc),
	.w5(32'hbc37d4d8),
	.w6(32'hb7a66fe2),
	.w7(32'hba0644c8),
	.w8(32'hbc04217c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc492435),
	.w1(32'hbb130d42),
	.w2(32'h3bcef5c9),
	.w3(32'hbc02fb60),
	.w4(32'hbbb090ce),
	.w5(32'hbb048cc0),
	.w6(32'hbc072a3c),
	.w7(32'h3adb1d3b),
	.w8(32'h3b98dbab),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11842f),
	.w1(32'h3c0a21b5),
	.w2(32'h3a623519),
	.w3(32'h3c7984f5),
	.w4(32'h3c72c371),
	.w5(32'hb603e604),
	.w6(32'h3c4ee5b6),
	.w7(32'h3b89ed5f),
	.w8(32'h3a8d63ac),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66646),
	.w1(32'h3b3732f4),
	.w2(32'h3aff5e80),
	.w3(32'hbb69306e),
	.w4(32'h3aaad21e),
	.w5(32'h3c232132),
	.w6(32'hba2d8d90),
	.w7(32'h3aeadbf9),
	.w8(32'h3c079183),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1a6d5),
	.w1(32'h3c15caf1),
	.w2(32'hbbd83f37),
	.w3(32'h3b9f5e35),
	.w4(32'h3c66a0a0),
	.w5(32'h3cb3f16e),
	.w6(32'hbb6bb871),
	.w7(32'h3b977cf6),
	.w8(32'h3c86261d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94dd94),
	.w1(32'h3c02ea74),
	.w2(32'hbad41916),
	.w3(32'hbbe83291),
	.w4(32'hbc8aac75),
	.w5(32'h3b26398d),
	.w6(32'h3cf1d9fe),
	.w7(32'h3cb92f7a),
	.w8(32'h3b27d561),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf5915),
	.w1(32'hbb864381),
	.w2(32'hbbda0dd0),
	.w3(32'h3b6423af),
	.w4(32'h3a9fa671),
	.w5(32'hbb7b288b),
	.w6(32'h3b4d6f0b),
	.w7(32'h3a9813db),
	.w8(32'h3aadcbd9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e9a1),
	.w1(32'hba4cce5a),
	.w2(32'h3c17330e),
	.w3(32'h3bc0c601),
	.w4(32'h3c1492eb),
	.w5(32'hbbba3c04),
	.w6(32'h3bc7d21f),
	.w7(32'h3b8b4067),
	.w8(32'hbbd3bd0c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb81f47),
	.w1(32'h3c853c1e),
	.w2(32'hb9dc1d36),
	.w3(32'h3c651273),
	.w4(32'h3c3615e3),
	.w5(32'hbc104975),
	.w6(32'hbbdc847e),
	.w7(32'hba32aed9),
	.w8(32'hbc675c9f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb69a61),
	.w1(32'h3b9bdae6),
	.w2(32'hbab8e843),
	.w3(32'hbabc838d),
	.w4(32'hbac929ec),
	.w5(32'h3b85f625),
	.w6(32'hbbff47a5),
	.w7(32'hbbf1b6b8),
	.w8(32'hbb77ddde),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993b102),
	.w1(32'h3c35066d),
	.w2(32'h3b921396),
	.w3(32'hbbbe29db),
	.w4(32'h3ae95118),
	.w5(32'hbbbff759),
	.w6(32'hbbc990e8),
	.w7(32'hbc459fc9),
	.w8(32'hbbbc7f44),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9138aa),
	.w1(32'h3bbda6c0),
	.w2(32'hbc3c2db1),
	.w3(32'hbb62df65),
	.w4(32'hbb174376),
	.w5(32'hba3bb992),
	.w6(32'hbc209eed),
	.w7(32'hbc029147),
	.w8(32'h3c49c033),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e460c),
	.w1(32'hbc080a19),
	.w2(32'h3c063407),
	.w3(32'hbc56fec0),
	.w4(32'hbca7fc86),
	.w5(32'h3abcb7fd),
	.w6(32'h3b851dfe),
	.w7(32'hbba7fe0e),
	.w8(32'hba9b922b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec90b0),
	.w1(32'h3ba0e43f),
	.w2(32'hbc34727a),
	.w3(32'h3baa21fe),
	.w4(32'h3ab19eaf),
	.w5(32'hbaa06135),
	.w6(32'h3b192259),
	.w7(32'h38d6e9d8),
	.w8(32'h3c050892),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f3b94),
	.w1(32'hbc8b2032),
	.w2(32'h3bbdef01),
	.w3(32'hbcaed2fd),
	.w4(32'hbc825b51),
	.w5(32'hb9a532c9),
	.w6(32'h3cae7326),
	.w7(32'h3c205e76),
	.w8(32'hbc6c2d3e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc057908),
	.w1(32'hbaa23138),
	.w2(32'h3a9bd138),
	.w3(32'h3ba8dbec),
	.w4(32'h3c034861),
	.w5(32'hba2ab160),
	.w6(32'hbc008ac3),
	.w7(32'h3c3727b9),
	.w8(32'h3b8fea4c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6876f),
	.w1(32'h3c04e0ab),
	.w2(32'hbbf084e3),
	.w3(32'hbb5e2d1b),
	.w4(32'hba4fe313),
	.w5(32'hbc1d356b),
	.w6(32'hbb6754c7),
	.w7(32'hbc33de44),
	.w8(32'hbc1d3b14),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc519394),
	.w1(32'hbbaff9de),
	.w2(32'hbba73fae),
	.w3(32'hbc3e838e),
	.w4(32'hbc03fb3e),
	.w5(32'h3bb77231),
	.w6(32'h3c2b2572),
	.w7(32'h3c1d09ec),
	.w8(32'h3be457e2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bb68b),
	.w1(32'hbc2d8da6),
	.w2(32'h3b96487b),
	.w3(32'hbb9e82b2),
	.w4(32'hbb57d01d),
	.w5(32'hbb2a2ab0),
	.w6(32'h3a32a7d1),
	.w7(32'h3c33c59c),
	.w8(32'h3b5fcba5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c48c7),
	.w1(32'h3b05080e),
	.w2(32'hbc646c24),
	.w3(32'hb8d7db7a),
	.w4(32'hba2ddeff),
	.w5(32'hbb7c6b71),
	.w6(32'hba973116),
	.w7(32'hba10c255),
	.w8(32'hbb719126),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b4bfb),
	.w1(32'hbc69bfac),
	.w2(32'hbcb33921),
	.w3(32'hbb8f82a9),
	.w4(32'hbc1eb4a0),
	.w5(32'hbc376746),
	.w6(32'h3b955258),
	.w7(32'hbbafb4bd),
	.w8(32'hbc758b3d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88abb2),
	.w1(32'h3c2a2bac),
	.w2(32'hbc075b7a),
	.w3(32'hbb2d460e),
	.w4(32'h3c06400a),
	.w5(32'hbbee3a6a),
	.w6(32'h3b8a110c),
	.w7(32'hbaed4d48),
	.w8(32'hbbd5ea79),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c879809),
	.w1(32'hbb52d1f0),
	.w2(32'hbc852bef),
	.w3(32'hbb6e146f),
	.w4(32'hbc133c32),
	.w5(32'h3b9ec317),
	.w6(32'hbc2864c9),
	.w7(32'hbc342e78),
	.w8(32'h3c6fa4d4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ee514),
	.w1(32'hbc82d588),
	.w2(32'h3ad4f8b8),
	.w3(32'hbc45ac51),
	.w4(32'hbc1e9bf6),
	.w5(32'h3b8cbaa7),
	.w6(32'h3c964fa8),
	.w7(32'hbad169d2),
	.w8(32'h3b185a9b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c47ba),
	.w1(32'hbb7a9c40),
	.w2(32'h3b670eb2),
	.w3(32'h3af48713),
	.w4(32'h3a7be371),
	.w5(32'hbbd5028f),
	.w6(32'h3a8af1fa),
	.w7(32'hba4cacc9),
	.w8(32'hbc7cf0e8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c13ae),
	.w1(32'h3be8220e),
	.w2(32'hba941993),
	.w3(32'h3c9fa3eb),
	.w4(32'h3c7fa3ab),
	.w5(32'hbbc8042a),
	.w6(32'hbc5a1679),
	.w7(32'hbc2f128c),
	.w8(32'hbc082a49),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e695),
	.w1(32'hbab3226c),
	.w2(32'hbcc459a3),
	.w3(32'hbc441947),
	.w4(32'h3a941d91),
	.w5(32'hbc7a9c86),
	.w6(32'hbc48a62d),
	.w7(32'h3a17903e),
	.w8(32'h3b5b38d1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa623c),
	.w1(32'hbba20ffa),
	.w2(32'hba58dc83),
	.w3(32'hbcad438d),
	.w4(32'hbbe7ccbf),
	.w5(32'hbafb2274),
	.w6(32'hb9affe80),
	.w7(32'hbaeb5e3a),
	.w8(32'hba9f704f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c894856),
	.w1(32'h3b88ee8f),
	.w2(32'hbc1b7d45),
	.w3(32'h3b3956a9),
	.w4(32'h3c0cd2b5),
	.w5(32'hbc096b2e),
	.w6(32'hbbb0b29a),
	.w7(32'hba2757e5),
	.w8(32'hbb5bbdab),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c815),
	.w1(32'hbb321447),
	.w2(32'hbc88c98a),
	.w3(32'hbc7c5a2e),
	.w4(32'hbc13a090),
	.w5(32'h3c32b2f9),
	.w6(32'hbb16ec4a),
	.w7(32'h379803e0),
	.w8(32'h3c27a849),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff16ae),
	.w1(32'hbbf42301),
	.w2(32'hbb906594),
	.w3(32'hbb2e7f6c),
	.w4(32'hbc362b31),
	.w5(32'h3a417058),
	.w6(32'h3c9ea959),
	.w7(32'h3c63af16),
	.w8(32'hbbea6a66),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4fc4f),
	.w1(32'hb88b8304),
	.w2(32'hba2b19ab),
	.w3(32'h3bf00dde),
	.w4(32'h3c317a89),
	.w5(32'hbc3fe2aa),
	.w6(32'hbc02caa8),
	.w7(32'h3acf48c5),
	.w8(32'hbc2d16ff),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b41d1d),
	.w1(32'hbc19a563),
	.w2(32'hbc164f23),
	.w3(32'hbb1a38f3),
	.w4(32'hbc03344b),
	.w5(32'hbc3c9d37),
	.w6(32'hbb958c05),
	.w7(32'hbbdd80f2),
	.w8(32'hbc6a17e1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f2e10),
	.w1(32'h3ba5b689),
	.w2(32'hbb423ec6),
	.w3(32'h3a7f1cb5),
	.w4(32'h3c0cd262),
	.w5(32'hbb50ced7),
	.w6(32'h3a4f6367),
	.w7(32'hba8f7cd1),
	.w8(32'hbc0ec47e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab24e6b),
	.w1(32'h3b14c3b6),
	.w2(32'h3ba0f054),
	.w3(32'hbb787110),
	.w4(32'hbb6b4642),
	.w5(32'hba39e548),
	.w6(32'hbbe4c8f6),
	.w7(32'hbc0cf7bd),
	.w8(32'h3af347cc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34bdbf),
	.w1(32'hba773a86),
	.w2(32'hbc986e90),
	.w3(32'h3aed2a2e),
	.w4(32'hbb9c6c95),
	.w5(32'hbc99fb2a),
	.w6(32'h3bbb875a),
	.w7(32'hbc2e4404),
	.w8(32'hbc944571),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4559c8),
	.w1(32'hb9c202c7),
	.w2(32'hbc32cc0c),
	.w3(32'h3a341f7d),
	.w4(32'h3bbcdb16),
	.w5(32'hbb1d34e5),
	.w6(32'h3ac5adc0),
	.w7(32'h3c65fecb),
	.w8(32'h3c4113a4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04c27a),
	.w1(32'hbc17b1dd),
	.w2(32'h3b3dc9b6),
	.w3(32'h3bbc5ca4),
	.w4(32'hbb8de777),
	.w5(32'hba1a5b8a),
	.w6(32'h3c222808),
	.w7(32'h3adf8c61),
	.w8(32'hbc256201),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92bb15),
	.w1(32'h3b82718a),
	.w2(32'hbbe5a882),
	.w3(32'h3b278144),
	.w4(32'h3bee9fcb),
	.w5(32'hbc26e85b),
	.w6(32'hbadc58ff),
	.w7(32'h3b2ea515),
	.w8(32'h3b60d4ad),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6f0b3),
	.w1(32'hbbba8b78),
	.w2(32'hbba49854),
	.w3(32'hbc584e97),
	.w4(32'hbc7f591b),
	.w5(32'hbc33ee86),
	.w6(32'hb944b6b3),
	.w7(32'hbbcbc428),
	.w8(32'hbc433bb3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37b5f2),
	.w1(32'hbc1db2fb),
	.w2(32'hbb1aaee4),
	.w3(32'hbc516de8),
	.w4(32'hbc1da709),
	.w5(32'hbb4864cb),
	.w6(32'hbc755f21),
	.w7(32'hbc29f75f),
	.w8(32'h3b5dda9d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49e4c5),
	.w1(32'h3b947fee),
	.w2(32'h3b7bf8d5),
	.w3(32'h3a9cd505),
	.w4(32'hba36eaed),
	.w5(32'hbaab78a2),
	.w6(32'h3b15cb21),
	.w7(32'hbab9f7e5),
	.w8(32'h3b459666),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5b7c2),
	.w1(32'h3b69124e),
	.w2(32'h3bb21772),
	.w3(32'h3b1e3147),
	.w4(32'h3b8a5ac7),
	.w5(32'hbad7e119),
	.w6(32'h3b463fd8),
	.w7(32'h3b28b14b),
	.w8(32'hbc280daf),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cf7d1),
	.w1(32'h3c973f3f),
	.w2(32'h3b9e18b5),
	.w3(32'hbbd629a1),
	.w4(32'h3b9feea6),
	.w5(32'hbc388233),
	.w6(32'hbb8d04e7),
	.w7(32'hbb09c57d),
	.w8(32'h3aca589b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc3e62),
	.w1(32'h3bf48762),
	.w2(32'hbbb867df),
	.w3(32'hbbd728d4),
	.w4(32'hba2afc78),
	.w5(32'h3b6ef0bf),
	.w6(32'hbb46b27b),
	.w7(32'hba45f502),
	.w8(32'h3b1819cf),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88926c),
	.w1(32'hbbe607f3),
	.w2(32'hbade6d49),
	.w3(32'h3bdbf5e2),
	.w4(32'h3b1a9a2d),
	.w5(32'h3b9f1cfb),
	.w6(32'h3b6f497f),
	.w7(32'hbab5c80c),
	.w8(32'hbbe7f368),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76cf12),
	.w1(32'hbac3cb14),
	.w2(32'hbc21d2e6),
	.w3(32'hbb0cc742),
	.w4(32'hbb3ebbb4),
	.w5(32'hbbfcd54a),
	.w6(32'hbb1e41b8),
	.w7(32'hba3c7623),
	.w8(32'hbb07a9d8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc37b1d),
	.w1(32'hb9206bb1),
	.w2(32'h3c3fc82d),
	.w3(32'hbc0a3b9c),
	.w4(32'hbb1fefdf),
	.w5(32'hbbdbc1b1),
	.w6(32'hbabf1c14),
	.w7(32'hbaaf7751),
	.w8(32'hbc25424d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caaa64a),
	.w1(32'h3c9afb42),
	.w2(32'hbcdb5c49),
	.w3(32'hbc5d370c),
	.w4(32'hbb1d7e8d),
	.w5(32'hbb3ebfc8),
	.w6(32'hbcabc7fa),
	.w7(32'hbc9f2108),
	.w8(32'hbb3d687c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9d587),
	.w1(32'hbcc0ee75),
	.w2(32'hbb67d8a6),
	.w3(32'h3c310cc5),
	.w4(32'h3c63cca5),
	.w5(32'h3b81da39),
	.w6(32'h3bd8fba7),
	.w7(32'h3c371808),
	.w8(32'h3baa4f75),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc7439),
	.w1(32'hbb81b89d),
	.w2(32'hbb266ce3),
	.w3(32'h3b7c6071),
	.w4(32'h3b9a8511),
	.w5(32'hbc9798c4),
	.w6(32'h3bdb75c2),
	.w7(32'h3bf85d40),
	.w8(32'hbcabc132),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4c733),
	.w1(32'h3c32360a),
	.w2(32'h3b63e285),
	.w3(32'hbc8f4f5b),
	.w4(32'hbb43690d),
	.w5(32'hbbff9a61),
	.w6(32'hbcbb2d93),
	.w7(32'hbc5384fc),
	.w8(32'hbbe12408),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb582f14),
	.w1(32'h3bcf5e30),
	.w2(32'hbc642067),
	.w3(32'hbb9fc6c5),
	.w4(32'hbb232b62),
	.w5(32'hbc56e617),
	.w6(32'hba18dee0),
	.w7(32'hbc18f118),
	.w8(32'hbbd453d0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8782c),
	.w1(32'hba848586),
	.w2(32'hbc694387),
	.w3(32'hbc5b6beb),
	.w4(32'hbbdb978a),
	.w5(32'h3b7caa1a),
	.w6(32'hbc098f4c),
	.w7(32'hbbf5b798),
	.w8(32'h3ad2510a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc05a6),
	.w1(32'hbc23b37a),
	.w2(32'hbb23fb1e),
	.w3(32'hbc83bf04),
	.w4(32'hbc8678ec),
	.w5(32'h3adc793b),
	.w6(32'h3c0cb47f),
	.w7(32'hbb513fe7),
	.w8(32'h3b128f42),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446f61),
	.w1(32'h394c69e5),
	.w2(32'hbaf56d20),
	.w3(32'h3ba96b62),
	.w4(32'h3bd834b4),
	.w5(32'h3b4422cd),
	.w6(32'hb9a95f1c),
	.w7(32'h3aa8e4b8),
	.w8(32'hb870cd08),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63f5a3),
	.w1(32'hbaa71803),
	.w2(32'hbb6b9837),
	.w3(32'hb8339f6e),
	.w4(32'h3aa4e741),
	.w5(32'hbc18d5f4),
	.w6(32'h3be6ebf1),
	.w7(32'h3b5ff882),
	.w8(32'hbbfc3474),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cc12c),
	.w1(32'h3b113272),
	.w2(32'h3c01fcc4),
	.w3(32'hbae874c1),
	.w4(32'h3ac062b4),
	.w5(32'h3ac91157),
	.w6(32'hbb0dd8fb),
	.w7(32'hba82f084),
	.w8(32'hbc39b95c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c283c22),
	.w1(32'hb91475e7),
	.w2(32'hbbb58e8e),
	.w3(32'h3baf9f68),
	.w4(32'h3b8dfb6f),
	.w5(32'hbb680f2a),
	.w6(32'hbc3eb258),
	.w7(32'h3b812be9),
	.w8(32'h3b6654cd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32874b),
	.w1(32'hbc8394d9),
	.w2(32'h3be2dade),
	.w3(32'hbc63a865),
	.w4(32'hbc96d149),
	.w5(32'hbbb1fc33),
	.w6(32'h3bd133ae),
	.w7(32'h3ad647de),
	.w8(32'hbc01fba3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8e61d),
	.w1(32'h3c492d9a),
	.w2(32'hbb11661d),
	.w3(32'hbc2a7dd9),
	.w4(32'hbb50df06),
	.w5(32'hbc916698),
	.w6(32'hbb875e27),
	.w7(32'hbcbb315a),
	.w8(32'hbc7066a6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b511390),
	.w1(32'h3b8d9adf),
	.w2(32'hba16ef3c),
	.w3(32'hbc87339e),
	.w4(32'hbb398cbc),
	.w5(32'hba276f8a),
	.w6(32'hbc280e93),
	.w7(32'h3b9198c3),
	.w8(32'h3b6338fd),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd9856),
	.w1(32'hb9e32178),
	.w2(32'hbc3577d3),
	.w3(32'h3c5fb1e3),
	.w4(32'h3bdedead),
	.w5(32'hbb2195e3),
	.w6(32'h3ac72ae6),
	.w7(32'hbab0f64f),
	.w8(32'hbb3e076c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb678ae5),
	.w1(32'hbb04b70a),
	.w2(32'hbb1b69f9),
	.w3(32'hbb757fa0),
	.w4(32'hb8a9d7c2),
	.w5(32'hbc1f0c6f),
	.w6(32'hbb11b472),
	.w7(32'hba692fbb),
	.w8(32'hbb69e3fc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0262b4),
	.w1(32'h3b6322d6),
	.w2(32'hbaa78126),
	.w3(32'hbbb0bd66),
	.w4(32'hb9c0f7cd),
	.w5(32'h3a4c8856),
	.w6(32'hbc1554a8),
	.w7(32'hbb6a3115),
	.w8(32'h3b16cdf0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb704ae),
	.w1(32'h3c4ab5c7),
	.w2(32'h3c3547e9),
	.w3(32'h3b5cd018),
	.w4(32'hbb184635),
	.w5(32'hbc1c4611),
	.w6(32'h3c86f112),
	.w7(32'h3bf281a5),
	.w8(32'h3b7b5b03),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd18b7d),
	.w1(32'h3c51d7da),
	.w2(32'hbae2e676),
	.w3(32'h3b8aebf0),
	.w4(32'hbbbc13b5),
	.w5(32'h3be811bf),
	.w6(32'hbb2e89c9),
	.w7(32'hbc347db9),
	.w8(32'hbb2d4697),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a9fdd),
	.w1(32'h3c5cf8f1),
	.w2(32'hbc39213b),
	.w3(32'h3cc83fe2),
	.w4(32'h3cababa8),
	.w5(32'hbb8785b3),
	.w6(32'h3c6809a8),
	.w7(32'h3c172b36),
	.w8(32'hbc3ac089),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc38315),
	.w1(32'h3acc41da),
	.w2(32'hb99d26f5),
	.w3(32'hbb88055d),
	.w4(32'h3b4d238b),
	.w5(32'h3b64a262),
	.w6(32'hbbc381e5),
	.w7(32'h3a743b1e),
	.w8(32'h3be15d97),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d7a1a),
	.w1(32'hbb7c13a5),
	.w2(32'h3baa79bf),
	.w3(32'hbbe9d2b7),
	.w4(32'h3bb635ce),
	.w5(32'hba839740),
	.w6(32'hbb5f5bf5),
	.w7(32'h3be0ee1a),
	.w8(32'hb9f00b5c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c014ddd),
	.w1(32'h3c12797d),
	.w2(32'h3c95ed54),
	.w3(32'hbaed8feb),
	.w4(32'h3bdca7d5),
	.w5(32'h3cb22c48),
	.w6(32'hbbd80b2e),
	.w7(32'hbb86ce08),
	.w8(32'hbb94f9c2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d23a4fa),
	.w1(32'h3ce4bbc0),
	.w2(32'h3b9b586b),
	.w3(32'h3d56a692),
	.w4(32'h3d6081a1),
	.w5(32'hbc2ec622),
	.w6(32'hb9955c09),
	.w7(32'h3bad7440),
	.w8(32'hbc0b24a2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b04af),
	.w1(32'h3bd8e184),
	.w2(32'hb9a1d716),
	.w3(32'hbc34b1c6),
	.w4(32'hbc336e1c),
	.w5(32'h3baf6a9c),
	.w6(32'hbc0dd077),
	.w7(32'hbbcba3c4),
	.w8(32'h3a341d1f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe39a42),
	.w1(32'hba517f53),
	.w2(32'hbac75212),
	.w3(32'h3a310a4f),
	.w4(32'hbb8b6876),
	.w5(32'hbc5d53cb),
	.w6(32'hba64156f),
	.w7(32'hbb1be11f),
	.w8(32'hbb0ad222),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10aa8f),
	.w1(32'hbc0d3caa),
	.w2(32'h3bf44a92),
	.w3(32'hbbe6ef56),
	.w4(32'hbbfb42c0),
	.w5(32'h3bd64bd8),
	.w6(32'hbc4c2e9b),
	.w7(32'hbc9b77b0),
	.w8(32'h3ae44e00),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4042b7),
	.w1(32'h3b0a7e4a),
	.w2(32'hbc607b36),
	.w3(32'hbaf535ac),
	.w4(32'h37d6e834),
	.w5(32'hbc47bcd4),
	.w6(32'h39b00cc8),
	.w7(32'hbc091917),
	.w8(32'hbbb53bdd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5967b9),
	.w1(32'hbb1830f4),
	.w2(32'hbbfb4444),
	.w3(32'hbba8ac16),
	.w4(32'hbab0b7ec),
	.w5(32'hbc7395bd),
	.w6(32'h3b41179b),
	.w7(32'hbb81cbcf),
	.w8(32'hbad54b8b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b460),
	.w1(32'hbb5b78b3),
	.w2(32'hbb647128),
	.w3(32'hbb2beb23),
	.w4(32'h3bd809d1),
	.w5(32'hbbcc676c),
	.w6(32'hbc1c46ac),
	.w7(32'hb96ebc3b),
	.w8(32'h3ad60acf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31a600),
	.w1(32'h3be6f3f1),
	.w2(32'hbc12ca4a),
	.w3(32'h3aca0106),
	.w4(32'hbbf6bca3),
	.w5(32'hbc435875),
	.w6(32'h3b4bf792),
	.w7(32'hbb89c76e),
	.w8(32'hbad591f4),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9938449),
	.w1(32'hbc143a68),
	.w2(32'hba09dbcb),
	.w3(32'hbc07fae1),
	.w4(32'hbc6cd4c2),
	.w5(32'hbc21bfa8),
	.w6(32'h3b9fd832),
	.w7(32'h3afcbb0a),
	.w8(32'hbb93b688),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82b759),
	.w1(32'hbbbb5719),
	.w2(32'hbb7b9582),
	.w3(32'hbc3b5fc1),
	.w4(32'hbbff0943),
	.w5(32'h398942ee),
	.w6(32'hbb814c8f),
	.w7(32'hbbcf71e1),
	.w8(32'h3b399e11),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb36640),
	.w1(32'h3a4aabbf),
	.w2(32'hbbc12a18),
	.w3(32'h39afc7cf),
	.w4(32'hba85c917),
	.w5(32'hbab08cbd),
	.w6(32'hb90d7674),
	.w7(32'hbb56511b),
	.w8(32'h3a53d90d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78eeb9),
	.w1(32'h3ad60cb6),
	.w2(32'hbc00651b),
	.w3(32'hbb07e347),
	.w4(32'h3b81f0a5),
	.w5(32'hba93818c),
	.w6(32'h3aa7b0f0),
	.w7(32'h3b01061c),
	.w8(32'h3bda5c89),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41e371),
	.w1(32'hbc19709f),
	.w2(32'h3c59b6cc),
	.w3(32'hbb8a7990),
	.w4(32'hbb87e27c),
	.w5(32'hbb88b1ed),
	.w6(32'h3bcda3bb),
	.w7(32'h3bf1e66d),
	.w8(32'hba3b4f46),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51d639),
	.w1(32'h3b2acab0),
	.w2(32'h3b75e80c),
	.w3(32'hbc293c06),
	.w4(32'hbb73d5bf),
	.w5(32'hbbbd779f),
	.w6(32'hbc863c38),
	.w7(32'hbc1e6e10),
	.w8(32'h3bcbf1f4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2cb86),
	.w1(32'hbc39878e),
	.w2(32'h3c191321),
	.w3(32'h3bcc2053),
	.w4(32'h3b6ba21b),
	.w5(32'h3c2dfebb),
	.w6(32'h3c08dd09),
	.w7(32'h3bef6a1a),
	.w8(32'h3879f450),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a860f),
	.w1(32'h3c123327),
	.w2(32'h3c0765df),
	.w3(32'h3b68f662),
	.w4(32'h3b14f4a6),
	.w5(32'h3ac53caf),
	.w6(32'h3b607300),
	.w7(32'h3af96cd1),
	.w8(32'hba90fb4a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0860e8),
	.w1(32'hbc4d1335),
	.w2(32'hbb8e7ec7),
	.w3(32'h3a7f7282),
	.w4(32'hba092ffa),
	.w5(32'hbba34afe),
	.w6(32'hbb254973),
	.w7(32'hbb988df0),
	.w8(32'hbc272a31),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab5b10),
	.w1(32'h3c944909),
	.w2(32'hbc713eae),
	.w3(32'h3c373759),
	.w4(32'h3c128bdd),
	.w5(32'h3c01ff69),
	.w6(32'hbc27efb5),
	.w7(32'hb9981b3b),
	.w8(32'hbb6d53a0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fde81),
	.w1(32'hbc0acd38),
	.w2(32'h3c872347),
	.w3(32'h3c4db328),
	.w4(32'hbb8b7e0e),
	.w5(32'h3bc87c64),
	.w6(32'h3b53caa7),
	.w7(32'h3ba36b33),
	.w8(32'hbc9b6025),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7a83a),
	.w1(32'h3c465038),
	.w2(32'hbb12797e),
	.w3(32'h3c7b407a),
	.w4(32'h3c8a69ce),
	.w5(32'h3b695f89),
	.w6(32'hbc077384),
	.w7(32'hbbca060a),
	.w8(32'h3b97b3d6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec33d),
	.w1(32'hbb91abf7),
	.w2(32'hbbee9c3d),
	.w3(32'hba670892),
	.w4(32'hba9953ee),
	.w5(32'hbbe9cc77),
	.w6(32'h3bd163b9),
	.w7(32'h3a8a4243),
	.w8(32'h394b68ed),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46c0b2),
	.w1(32'hbb031396),
	.w2(32'hb9d706a7),
	.w3(32'hbc197ba5),
	.w4(32'hbbc53d63),
	.w5(32'h3b03742b),
	.w6(32'h3b1771b0),
	.w7(32'h3c09fc9a),
	.w8(32'h3b379aef),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8487b4),
	.w1(32'hba3b91aa),
	.w2(32'hbb397c04),
	.w3(32'hbb26b35e),
	.w4(32'hbac1729f),
	.w5(32'hbb3fbc43),
	.w6(32'h3b1ec5e4),
	.w7(32'hbb39ad0d),
	.w8(32'h3b9d1844),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0229a),
	.w1(32'hbb1e9595),
	.w2(32'hbcbb8b4d),
	.w3(32'hbc13550b),
	.w4(32'h3a976259),
	.w5(32'hbc9a944f),
	.w6(32'h3b931d9e),
	.w7(32'hbbed5dda),
	.w8(32'hbc70528a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44ec79),
	.w1(32'h3ab62653),
	.w2(32'h3b732255),
	.w3(32'hbb91bf5c),
	.w4(32'hbb2ae6c4),
	.w5(32'hbb33e2a7),
	.w6(32'hbc0bba9c),
	.w7(32'hbb86aa60),
	.w8(32'h3b3e7827),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdf085),
	.w1(32'h3bd73a80),
	.w2(32'hbb30acd9),
	.w3(32'hbb8060c0),
	.w4(32'h3b2d1691),
	.w5(32'hba6b0b65),
	.w6(32'hbbbf240e),
	.w7(32'hbc1337a7),
	.w8(32'hba818ac9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfc587),
	.w1(32'hbb89f354),
	.w2(32'hb99bdbd4),
	.w3(32'hbabdb2a8),
	.w4(32'hbb415678),
	.w5(32'hbba1e6c9),
	.w6(32'hba532f18),
	.w7(32'hbab133f6),
	.w8(32'hbbb680cd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98dedb),
	.w1(32'h3b8b27a2),
	.w2(32'hbc5bd9be),
	.w3(32'hbb2ca861),
	.w4(32'hbb13dfa5),
	.w5(32'h3a78a1ac),
	.w6(32'hbaf386d1),
	.w7(32'hbb36af58),
	.w8(32'h3c36e07b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80e398),
	.w1(32'hbaac4ff5),
	.w2(32'hbb00d778),
	.w3(32'hbc610b9f),
	.w4(32'hbccb51f7),
	.w5(32'h3b26e777),
	.w6(32'h3c563e14),
	.w7(32'hbc1304e6),
	.w8(32'h3b08fbef),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf4441),
	.w1(32'hbbfc0aee),
	.w2(32'hbb989f52),
	.w3(32'h3a1b8ead),
	.w4(32'h3a58050e),
	.w5(32'hbc50c9f0),
	.w6(32'h3a89c137),
	.w7(32'h3b160c1e),
	.w8(32'hbbe175de),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5d7d8),
	.w1(32'hbbdfe32b),
	.w2(32'hbcbf248b),
	.w3(32'hbc346a11),
	.w4(32'hbbdad04f),
	.w5(32'hbc94ad56),
	.w6(32'hbc875cef),
	.w7(32'hbc550d19),
	.w8(32'hbc84828b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a515e),
	.w1(32'h3c275847),
	.w2(32'h3c7e08c8),
	.w3(32'hbc81f094),
	.w4(32'hbc1351f6),
	.w5(32'hbbf533be),
	.w6(32'hbc621075),
	.w7(32'hbc69bd94),
	.w8(32'hbb4a6eee),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6fea4),
	.w1(32'h3cd02ea8),
	.w2(32'h3c04b141),
	.w3(32'hbc91941e),
	.w4(32'hbbb46b22),
	.w5(32'h3a71d5cb),
	.w6(32'hbccf50a2),
	.w7(32'hbc501d33),
	.w8(32'hbbd19e56),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule