module layer_10_featuremap_185(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f0931b),
	.w1(32'hb5bdd883),
	.w2(32'hb619f4a0),
	.w3(32'h354b3557),
	.w4(32'h3610ce92),
	.w5(32'h35cc2758),
	.w6(32'h34c31fda),
	.w7(32'hb5d61565),
	.w8(32'h369cac10),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836fb86),
	.w1(32'hb84a3207),
	.w2(32'hb8823c12),
	.w3(32'hb796cd8d),
	.w4(32'hb7c3330f),
	.w5(32'hb864afef),
	.w6(32'hb821b307),
	.w7(32'hb7bc9dec),
	.w8(32'hb7c91c80),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b13e3d),
	.w1(32'h34f449c6),
	.w2(32'h3558ad3b),
	.w3(32'hb62f80fd),
	.w4(32'h35b8331e),
	.w5(32'h34ea23ab),
	.w6(32'h35c66810),
	.w7(32'h360c4ea0),
	.w8(32'h35b9a8ea),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37282a35),
	.w1(32'hb7089252),
	.w2(32'hb71c385d),
	.w3(32'hb698563f),
	.w4(32'hb7d527ba),
	.w5(32'h364a5eb3),
	.w6(32'h36253038),
	.w7(32'hb724dc5a),
	.w8(32'hb61f2171),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68a5350),
	.w1(32'hb5a8b907),
	.w2(32'h3659b5dc),
	.w3(32'hb6dba7c6),
	.w4(32'hb6884e25),
	.w5(32'hb520ac18),
	.w6(32'hb6444ff1),
	.w7(32'hb5eec6c3),
	.w8(32'hb669fdf6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358c4ba4),
	.w1(32'h358c3847),
	.w2(32'h3591e3d7),
	.w3(32'h35607eeb),
	.w4(32'h362cf840),
	.w5(32'h3624923d),
	.w6(32'h35fcdee9),
	.w7(32'h361d48c6),
	.w8(32'h358565ae),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc981d),
	.w1(32'hb73a01ce),
	.w2(32'h39428d93),
	.w3(32'hb8f69b0b),
	.w4(32'hb8d300b7),
	.w5(32'h390fadd9),
	.w6(32'hb915335a),
	.w7(32'h3841d320),
	.w8(32'h391003a0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ecd17b),
	.w1(32'h3a0a3f94),
	.w2(32'h39c2704e),
	.w3(32'h386aff97),
	.w4(32'h38be416c),
	.w5(32'h39af4112),
	.w6(32'hb805f38c),
	.w7(32'h38b5a39c),
	.w8(32'h38044436),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81231ca),
	.w1(32'hb7bff259),
	.w2(32'hb8122557),
	.w3(32'hb756595b),
	.w4(32'hb7991dcb),
	.w5(32'hb54e62fc),
	.w6(32'h37a88219),
	.w7(32'hb7eb91f2),
	.w8(32'hb7381663),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812a21b),
	.w1(32'h38854997),
	.w2(32'h38f3f75e),
	.w3(32'hb80dc389),
	.w4(32'h388693fc),
	.w5(32'h38fbf1e1),
	.w6(32'h38a4b7f3),
	.w7(32'h36ca7898),
	.w8(32'h378a344a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba68e9),
	.w1(32'hb786557c),
	.w2(32'hb704ad4b),
	.w3(32'hb723ca68),
	.w4(32'h35abb682),
	.w5(32'h36d74a2a),
	.w6(32'hb696aea0),
	.w7(32'hb6c8a2ba),
	.w8(32'h37259efb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884ebe2),
	.w1(32'hb82914fd),
	.w2(32'h3941a12f),
	.w3(32'hb900f8a1),
	.w4(32'hb928c5fb),
	.w5(32'h391ca041),
	.w6(32'hb93bc762),
	.w7(32'hb70c5309),
	.w8(32'h391eb844),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36eff498),
	.w1(32'h38cf4688),
	.w2(32'h39284247),
	.w3(32'hb85af4c0),
	.w4(32'h38a3a8cc),
	.w5(32'h38e8d48b),
	.w6(32'h36c42130),
	.w7(32'h37269ddb),
	.w8(32'h3815a851),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7abdb12),
	.w1(32'h387a67fe),
	.w2(32'h38df4528),
	.w3(32'hb831fb93),
	.w4(32'h388ee6cb),
	.w5(32'h38a21df6),
	.w6(32'hb8b5adda),
	.w7(32'hb6fabaa2),
	.w8(32'h38059d10),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891f246),
	.w1(32'hb87dd2ce),
	.w2(32'hb7a95b29),
	.w3(32'hb724b2d3),
	.w4(32'hb88df5ac),
	.w5(32'hb816dde3),
	.w6(32'hb6a0d4f9),
	.w7(32'hb880c7d9),
	.w8(32'hb81c4331),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382e57c8),
	.w1(32'h38d5a0a3),
	.w2(32'hb75fc738),
	.w3(32'hb866fc1d),
	.w4(32'h38e2d374),
	.w5(32'hb7ce8621),
	.w6(32'hb6281c9a),
	.w7(32'h381a9f57),
	.w8(32'hb7e2be4b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76bfed1),
	.w1(32'hb6c1388f),
	.w2(32'h36ad9f6d),
	.w3(32'h37afa70d),
	.w4(32'h37eaee1d),
	.w5(32'h37e1b109),
	.w6(32'h37f33b55),
	.w7(32'h37a8af96),
	.w8(32'h37b2514c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3702c663),
	.w1(32'h39942072),
	.w2(32'h396bfb78),
	.w3(32'hb85650e0),
	.w4(32'h3964ba78),
	.w5(32'h39818d51),
	.w6(32'h38ee8b13),
	.w7(32'h3912fee1),
	.w8(32'h38a98598),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37707929),
	.w1(32'h391e0b13),
	.w2(32'h38f9f91f),
	.w3(32'hb79e1a9d),
	.w4(32'h38c52cf2),
	.w5(32'h39015c47),
	.w6(32'h38791ecc),
	.w7(32'h389c6b13),
	.w8(32'h38307413),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59bf293),
	.w1(32'hb5b3f6a0),
	.w2(32'hb5d9d008),
	.w3(32'hb5b7223d),
	.w4(32'hb5d19c34),
	.w5(32'hb5562dab),
	.w6(32'hb5fd3a80),
	.w7(32'hb4e30a3e),
	.w8(32'hb5c1c57d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36117ef6),
	.w1(32'h367114c4),
	.w2(32'h368c9a96),
	.w3(32'hb5e33b77),
	.w4(32'h35f89c0b),
	.w5(32'h36413c7f),
	.w6(32'hb5a187a0),
	.w7(32'hb4143b4f),
	.w8(32'h35f2b593),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64c7a1a),
	.w1(32'hb7a06de4),
	.w2(32'hb7e16f27),
	.w3(32'hb76e2c6b),
	.w4(32'hb795374f),
	.w5(32'hb7a2cc65),
	.w6(32'hb7a55b5f),
	.w7(32'hb525bc32),
	.w8(32'hb5743e68),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371db51d),
	.w1(32'hb844bbd8),
	.w2(32'h39a00bcf),
	.w3(32'hb808f17a),
	.w4(32'h394af198),
	.w5(32'h392f7cf8),
	.w6(32'h3651d4b9),
	.w7(32'h388dd836),
	.w8(32'h38e6b02a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8593308),
	.w1(32'hb7ee2da6),
	.w2(32'h380ab52c),
	.w3(32'hb834774a),
	.w4(32'hb82c4fb8),
	.w5(32'h37469778),
	.w6(32'hb57eda01),
	.w7(32'hb80a0965),
	.w8(32'hb78cc5cc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0abab),
	.w1(32'hb87e2de8),
	.w2(32'hb89a9093),
	.w3(32'h385f498e),
	.w4(32'hb8792385),
	.w5(32'hb8bbdf6c),
	.w6(32'h37ad6243),
	.w7(32'hb82ad2d2),
	.w8(32'hb81a01bb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80971aa),
	.w1(32'hb8253b55),
	.w2(32'hb782812c),
	.w3(32'hb6f03eda),
	.w4(32'hb7ed72ad),
	.w5(32'hb78aa5ad),
	.w6(32'h35eb2989),
	.w7(32'hb7e4e80a),
	.w8(32'hb81fd0bf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e393f9),
	.w1(32'hb31580c8),
	.w2(32'hb6861754),
	.w3(32'h35ae5a96),
	.w4(32'h35c4efda),
	.w5(32'hb629b37d),
	.w6(32'hb5fe52f8),
	.w7(32'hb504875f),
	.w8(32'hb66f0d5f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e821b),
	.w1(32'h38fde1ab),
	.w2(32'hb8d5a935),
	.w3(32'h38db47d4),
	.w4(32'h391ea7b5),
	.w5(32'hb8760b2d),
	.w6(32'h389619c8),
	.w7(32'h37aa6110),
	.w8(32'hb8784fa4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb698d7d7),
	.w1(32'hb78a1e78),
	.w2(32'hb7eb9818),
	.w3(32'hb78f55aa),
	.w4(32'hb7936888),
	.w5(32'hb7a9ff98),
	.w6(32'hb74489c6),
	.w7(32'hb6ee3d8a),
	.w8(32'hb7943e27),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3720bc1d),
	.w1(32'hb8355cad),
	.w2(32'hb86c3ea2),
	.w3(32'h3783b019),
	.w4(32'hb84f2766),
	.w5(32'hb8fa15fd),
	.w6(32'hb7a8c046),
	.w7(32'hb8beeb45),
	.w8(32'hb8c310d4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb2d7a71f),
	.w1(32'hb4f95ef0),
	.w2(32'hb42ab2d1),
	.w3(32'h35050666),
	.w4(32'h34b1cb45),
	.w5(32'h349bd955),
	.w6(32'hb54a1744),
	.w7(32'h33e7b909),
	.w8(32'h3462239c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362191c4),
	.w1(32'hb507ff48),
	.w2(32'hb5eb77d2),
	.w3(32'h35d890cb),
	.w4(32'hb598dbe5),
	.w5(32'hb5e547cc),
	.w6(32'hb547ea35),
	.w7(32'hb6006faf),
	.w8(32'hb624da70),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f0027c),
	.w1(32'h38144cb0),
	.w2(32'h389ab262),
	.w3(32'hb8260718),
	.w4(32'h368dbd14),
	.w5(32'h3876a791),
	.w6(32'hb5a45e6a),
	.w7(32'hb6237f9e),
	.w8(32'hb645bfd5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ba08df),
	.w1(32'hb826f190),
	.w2(32'hb80ace73),
	.w3(32'h37eee507),
	.w4(32'hb7a716f1),
	.w5(32'hb7a53dd4),
	.w6(32'h371393c0),
	.w7(32'hb78747b4),
	.w8(32'hb79089ab),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3699c645),
	.w1(32'h382d7150),
	.w2(32'h37d09924),
	.w3(32'hb7111663),
	.w4(32'h3791ace4),
	.w5(32'h380feacc),
	.w6(32'h370e634f),
	.w7(32'h37bfd287),
	.w8(32'hb41d4d94),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86bcf1f),
	.w1(32'hb7b720a8),
	.w2(32'h391dd24f),
	.w3(32'hb856751c),
	.w4(32'hb8a95a4b),
	.w5(32'h38d8e467),
	.w6(32'hb8413672),
	.w7(32'h371056ba),
	.w8(32'h3880a567),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8967218),
	.w1(32'hb95cc1a1),
	.w2(32'h39bf497f),
	.w3(32'hb78f2fdc),
	.w4(32'hb946ffb1),
	.w5(32'h3a0eddf0),
	.w6(32'hb8f4c966),
	.w7(32'hb88f20ec),
	.w8(32'h39bc198b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a07a49),
	.w1(32'hb8f57b1f),
	.w2(32'hb936e5c8),
	.w3(32'h3917b50a),
	.w4(32'hb7b0dd4d),
	.w5(32'hb8d31463),
	.w6(32'hb8242483),
	.w7(32'hb81a4044),
	.w8(32'h36b9bdf0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36126f42),
	.w1(32'hb883c935),
	.w2(32'hb919936d),
	.w3(32'hb73b3e86),
	.w4(32'hb7676d02),
	.w5(32'hb8b5fda9),
	.w6(32'hb90726ae),
	.w7(32'hb891d120),
	.w8(32'hb8803977),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb635498e),
	.w1(32'hb78d70b6),
	.w2(32'hb713573d),
	.w3(32'h36e03913),
	.w4(32'hb7a5dac8),
	.w5(32'hb73824bc),
	.w6(32'h353a92af),
	.w7(32'hb756378a),
	.w8(32'hb759a75e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354a9d7b),
	.w1(32'hb5cdefe1),
	.w2(32'h36d2a9e6),
	.w3(32'h3562d2fb),
	.w4(32'hb29ec967),
	.w5(32'h37015c2e),
	.w6(32'hb61fe937),
	.w7(32'h3695956b),
	.w8(32'hb634dba3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36079d6e),
	.w1(32'h35795dab),
	.w2(32'hb6b87442),
	.w3(32'h35a2ac46),
	.w4(32'h351ac1bd),
	.w5(32'hb6ac8614),
	.w6(32'hb65981a6),
	.w7(32'hb643d1bc),
	.w8(32'hb690da67),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722ef5d),
	.w1(32'hb78e2a3f),
	.w2(32'hb7df6050),
	.w3(32'hb663b69f),
	.w4(32'hb6a868f5),
	.w5(32'hb703eef5),
	.w6(32'h359a2b6a),
	.w7(32'hb6fa77f3),
	.w8(32'hb7d8e9f1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39020159),
	.w1(32'h398b7e49),
	.w2(32'h37f68f16),
	.w3(32'h38c60c5d),
	.w4(32'h39a0fc42),
	.w5(32'hb761e551),
	.w6(32'h3903bfbe),
	.w7(32'h38e37698),
	.w8(32'hb8d63aa3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb770a98b),
	.w1(32'hb880205e),
	.w2(32'hb835b8ef),
	.w3(32'h37b369a4),
	.w4(32'hb8199c7a),
	.w5(32'hb87c7cc1),
	.w6(32'h367523c1),
	.w7(32'hb8b98958),
	.w8(32'hb880f01a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0ee5e),
	.w1(32'hb88f98ff),
	.w2(32'h385b6de3),
	.w3(32'hb7435305),
	.w4(32'hb88eb518),
	.w5(32'hb838c313),
	.w6(32'hb74e9bb1),
	.w7(32'hb88693a9),
	.w8(32'hb883009f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371bdae6),
	.w1(32'h37a423db),
	.w2(32'h37c643f5),
	.w3(32'h35cc3322),
	.w4(32'hb781debb),
	.w5(32'hb78c2dcf),
	.w6(32'h34c61750),
	.w7(32'hb7c330e7),
	.w8(32'hb7afba5c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a2c4cf),
	.w1(32'h39296de2),
	.w2(32'h39a3be74),
	.w3(32'hb902d223),
	.w4(32'h378b747a),
	.w5(32'h3958142c),
	.w6(32'hb686499b),
	.w7(32'h38ce5fe0),
	.w8(32'h39074af4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360f4700),
	.w1(32'h3608e6c6),
	.w2(32'h362080c8),
	.w3(32'h3645a2b9),
	.w4(32'hb64015fb),
	.w5(32'h3651dd85),
	.w6(32'hb66382c9),
	.w7(32'hb6f83ba3),
	.w8(32'hb5b7cdc6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7699a27),
	.w1(32'h37035e49),
	.w2(32'h37d4ab6d),
	.w3(32'hb74e88ed),
	.w4(32'hb7a85ece),
	.w5(32'hb5d1cb96),
	.w6(32'h37ae0808),
	.w7(32'hb7b328ec),
	.w8(32'hb6c38349),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb691a956),
	.w1(32'h35c0ad5a),
	.w2(32'h36f0f75d),
	.w3(32'hb6cbfde2),
	.w4(32'hb6ec1c1f),
	.w5(32'hb5fb7dde),
	.w6(32'hb6d1ec79),
	.w7(32'hb7223fd3),
	.w8(32'hb6c9fbbd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389283ce),
	.w1(32'h386c63d8),
	.w2(32'h38a36519),
	.w3(32'h381aeb1c),
	.w4(32'h38bf4e7d),
	.w5(32'h372b4285),
	.w6(32'h365417fa),
	.w7(32'h37988f35),
	.w8(32'hb661817c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37420ef3),
	.w1(32'h380a0277),
	.w2(32'h37c24d03),
	.w3(32'h35a9ad53),
	.w4(32'h37540803),
	.w5(32'h37a50237),
	.w6(32'hb5e986d2),
	.w7(32'h37541abc),
	.w8(32'h37407056),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aa647e),
	.w1(32'h394a5f84),
	.w2(32'h393f3c93),
	.w3(32'hb8a84518),
	.w4(32'h382d398a),
	.w5(32'h39010386),
	.w6(32'h38f22dae),
	.w7(32'h3851e7c7),
	.w8(32'hb7829fce),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381bb37c),
	.w1(32'h38c1adbe),
	.w2(32'h370405a7),
	.w3(32'h382f8b7d),
	.w4(32'h38c11910),
	.w5(32'hb682fe73),
	.w6(32'h382e0c90),
	.w7(32'h3846b85e),
	.w8(32'hb7cd6c71),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a56c90),
	.w1(32'hb746c489),
	.w2(32'hb6e96cc5),
	.w3(32'hb5bcc43d),
	.w4(32'hb745a2ee),
	.w5(32'hb7122967),
	.w6(32'hb6d28d31),
	.w7(32'hb7334b6f),
	.w8(32'hb7197c04),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb628ba62),
	.w1(32'hb6363d3c),
	.w2(32'h3597ce71),
	.w3(32'hb6120b22),
	.w4(32'hb5b17b1e),
	.w5(32'h35ee7664),
	.w6(32'hb5aefe27),
	.w7(32'h362cd2f5),
	.w8(32'h356b75cf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366b42ee),
	.w1(32'hb57e26a6),
	.w2(32'h3646d93c),
	.w3(32'h36c8ab25),
	.w4(32'hb6594eaa),
	.w5(32'hb627fcef),
	.w6(32'hb66ba4d7),
	.w7(32'hb6568080),
	.w8(32'hb7193731),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb762e205),
	.w1(32'hb79cb187),
	.w2(32'hb7a9faed),
	.w3(32'hb7156982),
	.w4(32'hb73e44bb),
	.w5(32'hb73b7534),
	.w6(32'hb6720383),
	.w7(32'hb60c0a84),
	.w8(32'hb50b2ff0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71c35f3),
	.w1(32'hb6ba4fd1),
	.w2(32'hb728f192),
	.w3(32'hb7234dcf),
	.w4(32'hb69c4bc9),
	.w5(32'hb73b36a3),
	.w6(32'hb7089e0c),
	.w7(32'h372b7e63),
	.w8(32'hb67a8696),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b20bff),
	.w1(32'h38eaae93),
	.w2(32'h38b43fc0),
	.w3(32'hb7837639),
	.w4(32'h38abf705),
	.w5(32'h3880f40c),
	.w6(32'hb61902aa),
	.w7(32'h384d5ef5),
	.w8(32'h3831deb7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392bdbc0),
	.w1(32'h393213f0),
	.w2(32'hb825495a),
	.w3(32'h38e39288),
	.w4(32'h396b431a),
	.w5(32'hb800affe),
	.w6(32'h38e7e876),
	.w7(32'h3900656d),
	.w8(32'hb815e4cf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb2fbef98),
	.w1(32'h3623c5d8),
	.w2(32'hb5f10e32),
	.w3(32'h36152fdf),
	.w4(32'h3675e2df),
	.w5(32'hb64ae886),
	.w6(32'h368052c2),
	.w7(32'hb6a6d716),
	.w8(32'hb65ce3ca),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34730bca),
	.w1(32'h35c7a430),
	.w2(32'h355d7ee5),
	.w3(32'hb6087bda),
	.w4(32'h35c99fa8),
	.w5(32'h3465040d),
	.w6(32'h3652b520),
	.w7(32'h35b72589),
	.w8(32'hb59ef5d6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb658e0dd),
	.w1(32'hb5970693),
	.w2(32'hb5a58a03),
	.w3(32'hb662fbf4),
	.w4(32'hb5c29691),
	.w5(32'hb60f5884),
	.w6(32'hb5fb4891),
	.w7(32'hb56a0915),
	.w8(32'hb5ced698),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356aca3c),
	.w1(32'h3570745d),
	.w2(32'hb62d5b5f),
	.w3(32'h338085bf),
	.w4(32'h3402507b),
	.w5(32'hb647698b),
	.w6(32'hb408142b),
	.w7(32'hb552c58e),
	.w8(32'hb6e4798a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f8898),
	.w1(32'h39c62045),
	.w2(32'h388a04b9),
	.w3(32'hb882d789),
	.w4(32'h3940e6a3),
	.w5(32'h391b335e),
	.w6(32'h37d408b2),
	.w7(32'h38ad2dd7),
	.w8(32'hb8562875),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927fe98),
	.w1(32'h3925aea8),
	.w2(32'h3989c03a),
	.w3(32'hb862b06b),
	.w4(32'h356a4fb0),
	.w5(32'h372bcde3),
	.w6(32'hb78ec2dc),
	.w7(32'h38e53cdc),
	.w8(32'h38642dfb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38928a85),
	.w1(32'h38fb7e99),
	.w2(32'h38d987cc),
	.w3(32'h37f9f45c),
	.w4(32'h395c5d3c),
	.w5(32'h3891723a),
	.w6(32'h38618520),
	.w7(32'h38f6b6cc),
	.w8(32'h38a49510),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b5cf33),
	.w1(32'hb8bc4e30),
	.w2(32'hb897131e),
	.w3(32'h38171c11),
	.w4(32'hb8b608d3),
	.w5(32'hb8e39a06),
	.w6(32'hb622eef6),
	.w7(32'hb88a24e0),
	.w8(32'hb7dafc82),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb651a0e8),
	.w1(32'hb4f7b038),
	.w2(32'h34045446),
	.w3(32'hb52e98a2),
	.w4(32'hb5d3f6e6),
	.w5(32'hb5e353cb),
	.w6(32'hb3ba0950),
	.w7(32'hb5bdb323),
	.w8(32'hb5939d78),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34eaa8c4),
	.w1(32'hb5cf5291),
	.w2(32'hb60b6a1c),
	.w3(32'hb5a6885f),
	.w4(32'hb5562f86),
	.w5(32'hb607bf8f),
	.w6(32'hb61ea505),
	.w7(32'hb631f6ec),
	.w8(32'hb65bccaf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360d0434),
	.w1(32'h36074363),
	.w2(32'hb596f6e8),
	.w3(32'h360bdb5c),
	.w4(32'h3635a045),
	.w5(32'h3175a68c),
	.w6(32'hb446855a),
	.w7(32'hb50d0b06),
	.w8(32'hb624f200),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74ccb62),
	.w1(32'h3890db26),
	.w2(32'h373de429),
	.w3(32'hb75d2b7b),
	.w4(32'h384686fb),
	.w5(32'hb6a6aa2e),
	.w6(32'h3726945d),
	.w7(32'h381c7336),
	.w8(32'hb6dda7c4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356cf743),
	.w1(32'h34aac752),
	.w2(32'hb5a539a0),
	.w3(32'h35858023),
	.w4(32'hb57ef81c),
	.w5(32'hb620af97),
	.w6(32'hb5d96186),
	.w7(32'hb672bdc7),
	.w8(32'hb63b2aad),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361d2526),
	.w1(32'h38fc33e0),
	.w2(32'h391b0029),
	.w3(32'hb7c76b49),
	.w4(32'h37f1aa80),
	.w5(32'h392455b1),
	.w6(32'hb870c2bd),
	.w7(32'hb75dc2f5),
	.w8(32'h38bb9e80),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa41d6),
	.w1(32'h38ea5dc3),
	.w2(32'h3971a412),
	.w3(32'hb8857d06),
	.w4(32'hb7e39715),
	.w5(32'h398e5d12),
	.w6(32'hb8b81fc9),
	.w7(32'h37836c15),
	.w8(32'h38f4b1e2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73a95c2),
	.w1(32'hb8a1aa9d),
	.w2(32'hb81625b3),
	.w3(32'h3785aa66),
	.w4(32'hb8802808),
	.w5(32'hb8364a91),
	.w6(32'h377491e1),
	.w7(32'hb895aaad),
	.w8(32'hb850d965),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ec7aec),
	.w1(32'h38ad835e),
	.w2(32'h381efc2a),
	.w3(32'hb5ad21fe),
	.w4(32'h38a9e6ee),
	.w5(32'h3810c320),
	.w6(32'h37e0ac17),
	.w7(32'h37f62b2b),
	.w8(32'hb74ee914),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b0b55e),
	.w1(32'h389ce438),
	.w2(32'h38dd9431),
	.w3(32'hb839ba28),
	.w4(32'hb855a170),
	.w5(32'h38c17fb5),
	.w6(32'hb89feca4),
	.w7(32'hb714866b),
	.w8(32'h389ed1b4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f2e5f7),
	.w1(32'h37b51652),
	.w2(32'hb7c1c2b0),
	.w3(32'h376c681c),
	.w4(32'h37fac176),
	.w5(32'hb7bb6f66),
	.w6(32'h3802f06d),
	.w7(32'h35389826),
	.w8(32'hb7cb79e0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ac4c1),
	.w1(32'h386e0364),
	.w2(32'h38d5b6e8),
	.w3(32'hb7a56f6f),
	.w4(32'h37f549d6),
	.w5(32'h38d6c562),
	.w6(32'hb7067f45),
	.w7(32'h38289c55),
	.w8(32'h38b8a350),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369088ab),
	.w1(32'h3630424f),
	.w2(32'hb5153f46),
	.w3(32'h3587c605),
	.w4(32'h3610eae4),
	.w5(32'hb40b2957),
	.w6(32'hb531323d),
	.w7(32'hb57a58a1),
	.w8(32'hb68270c3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb623a61b),
	.w1(32'hb6141130),
	.w2(32'hb64e3b21),
	.w3(32'hb5fd68be),
	.w4(32'hb5d5ee12),
	.w5(32'hb6229424),
	.w6(32'hb60c97b6),
	.w7(32'hb625a307),
	.w8(32'hb454eb98),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5aef5cb),
	.w1(32'hb6ee4297),
	.w2(32'h35a87374),
	.w3(32'hb64b692a),
	.w4(32'hb6eed6e3),
	.w5(32'hb564739e),
	.w6(32'hb6e04370),
	.w7(32'h35018de6),
	.w8(32'hb4bfd753),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3599479b),
	.w1(32'hb715e2d5),
	.w2(32'hb6d89d44),
	.w3(32'h3629fbc0),
	.w4(32'hb6ba5fd8),
	.w5(32'hb65ef464),
	.w6(32'hb61ca563),
	.w7(32'hb6b17577),
	.w8(32'hb6d2bf1e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37207ec9),
	.w1(32'hb889ddb9),
	.w2(32'hb87ca432),
	.w3(32'h387365d8),
	.w4(32'hb7d5cec6),
	.w5(32'hb87de73a),
	.w6(32'h38207e28),
	.w7(32'hb8398b71),
	.w8(32'hb7e255c6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362a7985),
	.w1(32'hb6c5e4ba),
	.w2(32'hb730fa9e),
	.w3(32'h369b1361),
	.w4(32'hb67e4228),
	.w5(32'hb6d9ce5c),
	.w6(32'h35d95674),
	.w7(32'hb6d50195),
	.w8(32'hb750d139),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ba80f),
	.w1(32'hb8182aa0),
	.w2(32'hb75c306b),
	.w3(32'hb8177530),
	.w4(32'hb8c7f606),
	.w5(32'hb91d9063),
	.w6(32'h36afecbd),
	.w7(32'hb8bb8a26),
	.w8(32'hb8c0f6aa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385385ee),
	.w1(32'h394cf2e9),
	.w2(32'h39551469),
	.w3(32'h379a0a5f),
	.w4(32'h38fa93b4),
	.w5(32'h3948f7a4),
	.w6(32'h38813fd1),
	.w7(32'h39078060),
	.w8(32'h38fdf0dc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381c1911),
	.w1(32'hb7b31fe0),
	.w2(32'hb8825d4a),
	.w3(32'h383053ab),
	.w4(32'hb7bd02d4),
	.w5(32'hb7e10b16),
	.w6(32'hb7644e51),
	.w7(32'hb8099f64),
	.w8(32'hb81cfd1b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb798bc00),
	.w1(32'hb88c38dc),
	.w2(32'h394eaf79),
	.w3(32'hb9302d90),
	.w4(32'hb6eff4f1),
	.w5(32'h394b9486),
	.w6(32'hb96ced25),
	.w7(32'hb8b1bb17),
	.w8(32'h39116680),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ae9d04),
	.w1(32'hb7dc3220),
	.w2(32'hb7b952a3),
	.w3(32'h37e54e35),
	.w4(32'hb844b79d),
	.w5(32'hb7370f8f),
	.w6(32'h36c3a224),
	.w7(32'hb7716251),
	.w8(32'hb71b0e7c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d82cf1),
	.w1(32'h398a17cb),
	.w2(32'h38d057ab),
	.w3(32'hb8272cc6),
	.w4(32'h38e0fde0),
	.w5(32'hb84f20b8),
	.w6(32'h389f8e54),
	.w7(32'h3872db8f),
	.w8(32'hb84bb637),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb770b36a),
	.w1(32'h35a3c0ab),
	.w2(32'hb7adeb80),
	.w3(32'hb8a6b487),
	.w4(32'hb882cec8),
	.w5(32'hb7f84dfe),
	.w6(32'hb866c205),
	.w7(32'hb845325c),
	.w8(32'h3398e1a0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803b21b),
	.w1(32'h37769c84),
	.w2(32'hb80f93d4),
	.w3(32'h38482284),
	.w4(32'h37aaad63),
	.w5(32'hb7b9b6b9),
	.w6(32'h363b88b4),
	.w7(32'hb7c231e3),
	.w8(32'hb835a3c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73f3046),
	.w1(32'hb6cc5f22),
	.w2(32'h37be14a3),
	.w3(32'hb70f44f7),
	.w4(32'h37484cae),
	.w5(32'h37d04d22),
	.w6(32'hb5483745),
	.w7(32'h372d9cea),
	.w8(32'hb5700012),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d33c0a),
	.w1(32'h3897dbd6),
	.w2(32'h39123166),
	.w3(32'hb8298dd3),
	.w4(32'h38310626),
	.w5(32'h39001ee6),
	.w6(32'h383c86dd),
	.w7(32'h380c7a8d),
	.w8(32'h3819a741),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbbb51),
	.w1(32'h38879eef),
	.w2(32'h3898da2d),
	.w3(32'hb7f44d36),
	.w4(32'hb8c5d8da),
	.w5(32'h38e5fd20),
	.w6(32'hb8173487),
	.w7(32'hb86466d6),
	.w8(32'h38cdf927),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882f0d1),
	.w1(32'hb8f7cc53),
	.w2(32'h39e3bc0a),
	.w3(32'hb832afec),
	.w4(32'h369c333f),
	.w5(32'h39ed0793),
	.w6(32'hb8b37351),
	.w7(32'h386b0f5f),
	.w8(32'h399a2897),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382d651e),
	.w1(32'hb8db4193),
	.w2(32'hb7558ecb),
	.w3(32'h38c3bb84),
	.w4(32'hb904eec7),
	.w5(32'hb8ef65e7),
	.w6(32'h37a76bd7),
	.w7(32'hb96fd3ba),
	.w8(32'hb9486d2c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba2ba9),
	.w1(32'hb8c66ad8),
	.w2(32'hb832b33a),
	.w3(32'h36de9f8e),
	.w4(32'hb8cf6977),
	.w5(32'hb8b9260f),
	.w6(32'h3785878a),
	.w7(32'hb8ca4e7a),
	.w8(32'hb8d4e33d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859af71),
	.w1(32'hb841e1fa),
	.w2(32'h398b8557),
	.w3(32'hb7086109),
	.w4(32'hb89ca183),
	.w5(32'h39697715),
	.w6(32'hb8d82a33),
	.w7(32'h36089a93),
	.w8(32'h3950714f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ae35be),
	.w1(32'hb6f02a89),
	.w2(32'hb759e72c),
	.w3(32'hb6cd12e4),
	.w4(32'hb78db960),
	.w5(32'hb6b429d7),
	.w6(32'hb74e075e),
	.w7(32'hb7ec2320),
	.w8(32'hb776d55f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8916fa3),
	.w1(32'h38ec6e80),
	.w2(32'h3a047023),
	.w3(32'h38a446bd),
	.w4(32'h3873d8fa),
	.w5(32'h3a072158),
	.w6(32'hb834e86f),
	.w7(32'h37842394),
	.w8(32'h39c0d6b9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364a338a),
	.w1(32'hb8867d3f),
	.w2(32'hb623d5bc),
	.w3(32'hb8126514),
	.w4(32'hb8b6d0a4),
	.w5(32'h37769947),
	.w6(32'hb82d1a49),
	.w7(32'hb8e53466),
	.w8(32'h37b78d05),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65af585),
	.w1(32'hb5b5be5a),
	.w2(32'hb60a23cf),
	.w3(32'hb6c159a9),
	.w4(32'hb614ddd4),
	.w5(32'hb635a9cb),
	.w6(32'hb5a97905),
	.w7(32'h35c72b23),
	.w8(32'h3672a560),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381446b8),
	.w1(32'h3618301e),
	.w2(32'h376bbe78),
	.w3(32'h36a08692),
	.w4(32'h3857c41d),
	.w5(32'hb82452f0),
	.w6(32'hb7951ebd),
	.w7(32'h38354971),
	.w8(32'hb7e10bc8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7945367),
	.w1(32'h37c0c84f),
	.w2(32'h386cbd00),
	.w3(32'hb82735f5),
	.w4(32'h36931510),
	.w5(32'h36df39e4),
	.w6(32'hb639aa3a),
	.w7(32'hb7b182b7),
	.w8(32'hb8034a69),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818c8b9),
	.w1(32'hb8a9b918),
	.w2(32'hb7dcd605),
	.w3(32'hb6f6a5ed),
	.w4(32'hb8c11502),
	.w5(32'hb85e655c),
	.w6(32'hb7acfa74),
	.w7(32'hb8e0d648),
	.w8(32'hb8acb674),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3862213d),
	.w1(32'hb4e6b6ce),
	.w2(32'hb785a48c),
	.w3(32'h38a12232),
	.w4(32'h38507326),
	.w5(32'hb7a13c7d),
	.w6(32'hb702828a),
	.w7(32'hb88c2c2c),
	.w8(32'hb84a0f7a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d852a2),
	.w1(32'h3687a608),
	.w2(32'hb82bc24c),
	.w3(32'h388058c2),
	.w4(32'h38257f99),
	.w5(32'hb857c266),
	.w6(32'h38328111),
	.w7(32'h36339592),
	.w8(32'hb82533ef),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d0716),
	.w1(32'hb8ae27e0),
	.w2(32'h38a14ef9),
	.w3(32'hb830c46d),
	.w4(32'hb94ee810),
	.w5(32'h37cefc30),
	.w6(32'hb8169ba5),
	.w7(32'hb8646cf3),
	.w8(32'hb4f54770),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0a127),
	.w1(32'h391fef9a),
	.w2(32'h37c3d25d),
	.w3(32'hb8a113d5),
	.w4(32'h3903f883),
	.w5(32'hb7c8ea9c),
	.w6(32'h36340b46),
	.w7(32'h3685f884),
	.w8(32'hb81190f1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb780ac11),
	.w1(32'hb823db81),
	.w2(32'hb7ffbaba),
	.w3(32'h37216a74),
	.w4(32'hb8150483),
	.w5(32'hb83cedc9),
	.w6(32'h37e4de11),
	.w7(32'hb8221819),
	.w8(32'hb846100a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b9af50),
	.w1(32'h36339c28),
	.w2(32'h366c3e81),
	.w3(32'h357c0d40),
	.w4(32'h36e31651),
	.w5(32'h3725c2a0),
	.w6(32'h3600f6c2),
	.w7(32'h34e9931c),
	.w8(32'h3502688e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b5aa49),
	.w1(32'h36d8f770),
	.w2(32'hb794929d),
	.w3(32'h3614aeea),
	.w4(32'h36f54344),
	.w5(32'hb7925528),
	.w6(32'h36e934ab),
	.w7(32'hb6968409),
	.w8(32'hb7560e36),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb054b920),
	.w1(32'h34e0e90a),
	.w2(32'h351b8fc6),
	.w3(32'h350ee231),
	.w4(32'h35e54f32),
	.w5(32'h35fa6836),
	.w6(32'h358dd70b),
	.w7(32'h358b46c3),
	.w8(32'hb51f91fb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62d1897),
	.w1(32'hb65dd337),
	.w2(32'hb69e099b),
	.w3(32'hb740f1bc),
	.w4(32'hb706efd2),
	.w5(32'h3689640b),
	.w6(32'hb71bc5d7),
	.w7(32'hb648ec70),
	.w8(32'h360c914a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d0a13),
	.w1(32'hb80bb5e7),
	.w2(32'hb72533f6),
	.w3(32'hb7bbea13),
	.w4(32'hb87d1c34),
	.w5(32'hb867faf0),
	.w6(32'hb7cbc608),
	.w7(32'hb8a7cab5),
	.w8(32'hb83dff07),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb754201b),
	.w1(32'h3698c33d),
	.w2(32'hb6d982f8),
	.w3(32'hb75a1070),
	.w4(32'hb71a6609),
	.w5(32'h366cc9d5),
	.w6(32'hb4714f79),
	.w7(32'hb7479372),
	.w8(32'h36c0c386),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ac44cb),
	.w1(32'h3883ce0f),
	.w2(32'h3916e4b2),
	.w3(32'hb7f4fc37),
	.w4(32'h35862dc4),
	.w5(32'h38dff457),
	.w6(32'hb8204dc3),
	.w7(32'h3761b3f2),
	.w8(32'h38c8a466),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ac9262),
	.w1(32'hb870bee7),
	.w2(32'hb8adbb8f),
	.w3(32'h380fe79e),
	.w4(32'hb7e40915),
	.w5(32'hb8adcad7),
	.w6(32'hb739cc78),
	.w7(32'hb7725ad0),
	.w8(32'hb74330f4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6112897),
	.w1(32'hb680d5dd),
	.w2(32'hb69cf00b),
	.w3(32'hb44cade8),
	.w4(32'h358dd985),
	.w5(32'h35b074e4),
	.w6(32'h35bb4bb6),
	.w7(32'h3660c006),
	.w8(32'h35771f01),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f4ca37),
	.w1(32'hb68dcb23),
	.w2(32'hb6bc62c1),
	.w3(32'h35898748),
	.w4(32'hb5a12bea),
	.w5(32'hb5552151),
	.w6(32'hb5fd6e93),
	.w7(32'h3466918c),
	.w8(32'h2f661b80),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb059f81a),
	.w1(32'hb3b7432c),
	.w2(32'hb1aec879),
	.w3(32'h3518b0ed),
	.w4(32'h358f4dcf),
	.w5(32'h349e8c3e),
	.w6(32'hb5b2192a),
	.w7(32'h349d5343),
	.w8(32'h35864388),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb751dbc1),
	.w1(32'hbaf8046d),
	.w2(32'hbb97e70f),
	.w3(32'hb676b4d2),
	.w4(32'hba22d599),
	.w5(32'hbb3ea100),
	.w6(32'hbb06bf11),
	.w7(32'hbb4dbcb3),
	.w8(32'hba96153e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae68111),
	.w1(32'hb8eac8f1),
	.w2(32'hb9d251bb),
	.w3(32'hbb3933ea),
	.w4(32'hb8e99fba),
	.w5(32'h3a5d28d3),
	.w6(32'hba45875e),
	.w7(32'hbab1bf52),
	.w8(32'hbae1f038),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc5df2),
	.w1(32'hbb5c26b2),
	.w2(32'hbba11326),
	.w3(32'hba1c1c11),
	.w4(32'h3a63eb7d),
	.w5(32'h3b2ac307),
	.w6(32'hb98084fc),
	.w7(32'h3a31b4d7),
	.w8(32'h3b6e7a15),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79cad1),
	.w1(32'h39ab8ae2),
	.w2(32'hb955a041),
	.w3(32'h3b060e68),
	.w4(32'h39a639b4),
	.w5(32'hba322e89),
	.w6(32'h3a7c04ee),
	.w7(32'h3aab85f1),
	.w8(32'h3a98fe07),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b3d920),
	.w1(32'hb9de0215),
	.w2(32'hb9a8cc97),
	.w3(32'hb980fef1),
	.w4(32'hb91489ca),
	.w5(32'hba1e6439),
	.w6(32'hba328569),
	.w7(32'h37e06b0c),
	.w8(32'hba95fd92),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48ee5e),
	.w1(32'h3b1b7015),
	.w2(32'h39f2d58d),
	.w3(32'hba7f34fa),
	.w4(32'hb84e5213),
	.w5(32'hbb7e23c3),
	.w6(32'hb56d9903),
	.w7(32'hbaef63c6),
	.w8(32'hbb65b194),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aace753),
	.w1(32'hb9a3d1a3),
	.w2(32'h3a91c2ae),
	.w3(32'hbb1745fb),
	.w4(32'h3aaa098f),
	.w5(32'h3a90c725),
	.w6(32'hba515553),
	.w7(32'h3a40d03a),
	.w8(32'hba5eca68),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac687b9),
	.w1(32'h39bc95a9),
	.w2(32'hba7c6c92),
	.w3(32'h3a91a9dc),
	.w4(32'hb8c18f58),
	.w5(32'hb9ecf467),
	.w6(32'h3ac60b35),
	.w7(32'h3ab9d7d4),
	.w8(32'h3a9686ca),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c0a37),
	.w1(32'h39fa381b),
	.w2(32'h39a146f4),
	.w3(32'hbac7b028),
	.w4(32'h3918ca22),
	.w5(32'h38b19839),
	.w6(32'h3af5261d),
	.w7(32'h3adee66e),
	.w8(32'hb9f4574c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba279717),
	.w1(32'hb9d36884),
	.w2(32'hba3059bf),
	.w3(32'h3aa13f47),
	.w4(32'h3a790859),
	.w5(32'h3a8523ba),
	.w6(32'hb890cf07),
	.w7(32'hba1feb9f),
	.w8(32'hba8471de),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace8fb7),
	.w1(32'hb9d69456),
	.w2(32'hbb108c2f),
	.w3(32'h399ee667),
	.w4(32'hba049828),
	.w5(32'hbaded7dc),
	.w6(32'h38a8dcaf),
	.w7(32'hbae235f0),
	.w8(32'hbb331f06),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb374311),
	.w1(32'hb9b46ced),
	.w2(32'hba61806c),
	.w3(32'hbb1ec8f3),
	.w4(32'hb96a9635),
	.w5(32'hba951a77),
	.w6(32'h3ad5b517),
	.w7(32'h3b53fd6f),
	.w8(32'h3b0754d4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba721ad4),
	.w1(32'h3c4db37e),
	.w2(32'h3c879774),
	.w3(32'hba883b7c),
	.w4(32'h3a3f71e4),
	.w5(32'h3b8258e9),
	.w6(32'h3bc9e855),
	.w7(32'h3bc201b2),
	.w8(32'h3be3471b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87b7a2),
	.w1(32'h3a76001f),
	.w2(32'h3952c244),
	.w3(32'h3bfadb26),
	.w4(32'h3b01bd7c),
	.w5(32'h3aeab9d2),
	.w6(32'h3b512c79),
	.w7(32'h3b271e6f),
	.w8(32'h3aa023b1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abd39c),
	.w1(32'h3a791ac0),
	.w2(32'h3a357899),
	.w3(32'h3b09148e),
	.w4(32'hb9535428),
	.w5(32'h3977931f),
	.w6(32'hba762d49),
	.w7(32'hbb0523ba),
	.w8(32'hba4430eb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaeb87),
	.w1(32'h3a4a5e4c),
	.w2(32'h3965a439),
	.w3(32'h3a200c66),
	.w4(32'h3b27534c),
	.w5(32'h3ac85504),
	.w6(32'h3b4920dd),
	.w7(32'h3b593227),
	.w8(32'h3b122363),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998b29b),
	.w1(32'hb970a630),
	.w2(32'h3b6c20e2),
	.w3(32'h3a7d19fd),
	.w4(32'hb9a24716),
	.w5(32'h3aa9e8de),
	.w6(32'h3b1e7e6c),
	.w7(32'h3b721018),
	.w8(32'h3aa6df59),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87d24f),
	.w1(32'hb94823ea),
	.w2(32'hb9a89bc2),
	.w3(32'h3b2f0ad9),
	.w4(32'h3894e77e),
	.w5(32'h3a2e3843),
	.w6(32'h3942e417),
	.w7(32'hb947ddc3),
	.w8(32'hba789c15),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51f42d),
	.w1(32'hbae8c4d0),
	.w2(32'h39f2fc32),
	.w3(32'hb79c0769),
	.w4(32'hbac7e2af),
	.w5(32'hba2332c3),
	.w6(32'hbb885c96),
	.w7(32'hb9df3e23),
	.w8(32'hbb247991),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070259),
	.w1(32'h3a5032b7),
	.w2(32'h39010a5d),
	.w3(32'hbb1b6c95),
	.w4(32'hba0a345e),
	.w5(32'hbada840f),
	.w6(32'h3a80aeb3),
	.w7(32'h3a74525a),
	.w8(32'hb99d0a81),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c3338),
	.w1(32'h39782079),
	.w2(32'hb9cc86a6),
	.w3(32'hba257cae),
	.w4(32'hba1ded48),
	.w5(32'hba2b3645),
	.w6(32'hb9f12746),
	.w7(32'hba5583a7),
	.w8(32'hbae902c0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b340c),
	.w1(32'hba60865f),
	.w2(32'hbb05b4f9),
	.w3(32'hba85eb1e),
	.w4(32'hba9708c0),
	.w5(32'hbaf8172f),
	.w6(32'hb9d14c43),
	.w7(32'hba4ebde9),
	.w8(32'hbaeb8e76),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1cd09),
	.w1(32'hba515556),
	.w2(32'hbb3f719f),
	.w3(32'hbad75230),
	.w4(32'h3a828e9a),
	.w5(32'h39f4032e),
	.w6(32'h3a2c68ed),
	.w7(32'h3a2066a3),
	.w8(32'hba80cd84),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf41a7f),
	.w1(32'h3a16a58c),
	.w2(32'h3b23cea8),
	.w3(32'hb9f378f2),
	.w4(32'hbad2e0cb),
	.w5(32'h3a7a4f9f),
	.w6(32'h3aef190c),
	.w7(32'h3b319c7c),
	.w8(32'h3b3185f1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5cb72),
	.w1(32'h3c097dc0),
	.w2(32'h3c1ab620),
	.w3(32'h3b5a4aa8),
	.w4(32'h3b7ca1b2),
	.w5(32'h3bb7da1c),
	.w6(32'h3c30eaa8),
	.w7(32'h3c65f8ab),
	.w8(32'h3c3077c7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0244fd),
	.w1(32'hb939bac1),
	.w2(32'h38fdbed1),
	.w3(32'h3b59efbc),
	.w4(32'h393791c6),
	.w5(32'h3a864c36),
	.w6(32'hb7f4b465),
	.w7(32'hb9fe0cdf),
	.w8(32'hba6c78d8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f3157),
	.w1(32'h3a9c7c4c),
	.w2(32'h3a40f07a),
	.w3(32'h39571c9d),
	.w4(32'h39a85248),
	.w5(32'h3a0c82ec),
	.w6(32'h3a29dfc7),
	.w7(32'h394fbde7),
	.w8(32'hba6befe5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb855a068),
	.w1(32'hbb97e533),
	.w2(32'hbb55a78b),
	.w3(32'hba3843fb),
	.w4(32'hba5db52e),
	.w5(32'hbb25fbc1),
	.w6(32'hb9eff839),
	.w7(32'h3b5dec9f),
	.w8(32'h39a63211),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ab4c),
	.w1(32'hbabcbab9),
	.w2(32'hbb06dcd4),
	.w3(32'hbb2299cb),
	.w4(32'hbaef4021),
	.w5(32'hbb1544cb),
	.w6(32'hba3ee163),
	.w7(32'hb9b52205),
	.w8(32'hbaae12b2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6da93),
	.w1(32'hbadce2d7),
	.w2(32'hbae9ff66),
	.w3(32'hbab87795),
	.w4(32'hbb0b180f),
	.w5(32'hbb3188e5),
	.w6(32'hbaecbe4e),
	.w7(32'hba9d93cd),
	.w8(32'hbb381c3b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be2d1),
	.w1(32'h3b6b0f0b),
	.w2(32'h3b1b2166),
	.w3(32'hbb831612),
	.w4(32'h39e6893f),
	.w5(32'h3b2cbf9e),
	.w6(32'h3c278eb7),
	.w7(32'h3c51af8c),
	.w8(32'h3bf78b53),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac32210),
	.w1(32'h3aface7e),
	.w2(32'h3b353331),
	.w3(32'h39cf461c),
	.w4(32'h3b5513a8),
	.w5(32'h3b93422a),
	.w6(32'h3ad463fa),
	.w7(32'h3a81a90a),
	.w8(32'hbb5fdd81),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84d04e),
	.w1(32'hb9c25365),
	.w2(32'hba872444),
	.w3(32'hbb082abe),
	.w4(32'hba03e4fa),
	.w5(32'hb9d65845),
	.w6(32'hb9f8e16a),
	.w7(32'hb9ac9674),
	.w8(32'hb9db8de1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa3e87),
	.w1(32'hb8c1d696),
	.w2(32'hb83adde7),
	.w3(32'hba182e89),
	.w4(32'h3a155f32),
	.w5(32'h3a3bb2f1),
	.w6(32'h399c667d),
	.w7(32'h388cca84),
	.w8(32'hb9875f94),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a21f9f),
	.w1(32'hb79d42e4),
	.w2(32'h3ab3cca7),
	.w3(32'h3a0c8d66),
	.w4(32'hba54880a),
	.w5(32'h3a485020),
	.w6(32'h39b506fc),
	.w7(32'h3b62bfc8),
	.w8(32'h399f0436),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f8356),
	.w1(32'hbc168416),
	.w2(32'hbc0851eb),
	.w3(32'hbaebdc46),
	.w4(32'hbbcd1164),
	.w5(32'hbba57bbb),
	.w6(32'hbc010d1c),
	.w7(32'hbc0b3e4e),
	.w8(32'hb9dd227b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153783),
	.w1(32'h39dea1d5),
	.w2(32'hba5daec3),
	.w3(32'h3ac4f18a),
	.w4(32'hb9173069),
	.w5(32'hbb051fa2),
	.w6(32'h399f5485),
	.w7(32'h3a55bd7c),
	.w8(32'h39aa7a38),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c44170),
	.w1(32'hb975425b),
	.w2(32'hba76d374),
	.w3(32'hbac0d2b3),
	.w4(32'hbab5ae1b),
	.w5(32'hbaa37e89),
	.w6(32'h39d56b18),
	.w7(32'hb9f77658),
	.w8(32'hba0c8f67),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fcca3),
	.w1(32'h3a865473),
	.w2(32'h3af081a7),
	.w3(32'hb9d7e639),
	.w4(32'hbb0a5a1e),
	.w5(32'hbafdad52),
	.w6(32'hb9d72088),
	.w7(32'hb9b7d062),
	.w8(32'hbae5c6cf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a279dc),
	.w1(32'hb94fb01a),
	.w2(32'hba0018b5),
	.w3(32'hba2e784f),
	.w4(32'hb965aa68),
	.w5(32'hba3c86b1),
	.w6(32'h3af97148),
	.w7(32'h3b277e8e),
	.w8(32'h3b0bce72),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927a545),
	.w1(32'h37b2e9f6),
	.w2(32'hb8bd3744),
	.w3(32'h39ebe639),
	.w4(32'h39cc862b),
	.w5(32'h3a991228),
	.w6(32'hb7823f4d),
	.w7(32'hb9eb7fcb),
	.w8(32'hba9c2cb5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c93fb),
	.w1(32'hb8be8d7a),
	.w2(32'h39d23775),
	.w3(32'h395703a2),
	.w4(32'hb9ead295),
	.w5(32'hb967f648),
	.w6(32'h39fcbe97),
	.w7(32'h39225c36),
	.w8(32'hba5f312d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a976f),
	.w1(32'h3aa438c7),
	.w2(32'h3ba25d54),
	.w3(32'h39888f2f),
	.w4(32'h3b662c05),
	.w5(32'h3c0fa8ed),
	.w6(32'h3c07dcc6),
	.w7(32'h3c1f1fdf),
	.w8(32'h3adfb435),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920066),
	.w1(32'h3aa63b08),
	.w2(32'h3af929af),
	.w3(32'hba68780a),
	.w4(32'hb9f8a668),
	.w5(32'hba8abb70),
	.w6(32'h3b00222f),
	.w7(32'h3a602ef6),
	.w8(32'h39286fe9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eafca),
	.w1(32'hb84379bf),
	.w2(32'h389194fd),
	.w3(32'h3a0a2aa7),
	.w4(32'h3898e570),
	.w5(32'h39168a93),
	.w6(32'h3a66193b),
	.w7(32'h3a31a1e5),
	.w8(32'hba4acee5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39409966),
	.w1(32'h3a46c18c),
	.w2(32'hb9ad8efd),
	.w3(32'hb9098db5),
	.w4(32'hb8c7bc4d),
	.w5(32'hbb07ec56),
	.w6(32'h3b85deba),
	.w7(32'h3b77277b),
	.w8(32'h3b47c49d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b80b6),
	.w1(32'h3b1a396f),
	.w2(32'hbaa558f9),
	.w3(32'hba677891),
	.w4(32'h3a92ff25),
	.w5(32'hbb040e3e),
	.w6(32'h3a79aa36),
	.w7(32'h3a20a175),
	.w8(32'h3a47bc9d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd3ce1),
	.w1(32'hb9fdcbb9),
	.w2(32'hbb22196a),
	.w3(32'hb99b3f7e),
	.w4(32'hbaf8ed38),
	.w5(32'hbb2a45d0),
	.w6(32'hb9bc9ef4),
	.w7(32'hbab912fa),
	.w8(32'hbb26751b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae896ca),
	.w1(32'hbabfdb75),
	.w2(32'h3b21d359),
	.w3(32'hbaa998dc),
	.w4(32'h3ac59040),
	.w5(32'h3b05f86e),
	.w6(32'h3ad7cd8e),
	.w7(32'h3ae95f5a),
	.w8(32'hb9eac36b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc78b3),
	.w1(32'h3b78818f),
	.w2(32'hba538bd6),
	.w3(32'h3b2e2eb8),
	.w4(32'hb9990130),
	.w5(32'hbaeb65cc),
	.w6(32'h3b8e3ab8),
	.w7(32'h3aa4023d),
	.w8(32'h3b20f90f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192d23),
	.w1(32'hba155e7f),
	.w2(32'hb91a6d0d),
	.w3(32'hbb0d2efd),
	.w4(32'hba0d4575),
	.w5(32'hb9fb2d3c),
	.w6(32'h3a2dfff1),
	.w7(32'h3ac1119a),
	.w8(32'h3915d25b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3510f),
	.w1(32'h3990b495),
	.w2(32'h3a03ae54),
	.w3(32'h39334cf4),
	.w4(32'h3ab153e6),
	.w5(32'h3adf621d),
	.w6(32'h3a19981c),
	.w7(32'h39a21705),
	.w8(32'hb6a187e6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f09be7),
	.w1(32'h3a9d4134),
	.w2(32'h3af6c360),
	.w3(32'h3a9a478f),
	.w4(32'h3a99b51e),
	.w5(32'h394b3d7a),
	.w6(32'h3b130c54),
	.w7(32'h3b23081e),
	.w8(32'h3aea3776),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80a9e2),
	.w1(32'h3a152fd8),
	.w2(32'h3b00a380),
	.w3(32'h3ad91545),
	.w4(32'h3b095cd3),
	.w5(32'h3b94ea0f),
	.w6(32'h3a9b9199),
	.w7(32'hbac63cd0),
	.w8(32'h39ca053d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad03984),
	.w1(32'hb9074e06),
	.w2(32'hba457d25),
	.w3(32'h3ac106a0),
	.w4(32'hb989827b),
	.w5(32'hba044800),
	.w6(32'h3b5f02d7),
	.w7(32'h3b8bc33f),
	.w8(32'h3b735496),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1418ce),
	.w1(32'h388a6f7b),
	.w2(32'h399e8f36),
	.w3(32'hb91b504d),
	.w4(32'hb951dc06),
	.w5(32'hb8673f43),
	.w6(32'h3a265b50),
	.w7(32'h3a197166),
	.w8(32'hba821271),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf59fb),
	.w1(32'h3a855a2b),
	.w2(32'h3b27127f),
	.w3(32'h3aa23224),
	.w4(32'h3a79c12a),
	.w5(32'h3a887247),
	.w6(32'h3a98030b),
	.w7(32'h3ba34d6e),
	.w8(32'h3b7602d9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b5d0),
	.w1(32'h3b602a82),
	.w2(32'h3b1f8f9d),
	.w3(32'h39ab1e87),
	.w4(32'h3ba7681a),
	.w5(32'h3bf8c6fa),
	.w6(32'h3c659587),
	.w7(32'h3c24efa3),
	.w8(32'h3ba027b9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13122a),
	.w1(32'hbae93139),
	.w2(32'hb9efe891),
	.w3(32'h3af8b6c1),
	.w4(32'hb8bbbff8),
	.w5(32'hb8ef6d4d),
	.w6(32'h3b457e3a),
	.w7(32'h3bceea02),
	.w8(32'h3bb91bdb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1605f3),
	.w1(32'hbb0612b9),
	.w2(32'hb9fc98ed),
	.w3(32'hbaafbc3d),
	.w4(32'h3917c618),
	.w5(32'h3a57a2e1),
	.w6(32'hbaa6d22f),
	.w7(32'h39e7c183),
	.w8(32'h39f64231),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba755f42),
	.w1(32'h38a1e04e),
	.w2(32'hba26cd5b),
	.w3(32'h3a005bae),
	.w4(32'h3a034591),
	.w5(32'hb991fc24),
	.w6(32'h38d58ae0),
	.w7(32'h39ff213f),
	.w8(32'h3a1ae582),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12737a),
	.w1(32'h38e29c20),
	.w2(32'h37202549),
	.w3(32'hba563a2a),
	.w4(32'h3a11d99e),
	.w5(32'h3a9be529),
	.w6(32'hb928f2b2),
	.w7(32'hba29c67a),
	.w8(32'hbac6bfe7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9675f7),
	.w1(32'h3a37d87d),
	.w2(32'hb856e298),
	.w3(32'h3947df6b),
	.w4(32'h3a32ca44),
	.w5(32'hb9d20429),
	.w6(32'hb899ca0d),
	.w7(32'hb959ed71),
	.w8(32'hba77080d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1da030),
	.w1(32'h3a4a0bcc),
	.w2(32'h3ab89844),
	.w3(32'hba2caef6),
	.w4(32'h3a3beb1b),
	.w5(32'h3acf9dd0),
	.w6(32'h3a69266a),
	.w7(32'h3895fb17),
	.w8(32'hb9ff51ad),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9109da9),
	.w1(32'h3a3d4da6),
	.w2(32'hb97d8604),
	.w3(32'h3aae0aa8),
	.w4(32'hbac67041),
	.w5(32'hba6a1e3f),
	.w6(32'h3ae8d21b),
	.w7(32'h3b0648da),
	.w8(32'hba7441f0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e838),
	.w1(32'h3a1eee34),
	.w2(32'hb9107ea1),
	.w3(32'hbb706352),
	.w4(32'hb9c12225),
	.w5(32'hbad0e633),
	.w6(32'h3b21756a),
	.w7(32'h3b0e6c03),
	.w8(32'h3ae4f8b7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecee5d),
	.w1(32'hb9ef21d2),
	.w2(32'hb98851ca),
	.w3(32'hba567fc0),
	.w4(32'hbabf3525),
	.w5(32'hbaa4d110),
	.w6(32'hba3c5fca),
	.w7(32'hb8dc3195),
	.w8(32'hba77a189),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c7a3e),
	.w1(32'hbb6338d3),
	.w2(32'hbb34fa96),
	.w3(32'hbaf94f17),
	.w4(32'hba983cc3),
	.w5(32'hba916931),
	.w6(32'hbb9aabd6),
	.w7(32'hbb99ce2a),
	.w8(32'hbaa9ddb2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9831ed),
	.w1(32'hbad2c55a),
	.w2(32'h39964b8c),
	.w3(32'hb96e7724),
	.w4(32'h3a1c7d5e),
	.w5(32'h391224dd),
	.w6(32'h3b7eb439),
	.w7(32'h3b3cbb23),
	.w8(32'h3a97037a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb861080),
	.w1(32'hb8594398),
	.w2(32'h39b26f97),
	.w3(32'hbb58b549),
	.w4(32'h3a9c81f7),
	.w5(32'h3ba62d12),
	.w6(32'h3c421db2),
	.w7(32'h3c5119c8),
	.w8(32'h3c181150),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981f120),
	.w1(32'hb9df5e44),
	.w2(32'hba25b7af),
	.w3(32'h3b0a4d6a),
	.w4(32'hb8d61dfc),
	.w5(32'h3a046925),
	.w6(32'h3a249cd9),
	.w7(32'h3a52c1ed),
	.w8(32'hba87fbd8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa50959),
	.w1(32'hba26d4aa),
	.w2(32'hb86e64d4),
	.w3(32'hb9759650),
	.w4(32'hb8ca20d5),
	.w5(32'hba7d163f),
	.w6(32'hbb0712d7),
	.w7(32'hbb048b68),
	.w8(32'hbb112981),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfaa73),
	.w1(32'h3a301ace),
	.w2(32'hba019d4c),
	.w3(32'h3a2c3fd9),
	.w4(32'hba536075),
	.w5(32'hbb168f9b),
	.w6(32'h3a95386d),
	.w7(32'h3a18bcf0),
	.w8(32'h39732c38),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a9986),
	.w1(32'h39b36446),
	.w2(32'hb9fbf8d0),
	.w3(32'hbab35ae1),
	.w4(32'hb98ef2a2),
	.w5(32'hba0bf11b),
	.w6(32'h3a1252f9),
	.w7(32'h393b95df),
	.w8(32'hb97de697),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26a14a),
	.w1(32'h38907edb),
	.w2(32'hb941c2a1),
	.w3(32'hbaa89dca),
	.w4(32'h3979b4cc),
	.w5(32'h3a66dbaa),
	.w6(32'hb7d58203),
	.w7(32'hba08e1b9),
	.w8(32'hbaccb6df),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c714a),
	.w1(32'h3a377027),
	.w2(32'h383ed674),
	.w3(32'hb94836ac),
	.w4(32'hb9c65d65),
	.w5(32'hb8c5d19d),
	.w6(32'h3ac26971),
	.w7(32'h3a846810),
	.w8(32'h393c9445),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a563e),
	.w1(32'h37a300dc),
	.w2(32'h39f0f088),
	.w3(32'h39b53bd0),
	.w4(32'h3a03ccc6),
	.w5(32'hb8778126),
	.w6(32'hba7c4c0a),
	.w7(32'hba40d690),
	.w8(32'hba496f53),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b824d0),
	.w1(32'hbb6881bd),
	.w2(32'hbb65ce13),
	.w3(32'hba20e23a),
	.w4(32'hba962a96),
	.w5(32'hbac873b1),
	.w6(32'h3b2d63fa),
	.w7(32'h3af1b473),
	.w8(32'hbaf08a75),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77283d),
	.w1(32'hb9fbe459),
	.w2(32'hba6b5812),
	.w3(32'hba763e02),
	.w4(32'h39f82971),
	.w5(32'h3a675436),
	.w6(32'h3a6396ef),
	.w7(32'h3a3190a2),
	.w8(32'hb9aa9e7d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e5e4),
	.w1(32'h3a919e81),
	.w2(32'hbadb8087),
	.w3(32'hb94df825),
	.w4(32'h3a823d5d),
	.w5(32'hba9a5db0),
	.w6(32'hba07fc46),
	.w7(32'hbaf43076),
	.w8(32'hbaf4b708),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb709),
	.w1(32'h3a10dfb2),
	.w2(32'h3b1522ac),
	.w3(32'hbb2d9c99),
	.w4(32'h3a9189b1),
	.w5(32'h3ab0e682),
	.w6(32'hbb00fcb7),
	.w7(32'h3b652bdc),
	.w8(32'h3b17c8bf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9a1b9),
	.w1(32'hbb22404c),
	.w2(32'hbb8b06d7),
	.w3(32'h3b01d722),
	.w4(32'hbaca3b8a),
	.w5(32'hbb179417),
	.w6(32'hbaf3f750),
	.w7(32'hbae080fe),
	.w8(32'hbabfc79b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb088b6f),
	.w1(32'hbb357fa0),
	.w2(32'hbb012dd6),
	.w3(32'hbb1d0465),
	.w4(32'hb8da8a2b),
	.w5(32'h3b5498b0),
	.w6(32'h3c465d1d),
	.w7(32'h3c3c6933),
	.w8(32'h3c3ca21c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4f5d7),
	.w1(32'hba7f7635),
	.w2(32'hbaabc2eb),
	.w3(32'h3b1e4416),
	.w4(32'hb8b127d6),
	.w5(32'hbaac95b1),
	.w6(32'hb910f1c8),
	.w7(32'h3a0e0ba1),
	.w8(32'hb69a394e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82055a),
	.w1(32'h3b0d6abc),
	.w2(32'h3ac8ac5f),
	.w3(32'hba56c8da),
	.w4(32'h3924f56a),
	.w5(32'h39a5c938),
	.w6(32'h3b6a25bd),
	.w7(32'h3b490972),
	.w8(32'h3a5579aa),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb751bf7f),
	.w1(32'hba0700dc),
	.w2(32'hba91e2a3),
	.w3(32'hbab903e2),
	.w4(32'hb94a7737),
	.w5(32'hb9f1052d),
	.w6(32'h389c9ef0),
	.w7(32'h3a5d4982),
	.w8(32'h3a873e91),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba865d79),
	.w1(32'h3c4a77cc),
	.w2(32'h3c320081),
	.w3(32'hb9e4a715),
	.w4(32'hbb164f06),
	.w5(32'hba06fca5),
	.w6(32'h3c336942),
	.w7(32'h3c0e30b0),
	.w8(32'h3c91820a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4b32a),
	.w1(32'hbaa493eb),
	.w2(32'hbaa9d3af),
	.w3(32'h3bb87896),
	.w4(32'h3a978a59),
	.w5(32'h3918018d),
	.w6(32'hba41bcdd),
	.w7(32'h39511815),
	.w8(32'h3a55d355),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63682f),
	.w1(32'hb949a606),
	.w2(32'hbad6a9a8),
	.w3(32'h3a09fec0),
	.w4(32'h3a783c55),
	.w5(32'hba227778),
	.w6(32'h3aa03a1c),
	.w7(32'hba90e83e),
	.w8(32'hbabb8a73),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040a6f),
	.w1(32'hba144522),
	.w2(32'hbaa8abd0),
	.w3(32'hbaaf0f93),
	.w4(32'h390e0998),
	.w5(32'h3967a06f),
	.w6(32'hb7bd406f),
	.w7(32'h39518712),
	.w8(32'hba14aef5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71cec3),
	.w1(32'h3aff8add),
	.w2(32'h3b504e2c),
	.w3(32'hb9b6834e),
	.w4(32'h3abaa25c),
	.w5(32'h3aded664),
	.w6(32'h3b5a71df),
	.w7(32'h3bd2c992),
	.w8(32'h3bae0671),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48a1c1),
	.w1(32'hba7ebefd),
	.w2(32'hbac4bbb7),
	.w3(32'h3a670b15),
	.w4(32'h3a11bf35),
	.w5(32'h3a6e6276),
	.w6(32'h3a2fae35),
	.w7(32'h3a076cf4),
	.w8(32'hb8151fe8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba998d79),
	.w1(32'h3b19d71a),
	.w2(32'h3b1e47c8),
	.w3(32'hba564e45),
	.w4(32'h3adb1b64),
	.w5(32'h3b16055e),
	.w6(32'h3a6901cb),
	.w7(32'h3a6da6b1),
	.w8(32'hb96dc607),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f6ce),
	.w1(32'h399f825b),
	.w2(32'hb8a38878),
	.w3(32'h3aecadc4),
	.w4(32'hba7653cf),
	.w5(32'hbb089b63),
	.w6(32'h3b580541),
	.w7(32'h3b97bea9),
	.w8(32'h3b8a8451),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab0893),
	.w1(32'hba8d0e02),
	.w2(32'hbb04b223),
	.w3(32'hb966dd75),
	.w4(32'hbade07bc),
	.w5(32'hbb346e83),
	.w6(32'h3a49dd67),
	.w7(32'h3b01092d),
	.w8(32'h3b1b24db),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d0c5f),
	.w1(32'hbb2d5d3e),
	.w2(32'h3a14693b),
	.w3(32'hbb3afc44),
	.w4(32'hb8691c11),
	.w5(32'h3bd76c56),
	.w6(32'h3c830070),
	.w7(32'h3c9bafd2),
	.w8(32'h3c61133f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb5fec),
	.w1(32'h386887b0),
	.w2(32'h3a59a0fc),
	.w3(32'h3b464ba1),
	.w4(32'h3a1c5d6c),
	.w5(32'h3a2a1ee5),
	.w6(32'h39a80233),
	.w7(32'h3a800977),
	.w8(32'h37d37e72),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e4bae2),
	.w1(32'h3ab649eb),
	.w2(32'h398a100a),
	.w3(32'h39df4e4a),
	.w4(32'h3a8f7368),
	.w5(32'h3a9517fd),
	.w6(32'h3b37d595),
	.w7(32'h3a2a02d5),
	.w8(32'h3a6a3150),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38884aea),
	.w1(32'hb9939d35),
	.w2(32'h3a596b44),
	.w3(32'h3aacf3cf),
	.w4(32'h3af3ac7c),
	.w5(32'h3a842beb),
	.w6(32'hbae994d2),
	.w7(32'h3a3640db),
	.w8(32'h3a132ff6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acce53),
	.w1(32'hba8c32eb),
	.w2(32'hbb8df5b0),
	.w3(32'h3b15b4f0),
	.w4(32'hba002f5f),
	.w5(32'hbb49d2eb),
	.w6(32'hba953a7a),
	.w7(32'hbb53b2c5),
	.w8(32'hbb9eb4f9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e78b2),
	.w1(32'h3a171f16),
	.w2(32'h39698b91),
	.w3(32'hbbb72fdf),
	.w4(32'h39abce5b),
	.w5(32'hba0748e6),
	.w6(32'hba2ae9ec),
	.w7(32'hba038b55),
	.w8(32'hbaad5fe5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aef671),
	.w1(32'hba6483ee),
	.w2(32'hbb4b3b12),
	.w3(32'hba2377f6),
	.w4(32'hba870ca9),
	.w5(32'hbb366b8d),
	.w6(32'h3a4187bf),
	.w7(32'hb8c6e027),
	.w8(32'hb989ff05),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12849a),
	.w1(32'hbb469a5a),
	.w2(32'h3b0e057a),
	.w3(32'hbb594243),
	.w4(32'hbb6ccee2),
	.w5(32'hba985245),
	.w6(32'hba8f7445),
	.w7(32'h3b342586),
	.w8(32'hbaa95db2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aa7af),
	.w1(32'h3a9b74ff),
	.w2(32'h3b2231ea),
	.w3(32'hbb3ae7f8),
	.w4(32'h3ba431c6),
	.w5(32'h3ba45c98),
	.w6(32'hb9e5d29d),
	.w7(32'h3a84dab2),
	.w8(32'hba3df813),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5bd1),
	.w1(32'hba344214),
	.w2(32'hba86ff6b),
	.w3(32'h3b5af9e0),
	.w4(32'h3a4ed9ef),
	.w5(32'h3add23c3),
	.w6(32'h3a9bb84e),
	.w7(32'h3a9980c9),
	.w8(32'hb9478e8e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d7305),
	.w1(32'hba8b99f9),
	.w2(32'hbae0ae8d),
	.w3(32'hb98952bb),
	.w4(32'hb9854c7a),
	.w5(32'hba2ca19e),
	.w6(32'h39b29e71),
	.w7(32'h3a2ce82e),
	.w8(32'hb339d3e8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46387),
	.w1(32'hb93c291b),
	.w2(32'hba112b0a),
	.w3(32'hbaf4a99f),
	.w4(32'h399634f8),
	.w5(32'h3a2c9be1),
	.w6(32'h3a1cd4ac),
	.w7(32'h39c661ce),
	.w8(32'hb9d1895a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0edfe),
	.w1(32'hba74e26e),
	.w2(32'hbb300576),
	.w3(32'hb9a04450),
	.w4(32'hbae9064f),
	.w5(32'hbb240760),
	.w6(32'hb9339271),
	.w7(32'hba74a725),
	.w8(32'hbaf71a58),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17fcb9),
	.w1(32'h3aae0d58),
	.w2(32'h3ab9ff48),
	.w3(32'hbb0fbd7c),
	.w4(32'h3980281f),
	.w5(32'h39b54008),
	.w6(32'h37dba05d),
	.w7(32'h38ee2498),
	.w8(32'h392aa32c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfcd5e),
	.w1(32'h3b1549a3),
	.w2(32'h3acd6deb),
	.w3(32'h3a749e09),
	.w4(32'h3b028b03),
	.w5(32'h3b1138f0),
	.w6(32'h3a566bda),
	.w7(32'h3a994adf),
	.w8(32'hba2e5d5e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a970ebf),
	.w1(32'hb9d0e902),
	.w2(32'hba4be27b),
	.w3(32'h3ac95060),
	.w4(32'h3a01bacf),
	.w5(32'h3a3bf352),
	.w6(32'h3a407fce),
	.w7(32'h3a21aad1),
	.w8(32'hb94185ac),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8cfac),
	.w1(32'h3ac8aa47),
	.w2(32'h397cfa44),
	.w3(32'hb7a5572a),
	.w4(32'h3ac67044),
	.w5(32'hb99cae17),
	.w6(32'hb91c9f94),
	.w7(32'h3ab211d1),
	.w8(32'h3acda25d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cf4d2),
	.w1(32'hba81a50c),
	.w2(32'hba17daa0),
	.w3(32'h390d8bd1),
	.w4(32'hb98e93ee),
	.w5(32'h3aab73e8),
	.w6(32'h3a0d4286),
	.w7(32'hb9b535ae),
	.w8(32'hbaf1acbe),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc05f1),
	.w1(32'hba68b6cc),
	.w2(32'hbb08cedd),
	.w3(32'h39da3b04),
	.w4(32'h3a0a39a5),
	.w5(32'h3b3494cf),
	.w6(32'h3904a0a3),
	.w7(32'hba1d6151),
	.w8(32'hba714477),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022722),
	.w1(32'hb9815a73),
	.w2(32'hb90956fd),
	.w3(32'hba73651c),
	.w4(32'hb99465ad),
	.w5(32'h3a5d78b8),
	.w6(32'h39553309),
	.w7(32'hba56fcc7),
	.w8(32'hba846d63),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12686f),
	.w1(32'h3ac14acf),
	.w2(32'h3aead695),
	.w3(32'h38c3b58d),
	.w4(32'h3a82292a),
	.w5(32'h394e84da),
	.w6(32'hb90db24a),
	.w7(32'hb9887baa),
	.w8(32'hb790aaf8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6826e),
	.w1(32'hbacb22ea),
	.w2(32'hba11b19b),
	.w3(32'hba12b9fa),
	.w4(32'hba9f2bbd),
	.w5(32'hb9fd4ac6),
	.w6(32'h3ab61405),
	.w7(32'h3b0a3a3a),
	.w8(32'h3ab12da4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39709d92),
	.w1(32'hb9f9a941),
	.w2(32'hba804bbd),
	.w3(32'h3904760b),
	.w4(32'h3a1b46b2),
	.w5(32'h3a8affd6),
	.w6(32'h3a7b1873),
	.w7(32'h3a592523),
	.w8(32'hb9b548e1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14bccf),
	.w1(32'h3a4c48c1),
	.w2(32'h37782413),
	.w3(32'hb9627267),
	.w4(32'hb8b14257),
	.w5(32'hb91db904),
	.w6(32'h395d5529),
	.w7(32'hba0724f9),
	.w8(32'hba9cebd5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af4215),
	.w1(32'h3a329144),
	.w2(32'hb9fd13e4),
	.w3(32'hba487c26),
	.w4(32'hb7f27ee9),
	.w5(32'hb903402c),
	.w6(32'hb9c7b6d1),
	.w7(32'hba9c1ab1),
	.w8(32'hbad67fc3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ecd40),
	.w1(32'h3b1ca208),
	.w2(32'h3abd9445),
	.w3(32'hba4a81c6),
	.w4(32'h3973d930),
	.w5(32'h38ecfb75),
	.w6(32'hbab962ba),
	.w7(32'hbb06a257),
	.w8(32'hbafd8573),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a3e99),
	.w1(32'hba7ecd6e),
	.w2(32'hbb64c5f6),
	.w3(32'h3a3808d3),
	.w4(32'hbb365733),
	.w5(32'hbb7b3c45),
	.w6(32'hba0e3e9c),
	.w7(32'hbb375620),
	.w8(32'hbb8da44e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e0c8),
	.w1(32'h3a345cbf),
	.w2(32'hba885cf8),
	.w3(32'hbb2d5b12),
	.w4(32'hbab46e3b),
	.w5(32'hbb2cbd2d),
	.w6(32'h3ac98fce),
	.w7(32'h383e6610),
	.w8(32'h3a3b94de),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa94f3e),
	.w1(32'h3a581ef8),
	.w2(32'hba29c374),
	.w3(32'hba7b417b),
	.w4(32'h38e72556),
	.w5(32'hba837eb6),
	.w6(32'h39e1f605),
	.w7(32'hbad54966),
	.w8(32'hbaf78526),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba498e92),
	.w1(32'hb9049315),
	.w2(32'h3782d341),
	.w3(32'hba1c4cac),
	.w4(32'h39cde1dc),
	.w5(32'h3a835022),
	.w6(32'hb918dd44),
	.w7(32'hba12c4c5),
	.w8(32'hba918165),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9632fa),
	.w1(32'hbaae6418),
	.w2(32'hbb66dee4),
	.w3(32'h38fea6fd),
	.w4(32'h3b211114),
	.w5(32'h3a976c8a),
	.w6(32'h3a612095),
	.w7(32'h3ae5ee46),
	.w8(32'h3af131bf),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934e9c),
	.w1(32'hba3a5609),
	.w2(32'hbb246d91),
	.w3(32'h3b26a11e),
	.w4(32'hbae4cd24),
	.w5(32'hbb5174c7),
	.w6(32'h3b30f9ca),
	.w7(32'h3b3c629a),
	.w8(32'h3b7cf417),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83894bf),
	.w1(32'hb8447948),
	.w2(32'hbb2fc370),
	.w3(32'hbaf07693),
	.w4(32'hba6817b6),
	.w5(32'hbb00ac08),
	.w6(32'hba434152),
	.w7(32'hbb058a07),
	.w8(32'hbb0e9750),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27c2b3),
	.w1(32'h37591c5d),
	.w2(32'h372f9fea),
	.w3(32'hba471a83),
	.w4(32'h37262adc),
	.w5(32'h36eec725),
	.w6(32'hb566ebe6),
	.w7(32'h371647ab),
	.w8(32'h34a2924c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d1f4b5),
	.w1(32'hb86dccae),
	.w2(32'h38d3a3ed),
	.w3(32'h3807bbc2),
	.w4(32'hb902aace),
	.w5(32'hb897c795),
	.w6(32'h38acd68a),
	.w7(32'h368c204e),
	.w8(32'hb8755e4a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule