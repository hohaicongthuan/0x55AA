module layer_10_featuremap_49(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d11b59a),
	.w1(32'hba4dcf6d),
	.w2(32'h3b85af21),
	.w3(32'h3d127571),
	.w4(32'h3d031643),
	.w5(32'h3c622d2d),
	.w6(32'h3c0cbbd0),
	.w7(32'h3d04da25),
	.w8(32'h3c145787),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60c149),
	.w1(32'h3c985e25),
	.w2(32'hbb461bf0),
	.w3(32'h3c0de2af),
	.w4(32'h3af2515e),
	.w5(32'hbb7d6ce3),
	.w6(32'h3c653361),
	.w7(32'h39afb65a),
	.w8(32'h3a4eb7d6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58c23f),
	.w1(32'h3b1451ae),
	.w2(32'hbc79af6e),
	.w3(32'hbc0ba9bf),
	.w4(32'hbba42b2c),
	.w5(32'hbc0eac43),
	.w6(32'hbba6f686),
	.w7(32'hbbb16d41),
	.w8(32'hbc05ba78),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc438e20),
	.w1(32'hbb34ddc2),
	.w2(32'hbb885d31),
	.w3(32'hbc8e65d2),
	.w4(32'hbc71f925),
	.w5(32'hb9f04072),
	.w6(32'hbb55903a),
	.w7(32'hbb76b266),
	.w8(32'hbaccc97d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8475ba),
	.w1(32'h3b874c49),
	.w2(32'hbc086ba5),
	.w3(32'hbb8d2337),
	.w4(32'hbbdbaec6),
	.w5(32'hbc329e90),
	.w6(32'h3ac6f5a1),
	.w7(32'h39655145),
	.w8(32'hbbf4deba),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8405c9),
	.w1(32'hb9f6395a),
	.w2(32'h3a4aa79f),
	.w3(32'hbc81f2bb),
	.w4(32'hbba30e91),
	.w5(32'hb94bd3b3),
	.w6(32'hbc9123b8),
	.w7(32'hbbaa6650),
	.w8(32'h39da52eb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ead8),
	.w1(32'hbc06822b),
	.w2(32'hbb2f3908),
	.w3(32'hbbe44d25),
	.w4(32'hbbe9c841),
	.w5(32'h3a0eed9d),
	.w6(32'hba3d17ec),
	.w7(32'hbb04835c),
	.w8(32'h3ba210c5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab226c),
	.w1(32'h3b42c103),
	.w2(32'h3c2faded),
	.w3(32'h3c1f1587),
	.w4(32'h3c2f2bbb),
	.w5(32'hbc2e0389),
	.w6(32'h3ca0ac71),
	.w7(32'hba3ee51c),
	.w8(32'h3b6e381c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147604),
	.w1(32'hbb48d203),
	.w2(32'h3c312315),
	.w3(32'h3b553947),
	.w4(32'h3c1fe965),
	.w5(32'h3c7982c3),
	.w6(32'hbcabfd41),
	.w7(32'hbb494363),
	.w8(32'h3c5a5360),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2951c3),
	.w1(32'h3c228a9f),
	.w2(32'hbb27c3ff),
	.w3(32'h3c9fb557),
	.w4(32'h3c536209),
	.w5(32'hbb7cf87c),
	.w6(32'h3cc83aee),
	.w7(32'h3cd8d386),
	.w8(32'h3b92794d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fabfe),
	.w1(32'h3b47ecf1),
	.w2(32'hbc0bd1fb),
	.w3(32'hbacb21b4),
	.w4(32'h3a4fdcb2),
	.w5(32'hbc17d126),
	.w6(32'h3b280b4c),
	.w7(32'h3ab0c122),
	.w8(32'h3bd5196d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10509d),
	.w1(32'h3b303681),
	.w2(32'hbc1da631),
	.w3(32'hbc5a58fe),
	.w4(32'hbb404ff7),
	.w5(32'hbc2a060e),
	.w6(32'hbb58c0a6),
	.w7(32'hbb823a2c),
	.w8(32'h38631467),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b3cb5),
	.w1(32'hbae6b6ec),
	.w2(32'h3c423043),
	.w3(32'hbbf4be1c),
	.w4(32'hbb9afae7),
	.w5(32'h3c40e607),
	.w6(32'hb94cb299),
	.w7(32'hbb4359f3),
	.w8(32'h3c7eef5b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe421d),
	.w1(32'h3b544bdf),
	.w2(32'hba610d05),
	.w3(32'h3c10f352),
	.w4(32'h3c0d5869),
	.w5(32'hbb41fa86),
	.w6(32'h3c735a86),
	.w7(32'h3c3cfc27),
	.w8(32'h3bf4dc12),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29bd4e),
	.w1(32'h3b635e23),
	.w2(32'hb9796533),
	.w3(32'hbc8025a4),
	.w4(32'hbc72826d),
	.w5(32'h3be31f64),
	.w6(32'hbb88596c),
	.w7(32'hbb9798c9),
	.w8(32'h38b5f731),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aba1e),
	.w1(32'h3bd65263),
	.w2(32'hbaa47b10),
	.w3(32'hba24ecdc),
	.w4(32'hbc19d49d),
	.w5(32'h3ae76176),
	.w6(32'h3c230a06),
	.w7(32'h3b54c1e6),
	.w8(32'h3b8748ca),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b145811),
	.w1(32'h3b8f9338),
	.w2(32'hbc25519c),
	.w3(32'h38cdc5c3),
	.w4(32'h3b4018c4),
	.w5(32'hbc22bc39),
	.w6(32'h3b20fd44),
	.w7(32'h3a9b9f07),
	.w8(32'hb96d91bc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae20e4),
	.w1(32'hbba19ef2),
	.w2(32'h3be7c909),
	.w3(32'hbbc92998),
	.w4(32'hbb2bd8c4),
	.w5(32'h3b40f24c),
	.w6(32'h39c46a9a),
	.w7(32'h3be8cbc8),
	.w8(32'h3c166184),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7df18),
	.w1(32'h3b532185),
	.w2(32'hbb6002a0),
	.w3(32'h3b924c64),
	.w4(32'h3b8017e4),
	.w5(32'h3c86a5e0),
	.w6(32'hba3d9fe3),
	.w7(32'h3bed862a),
	.w8(32'h3cf63391),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f37e2),
	.w1(32'h3ce1000e),
	.w2(32'hbc050bda),
	.w3(32'h3babea4d),
	.w4(32'h3c8f9071),
	.w5(32'hbb9a4a56),
	.w6(32'h3cd2d113),
	.w7(32'h3a732a68),
	.w8(32'h3a6af9c7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f1f31),
	.w1(32'h3bd33b0b),
	.w2(32'h399c0e62),
	.w3(32'hbad46110),
	.w4(32'h3b0a61ab),
	.w5(32'h3c0ffd52),
	.w6(32'h3b91d857),
	.w7(32'h3aad66cb),
	.w8(32'hbbc55fe0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a06d),
	.w1(32'h3c00429e),
	.w2(32'hbb78674d),
	.w3(32'h3c0805d0),
	.w4(32'h3b145de7),
	.w5(32'hbb5713b5),
	.w6(32'h3c0e234d),
	.w7(32'h3bc85ca9),
	.w8(32'h3a961287),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06718),
	.w1(32'h3bd3d4f7),
	.w2(32'hbc21778e),
	.w3(32'h3ae3fbf9),
	.w4(32'h3a9031a1),
	.w5(32'hba8b0e40),
	.w6(32'h3b3a55ee),
	.w7(32'hbb7d88ec),
	.w8(32'hbb8c5845),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bf4d8),
	.w1(32'h3b846903),
	.w2(32'h3c0ae86b),
	.w3(32'hbc5d5d22),
	.w4(32'hbbc27d20),
	.w5(32'h3c024492),
	.w6(32'hbb851931),
	.w7(32'hbb3f4f63),
	.w8(32'h3c35b844),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8e2d),
	.w1(32'h3c3eae72),
	.w2(32'hbc037c26),
	.w3(32'h3bb516d7),
	.w4(32'h3c218c78),
	.w5(32'hbc982d91),
	.w6(32'hbb8d1905),
	.w7(32'h3c31326c),
	.w8(32'hbc7029d8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e26971),
	.w1(32'h3c02652f),
	.w2(32'hba66958e),
	.w3(32'h3b2a57d2),
	.w4(32'h3ba73c8b),
	.w5(32'hbbf6de74),
	.w6(32'hbcca5d2e),
	.w7(32'h3a98b871),
	.w8(32'hbb0d7c72),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae2d62),
	.w1(32'hba90f7bb),
	.w2(32'hbb0a95fc),
	.w3(32'hbbb3e8b7),
	.w4(32'hbbef99a0),
	.w5(32'h39b9145d),
	.w6(32'h3b3169a2),
	.w7(32'hbb15ba60),
	.w8(32'hbad7de47),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391af592),
	.w1(32'h3b394e4c),
	.w2(32'h3bc4b2ee),
	.w3(32'hba031a9c),
	.w4(32'h3b17046d),
	.w5(32'h3c11ee0b),
	.w6(32'hba2d90dd),
	.w7(32'h3be3e5a0),
	.w8(32'h3c0bd838),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98dbbd),
	.w1(32'h3a8e83e4),
	.w2(32'h3a84702b),
	.w3(32'hbc001fe2),
	.w4(32'hbb732c1b),
	.w5(32'hbae8a80e),
	.w6(32'hbbc3b0c8),
	.w7(32'h3b190a7a),
	.w8(32'h3bca53e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c3ed1),
	.w1(32'h3b011681),
	.w2(32'h3c8af333),
	.w3(32'hbb9795db),
	.w4(32'h3a4f0673),
	.w5(32'h3ae53afa),
	.w6(32'hbb74ad10),
	.w7(32'hbad5f321),
	.w8(32'h3c122668),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9500f),
	.w1(32'h3c2d0db0),
	.w2(32'hbb5e489c),
	.w3(32'hbc4f35d3),
	.w4(32'hbb9e5a45),
	.w5(32'hbac5f427),
	.w6(32'hbb1284f5),
	.w7(32'h3b9272b8),
	.w8(32'h3b555e62),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc274e),
	.w1(32'h3aef1744),
	.w2(32'hbb0fa969),
	.w3(32'h3bcbe083),
	.w4(32'hba3da0f5),
	.w5(32'h3a742d39),
	.w6(32'h3b5bb1d9),
	.w7(32'hbbcda528),
	.w8(32'h3c028bc2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6278df),
	.w1(32'h3b63a952),
	.w2(32'hbc3834ac),
	.w3(32'h3b3641cf),
	.w4(32'h3b80d652),
	.w5(32'hbd121386),
	.w6(32'h3c4a87c6),
	.w7(32'h3c2cfa5a),
	.w8(32'hbcb1a63d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1441d6),
	.w1(32'hbc921596),
	.w2(32'hb93a1bb6),
	.w3(32'hbd9b78f8),
	.w4(32'hbd53409b),
	.w5(32'hbb333f17),
	.w6(32'hbd7019fe),
	.w7(32'hbd1a529e),
	.w8(32'hbbb1c391),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59dce5),
	.w1(32'h3a899475),
	.w2(32'hbbfbf4c2),
	.w3(32'hbc0db186),
	.w4(32'hb9524ac9),
	.w5(32'hbb88bc5f),
	.w6(32'hbc0d00db),
	.w7(32'h3aef9f59),
	.w8(32'hbbb720d2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64a08e),
	.w1(32'hbc2f8c2e),
	.w2(32'hbbd04afa),
	.w3(32'h3c0b54f8),
	.w4(32'hbb07fa63),
	.w5(32'h3b137fc0),
	.w6(32'h3ba07dde),
	.w7(32'hbba999a9),
	.w8(32'h3bb5324c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2931),
	.w1(32'h3bc5d4aa),
	.w2(32'hbcfabf6b),
	.w3(32'hbc605756),
	.w4(32'hb9425b1d),
	.w5(32'hbd7a272a),
	.w6(32'hb81a77f4),
	.w7(32'hbc980098),
	.w8(32'hbd2e9f23),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd31c404),
	.w1(32'hbc9eb6e6),
	.w2(32'h3c42ea3e),
	.w3(32'hbdb10e2f),
	.w4(32'hbd58c8d0),
	.w5(32'h3ab812b7),
	.w6(32'hbd8edecf),
	.w7(32'hbd27836a),
	.w8(32'h3c022864),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7838fc),
	.w1(32'h3c1d7484),
	.w2(32'h3b80c759),
	.w3(32'hbc1ad436),
	.w4(32'h39f3a779),
	.w5(32'h3b5c0ce0),
	.w6(32'hbc27cb69),
	.w7(32'h3bb476a4),
	.w8(32'h3b0e35e4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc747e4),
	.w1(32'h3b244c05),
	.w2(32'h395d560c),
	.w3(32'h3c2100c1),
	.w4(32'h3b522413),
	.w5(32'h3b2ca93a),
	.w6(32'h3bc5630b),
	.w7(32'h3b1995d2),
	.w8(32'h395de181),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb083441),
	.w1(32'hbb9349b9),
	.w2(32'hbbe58680),
	.w3(32'h3b229964),
	.w4(32'hbb24209a),
	.w5(32'hba28a384),
	.w6(32'h3a227571),
	.w7(32'hbac41774),
	.w8(32'hbb165062),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b029025),
	.w1(32'h3b65371c),
	.w2(32'h38055709),
	.w3(32'hba9615ec),
	.w4(32'h3b0c6e3d),
	.w5(32'h399e49ff),
	.w6(32'hbbed2b14),
	.w7(32'hbacd9cfd),
	.w8(32'h3a645790),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37cef6),
	.w1(32'h39fa4a51),
	.w2(32'hbc8e39ff),
	.w3(32'h3afac846),
	.w4(32'h38f2c449),
	.w5(32'hbb87674a),
	.w6(32'h3a771348),
	.w7(32'h3ba94849),
	.w8(32'hbc3b27c9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9eef0),
	.w1(32'hbca1581b),
	.w2(32'h3bfd5f9b),
	.w3(32'h3c83b637),
	.w4(32'h3b9f117c),
	.w5(32'h3c246dbe),
	.w6(32'h3bebcffe),
	.w7(32'hbab9272d),
	.w8(32'h3a915a7a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dc0a5),
	.w1(32'h3bb313f3),
	.w2(32'h3afa337d),
	.w3(32'hbaeab923),
	.w4(32'h3c4d4c4d),
	.w5(32'h3bc27fbe),
	.w6(32'h3ad459a8),
	.w7(32'h3bd48e25),
	.w8(32'h3b941978),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0cd54),
	.w1(32'h3c0d5d09),
	.w2(32'h3c18e1f2),
	.w3(32'h3ba73bca),
	.w4(32'h3c2351d9),
	.w5(32'h3c201bc6),
	.w6(32'hbab2a61e),
	.w7(32'h3ba28e0f),
	.w8(32'h3a9361e3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b136f81),
	.w1(32'h3be218e7),
	.w2(32'h3c4379cf),
	.w3(32'h3b578a81),
	.w4(32'h3c0d8aeb),
	.w5(32'h3c22ac9f),
	.w6(32'h3bac5c6a),
	.w7(32'h3c22e4f0),
	.w8(32'h3bcc85fe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5192d),
	.w1(32'h3b73e19b),
	.w2(32'hbd073ea1),
	.w3(32'h3c5618f1),
	.w4(32'h3c09d88d),
	.w5(32'hbca458a1),
	.w6(32'h3ca3140a),
	.w7(32'h3c3e0456),
	.w8(32'hbcbe5f55),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc815e84),
	.w1(32'hbcc7bb3a),
	.w2(32'hba05adc7),
	.w3(32'h3b6a9ecc),
	.w4(32'hbc0d6176),
	.w5(32'hba3db2c1),
	.w6(32'hbc0aa12f),
	.w7(32'hbca22d24),
	.w8(32'h3b96892f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891399),
	.w1(32'hb992b44b),
	.w2(32'h3a9c34c0),
	.w3(32'hbb9e803c),
	.w4(32'hbbffff63),
	.w5(32'hba89548b),
	.w6(32'hbb881707),
	.w7(32'hbb915fda),
	.w8(32'h3b80d552),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a4d48),
	.w1(32'h3b332952),
	.w2(32'h3b2d45f1),
	.w3(32'hba3ed68a),
	.w4(32'hba18a6ad),
	.w5(32'hb85b5b66),
	.w6(32'hbb044ee8),
	.w7(32'h3b3d653d),
	.w8(32'h3b5d5f6e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12032a),
	.w1(32'h3b7d0c25),
	.w2(32'hbb7e0bbd),
	.w3(32'h3bf93e7e),
	.w4(32'h3b768f87),
	.w5(32'hbad34cd2),
	.w6(32'h3b5be9bc),
	.w7(32'h39d94e94),
	.w8(32'h3a915b97),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1192ce),
	.w1(32'hbb7caa10),
	.w2(32'h3b4ac3da),
	.w3(32'h3ac7933b),
	.w4(32'h3bfa6ed6),
	.w5(32'h3bb6d785),
	.w6(32'h3baeb695),
	.w7(32'hbb83588d),
	.w8(32'h3be52687),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ead11),
	.w1(32'hbb4d61f0),
	.w2(32'hbabdd129),
	.w3(32'h3b224995),
	.w4(32'h3b5a72b5),
	.w5(32'hbae6558f),
	.w6(32'h3c6da0ef),
	.w7(32'h3c6a8c35),
	.w8(32'h3bf0d841),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29b681),
	.w1(32'hbb4ead83),
	.w2(32'hb9f0d1fa),
	.w3(32'hbb963fbe),
	.w4(32'hb99f257e),
	.w5(32'hbad33233),
	.w6(32'h3b51b237),
	.w7(32'h3b179778),
	.w8(32'h3a4798a8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00fd37),
	.w1(32'hbb02d46d),
	.w2(32'hbb5082f4),
	.w3(32'hba3f6c20),
	.w4(32'h3b6467c2),
	.w5(32'h3be3cad4),
	.w6(32'h3b6b531b),
	.w7(32'h3a9888aa),
	.w8(32'h3c39f95d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b378072),
	.w1(32'h3bfd787c),
	.w2(32'h3bc5718e),
	.w3(32'h3997128c),
	.w4(32'hb9f97dc6),
	.w5(32'h3bf7491d),
	.w6(32'h3b89cc6a),
	.w7(32'h3b49939b),
	.w8(32'h3b9ad8ed),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f60f51),
	.w1(32'hbbe2a5c1),
	.w2(32'hba9da687),
	.w3(32'hba81b405),
	.w4(32'hbc2011ee),
	.w5(32'hbb4d3bf3),
	.w6(32'hba9239a0),
	.w7(32'hbbf9fefd),
	.w8(32'hbb599223),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20523),
	.w1(32'h3b245a52),
	.w2(32'h3aa3881a),
	.w3(32'hbb7dbdc7),
	.w4(32'h3a94d396),
	.w5(32'h3b2cd0f8),
	.w6(32'h3a6a88cc),
	.w7(32'h3bb835f3),
	.w8(32'h3ab77180),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc03329),
	.w1(32'h3adc1fe0),
	.w2(32'h3b6aa459),
	.w3(32'h3b80e94c),
	.w4(32'h3b5076f7),
	.w5(32'h3a7c7197),
	.w6(32'hbb2da50a),
	.w7(32'hbb444015),
	.w8(32'hbb2b429a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54d9d7),
	.w1(32'hbbb37f03),
	.w2(32'h3a98255f),
	.w3(32'h3b0edcd2),
	.w4(32'hbbc93173),
	.w5(32'hb99a55f4),
	.w6(32'hbbaf8ec7),
	.w7(32'hbbca88de),
	.w8(32'h3b04a7d4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48e32),
	.w1(32'h3b64d519),
	.w2(32'h3a583a29),
	.w3(32'hbb4d068c),
	.w4(32'hba587cf5),
	.w5(32'hbbc362fa),
	.w6(32'hbb70b86f),
	.w7(32'hb985cc2c),
	.w8(32'hbb88fc60),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a33a),
	.w1(32'hba92bf64),
	.w2(32'h3abc2292),
	.w3(32'hbc12372d),
	.w4(32'hba921a02),
	.w5(32'hbb10638f),
	.w6(32'hbbbf597d),
	.w7(32'hbb8e905f),
	.w8(32'h3992fd47),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389623a9),
	.w1(32'h3ad1fcd5),
	.w2(32'h3af2f0c1),
	.w3(32'hbb339521),
	.w4(32'hbb25bdae),
	.w5(32'h3b8accbe),
	.w6(32'hbae28312),
	.w7(32'h3a40f7ea),
	.w8(32'h3b5c171d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c0d0),
	.w1(32'hbb3daec9),
	.w2(32'hb9ad493a),
	.w3(32'h3b56c1a1),
	.w4(32'h3ba359ea),
	.w5(32'h3b9acdf1),
	.w6(32'h3b12a102),
	.w7(32'hbb102f37),
	.w8(32'h3bbe6578),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5b4ca),
	.w1(32'hbbcaaa02),
	.w2(32'hbbf7d2db),
	.w3(32'hbb3c433e),
	.w4(32'hbb45781e),
	.w5(32'hbc476c23),
	.w6(32'h3a30ad3a),
	.w7(32'h38155fd1),
	.w8(32'hbbf952bb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592e19),
	.w1(32'hbc4f24c9),
	.w2(32'h3bf34c0e),
	.w3(32'hbcfb1a27),
	.w4(32'hbca76e9a),
	.w5(32'h3b23c5da),
	.w6(32'hbb6e2424),
	.w7(32'hbaa4e659),
	.w8(32'h3c3b1a7c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3571b1),
	.w1(32'h3b3e703c),
	.w2(32'hbb5daa74),
	.w3(32'h3c5ff309),
	.w4(32'h3c56896e),
	.w5(32'h3b8c19b7),
	.w6(32'h3c0444ac),
	.w7(32'h3b52e303),
	.w8(32'hbaed136b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe547a),
	.w1(32'hbb20bcc2),
	.w2(32'h3b9a10f7),
	.w3(32'hbbac9d3e),
	.w4(32'hbad7e282),
	.w5(32'h3c0a015e),
	.w6(32'hbb5a1e11),
	.w7(32'hbb2659e0),
	.w8(32'h3b8777a3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0cc67),
	.w1(32'h3c364493),
	.w2(32'h3b92098a),
	.w3(32'hbb3bd33b),
	.w4(32'h3c019046),
	.w5(32'hbad9546c),
	.w6(32'hbba79204),
	.w7(32'h3bad191b),
	.w8(32'hbbc6f527),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff268d),
	.w1(32'h3c173568),
	.w2(32'h3c17c46e),
	.w3(32'h3b87158c),
	.w4(32'h3c6df8bb),
	.w5(32'h3c648e30),
	.w6(32'h3ba6e465),
	.w7(32'h3c304371),
	.w8(32'h3bfa078d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c424dbd),
	.w1(32'h3be6f44c),
	.w2(32'h3a7460e1),
	.w3(32'h3c536a09),
	.w4(32'h3ba62a1e),
	.w5(32'hbae0c10c),
	.w6(32'h3c3f1afb),
	.w7(32'h3bffb95e),
	.w8(32'h3a57f8cb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443570),
	.w1(32'hbaed230d),
	.w2(32'hbb879c32),
	.w3(32'hbb37cec1),
	.w4(32'hba9c08ae),
	.w5(32'hbbbbfda9),
	.w6(32'hbac50903),
	.w7(32'h3b8f87fe),
	.w8(32'hbbbda899),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac90a4e),
	.w1(32'h3b047662),
	.w2(32'hbb8c0428),
	.w3(32'hba9f5c98),
	.w4(32'hbb872901),
	.w5(32'h3c39a38d),
	.w6(32'h3b3fcd86),
	.w7(32'hbb9b7a82),
	.w8(32'h3b5d9f4a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cace4e7),
	.w1(32'h3b11c0a0),
	.w2(32'h3c08f762),
	.w3(32'h3d356ba7),
	.w4(32'h3cc01645),
	.w5(32'h3c188f6b),
	.w6(32'h3d043d1c),
	.w7(32'h3c2ed238),
	.w8(32'h3bcff470),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c080caf),
	.w1(32'h3bd1437c),
	.w2(32'hbb31b8f0),
	.w3(32'h3c315eeb),
	.w4(32'h3b92e950),
	.w5(32'hbc2db457),
	.w6(32'h3c6c04c7),
	.w7(32'h3be9eb14),
	.w8(32'h3986114a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa528b),
	.w1(32'h3ac61bf0),
	.w2(32'h3b1d4c20),
	.w3(32'h3bab6327),
	.w4(32'h3b017ad7),
	.w5(32'hba505d7e),
	.w6(32'h3c37676e),
	.w7(32'hbad620fd),
	.w8(32'h3bfaca55),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59f552),
	.w1(32'h3bcfb366),
	.w2(32'h3bbe8f70),
	.w3(32'hbaf5be74),
	.w4(32'hb9d69884),
	.w5(32'h3b876f1b),
	.w6(32'h3b4a2e77),
	.w7(32'hba3ba7b4),
	.w8(32'h3b52504f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacea356),
	.w1(32'hbbb8c5bf),
	.w2(32'hbb43ae64),
	.w3(32'h3b77083d),
	.w4(32'hbb7370dd),
	.w5(32'hbaf30fa7),
	.w6(32'h3ba0bb16),
	.w7(32'h3b11c112),
	.w8(32'hbb425595),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83bb4e),
	.w1(32'hbb04df7e),
	.w2(32'h3b570704),
	.w3(32'h3a8efe3d),
	.w4(32'hbb0482c0),
	.w5(32'hbae51fd8),
	.w6(32'h3b8b200e),
	.w7(32'hb9903e3d),
	.w8(32'h3b04ef9a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0e95),
	.w1(32'h3bf69bc1),
	.w2(32'h3c074449),
	.w3(32'hbabc8db6),
	.w4(32'h3bd4dc9f),
	.w5(32'h3b810f57),
	.w6(32'h3a67b056),
	.w7(32'h3be93ffd),
	.w8(32'h3bc41e99),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12a3d1),
	.w1(32'h3bed7418),
	.w2(32'hbb92aa48),
	.w3(32'h3be60701),
	.w4(32'h3bc878b0),
	.w5(32'h3b429921),
	.w6(32'h3c93ef39),
	.w7(32'h3c5822d4),
	.w8(32'hb8483df0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d717b),
	.w1(32'hb9317d86),
	.w2(32'h3b427672),
	.w3(32'hbb85e437),
	.w4(32'hbb31674b),
	.w5(32'h3b86676d),
	.w6(32'hbb934c88),
	.w7(32'hba85fba1),
	.w8(32'h3a836c7f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed4672),
	.w1(32'h3baf06e3),
	.w2(32'h3b32ed32),
	.w3(32'h3b987da9),
	.w4(32'h3bc5e3f4),
	.w5(32'h3b288b6b),
	.w6(32'hba9644df),
	.w7(32'h3bdd8fcd),
	.w8(32'hb988f879),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc85db),
	.w1(32'h3b18c089),
	.w2(32'h3b87a7ae),
	.w3(32'h3bb3373c),
	.w4(32'h3ad84115),
	.w5(32'h3b8d45e8),
	.w6(32'hbafaba0e),
	.w7(32'h3b9928e3),
	.w8(32'h3b331016),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd42a1),
	.w1(32'h3a4de09e),
	.w2(32'h3b8eef9f),
	.w3(32'hbb88741c),
	.w4(32'hbb7b3541),
	.w5(32'h3c0983d0),
	.w6(32'hbb8254cd),
	.w7(32'h3a84ac73),
	.w8(32'h3bd7a715),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29dd8),
	.w1(32'hbadd2ff8),
	.w2(32'h3bfeae9f),
	.w3(32'hbbb624d9),
	.w4(32'hbbab2e20),
	.w5(32'h3c3f819b),
	.w6(32'hbba6eede),
	.w7(32'hbc1716b1),
	.w8(32'h3c1cdfb3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bfb1e),
	.w1(32'h3c12c5d4),
	.w2(32'hba1af9f8),
	.w3(32'h3c8cacf2),
	.w4(32'h3c851426),
	.w5(32'h3b8ee13b),
	.w6(32'h3c8f73ee),
	.w7(32'h3c7561d4),
	.w8(32'h3be9533f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617ad8),
	.w1(32'h3c070fac),
	.w2(32'h3c247fb1),
	.w3(32'h3ba07380),
	.w4(32'h3c23e165),
	.w5(32'h3bc47c1e),
	.w6(32'h3b89e83e),
	.w7(32'hbabe576b),
	.w8(32'h3b3e7588),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c0d6),
	.w1(32'h3aa952e2),
	.w2(32'hbbd622e1),
	.w3(32'h3a97c1da),
	.w4(32'h3b32b813),
	.w5(32'hbbb0ea91),
	.w6(32'h3c488cc7),
	.w7(32'h3c0abd99),
	.w8(32'hbaf8f410),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc842c34),
	.w1(32'hbc48a19b),
	.w2(32'h3bd3954b),
	.w3(32'hbc54b112),
	.w4(32'hbc0a1552),
	.w5(32'h3b8c0612),
	.w6(32'hbb9d82b9),
	.w7(32'hbb889da3),
	.w8(32'h3bb807cc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27ff2b),
	.w1(32'h3c02de11),
	.w2(32'hbc336891),
	.w3(32'h3b9f7c52),
	.w4(32'hba11e60f),
	.w5(32'hbc90893f),
	.w6(32'h3c58ca61),
	.w7(32'h3bfd80ce),
	.w8(32'hbc30f2d9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc427bb6),
	.w1(32'hbc1712e3),
	.w2(32'hbb9a3f92),
	.w3(32'hbcb1f389),
	.w4(32'hbc8453d1),
	.w5(32'h3b879958),
	.w6(32'hbc9eaa09),
	.w7(32'hbc5946da),
	.w8(32'hb9ba5868),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07edbc),
	.w1(32'hbc0d794f),
	.w2(32'h3ad67ab4),
	.w3(32'h3c7f23a8),
	.w4(32'h3b81bac5),
	.w5(32'hb9d31708),
	.w6(32'h3c4fff87),
	.w7(32'h3b93bfa1),
	.w8(32'h3a6cc553),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d5e39),
	.w1(32'h3b5459ea),
	.w2(32'hbab25ccd),
	.w3(32'hbb334a24),
	.w4(32'hbb995665),
	.w5(32'hbc14262e),
	.w6(32'hbac3f28b),
	.w7(32'h3afd2515),
	.w8(32'hbc2068af),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf54ebe),
	.w1(32'hbac8ac54),
	.w2(32'h3aa53f2c),
	.w3(32'hbc870618),
	.w4(32'hbc20e7e3),
	.w5(32'h39b3938f),
	.w6(32'hbaf65d4b),
	.w7(32'hbb3988ba),
	.w8(32'hba92c8db),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabefc39),
	.w1(32'hbae52342),
	.w2(32'h3b65298e),
	.w3(32'h3a5f9a22),
	.w4(32'hbb115cd5),
	.w5(32'h3b1f9308),
	.w6(32'hbb1d043b),
	.w7(32'hbb5e9ed0),
	.w8(32'hba6328b8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa48461),
	.w1(32'h3ae6aa29),
	.w2(32'h3b98144d),
	.w3(32'h3b77cf20),
	.w4(32'h39df538c),
	.w5(32'h3c10635c),
	.w6(32'h3b213b02),
	.w7(32'h3c0edba6),
	.w8(32'h3c145c6a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c369d23),
	.w1(32'h3b6b5566),
	.w2(32'hbc64baec),
	.w3(32'h3b479cd2),
	.w4(32'hbb508bc3),
	.w5(32'hbcc748ae),
	.w6(32'h3c75a43f),
	.w7(32'h3bb89e5c),
	.w8(32'hbcaf218d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1df0bd),
	.w1(32'h3c048bb2),
	.w2(32'hbb69b16c),
	.w3(32'h3af1a0d1),
	.w4(32'h3a2b41aa),
	.w5(32'h39b00906),
	.w6(32'hba38696d),
	.w7(32'hbc43580b),
	.w8(32'hbacb51e2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01e11b),
	.w1(32'h3ba1cc59),
	.w2(32'h3b81ea59),
	.w3(32'hbb5f2866),
	.w4(32'h3b76b66a),
	.w5(32'hbb0582d3),
	.w6(32'hbaae77a7),
	.w7(32'hbb5f91c2),
	.w8(32'h3b58aff4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda551b),
	.w1(32'hbab27157),
	.w2(32'h3beb92d9),
	.w3(32'hbb92a659),
	.w4(32'hbb0cc1fe),
	.w5(32'h3bf87dc9),
	.w6(32'hbba964b5),
	.w7(32'hbb41d50d),
	.w8(32'h3b8b0e3f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb640fa),
	.w1(32'h3bc958a3),
	.w2(32'hbc48eee4),
	.w3(32'h3a6bf171),
	.w4(32'hbb0da904),
	.w5(32'hbc5273bc),
	.w6(32'h3c3ab5c9),
	.w7(32'hbb402f18),
	.w8(32'hbbd5f8a5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e5cb),
	.w1(32'hba615ecf),
	.w2(32'h3a8a2dab),
	.w3(32'h3a307635),
	.w4(32'h3bca4e55),
	.w5(32'hbad9a10c),
	.w6(32'h3b9c6b46),
	.w7(32'h3b43a1b8),
	.w8(32'h3b6d4110),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c079359),
	.w1(32'h3c60c7ca),
	.w2(32'h3c299770),
	.w3(32'h3bcab332),
	.w4(32'h3b324994),
	.w5(32'h3b5a09bd),
	.w6(32'h3c798e6b),
	.w7(32'hba87a4ef),
	.w8(32'h3c53bb24),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc659a9),
	.w1(32'h3bd75206),
	.w2(32'h39babf17),
	.w3(32'h3bff5464),
	.w4(32'h3b3d3925),
	.w5(32'h3b34d7d1),
	.w6(32'h3c6d4927),
	.w7(32'h3bfe3dd8),
	.w8(32'h3bcee7f4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e5613),
	.w1(32'h3b81ad38),
	.w2(32'hbba5b9e1),
	.w3(32'hb97b7f94),
	.w4(32'h3a8ce8ae),
	.w5(32'hbab5ef06),
	.w6(32'h3b164265),
	.w7(32'h3b9514d0),
	.w8(32'hba23a37d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb09c7),
	.w1(32'hbae84020),
	.w2(32'h3b4b61f6),
	.w3(32'h3b41269a),
	.w4(32'h3b71bba5),
	.w5(32'h3b8f9aec),
	.w6(32'hbb26e694),
	.w7(32'h3ac1d0e1),
	.w8(32'hbab54e4d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7290c),
	.w1(32'h3a0c0a1e),
	.w2(32'h3ac6f6fd),
	.w3(32'h3be65d9e),
	.w4(32'h3b5f2814),
	.w5(32'h3a144d0e),
	.w6(32'h3bf18d36),
	.w7(32'h3bfc73f2),
	.w8(32'h3bfa021c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dfb12),
	.w1(32'h3bd8828c),
	.w2(32'h3af3f0c9),
	.w3(32'hbae049ef),
	.w4(32'h3b8012f7),
	.w5(32'h397f6f7f),
	.w6(32'h3a2a5f20),
	.w7(32'h3b84223d),
	.w8(32'hba9b31a1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a991b5e),
	.w1(32'h3bd22f0e),
	.w2(32'h3ba5251e),
	.w3(32'hba03d31e),
	.w4(32'h3bf9e515),
	.w5(32'h3bc61e63),
	.w6(32'h3ab33ad7),
	.w7(32'hba31354d),
	.w8(32'h3bcb790b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde272a),
	.w1(32'h3b1e8911),
	.w2(32'h3be4bd3a),
	.w3(32'h3b9a6836),
	.w4(32'h3b1e88b3),
	.w5(32'h39e73a73),
	.w6(32'hbba19c18),
	.w7(32'hbb4f4e8f),
	.w8(32'hb6fe3236),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97afb0),
	.w1(32'h3b2f897b),
	.w2(32'hbb25e37e),
	.w3(32'h3c1ed566),
	.w4(32'h3bf6008f),
	.w5(32'h3bbec4b1),
	.w6(32'h3baeb289),
	.w7(32'h3ba87f08),
	.w8(32'h3b93fdb0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3aafe),
	.w1(32'h3b8919f3),
	.w2(32'hbba24388),
	.w3(32'h3c247f3c),
	.w4(32'h3b9b78cf),
	.w5(32'h3aa2768f),
	.w6(32'h3ba28768),
	.w7(32'h3bd57740),
	.w8(32'hbb98f4e1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab33f6a),
	.w1(32'h39df7200),
	.w2(32'h3b889305),
	.w3(32'h3a8ebe5f),
	.w4(32'hba1ad2f4),
	.w5(32'hbb308df7),
	.w6(32'hbb80bacf),
	.w7(32'hbb9ba9ba),
	.w8(32'hbbc36c03),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be433e1),
	.w1(32'h3b6c84b8),
	.w2(32'hbaa254b4),
	.w3(32'hbb07d25c),
	.w4(32'hbacb1a6d),
	.w5(32'h3bbdd47e),
	.w6(32'hbb9c0d7e),
	.w7(32'hbb5f4f9e),
	.w8(32'h3b41f43d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18df16),
	.w1(32'hbc014e10),
	.w2(32'h3b6977d9),
	.w3(32'h3b936890),
	.w4(32'h3a1a0307),
	.w5(32'hbba378ac),
	.w6(32'h3b80a62c),
	.w7(32'h3b1b6069),
	.w8(32'hbbbe40df),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b3ef0),
	.w1(32'h3b26840f),
	.w2(32'h3b7a335d),
	.w3(32'hbb9d7922),
	.w4(32'hbadf9494),
	.w5(32'h3c096e76),
	.w6(32'hbbc1997d),
	.w7(32'hbb54ee17),
	.w8(32'h3bef217f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977199),
	.w1(32'h3b85e22d),
	.w2(32'hbb5460e0),
	.w3(32'h3bea8df8),
	.w4(32'h3bbeb39d),
	.w5(32'hbaaf43be),
	.w6(32'h3c113f29),
	.w7(32'h3bb4aeb5),
	.w8(32'h3a60fb58),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bf9b9),
	.w1(32'hbae97e2c),
	.w2(32'hbac5bae1),
	.w3(32'hbb081154),
	.w4(32'hba8ef7c1),
	.w5(32'hbb02e845),
	.w6(32'hbad79dcb),
	.w7(32'hbb89f5da),
	.w8(32'hbb09ac4b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f89f15),
	.w1(32'h3b338e83),
	.w2(32'h3c06eacd),
	.w3(32'hba614649),
	.w4(32'hbb108040),
	.w5(32'h3bef5db0),
	.w6(32'hbb52c646),
	.w7(32'h3b27c06a),
	.w8(32'h3beda15f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba521b6),
	.w1(32'h3bb8f7db),
	.w2(32'h3a6f5067),
	.w3(32'h386ea579),
	.w4(32'hb96cae99),
	.w5(32'hbb9d427f),
	.w6(32'h3be9ffeb),
	.w7(32'h3b7f57af),
	.w8(32'h3b25bc73),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9965),
	.w1(32'h38c2985c),
	.w2(32'h3c1b08e3),
	.w3(32'hbc80bf68),
	.w4(32'hbbf1741b),
	.w5(32'h3c536720),
	.w6(32'hbc3fbb08),
	.w7(32'hbbe85a5a),
	.w8(32'h3c1c9d0d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdebcc9),
	.w1(32'hbad1dc80),
	.w2(32'h3baae026),
	.w3(32'h3c40ea42),
	.w4(32'h3b1811c7),
	.w5(32'h3b5e5716),
	.w6(32'h3c585982),
	.w7(32'h3b5869e5),
	.w8(32'hb919d671),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba255f49),
	.w1(32'h3a4eace7),
	.w2(32'h3c0d3ca9),
	.w3(32'hbb2382d4),
	.w4(32'hbb3ff944),
	.w5(32'h3c4131d0),
	.w6(32'hbb377871),
	.w7(32'hbb66487b),
	.w8(32'h3c2698b7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc50641),
	.w1(32'h3bf86a91),
	.w2(32'hba671c6a),
	.w3(32'h3bff9a5f),
	.w4(32'h3c40352c),
	.w5(32'hb8c74d64),
	.w6(32'h3bd03a7f),
	.w7(32'h3c5014ee),
	.w8(32'hbab00f5b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013ce8),
	.w1(32'h3b149543),
	.w2(32'h3b8617d7),
	.w3(32'h39fad728),
	.w4(32'h3b034c93),
	.w5(32'h3ba68dcd),
	.w6(32'h3ae8b202),
	.w7(32'h3b954647),
	.w8(32'h3bc5d608),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e5e39),
	.w1(32'hbbbd6ad2),
	.w2(32'hbbc6b87e),
	.w3(32'h3c82638a),
	.w4(32'h3b90944f),
	.w5(32'h3b9669d9),
	.w6(32'h3c5c2158),
	.w7(32'hbb53b1b2),
	.w8(32'h3a162798),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbf864),
	.w1(32'h39c975a8),
	.w2(32'hba8b0b02),
	.w3(32'hbb2149b9),
	.w4(32'hbb340a30),
	.w5(32'hbb5409c8),
	.w6(32'hbb88532c),
	.w7(32'hbae0924d),
	.w8(32'h3bd9a614),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3815ab),
	.w1(32'h3b6211ee),
	.w2(32'hbb5b8228),
	.w3(32'hba81e409),
	.w4(32'hbb1c63ac),
	.w5(32'hbc0a582a),
	.w6(32'hbae6351b),
	.w7(32'h38d71dc2),
	.w8(32'hbbc324c2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b4674),
	.w1(32'hbb197eb7),
	.w2(32'h39a7b101),
	.w3(32'hbbaef8ad),
	.w4(32'hbb840eb9),
	.w5(32'hb8bb5284),
	.w6(32'hbbdd1763),
	.w7(32'hbc03796d),
	.w8(32'hbb6cb79b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af84080),
	.w1(32'hbaca070b),
	.w2(32'h3be89b4a),
	.w3(32'hbb8e236a),
	.w4(32'hbb56b45f),
	.w5(32'h3a2015db),
	.w6(32'h3b5aa24a),
	.w7(32'hbaace18e),
	.w8(32'h3be7c578),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f0233),
	.w1(32'h3b8391e2),
	.w2(32'h3bd6958b),
	.w3(32'hb9faa7d7),
	.w4(32'hbbd5b5da),
	.w5(32'h3b8b8533),
	.w6(32'h3817f49c),
	.w7(32'h3b70b548),
	.w8(32'h3b03a5a0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b56b9),
	.w1(32'h3aca147e),
	.w2(32'hbac31393),
	.w3(32'hbae510a8),
	.w4(32'hbb717470),
	.w5(32'h3ca9d33c),
	.w6(32'hbba1fe68),
	.w7(32'h3a77aebc),
	.w8(32'h3ba9ccd9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf27062),
	.w1(32'h3b885c33),
	.w2(32'hb965af78),
	.w3(32'h3d890b1e),
	.w4(32'h3d0c236a),
	.w5(32'hbc05625c),
	.w6(32'h3d71e097),
	.w7(32'h3cd9981e),
	.w8(32'h3abe4e6a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc6c0f),
	.w1(32'h3b3bb6af),
	.w2(32'h3b31152c),
	.w3(32'hbc05e0a9),
	.w4(32'h3acb26e1),
	.w5(32'h3c17aee6),
	.w6(32'hbbd4db7d),
	.w7(32'hbb0a1fa2),
	.w8(32'h3b9f5ebe),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6692ff),
	.w1(32'hbb39e845),
	.w2(32'h3b933762),
	.w3(32'h3aca1a74),
	.w4(32'h39b6a000),
	.w5(32'h3b0fc730),
	.w6(32'h3ab691b3),
	.w7(32'h3b55b4b8),
	.w8(32'h3b1b21a6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a4af0),
	.w1(32'h3b328d33),
	.w2(32'h3b975812),
	.w3(32'h3aff5bb2),
	.w4(32'hbb722e5b),
	.w5(32'hbb5178eb),
	.w6(32'h3c1a68c4),
	.w7(32'h3b86d955),
	.w8(32'h3ba84e51),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6241ea),
	.w1(32'h3c0b23c9),
	.w2(32'hbb1f1c74),
	.w3(32'hbbe79613),
	.w4(32'h3ae364b2),
	.w5(32'hba8c92b0),
	.w6(32'hbb59c1d7),
	.w7(32'h3b70e180),
	.w8(32'hbb4b3270),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba756904),
	.w1(32'hb88fa9ff),
	.w2(32'h3b99bb6f),
	.w3(32'hbb431cc7),
	.w4(32'h3ae6d2a4),
	.w5(32'h3c157bc1),
	.w6(32'h3b10e297),
	.w7(32'h3a4647d5),
	.w8(32'h3c38bc13),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ba412),
	.w1(32'h3c158f5b),
	.w2(32'hbc39be2b),
	.w3(32'h3cbf5247),
	.w4(32'h3c8a5202),
	.w5(32'hbc8212c6),
	.w6(32'h3ca851af),
	.w7(32'h3c70c16d),
	.w8(32'hbbf1b70b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79b9da),
	.w1(32'hbbc1fed4),
	.w2(32'h3bfad2d6),
	.w3(32'hbcc5266d),
	.w4(32'hbc363b66),
	.w5(32'h3ba4b130),
	.w6(32'hbcb3e5cc),
	.w7(32'hbc19a13b),
	.w8(32'h3b0ce06b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b711182),
	.w1(32'h3bcb954f),
	.w2(32'h39e95051),
	.w3(32'h3b723208),
	.w4(32'h3b1f2db9),
	.w5(32'hba24eec4),
	.w6(32'hb946d247),
	.w7(32'h3b2c815b),
	.w8(32'hbb9b8d2c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c844),
	.w1(32'h3b2a0578),
	.w2(32'h3ae6b37a),
	.w3(32'hba2ccbad),
	.w4(32'h3bb10c37),
	.w5(32'hba4f3f21),
	.w6(32'hbba6b0c2),
	.w7(32'h3a90065a),
	.w8(32'h3adc64fd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a0cf),
	.w1(32'h39e92439),
	.w2(32'h3b6e3c3c),
	.w3(32'hbbad6e98),
	.w4(32'hba9c5d0a),
	.w5(32'h3a3d747f),
	.w6(32'hbaaff6a8),
	.w7(32'h3adfb260),
	.w8(32'hbb15d6e3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1354),
	.w1(32'h3bcaac28),
	.w2(32'hbc05e0be),
	.w3(32'h3b59f9bc),
	.w4(32'h3bad41c8),
	.w5(32'hbc162520),
	.w6(32'h3a8e3f6b),
	.w7(32'h3b305290),
	.w8(32'hbc1721dd),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd5e79),
	.w1(32'hbaddc4a4),
	.w2(32'h3b1a7c5e),
	.w3(32'hbc28009d),
	.w4(32'hbbab2cb0),
	.w5(32'hbc066ffd),
	.w6(32'hbc3d6b8a),
	.w7(32'hbbfa9319),
	.w8(32'hba34d35b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc58027),
	.w1(32'hbb77bade),
	.w2(32'h3aea807b),
	.w3(32'h39b43489),
	.w4(32'hbbb05420),
	.w5(32'h3aad9738),
	.w6(32'h38cb87dc),
	.w7(32'h3af6b722),
	.w8(32'h3b8e08e4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227589),
	.w1(32'h3bd79cd6),
	.w2(32'hbab80bef),
	.w3(32'hba5587f4),
	.w4(32'h3bb489c3),
	.w5(32'hbbf6aac7),
	.w6(32'h3b1ade2b),
	.w7(32'h3ba13552),
	.w8(32'hbba9afc2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c317d),
	.w1(32'hb9d09c13),
	.w2(32'h3bb848ac),
	.w3(32'h3a9e2e2d),
	.w4(32'hbb37c17a),
	.w5(32'hbaa9126e),
	.w6(32'h3b85ecdd),
	.w7(32'h3a829cc9),
	.w8(32'h3ae528cf),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92627c),
	.w1(32'h3ba90dc9),
	.w2(32'hbaed77a1),
	.w3(32'h3bb247fb),
	.w4(32'h3baac483),
	.w5(32'hbc517083),
	.w6(32'hba10809e),
	.w7(32'h3b92ba9e),
	.w8(32'hbbef31ab),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56024f),
	.w1(32'hbc26d2e7),
	.w2(32'hbc5d810c),
	.w3(32'hbd0013ab),
	.w4(32'hbcf83e56),
	.w5(32'hbc4e49b1),
	.w6(32'hbc81a15b),
	.w7(32'hbc8a48bb),
	.w8(32'hbc26a417),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ec8b8),
	.w1(32'hb9f888ee),
	.w2(32'h3b884711),
	.w3(32'hbcbcfb0e),
	.w4(32'hbb9ffef8),
	.w5(32'h3c437414),
	.w6(32'hbca79fff),
	.w7(32'hbbb08656),
	.w8(32'h3ae68eb4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a5d87),
	.w1(32'h3b902766),
	.w2(32'hb96c1a4e),
	.w3(32'h3b56c73b),
	.w4(32'h3b1ff3f4),
	.w5(32'h3af86346),
	.w6(32'hba4b4a8d),
	.w7(32'h3a810fe2),
	.w8(32'hbbac15ce),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399602ed),
	.w1(32'h39b66489),
	.w2(32'hba41c902),
	.w3(32'hb8e69ce3),
	.w4(32'h3997e30a),
	.w5(32'hbac6bcab),
	.w6(32'h3966f061),
	.w7(32'h3b73da2c),
	.w8(32'h39947a5b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad72b2f),
	.w1(32'h3b5b1a06),
	.w2(32'hbb88b380),
	.w3(32'h3be85711),
	.w4(32'h3aa697be),
	.w5(32'hb9f8c5ab),
	.w6(32'hba27b419),
	.w7(32'h39c23310),
	.w8(32'hbb1adf55),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac8de),
	.w1(32'hbb52a48a),
	.w2(32'hbc5c520c),
	.w3(32'hbb295325),
	.w4(32'hbb981769),
	.w5(32'hbc33b78a),
	.w6(32'h3b1d55df),
	.w7(32'h3c1fd8db),
	.w8(32'hbbed1dfa),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7760e7),
	.w1(32'h3af7d25e),
	.w2(32'hb8f15c26),
	.w3(32'hbc86bea6),
	.w4(32'hbc661d5e),
	.w5(32'hba81b848),
	.w6(32'hbb911e04),
	.w7(32'h3aa0f224),
	.w8(32'h3a8b7222),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac91959),
	.w1(32'h3a716491),
	.w2(32'h3ae57dec),
	.w3(32'h3a557c36),
	.w4(32'hbaf4b206),
	.w5(32'hbc104af3),
	.w6(32'hbab57b5d),
	.w7(32'h3853fe7f),
	.w8(32'h3c3f7bd6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000fce),
	.w1(32'hba00f3f1),
	.w2(32'hbb44cf3a),
	.w3(32'hbb928205),
	.w4(32'hbb81491b),
	.w5(32'hbbf45f82),
	.w6(32'h3c227415),
	.w7(32'h3ba63afc),
	.w8(32'h3bb67a25),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8a3b5),
	.w1(32'hbc74a964),
	.w2(32'hbab32d7e),
	.w3(32'hbba00431),
	.w4(32'hbc089646),
	.w5(32'hbaafe950),
	.w6(32'h3c6518b7),
	.w7(32'h3bd15935),
	.w8(32'h3b02d738),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fa445),
	.w1(32'hba544d9e),
	.w2(32'hbaeffac8),
	.w3(32'hbb2e1a39),
	.w4(32'hbb090c42),
	.w5(32'h3cbf4c19),
	.w6(32'hb8b10053),
	.w7(32'h3ad02c34),
	.w8(32'h3c9350a1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bce19),
	.w1(32'h3c1ea692),
	.w2(32'h3b817e38),
	.w3(32'h3caeff3e),
	.w4(32'h3b1a17b3),
	.w5(32'hba28cc63),
	.w6(32'hbc0ed562),
	.w7(32'hbb8b00da),
	.w8(32'hbabf67f1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d70f3),
	.w1(32'hbb50a6ed),
	.w2(32'hbc8caaa2),
	.w3(32'h3a364abc),
	.w4(32'h3a73363b),
	.w5(32'h3c8fbd5a),
	.w6(32'h3b3c49cf),
	.w7(32'h388608bf),
	.w8(32'h3d042958),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63a41d),
	.w1(32'h3c88eef4),
	.w2(32'hba83b815),
	.w3(32'h3cd6b0f7),
	.w4(32'hbbbda2f7),
	.w5(32'hba207f9c),
	.w6(32'hbbb67d98),
	.w7(32'hbbad65de),
	.w8(32'hbb4dca6c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46676),
	.w1(32'hbbc2dabc),
	.w2(32'hba92cba7),
	.w3(32'hbaec7dd1),
	.w4(32'hbb9db3d6),
	.w5(32'h3a013c26),
	.w6(32'hbbad27d5),
	.w7(32'h3b040f84),
	.w8(32'hbb2052b7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb8e7),
	.w1(32'h3a443b25),
	.w2(32'h3c698b76),
	.w3(32'h3ba25368),
	.w4(32'h3a839f8b),
	.w5(32'hbab481cf),
	.w6(32'h3a9b38c1),
	.w7(32'hbb724cce),
	.w8(32'h3ae47d39),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac0b9),
	.w1(32'h3b413fff),
	.w2(32'hbb0c1090),
	.w3(32'h3a5a1cde),
	.w4(32'hbc19fdd8),
	.w5(32'hba0672d0),
	.w6(32'hbbd2ab77),
	.w7(32'hbc133794),
	.w8(32'h3c0b8134),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c9286),
	.w1(32'hba72f093),
	.w2(32'hbbc28763),
	.w3(32'h3bdcc1c0),
	.w4(32'h3baec96e),
	.w5(32'hbbc1bd72),
	.w6(32'h3c1f4edf),
	.w7(32'hbab5f728),
	.w8(32'h3b63f40a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf0500),
	.w1(32'h3aa83f4c),
	.w2(32'hbcbeb4d9),
	.w3(32'hba7fa30c),
	.w4(32'h3b83bb0b),
	.w5(32'hbba68a37),
	.w6(32'h3b01368a),
	.w7(32'hbb44afff),
	.w8(32'h3c22a962),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdc16b),
	.w1(32'hbc0f5bca),
	.w2(32'hbb28445f),
	.w3(32'hbb8adf1c),
	.w4(32'hbabdb81e),
	.w5(32'hbac8e1c0),
	.w6(32'h3c0ee22d),
	.w7(32'h3b542d04),
	.w8(32'hbb61821d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06c88),
	.w1(32'hbbb04373),
	.w2(32'h3c554b89),
	.w3(32'hba209305),
	.w4(32'h3aa14eb6),
	.w5(32'hbb86fc14),
	.w6(32'h3b488266),
	.w7(32'h3b4c3894),
	.w8(32'hbbf3d91f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23aebe),
	.w1(32'hbc849f5f),
	.w2(32'h3c1bc0c2),
	.w3(32'hbcb07ed0),
	.w4(32'hbc27e69e),
	.w5(32'h3ad3dc11),
	.w6(32'h39f7e227),
	.w7(32'h3b887f50),
	.w8(32'h3cbeeb3c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ef5b9),
	.w1(32'h3c796b3d),
	.w2(32'hbc28e342),
	.w3(32'h3c057757),
	.w4(32'hbbdeacf1),
	.w5(32'hbcafe474),
	.w6(32'h3c89ede3),
	.w7(32'hbbe6ae3c),
	.w8(32'hbbd39199),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c3cfb),
	.w1(32'h3bc907ad),
	.w2(32'hbaba9db1),
	.w3(32'h3bb88447),
	.w4(32'h3c881a5d),
	.w5(32'h3b925465),
	.w6(32'h3c6f60e4),
	.w7(32'h3c4a4347),
	.w8(32'h3b5a4dd0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d362e),
	.w1(32'h3b733a57),
	.w2(32'h3b51511d),
	.w3(32'hbaca77e8),
	.w4(32'h3babafbd),
	.w5(32'h3a631a7b),
	.w6(32'hbc9a3fda),
	.w7(32'hbb9c1d9a),
	.w8(32'hba1b1351),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9744524),
	.w1(32'hbb52cc77),
	.w2(32'h3bb2757e),
	.w3(32'hbabf1bb5),
	.w4(32'hbb7718e0),
	.w5(32'hbbb07614),
	.w6(32'hb98e3bfe),
	.w7(32'hbb2c7493),
	.w8(32'hbc0706f8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014611),
	.w1(32'h3a80f5b5),
	.w2(32'h3c0584a3),
	.w3(32'hbc2228f8),
	.w4(32'h3c18a300),
	.w5(32'h3cfd691a),
	.w6(32'hbb1591c0),
	.w7(32'hbb130011),
	.w8(32'h3c33a006),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9be43d),
	.w1(32'hbc89b093),
	.w2(32'h3bc9d7e3),
	.w3(32'h3b8762ae),
	.w4(32'hbcaaf08d),
	.w5(32'h3b4284c0),
	.w6(32'hbc3e0d17),
	.w7(32'hbc2fa28c),
	.w8(32'hbc26f49b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ce91b),
	.w1(32'hbc0cbb0e),
	.w2(32'h3c809c8b),
	.w3(32'hbb1178c8),
	.w4(32'hbc2a48f5),
	.w5(32'h3ce193f7),
	.w6(32'hbb92ce18),
	.w7(32'hbbed19b8),
	.w8(32'hbb0a6329),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c827d8a),
	.w1(32'hbbfe00cb),
	.w2(32'h3bf26d74),
	.w3(32'hbadfda8a),
	.w4(32'hbcf9c52b),
	.w5(32'h3b84a25a),
	.w6(32'hbc8cb129),
	.w7(32'hbc943bdf),
	.w8(32'hbbbac603),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08016c),
	.w1(32'hbbdaba4a),
	.w2(32'h3b6ea8e3),
	.w3(32'hbaf09f11),
	.w4(32'hbb83b98f),
	.w5(32'h3ca4e648),
	.w6(32'hbb954989),
	.w7(32'h3accb852),
	.w8(32'h3ad51c4c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1588e),
	.w1(32'h3ab8a41c),
	.w2(32'hbaa05445),
	.w3(32'h3c84b84d),
	.w4(32'hbc5be571),
	.w5(32'hbbc58d42),
	.w6(32'hb8f4e1cf),
	.w7(32'hbb3a76b8),
	.w8(32'hbb9a0adf),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76e591),
	.w1(32'h3c380a0c),
	.w2(32'h3a008aaf),
	.w3(32'h3b069699),
	.w4(32'hbb13fa92),
	.w5(32'hbae8bdd2),
	.w6(32'hbb51e9a0),
	.w7(32'hbc111f09),
	.w8(32'hbbf6dd6e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b852a81),
	.w1(32'h3b773604),
	.w2(32'h398963f0),
	.w3(32'h3a999799),
	.w4(32'hbc0a7a52),
	.w5(32'h3beaf54f),
	.w6(32'hbb075cc1),
	.w7(32'hbc53cb69),
	.w8(32'hbb48af37),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaaf51),
	.w1(32'hbb007463),
	.w2(32'hbba44345),
	.w3(32'hbae7a8ef),
	.w4(32'h3a4b7b42),
	.w5(32'hbb252077),
	.w6(32'h3b3479f1),
	.w7(32'hbbdd2f6b),
	.w8(32'hba7ff98f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4566f7),
	.w1(32'hbb42159e),
	.w2(32'hba608ba3),
	.w3(32'h3bbe9832),
	.w4(32'hbbac029e),
	.w5(32'h3b866722),
	.w6(32'hba9f9c98),
	.w7(32'hbb9ba1f5),
	.w8(32'hbae11494),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c1dec),
	.w1(32'hbba08a62),
	.w2(32'hbab69ce8),
	.w3(32'h3b930dce),
	.w4(32'hbb94b23f),
	.w5(32'h3b051470),
	.w6(32'h3bbabb6d),
	.w7(32'h3b0f2c31),
	.w8(32'hbb05869a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e6279),
	.w1(32'hbb45baf1),
	.w2(32'h3b564f76),
	.w3(32'hbc408746),
	.w4(32'h3b365052),
	.w5(32'hbc3e1bc5),
	.w6(32'h3a50c0a5),
	.w7(32'h3c404c9e),
	.w8(32'h3a297f9b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c2bb),
	.w1(32'hbb935770),
	.w2(32'hbbdc9c79),
	.w3(32'h3c25b173),
	.w4(32'hba8a186c),
	.w5(32'hbba80f12),
	.w6(32'h3af6ef18),
	.w7(32'hbbde44fb),
	.w8(32'hba9d5181),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06117b),
	.w1(32'hbb3bb2a6),
	.w2(32'hbac09525),
	.w3(32'h3ac980ec),
	.w4(32'hbc40ecb2),
	.w5(32'hbb868dc3),
	.w6(32'hbb55dc4b),
	.w7(32'hbc30b2d9),
	.w8(32'hb9de1b7d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed0c64),
	.w1(32'hbbbe31d7),
	.w2(32'hbb837c06),
	.w3(32'hba87cb4b),
	.w4(32'h3b8dc6da),
	.w5(32'h3a84c01d),
	.w6(32'h3b5a98b7),
	.w7(32'h3ba71110),
	.w8(32'h3b55248d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf95805),
	.w1(32'h3bcb1c15),
	.w2(32'h3bbc8ad9),
	.w3(32'h3c03fd5b),
	.w4(32'h3c4850e2),
	.w5(32'h3bb84cfd),
	.w6(32'h394e77bb),
	.w7(32'h3bc55256),
	.w8(32'hb9176141),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baada86),
	.w1(32'hbb8a41b6),
	.w2(32'hbbea2e6e),
	.w3(32'h3bac6cd0),
	.w4(32'hbac24f48),
	.w5(32'hbb3a8249),
	.w6(32'h3b4464bd),
	.w7(32'hbb6868a7),
	.w8(32'h3a451484),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71db35),
	.w1(32'hbba0b30c),
	.w2(32'h3bd5269b),
	.w3(32'h390e23c7),
	.w4(32'hbb5bc0ba),
	.w5(32'hbb9f4465),
	.w6(32'h3a31d48e),
	.w7(32'h3b002d41),
	.w8(32'h3a4b0f0e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e434),
	.w1(32'hbc3c5bac),
	.w2(32'h3c4dad12),
	.w3(32'hbc6e1b2a),
	.w4(32'h3b9f67da),
	.w5(32'h3c7e182f),
	.w6(32'hbaaa894a),
	.w7(32'h3c117bcc),
	.w8(32'hbc37a94d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96adb3),
	.w1(32'h3b9bef3b),
	.w2(32'h3bb3a26b),
	.w3(32'h3c2704b4),
	.w4(32'hbc9a3a34),
	.w5(32'h3b46e5cf),
	.w6(32'hbc940579),
	.w7(32'hbc558f9d),
	.w8(32'h3b8623be),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2154e),
	.w1(32'h3b12fd6f),
	.w2(32'hbc34aee2),
	.w3(32'hbb8332dd),
	.w4(32'hbb1d76ee),
	.w5(32'hbc2cb199),
	.w6(32'h39fa1c76),
	.w7(32'h3ac28852),
	.w8(32'hbb2c54e2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2818b6),
	.w1(32'h3b75f96a),
	.w2(32'hbb7e0b2c),
	.w3(32'h3b8f5858),
	.w4(32'h3bbe65dc),
	.w5(32'h3abde0e8),
	.w6(32'h3b16c5ae),
	.w7(32'h3ae57884),
	.w8(32'h3b4e7355),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e2c8e),
	.w1(32'hbac3ec87),
	.w2(32'hbc8b4b54),
	.w3(32'h3c1a96ab),
	.w4(32'hb9c87753),
	.w5(32'hbccd061d),
	.w6(32'h3ac83f3b),
	.w7(32'hbbe01139),
	.w8(32'hbbeac8d0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc432f36),
	.w1(32'h3cc6e268),
	.w2(32'h3c782559),
	.w3(32'h3b991bec),
	.w4(32'h3ceaaa4a),
	.w5(32'h3cc29f57),
	.w6(32'h3c1a1065),
	.w7(32'h3c83755d),
	.w8(32'h3bdd3298),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92d2ea),
	.w1(32'hbb7d3a1c),
	.w2(32'hbac5d873),
	.w3(32'h3c9f9f6b),
	.w4(32'hbc6577a7),
	.w5(32'hbbe48cf0),
	.w6(32'h3b564d8b),
	.w7(32'hbc87530c),
	.w8(32'hbba38a41),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf28420),
	.w1(32'hbb6c32be),
	.w2(32'hbb6a088c),
	.w3(32'hbbc92a3b),
	.w4(32'hbb08f87e),
	.w5(32'hbc21e87d),
	.w6(32'hbb763b5d),
	.w7(32'hbbe375a1),
	.w8(32'hbb35eabd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca226),
	.w1(32'hb9e5a866),
	.w2(32'h3c64b4b0),
	.w3(32'hbc6cb9ce),
	.w4(32'h3b607e73),
	.w5(32'h3c81c2f7),
	.w6(32'hbbeba851),
	.w7(32'hbb938f68),
	.w8(32'hbc61c1a3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabdc63),
	.w1(32'h3ccee0e1),
	.w2(32'hbb1b4b5c),
	.w3(32'h3cb9c0c2),
	.w4(32'hbc11d2f3),
	.w5(32'h3c1520eb),
	.w6(32'hbc9c156e),
	.w7(32'hbc5448c4),
	.w8(32'hbc5aa480),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f11c6),
	.w1(32'h3c758627),
	.w2(32'hbc12e707),
	.w3(32'h3c58742e),
	.w4(32'hbb868f6b),
	.w5(32'hbc5d7fe5),
	.w6(32'hbc442cc5),
	.w7(32'hbc937489),
	.w8(32'hbbae97e1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc532a17),
	.w1(32'h3c006962),
	.w2(32'h3a9124f9),
	.w3(32'hbc182970),
	.w4(32'h3c0ddd03),
	.w5(32'h3b43e593),
	.w6(32'hbb1b58ee),
	.w7(32'hbbcf7527),
	.w8(32'h3a26c83c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6788e),
	.w1(32'h39e18e04),
	.w2(32'h3b9a2af5),
	.w3(32'h3c8d6b6a),
	.w4(32'h395d72c8),
	.w5(32'h3c04215c),
	.w6(32'h3c3992c9),
	.w7(32'h3b1557ea),
	.w8(32'hbaf68f55),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c395b),
	.w1(32'h3bf1b5ca),
	.w2(32'hbacc2499),
	.w3(32'h3b03910d),
	.w4(32'h3b71dcba),
	.w5(32'hb9ab52b7),
	.w6(32'hbab9da3c),
	.w7(32'h3b74b91b),
	.w8(32'h3be43445),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb604211),
	.w1(32'h3ac7c610),
	.w2(32'hbc3e4a56),
	.w3(32'h3ae6af7c),
	.w4(32'h3b46788d),
	.w5(32'h3c4a837a),
	.w6(32'h3b93b444),
	.w7(32'h3bb9b92b),
	.w8(32'h3b33dbf1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e6a24),
	.w1(32'hbb99ab65),
	.w2(32'hbafb3a4c),
	.w3(32'hbb8e838c),
	.w4(32'hbbbb024d),
	.w5(32'hbb7d653d),
	.w6(32'hbc9288e5),
	.w7(32'h39aa308b),
	.w8(32'h3a10aec8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4c8a9),
	.w1(32'h3c175b20),
	.w2(32'hbc89dbea),
	.w3(32'h3c0b10b8),
	.w4(32'h3ca88f15),
	.w5(32'hbccb5f88),
	.w6(32'h3b25799d),
	.w7(32'h3ad7bd92),
	.w8(32'hbc2ed0f9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b4d05),
	.w1(32'h3c9444f4),
	.w2(32'hba2ca00a),
	.w3(32'h3b879a7d),
	.w4(32'h3c9d669b),
	.w5(32'h3b4695ca),
	.w6(32'h3aac4c04),
	.w7(32'h3ac1107b),
	.w8(32'hbba1fffe),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcabc6b),
	.w1(32'h39e04839),
	.w2(32'hba322ae3),
	.w3(32'hbb86f18b),
	.w4(32'h3ae975f2),
	.w5(32'h3b8a059f),
	.w6(32'hbb953d9d),
	.w7(32'hbc084fad),
	.w8(32'h3a3127a5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b871612),
	.w1(32'hbb7c6b2f),
	.w2(32'hba3e2a7c),
	.w3(32'hba563adf),
	.w4(32'hbc1fe3bf),
	.w5(32'hbbe6b748),
	.w6(32'h3c006f26),
	.w7(32'hbb28646f),
	.w8(32'h394d57f2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa150bc),
	.w1(32'h3b5acda7),
	.w2(32'h3c93e762),
	.w3(32'h3b531da9),
	.w4(32'h3b7b130e),
	.w5(32'h3cdcd9a4),
	.w6(32'h3b7e3798),
	.w7(32'h3ae03778),
	.w8(32'h3bb9dffa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8cfb8),
	.w1(32'hbc9a5c67),
	.w2(32'hbbf4a117),
	.w3(32'h3c181206),
	.w4(32'hbc98c94a),
	.w5(32'hbbac02fc),
	.w6(32'hbc6b1427),
	.w7(32'hbc250bab),
	.w8(32'h3a0026d3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47d789),
	.w1(32'h3c60689e),
	.w2(32'hbc2a82ec),
	.w3(32'h3c2e8e11),
	.w4(32'h3c358a38),
	.w5(32'hbc1fc16a),
	.w6(32'h3c4f46f9),
	.w7(32'h3afeddaf),
	.w8(32'hbb9e7418),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0347f),
	.w1(32'hbbeae387),
	.w2(32'hbbf19184),
	.w3(32'h3bd45202),
	.w4(32'h3ba5ff85),
	.w5(32'h3a4dc80b),
	.w6(32'h3c2b7333),
	.w7(32'h3be9039d),
	.w8(32'hbacce9f0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f327c),
	.w1(32'hbc16ecbf),
	.w2(32'h3b69e4b5),
	.w3(32'h3b88cb69),
	.w4(32'hba5a15b2),
	.w5(32'h3b7c1f0e),
	.w6(32'h3c3aafec),
	.w7(32'h3bb4af67),
	.w8(32'h3c25a51b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f3bc),
	.w1(32'h3c58f91d),
	.w2(32'h3b4bbf26),
	.w3(32'h3bc465fa),
	.w4(32'h3bc73be4),
	.w5(32'h3b69013d),
	.w6(32'h3b0cda9f),
	.w7(32'h3bae2bc1),
	.w8(32'h3b186108),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d5d57),
	.w1(32'h3b9b7150),
	.w2(32'h3be8d5ff),
	.w3(32'h3b717ff6),
	.w4(32'h3b5ab7b4),
	.w5(32'h3cd175b8),
	.w6(32'h3a2cea59),
	.w7(32'hb866b084),
	.w8(32'hba4da717),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e3802),
	.w1(32'hbb364acc),
	.w2(32'h3cc17d11),
	.w3(32'h3bcf9044),
	.w4(32'hbc2ab98e),
	.w5(32'hbabca36b),
	.w6(32'hbc7293db),
	.w7(32'hbc8dc9fd),
	.w8(32'hbc1d4216),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e33f6),
	.w1(32'hbb0fca04),
	.w2(32'hbc02bc9c),
	.w3(32'hbbaf470c),
	.w4(32'h3b87c275),
	.w5(32'h3aa855d5),
	.w6(32'hbb02c617),
	.w7(32'h3c14f316),
	.w8(32'hb907c8bb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06aba4),
	.w1(32'h3b2c1a05),
	.w2(32'hbb85a4e3),
	.w3(32'h3af9eb04),
	.w4(32'h3aa59d4e),
	.w5(32'hbc7a3e61),
	.w6(32'h3b0cb067),
	.w7(32'hbafb19ab),
	.w8(32'hba9df413),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb89543),
	.w1(32'hbbc80d41),
	.w2(32'h3c345f76),
	.w3(32'hbbbb19e9),
	.w4(32'hbcceab6a),
	.w5(32'h3b6ded9c),
	.w6(32'hbc37c199),
	.w7(32'hbcb45558),
	.w8(32'hbc5f61b2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d382c),
	.w1(32'hbad4d8c3),
	.w2(32'hbb2734e6),
	.w3(32'hbb6fe2e1),
	.w4(32'hbc8df68b),
	.w5(32'h3a864748),
	.w6(32'hbc409688),
	.w7(32'hbc1c79f4),
	.w8(32'h3b4a3aad),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4de765),
	.w1(32'hbbdc1e3d),
	.w2(32'hbcd55019),
	.w3(32'h3ad221fb),
	.w4(32'hbbaacbc3),
	.w5(32'hba78210e),
	.w6(32'h3b775b64),
	.w7(32'hba2e81ba),
	.w8(32'h3c938bcd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdff042),
	.w1(32'hbb844c98),
	.w2(32'hbc4a1658),
	.w3(32'h3b2a327b),
	.w4(32'h3c8706d4),
	.w5(32'hbc0d6ef0),
	.w6(32'h3cbbe0ca),
	.w7(32'h3c97b6c4),
	.w8(32'h3c0ca76e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44afc9),
	.w1(32'h3bdee05b),
	.w2(32'h3b42c579),
	.w3(32'h3c3b2749),
	.w4(32'h3cc80b59),
	.w5(32'hbb55ed93),
	.w6(32'h3c8b5d6e),
	.w7(32'h3c4b5484),
	.w8(32'hbb8c56f5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c463),
	.w1(32'hbb4b28d4),
	.w2(32'hbc0d1cef),
	.w3(32'h3b8c6726),
	.w4(32'hbbaf5a7f),
	.w5(32'hbc109044),
	.w6(32'h3c8e31cf),
	.w7(32'h3bd63527),
	.w8(32'hbbf5bb7e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace59a3),
	.w1(32'hba9ff159),
	.w2(32'h3b9ba5db),
	.w3(32'hbb2d55b1),
	.w4(32'h3ac17de2),
	.w5(32'h3b61b654),
	.w6(32'h3bddac37),
	.w7(32'h3bc870e0),
	.w8(32'hbaadccce),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89f6cf),
	.w1(32'hbb6142d0),
	.w2(32'h3c2aeda9),
	.w3(32'hbba23739),
	.w4(32'hba877813),
	.w5(32'h3c2a8e26),
	.w6(32'hb953254b),
	.w7(32'hba46d867),
	.w8(32'hbbb8bf83),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e3eab),
	.w1(32'h3ad18d64),
	.w2(32'hbb5b0d69),
	.w3(32'h3a79a3b8),
	.w4(32'hbb8e21c8),
	.w5(32'h3b9b404d),
	.w6(32'h3b372ba6),
	.w7(32'h3b2b091d),
	.w8(32'hb9f2da5a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7909dc),
	.w1(32'h3a478c11),
	.w2(32'hbbbe2732),
	.w3(32'hbaf34c7c),
	.w4(32'hba5e180e),
	.w5(32'hbbdc9ed9),
	.w6(32'hbba69c6c),
	.w7(32'hba9ce304),
	.w8(32'h3a588320),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd4dff),
	.w1(32'h39ef20e0),
	.w2(32'hbc4b9ced),
	.w3(32'h3ade4b15),
	.w4(32'hbb447d8e),
	.w5(32'hbc138245),
	.w6(32'hbab28418),
	.w7(32'hbb5210f3),
	.w8(32'hbaaef94d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59fadb),
	.w1(32'h3c5332c8),
	.w2(32'hbc4a93ea),
	.w3(32'h3c058eb5),
	.w4(32'h3bad2e8f),
	.w5(32'hbb951155),
	.w6(32'h3a578d02),
	.w7(32'h3bd142e2),
	.w8(32'h3c80e7cf),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc663e16),
	.w1(32'hbba04309),
	.w2(32'hbc581c4e),
	.w3(32'hb9b9f924),
	.w4(32'h3b49cc24),
	.w5(32'hbbbe8f47),
	.w6(32'h3c36879a),
	.w7(32'h3b6baf4f),
	.w8(32'hbaae273a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc747c1a),
	.w1(32'hbbca0484),
	.w2(32'h3b1200b8),
	.w3(32'hbbb276b7),
	.w4(32'hbc2ea4dd),
	.w5(32'hbab4a4ce),
	.w6(32'hbc3b52e0),
	.w7(32'hbc6941f7),
	.w8(32'hbb7d578c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac1fa),
	.w1(32'hba308bab),
	.w2(32'hbc006228),
	.w3(32'hbac8351d),
	.w4(32'hbb735b0c),
	.w5(32'h3c74efb8),
	.w6(32'h3b3af88d),
	.w7(32'h39cce2bb),
	.w8(32'h3cf5877e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8678f8),
	.w1(32'h3c23892d),
	.w2(32'hbc6b3ef0),
	.w3(32'h3d050cff),
	.w4(32'hb9f38daf),
	.w5(32'hbc54ad4a),
	.w6(32'h3c5f0619),
	.w7(32'hbb1e1237),
	.w8(32'h3c7962b3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41cca2),
	.w1(32'hbc328bde),
	.w2(32'hbbe6ba8f),
	.w3(32'hbbc34374),
	.w4(32'hbb76c857),
	.w5(32'h3b8f3b4d),
	.w6(32'h3c6fb36a),
	.w7(32'h3bec8304),
	.w8(32'h3c7b1a56),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcda0d),
	.w1(32'h3bb0f050),
	.w2(32'h3b1a465a),
	.w3(32'h3bb1d196),
	.w4(32'h3a23d98b),
	.w5(32'h3af01854),
	.w6(32'h3a8c19d3),
	.w7(32'hbb47dfd3),
	.w8(32'h3b199fd6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474bfa),
	.w1(32'hbb9266b4),
	.w2(32'hb829cb55),
	.w3(32'hbad9d850),
	.w4(32'hbc113f69),
	.w5(32'hbc0b18cb),
	.w6(32'hbb6451b0),
	.w7(32'hbb950560),
	.w8(32'hbc074160),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a2236),
	.w1(32'hbb113e7e),
	.w2(32'hbafac9aa),
	.w3(32'hbb096e9d),
	.w4(32'hbb29409e),
	.w5(32'h3bc6989f),
	.w6(32'hbba34fee),
	.w7(32'hba93e2cc),
	.w8(32'h37365899),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8f05c),
	.w1(32'h3aad12c4),
	.w2(32'h3b827ebf),
	.w3(32'h3b7aa742),
	.w4(32'hb9be224d),
	.w5(32'h3b845a46),
	.w6(32'hba03b6e3),
	.w7(32'hba4f6aee),
	.w8(32'h3ae1ab70),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b5815),
	.w1(32'h3b7b175c),
	.w2(32'hbc500c1b),
	.w3(32'h3b99a3fb),
	.w4(32'hbae6115a),
	.w5(32'hbc88a69f),
	.w6(32'hbc23d309),
	.w7(32'hbaeec8b2),
	.w8(32'h3c73c343),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafef1e),
	.w1(32'hbb82c867),
	.w2(32'hb99cc57d),
	.w3(32'hbc01ec04),
	.w4(32'h3c902d7c),
	.w5(32'hbbb23d2a),
	.w6(32'h3c8ff2e8),
	.w7(32'h3c58fdba),
	.w8(32'h3bd7cb26),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69a5d9),
	.w1(32'hbb8e7e5f),
	.w2(32'hbad8ddf1),
	.w3(32'h39f34a28),
	.w4(32'hbc160d21),
	.w5(32'hb985d314),
	.w6(32'h3a8de4fe),
	.w7(32'hbc18f4ea),
	.w8(32'h3876e3bd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28e97f),
	.w1(32'h3b39298d),
	.w2(32'hbb878d76),
	.w3(32'hb985db59),
	.w4(32'h3ac89536),
	.w5(32'hbb8ce48b),
	.w6(32'hba2722cb),
	.w7(32'h3a740c47),
	.w8(32'hbb2dfbd2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc0ff),
	.w1(32'hbb1a9f83),
	.w2(32'h3b520724),
	.w3(32'hbb923afc),
	.w4(32'hbaba3029),
	.w5(32'h3be153ca),
	.w6(32'hbbb96d75),
	.w7(32'hbba4be95),
	.w8(32'h3b992691),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc691e77),
	.w1(32'h3b36ba9d),
	.w2(32'hbbe35bf5),
	.w3(32'hbc4cc7cc),
	.w4(32'h3b212c25),
	.w5(32'hbab74467),
	.w6(32'hbc25e6cc),
	.w7(32'h3b9b99ab),
	.w8(32'h3a6d8673),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a48d2),
	.w1(32'h3b839ec1),
	.w2(32'h3c3fd63c),
	.w3(32'h398766cc),
	.w4(32'h3b5ab6d0),
	.w5(32'h3ca7456d),
	.w6(32'h3b89da0e),
	.w7(32'h3ba9fefe),
	.w8(32'h3ac643ef),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3982f3),
	.w1(32'hbc30006e),
	.w2(32'h3a8633ed),
	.w3(32'hbc593183),
	.w4(32'hbc659c3a),
	.w5(32'h3b8b3307),
	.w6(32'hbc36376c),
	.w7(32'h3c48ec3b),
	.w8(32'h3bf52acf),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb55c4d),
	.w1(32'h3b912f28),
	.w2(32'hbbae0154),
	.w3(32'hbc157b46),
	.w4(32'h3c568585),
	.w5(32'hbc8506dd),
	.w6(32'h3bb50683),
	.w7(32'h3c5835cb),
	.w8(32'h3b806340),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc209091),
	.w1(32'h3c03b132),
	.w2(32'h3ae0801e),
	.w3(32'h3b201df6),
	.w4(32'h3c9cf776),
	.w5(32'hbbdce100),
	.w6(32'h3c224a0f),
	.w7(32'h3c1d25a7),
	.w8(32'h3c1afa20),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule