module layer_10_featuremap_334(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77e9ca),
	.w1(32'hbb4b6f7d),
	.w2(32'hbb3c9eb3),
	.w3(32'hbafa43f7),
	.w4(32'hb9c2cf94),
	.w5(32'hba0b5cbf),
	.w6(32'hbc61c95a),
	.w7(32'hbc52ad4c),
	.w8(32'hb93849fa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30c7b6),
	.w1(32'hbaca1d03),
	.w2(32'hbb45e70e),
	.w3(32'hbbb1ff13),
	.w4(32'hbb8629af),
	.w5(32'hbb1388a3),
	.w6(32'h3c01d664),
	.w7(32'h3b904b04),
	.w8(32'h3c560f3e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefa0b7),
	.w1(32'h3bcc8504),
	.w2(32'h3a90b404),
	.w3(32'h3ba06e7f),
	.w4(32'hbb27dda8),
	.w5(32'hba90e2d3),
	.w6(32'h3c7e4b39),
	.w7(32'h3c768bc2),
	.w8(32'h3a0db753),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae23f50),
	.w1(32'hbaf8a650),
	.w2(32'hb9851222),
	.w3(32'hbb228bdb),
	.w4(32'hbb5680ca),
	.w5(32'h3abe0337),
	.w6(32'h3c38037b),
	.w7(32'h3ac60717),
	.w8(32'hba8cdd5b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fecdc),
	.w1(32'h3a3fa19c),
	.w2(32'hba4cc7c1),
	.w3(32'hbb5abb20),
	.w4(32'hbbd7a7bd),
	.w5(32'h3b14a2e0),
	.w6(32'h3b3a885c),
	.w7(32'hbb7b6bb9),
	.w8(32'h3a71ee80),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe5d95),
	.w1(32'h395c4dc6),
	.w2(32'hba82ad0b),
	.w3(32'h3aaa7c84),
	.w4(32'h3b3c375d),
	.w5(32'hbafda1e6),
	.w6(32'hb989af8c),
	.w7(32'hba2c7512),
	.w8(32'hbb129700),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695d0e),
	.w1(32'hba1c831d),
	.w2(32'h39e222a5),
	.w3(32'hbafdd9e4),
	.w4(32'hbb01bed5),
	.w5(32'hbaa78918),
	.w6(32'h3b4dc610),
	.w7(32'hbaa75803),
	.w8(32'hbb965cc5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b206),
	.w1(32'hbc38f078),
	.w2(32'hbc1ec42e),
	.w3(32'hbb1e106f),
	.w4(32'hbb15afc6),
	.w5(32'hbaf92f63),
	.w6(32'hbbc513e1),
	.w7(32'hbc159687),
	.w8(32'hbbd6a9b5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b9513),
	.w1(32'hbb80b334),
	.w2(32'hbb264943),
	.w3(32'hbb70c1b3),
	.w4(32'hba1968dc),
	.w5(32'h3b9fc283),
	.w6(32'hbc13610c),
	.w7(32'hbb9504fb),
	.w8(32'h3b572545),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d9fd6),
	.w1(32'h3ab6e9f7),
	.w2(32'h3abd7a0b),
	.w3(32'h3b5faa8e),
	.w4(32'h3b87d224),
	.w5(32'hb95486ac),
	.w6(32'h3aaafddd),
	.w7(32'h3a1a7104),
	.w8(32'hbace8e28),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cef28),
	.w1(32'h3b63b459),
	.w2(32'h3a7416af),
	.w3(32'hbb3dac10),
	.w4(32'hba8b60b3),
	.w5(32'h3b0ee4ee),
	.w6(32'h3b56bac3),
	.w7(32'hbb18772f),
	.w8(32'h3ae334a4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74fbf3),
	.w1(32'h3b5d23d5),
	.w2(32'h3bef019e),
	.w3(32'hba9c1f90),
	.w4(32'hba20d2c7),
	.w5(32'h3be97f54),
	.w6(32'h3c024a6a),
	.w7(32'h3bd8d6f6),
	.w8(32'hbc3e6ac2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10b593),
	.w1(32'hbb393c71),
	.w2(32'h38858b98),
	.w3(32'hbae57b06),
	.w4(32'h3b49556a),
	.w5(32'h39f9921a),
	.w6(32'h37c8aa56),
	.w7(32'hba416f9a),
	.w8(32'hbb41d378),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840398),
	.w1(32'hbbd47c37),
	.w2(32'h3a0a314f),
	.w3(32'h3a6f379e),
	.w4(32'h3a8dbb26),
	.w5(32'hbbf66173),
	.w6(32'hbb07fccb),
	.w7(32'h3a8950d6),
	.w8(32'hbb0b47e1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81088f),
	.w1(32'hbb4f4fd0),
	.w2(32'hb9028f92),
	.w3(32'hbb88671e),
	.w4(32'hbbb1ddde),
	.w5(32'hbb3f36fb),
	.w6(32'h3c0b51c0),
	.w7(32'h3a045c88),
	.w8(32'hbb17377f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fd244),
	.w1(32'hbb0093b5),
	.w2(32'hbbadbea6),
	.w3(32'hbb562b69),
	.w4(32'hbb15e937),
	.w5(32'h3a435c62),
	.w6(32'hba8f0a26),
	.w7(32'hbb9a24f1),
	.w8(32'hbc187dfd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9345fe),
	.w1(32'hbbfdc8f1),
	.w2(32'hbc0bd525),
	.w3(32'hbb93561f),
	.w4(32'hba661f6e),
	.w5(32'hbac13c24),
	.w6(32'hbbe7536b),
	.w7(32'hbbc2a0ef),
	.w8(32'hbb35f146),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc61602),
	.w1(32'h3a823a3d),
	.w2(32'hbb13e00c),
	.w3(32'hbb44b4e1),
	.w4(32'hbb5688d4),
	.w5(32'h3ac39a7b),
	.w6(32'h3b26797e),
	.w7(32'hbba613de),
	.w8(32'h3bbb841a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1529d),
	.w1(32'h3b8cff86),
	.w2(32'h39a8730b),
	.w3(32'h3b9ebb90),
	.w4(32'hba0b24aa),
	.w5(32'hba64bf26),
	.w6(32'h3ba832dd),
	.w7(32'h3ad4f1b3),
	.w8(32'hba5c55fb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baaada),
	.w1(32'hbba3aa22),
	.w2(32'hbabcdc21),
	.w3(32'h377b75de),
	.w4(32'hbbb1d41e),
	.w5(32'hbb9dbb70),
	.w6(32'h37f8703c),
	.w7(32'hbbcea258),
	.w8(32'hbb65f8cc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f9270),
	.w1(32'hbaef0171),
	.w2(32'hbbe0df8f),
	.w3(32'hbb91c4fa),
	.w4(32'hbb216c75),
	.w5(32'hba672b75),
	.w6(32'h39972481),
	.w7(32'hbad8032f),
	.w8(32'hbb240009),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4184cb),
	.w1(32'hbae20c54),
	.w2(32'h397c1573),
	.w3(32'hba638809),
	.w4(32'h3a1de776),
	.w5(32'h3a5f5106),
	.w6(32'hbb9937ea),
	.w7(32'hbb4b6ea4),
	.w8(32'h3aa4301f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7543c8),
	.w1(32'h3b4a3e99),
	.w2(32'h39ab9a95),
	.w3(32'hba80c53c),
	.w4(32'hbad34732),
	.w5(32'hbb9c600f),
	.w6(32'h3b073664),
	.w7(32'h3aaf0a07),
	.w8(32'hbb9ec5e6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124a20),
	.w1(32'hbb718f5d),
	.w2(32'hbb4ebe90),
	.w3(32'hbbd7958c),
	.w4(32'hbbbaaecc),
	.w5(32'hbb8cc999),
	.w6(32'hbbabca4e),
	.w7(32'hbbe416d7),
	.w8(32'h399a6ef5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3377d7),
	.w1(32'h3ba72968),
	.w2(32'h39af2e69),
	.w3(32'hb954d75f),
	.w4(32'hbadfae69),
	.w5(32'h3b290762),
	.w6(32'hbba1e61a),
	.w7(32'h3a02b786),
	.w8(32'hba9101bf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70b129),
	.w1(32'h3b88fa09),
	.w2(32'h3b913f9d),
	.w3(32'h3b226d22),
	.w4(32'h3b4accfa),
	.w5(32'h3c07b30a),
	.w6(32'hb997dc1e),
	.w7(32'hbb6c830b),
	.w8(32'h3b9b8e5f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2449),
	.w1(32'hba705624),
	.w2(32'hba3402f5),
	.w3(32'h3b05a3a8),
	.w4(32'h3bc51398),
	.w5(32'h3adabe22),
	.w6(32'hb9fe141d),
	.w7(32'h3c06c3e4),
	.w8(32'hbb9230ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b25f12),
	.w1(32'hbb3d8b5b),
	.w2(32'hbb1f3a1e),
	.w3(32'hba956618),
	.w4(32'h3a7c2dea),
	.w5(32'h3bcd5101),
	.w6(32'hbc4367d8),
	.w7(32'hbc00dd58),
	.w8(32'h3a1bca3f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e6c65),
	.w1(32'hbaa68b92),
	.w2(32'hbb5336a4),
	.w3(32'hbb24da4f),
	.w4(32'h3aa55fdd),
	.w5(32'hba88c4a9),
	.w6(32'h3aeacd56),
	.w7(32'h3a480483),
	.w8(32'hbb7bea71),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95455e),
	.w1(32'hbb6f5e31),
	.w2(32'hbbbd5af0),
	.w3(32'hbb10ab59),
	.w4(32'hba35cbcc),
	.w5(32'hbbfe07b9),
	.w6(32'hb9f253e8),
	.w7(32'hbb25510a),
	.w8(32'h3b94c28c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23609c),
	.w1(32'hba737e0c),
	.w2(32'hbb87ea6a),
	.w3(32'h3a16f080),
	.w4(32'hbc42cc66),
	.w5(32'h3a954e73),
	.w6(32'hbc2950f7),
	.w7(32'hbb771dcc),
	.w8(32'h3883a521),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851c5d),
	.w1(32'h3bbd3c1e),
	.w2(32'h3bd606e2),
	.w3(32'hbbd768f1),
	.w4(32'h3a97b7f1),
	.w5(32'h3b9a24ec),
	.w6(32'h3c06e28f),
	.w7(32'h39d68cf4),
	.w8(32'hbbb6a671),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae708d9),
	.w1(32'hb99f683d),
	.w2(32'h3abce3ae),
	.w3(32'h3ba92a36),
	.w4(32'hb9691c21),
	.w5(32'h394198a1),
	.w6(32'hbc240cdb),
	.w7(32'hbbf6703f),
	.w8(32'hbb30ae73),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37258e),
	.w1(32'h3b0c7e81),
	.w2(32'hbb92cd2b),
	.w3(32'hbbb9f517),
	.w4(32'hbbca317e),
	.w5(32'hba5a6208),
	.w6(32'h3b24a3fa),
	.w7(32'hbc0e44f6),
	.w8(32'hb8b5aa6d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0364e),
	.w1(32'h3a89ddc8),
	.w2(32'h3a83c820),
	.w3(32'h37ee876d),
	.w4(32'h3b3db983),
	.w5(32'hbbbb7346),
	.w6(32'h3ba23f62),
	.w7(32'hbaeacd8a),
	.w8(32'h3c190692),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b1dc0),
	.w1(32'h3bf80990),
	.w2(32'h3ad2185e),
	.w3(32'hbb58dcee),
	.w4(32'hbc09a969),
	.w5(32'h3bb51029),
	.w6(32'h3b9f05d3),
	.w7(32'hba108c6a),
	.w8(32'hbba798cc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d031),
	.w1(32'h3a8bbf15),
	.w2(32'h3a63d059),
	.w3(32'h3cbf5a09),
	.w4(32'h3c226a5d),
	.w5(32'h3ab3316d),
	.w6(32'hbc9273a4),
	.w7(32'hbb756684),
	.w8(32'h3b692b22),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64dd46),
	.w1(32'h3ae46978),
	.w2(32'h3a705db0),
	.w3(32'h3bbe2f28),
	.w4(32'h3c372985),
	.w5(32'h3b45c891),
	.w6(32'hbbe82e5a),
	.w7(32'h3c788fa5),
	.w8(32'h3bb8c9e3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d92a2b),
	.w1(32'h3ba2b2c9),
	.w2(32'h3b4b9530),
	.w3(32'h3b0fa53e),
	.w4(32'h3a7b37ea),
	.w5(32'h3b5ec6bd),
	.w6(32'h3bd228e2),
	.w7(32'h3c08a01b),
	.w8(32'h3a630a52),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabaec5),
	.w1(32'hbb3d5554),
	.w2(32'hbb90b8a6),
	.w3(32'hb8da4f89),
	.w4(32'hbb037161),
	.w5(32'h3add3351),
	.w6(32'hbc447c64),
	.w7(32'hbc0bad7e),
	.w8(32'hbb6eb0a6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b959a9a),
	.w1(32'hbaebb351),
	.w2(32'h3bb1feff),
	.w3(32'hb88f640e),
	.w4(32'h3bcdbae5),
	.w5(32'h3a9c49a8),
	.w6(32'h3bdd8414),
	.w7(32'h3b01ddc0),
	.w8(32'h3b0b0d9d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfd419),
	.w1(32'h3b17cd70),
	.w2(32'h3b6c21be),
	.w3(32'h3b82e3aa),
	.w4(32'h3b7e054b),
	.w5(32'h3a5921c2),
	.w6(32'h3b94f4e4),
	.w7(32'h3b93f2e9),
	.w8(32'h3bb6e321),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14cb91),
	.w1(32'hbb1397bf),
	.w2(32'h3ab699d0),
	.w3(32'h3bfaa6ec),
	.w4(32'h3b36f717),
	.w5(32'hbc19e8b4),
	.w6(32'h3cbc03c5),
	.w7(32'h3c7cc657),
	.w8(32'hbaac145c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cd9fb),
	.w1(32'h3a1efc48),
	.w2(32'hbbc747d3),
	.w3(32'hbbb90b3b),
	.w4(32'hbbe206d2),
	.w5(32'hbb4913d4),
	.w6(32'h3cb71d69),
	.w7(32'h3ab95add),
	.w8(32'hb9104a78),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eeb80),
	.w1(32'hba61f965),
	.w2(32'hb9a02d7d),
	.w3(32'hba6ecd6f),
	.w4(32'h3a90c6ee),
	.w5(32'hbb151b4b),
	.w6(32'hbc1d7f9a),
	.w7(32'hbc026e21),
	.w8(32'hbb376df8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5d00),
	.w1(32'h3b148b81),
	.w2(32'hbaf57fbf),
	.w3(32'hbb98da4b),
	.w4(32'hbbc44886),
	.w5(32'h3bafa9bc),
	.w6(32'hbba94e9e),
	.w7(32'hbb776708),
	.w8(32'hba97e86f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f6c77),
	.w1(32'h3c083218),
	.w2(32'h3b9cba22),
	.w3(32'h3aedf30a),
	.w4(32'h3aaefd0f),
	.w5(32'h3aaa64ce),
	.w6(32'hbb61e8a7),
	.w7(32'hbaea8728),
	.w8(32'hbb01a4a3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30241c),
	.w1(32'h38c77cf3),
	.w2(32'h3b7b527a),
	.w3(32'h394e9d00),
	.w4(32'h3b6e8914),
	.w5(32'h3b61fa50),
	.w6(32'hbb735a5b),
	.w7(32'h3b25f102),
	.w8(32'hba32611c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06efe7),
	.w1(32'h3a57c1e5),
	.w2(32'h3b081716),
	.w3(32'h3a01f7ee),
	.w4(32'hb9f625b6),
	.w5(32'hbb55d423),
	.w6(32'h3a8dbe88),
	.w7(32'h3b706059),
	.w8(32'hbb278df8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53bc61),
	.w1(32'hbad34451),
	.w2(32'h395fd5bb),
	.w3(32'h3abbda11),
	.w4(32'h3aa11f70),
	.w5(32'h3bd62cd4),
	.w6(32'hbb62e34f),
	.w7(32'hbb435548),
	.w8(32'h3a86bead),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a4aec),
	.w1(32'hba0ff32a),
	.w2(32'hbb989c59),
	.w3(32'h3b413ba6),
	.w4(32'hbbd28951),
	.w5(32'h3bde9d90),
	.w6(32'hbb94fadc),
	.w7(32'hbc3670af),
	.w8(32'h3bfb4c48),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f25fd),
	.w1(32'hbb892a51),
	.w2(32'hba9b8ae4),
	.w3(32'hbb77f481),
	.w4(32'h3b919526),
	.w5(32'hbb1ff4e6),
	.w6(32'h3cb62ba7),
	.w7(32'h3c2c9125),
	.w8(32'hbbc176a5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8c24),
	.w1(32'hba4b3919),
	.w2(32'hbb564bbd),
	.w3(32'hbabd241e),
	.w4(32'hbb1e9d22),
	.w5(32'h3aee3951),
	.w6(32'h3b4f1cea),
	.w7(32'hba6e5658),
	.w8(32'h3a9f3c4f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c161651),
	.w1(32'h3b6217e7),
	.w2(32'hbb90778d),
	.w3(32'hbbb8087f),
	.w4(32'hbbb80dd2),
	.w5(32'h39b5b62a),
	.w6(32'hbbd61a5d),
	.w7(32'hbc85bb6e),
	.w8(32'h3b581d1c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c948),
	.w1(32'h3b8dc4ef),
	.w2(32'hb98fd35f),
	.w3(32'hbad248fb),
	.w4(32'hba78bee9),
	.w5(32'hbb363306),
	.w6(32'h39c78ab5),
	.w7(32'hbba0d264),
	.w8(32'hbb089717),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5247a3),
	.w1(32'hba98e4b7),
	.w2(32'hba9763db),
	.w3(32'hbb23480e),
	.w4(32'h3a36a1df),
	.w5(32'hbb268f10),
	.w6(32'h3a3b4e43),
	.w7(32'hbc3066fc),
	.w8(32'hbb6ce013),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5ae2),
	.w1(32'hbab6012e),
	.w2(32'h3b763948),
	.w3(32'hba0a3d49),
	.w4(32'h3b2fe0c3),
	.w5(32'hbb2eaba7),
	.w6(32'hb9a0c5a1),
	.w7(32'hb9e603b1),
	.w8(32'hbb28d01a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b922941),
	.w1(32'hba912ed5),
	.w2(32'h3b0caf8e),
	.w3(32'hbbd73406),
	.w4(32'h3bb153af),
	.w5(32'hbb9cb189),
	.w6(32'hbb67e72f),
	.w7(32'hbbaca605),
	.w8(32'hbb0377ef),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fda12),
	.w1(32'hb9d0da4c),
	.w2(32'h3b553ce9),
	.w3(32'h396b22b0),
	.w4(32'h3a51fef2),
	.w5(32'h3c485a4b),
	.w6(32'hbb033791),
	.w7(32'hbb2c2498),
	.w8(32'h3b8b2367),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9feef3),
	.w1(32'h3c52792f),
	.w2(32'h3c35ecc7),
	.w3(32'h3b516924),
	.w4(32'h3c878e08),
	.w5(32'h3abaa879),
	.w6(32'hbc81f2b7),
	.w7(32'h3c4a8729),
	.w8(32'h3aa604a1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa76773),
	.w1(32'hbae60466),
	.w2(32'hbb023bdb),
	.w3(32'h38fc09f4),
	.w4(32'hbb43bcc5),
	.w5(32'hbb2354b7),
	.w6(32'h3b6344d5),
	.w7(32'h3b0c6fa3),
	.w8(32'hbb7f1edd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17bbe6),
	.w1(32'hbbb7ee3c),
	.w2(32'hbbcdfcbd),
	.w3(32'hbb07b682),
	.w4(32'hbbc7345c),
	.w5(32'hb974511e),
	.w6(32'h3ac2ea1b),
	.w7(32'hbbcbeeca),
	.w8(32'hbba491d1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3402),
	.w1(32'h3aa57106),
	.w2(32'hbabe32a1),
	.w3(32'h3b3285e9),
	.w4(32'h3bac1200),
	.w5(32'hbaec7433),
	.w6(32'h3b6d35db),
	.w7(32'h39bb7ac0),
	.w8(32'hbaa2343d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83767),
	.w1(32'h3a3a6b18),
	.w2(32'h3b90e626),
	.w3(32'h3ace092b),
	.w4(32'h3a66415a),
	.w5(32'hbb5de15a),
	.w6(32'h3bbe0b24),
	.w7(32'hbb080151),
	.w8(32'hbb4b27b4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac249a),
	.w1(32'hbbd3ca66),
	.w2(32'hbb6b5167),
	.w3(32'h3a6b072a),
	.w4(32'h398aee04),
	.w5(32'hbbad607a),
	.w6(32'h3b160b36),
	.w7(32'hbc3f63e6),
	.w8(32'h3b98eec4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95bfca),
	.w1(32'h3c2297a3),
	.w2(32'h3b9670e1),
	.w3(32'hbb799e76),
	.w4(32'h3b891e0d),
	.w5(32'hbb2a0af4),
	.w6(32'h3bd7af26),
	.w7(32'hbb10a115),
	.w8(32'hbb16507c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f719),
	.w1(32'hbbb21bf0),
	.w2(32'hbbd51fa6),
	.w3(32'hbba94160),
	.w4(32'hbbe3d2b2),
	.w5(32'h3b395f76),
	.w6(32'hba755ac2),
	.w7(32'hbbd96ae8),
	.w8(32'h3b5da053),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9df67),
	.w1(32'hbadbbcd0),
	.w2(32'h3aaa17ba),
	.w3(32'h3b21bdcd),
	.w4(32'h3aff449a),
	.w5(32'h3b995046),
	.w6(32'h3bb5141f),
	.w7(32'h3c0f6053),
	.w8(32'h3bc2e2e7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0efbfb),
	.w1(32'hbb370e58),
	.w2(32'hb9eb9eec),
	.w3(32'hb9b4e10d),
	.w4(32'hbb5a0baa),
	.w5(32'h3af9d914),
	.w6(32'hbba3092b),
	.w7(32'hbb6e5582),
	.w8(32'hbb097579),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37c62),
	.w1(32'h3b924501),
	.w2(32'h3a6b8ef9),
	.w3(32'hbaf7a6e8),
	.w4(32'h3b5f419e),
	.w5(32'h3b9575d8),
	.w6(32'h392831b4),
	.w7(32'hba95ac8e),
	.w8(32'h3b1602f5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bc47d),
	.w1(32'h3b7ce658),
	.w2(32'h3bb4611e),
	.w3(32'h3c79633a),
	.w4(32'h3c09a404),
	.w5(32'hbb414825),
	.w6(32'h3a28d68a),
	.w7(32'h3bf9a4b7),
	.w8(32'hbbbb94cb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63244e),
	.w1(32'hba626595),
	.w2(32'h3a79bcda),
	.w3(32'hbb79f8f1),
	.w4(32'hbadb492e),
	.w5(32'h3b837470),
	.w6(32'hbbcd04e6),
	.w7(32'h3a4ae358),
	.w8(32'h3b949468),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296c43),
	.w1(32'h3bf5a2f0),
	.w2(32'h3bcaa08b),
	.w3(32'h3bd435e5),
	.w4(32'h3b97a3b1),
	.w5(32'hb903a576),
	.w6(32'h3b674d27),
	.w7(32'h3b5dc038),
	.w8(32'hbb59069d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59c89d),
	.w1(32'h39e8b84c),
	.w2(32'hbb8e4ed2),
	.w3(32'hbb7754ef),
	.w4(32'hbb187fea),
	.w5(32'hbad57474),
	.w6(32'hba9c962a),
	.w7(32'hb9ae56ef),
	.w8(32'hbb1f4e0e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167ca0),
	.w1(32'hbb9665d8),
	.w2(32'hbb879776),
	.w3(32'hbb8f2475),
	.w4(32'hba9bc5bf),
	.w5(32'hbb33df24),
	.w6(32'h3b0b7f4b),
	.w7(32'hbb986fcf),
	.w8(32'hbaaf2639),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc4a6),
	.w1(32'hb91cdf48),
	.w2(32'h3a9e0af9),
	.w3(32'hbbdab132),
	.w4(32'hba9faeb7),
	.w5(32'hbb1c34f2),
	.w6(32'h3b578e54),
	.w7(32'h3b5eb36d),
	.w8(32'hbac3f6b7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b884dcd),
	.w1(32'h3b0642de),
	.w2(32'h3b497c62),
	.w3(32'hbb275b0b),
	.w4(32'h3b0e6d38),
	.w5(32'hbc0407f5),
	.w6(32'hb8ec087e),
	.w7(32'hbb38289d),
	.w8(32'h3bad2543),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba31727),
	.w1(32'hbb7f4d31),
	.w2(32'hbbe0a31d),
	.w3(32'hbbe1dd04),
	.w4(32'hbb976a68),
	.w5(32'hbb02a226),
	.w6(32'h3b295089),
	.w7(32'hbb979ecc),
	.w8(32'hba6318f9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa4dc),
	.w1(32'hbb3a7c4f),
	.w2(32'hbb8d4140),
	.w3(32'hbbe9a959),
	.w4(32'hbc17fbac),
	.w5(32'hbb0d42a4),
	.w6(32'hbb904501),
	.w7(32'hbb690129),
	.w8(32'hbba3579f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f11e5),
	.w1(32'hbbac7a01),
	.w2(32'hbbd31ed8),
	.w3(32'hbbda2847),
	.w4(32'hbbd6cdb9),
	.w5(32'hbb88b541),
	.w6(32'hbb4d2e1e),
	.w7(32'hbbb967e3),
	.w8(32'hbba3c814),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29d31c),
	.w1(32'hbb56ab5a),
	.w2(32'hb9aee100),
	.w3(32'hbbe65eac),
	.w4(32'hbc16417a),
	.w5(32'hb9f9439d),
	.w6(32'hbbb65e25),
	.w7(32'hbc02c6b0),
	.w8(32'h3abfbb0e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee1939),
	.w1(32'hbb190972),
	.w2(32'hbb4ddc2b),
	.w3(32'hbbc4a885),
	.w4(32'hbb924ad1),
	.w5(32'hbb58b44d),
	.w6(32'hba843363),
	.w7(32'h3a4dffa4),
	.w8(32'hbb4b2afb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d56b),
	.w1(32'hbb1279a5),
	.w2(32'hbb7f9f35),
	.w3(32'hba3db160),
	.w4(32'hbbb8ba7d),
	.w5(32'h3c603ebe),
	.w6(32'hbb5084c2),
	.w7(32'hbbc22ec6),
	.w8(32'h3c25750f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4474),
	.w1(32'h3bf83da9),
	.w2(32'h3bd35e30),
	.w3(32'hb9dff306),
	.w4(32'h3c18e68c),
	.w5(32'hbb27e65f),
	.w6(32'h3b5553be),
	.w7(32'h3c675194),
	.w8(32'hbbbf6e4d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b600849),
	.w1(32'h3b9b1624),
	.w2(32'h3accd48d),
	.w3(32'h39add716),
	.w4(32'hbb8c5939),
	.w5(32'h3ab07f1f),
	.w6(32'hbb1e4f71),
	.w7(32'hba9a7cd0),
	.w8(32'h3ad24ec7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f678a),
	.w1(32'hbb8c7e21),
	.w2(32'hbbab4d7e),
	.w3(32'h3be2b20a),
	.w4(32'hbb0bfe43),
	.w5(32'hbb2bb86e),
	.w6(32'h3c092e29),
	.w7(32'h395957f2),
	.w8(32'hbb1e37e6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3806a),
	.w1(32'h3aed88f2),
	.w2(32'h3b418756),
	.w3(32'h3b8bc1ce),
	.w4(32'hbb41f006),
	.w5(32'h3a971ac3),
	.w6(32'h3a2625a3),
	.w7(32'hbaf86533),
	.w8(32'h3b88d76f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51276b),
	.w1(32'h3b38a5f3),
	.w2(32'h3ae52b83),
	.w3(32'h3a6f84fb),
	.w4(32'hb98b1e5a),
	.w5(32'hbae00c56),
	.w6(32'h3bd0105d),
	.w7(32'h3be68cdf),
	.w8(32'hbbb04252),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2d06e),
	.w1(32'hbb744ba5),
	.w2(32'hbb85c04b),
	.w3(32'hbb9de9c8),
	.w4(32'hbb07edcf),
	.w5(32'h3a8a8704),
	.w6(32'hbae515c4),
	.w7(32'hbb9fd3fd),
	.w8(32'hbbabbda6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acab82b),
	.w1(32'hbb56db31),
	.w2(32'h3b3a6d41),
	.w3(32'hbc35c3a6),
	.w4(32'hbbcf6c3e),
	.w5(32'hbb0ddd9f),
	.w6(32'hbbb274c9),
	.w7(32'hbc0e7517),
	.w8(32'h39bb6cb1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b170198),
	.w1(32'h3b8260e9),
	.w2(32'h3b454930),
	.w3(32'hbb83429e),
	.w4(32'hbb6ce2a0),
	.w5(32'h3ab6e30c),
	.w6(32'hbb994274),
	.w7(32'hbb9fb8b7),
	.w8(32'h3b621136),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2efe3a),
	.w1(32'hbb2f0160),
	.w2(32'h3be38e2c),
	.w3(32'hbb2e7e12),
	.w4(32'h3bce3b6b),
	.w5(32'hbab44a61),
	.w6(32'h3bb489f8),
	.w7(32'hbb5d54b8),
	.w8(32'hbbbb7140),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42b78),
	.w1(32'hbbce2ad6),
	.w2(32'hbc1f5bc1),
	.w3(32'hbb2c072a),
	.w4(32'hbb323881),
	.w5(32'h3c227632),
	.w6(32'h3ba08948),
	.w7(32'hbb72b626),
	.w8(32'h3c6270d5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae269d),
	.w1(32'hbb756690),
	.w2(32'hbb127d3d),
	.w3(32'hbabe8520),
	.w4(32'hba2e937b),
	.w5(32'h3a47c9c4),
	.w6(32'h3c2ed51a),
	.w7(32'h3c380701),
	.w8(32'h3a45100b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95939),
	.w1(32'hba21fef4),
	.w2(32'h39b5fc82),
	.w3(32'h3ab15a3b),
	.w4(32'h3b19346d),
	.w5(32'hba0f9cef),
	.w6(32'hbc015cf3),
	.w7(32'hba334d49),
	.w8(32'h3c26d91a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60317c),
	.w1(32'hbc4b420d),
	.w2(32'hbbc302b1),
	.w3(32'hbc1e0d21),
	.w4(32'h3b081bb7),
	.w5(32'h3ad64518),
	.w6(32'h3d0142bf),
	.w7(32'h3c7b9a03),
	.w8(32'h3ba37289),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269e84),
	.w1(32'h3bb9ebd3),
	.w2(32'h3b8add51),
	.w3(32'hbb6aa828),
	.w4(32'hbaba20a1),
	.w5(32'h3befa185),
	.w6(32'hbbdab9e8),
	.w7(32'h3aada69e),
	.w8(32'hbc285e2e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba069131),
	.w1(32'hbbbcc69f),
	.w2(32'hba9622f3),
	.w3(32'h3b9d52d5),
	.w4(32'h3bacc5c9),
	.w5(32'h39ecb524),
	.w6(32'hbbb01e80),
	.w7(32'hbbecde4b),
	.w8(32'h3970818d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37de1ff9),
	.w1(32'hb85d0071),
	.w2(32'hb9e1d12d),
	.w3(32'hb9a8229d),
	.w4(32'hb9bbd1e4),
	.w5(32'h3a754a06),
	.w6(32'hba12d84a),
	.w7(32'hb9085ff6),
	.w8(32'hb984fb25),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42c5f),
	.w1(32'h3ac55757),
	.w2(32'h3a941e7f),
	.w3(32'h3a10566f),
	.w4(32'h3a64f53f),
	.w5(32'h3a6b4b1b),
	.w6(32'h3a59a5aa),
	.w7(32'h3a215255),
	.w8(32'h3a7793df),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376b489c),
	.w1(32'hb9582946),
	.w2(32'h39ccc881),
	.w3(32'h398ed3b3),
	.w4(32'h3a025ccd),
	.w5(32'h3a0ea8cc),
	.w6(32'hb9baf27e),
	.w7(32'h3a5259f9),
	.w8(32'h3a3e4cd1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef5e2f),
	.w1(32'hba283399),
	.w2(32'hba2d1983),
	.w3(32'h3aa13aab),
	.w4(32'h3a9eb3f8),
	.w5(32'hb9a4afa0),
	.w6(32'h3a822764),
	.w7(32'h39ef5a13),
	.w8(32'h390e5c95),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992790b),
	.w1(32'h38da69ae),
	.w2(32'hba249704),
	.w3(32'hba878e88),
	.w4(32'hba378517),
	.w5(32'hbb208750),
	.w6(32'hba59f233),
	.w7(32'hb9c4a445),
	.w8(32'hbb1069f8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a4897),
	.w1(32'hbb0648f3),
	.w2(32'hbaa8384d),
	.w3(32'hbb1db4ae),
	.w4(32'hbb187e21),
	.w5(32'h3afc3d61),
	.w6(32'hbb56df76),
	.w7(32'hbb085b45),
	.w8(32'h3b1561a0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2db332),
	.w1(32'h3a99cb8d),
	.w2(32'h39f473db),
	.w3(32'h3a00a675),
	.w4(32'h3a580256),
	.w5(32'h398c8849),
	.w6(32'h3a0f638b),
	.w7(32'h39e827a3),
	.w8(32'h394a1578),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8029515),
	.w1(32'h389002e0),
	.w2(32'hb8c8d219),
	.w3(32'h3a2f2d38),
	.w4(32'h39b03ecd),
	.w5(32'hb982071d),
	.w6(32'h3a0aee86),
	.w7(32'h394ec483),
	.w8(32'hba060687),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88fe80e),
	.w1(32'hb91ae3cb),
	.w2(32'hb880952c),
	.w3(32'hb803f153),
	.w4(32'hb963b9d9),
	.w5(32'h39a9ca3c),
	.w6(32'hba8f4e44),
	.w7(32'hba464b54),
	.w8(32'h39fb2d2c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6967f),
	.w1(32'h39b9ed29),
	.w2(32'hb9dc584f),
	.w3(32'h3a06ff8f),
	.w4(32'h39e03fff),
	.w5(32'h3ac91333),
	.w6(32'h3a16ef26),
	.w7(32'h3a135953),
	.w8(32'h3acbbe93),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad73794),
	.w1(32'h3a9aa79a),
	.w2(32'h3a9923dc),
	.w3(32'h3aac9978),
	.w4(32'h3ae08061),
	.w5(32'h3ab990cd),
	.w6(32'h3a46b981),
	.w7(32'h3ad6d0d9),
	.w8(32'h3a612c3c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d17fa6),
	.w1(32'h37932da2),
	.w2(32'h39c9f8ca),
	.w3(32'h3a30a38d),
	.w4(32'h3a7385e3),
	.w5(32'h39a29f8f),
	.w6(32'h39a23947),
	.w7(32'h3a3a3308),
	.w8(32'h38e613db),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b998f9),
	.w1(32'h3a29019d),
	.w2(32'h399da063),
	.w3(32'h39dbe82f),
	.w4(32'h39e87f71),
	.w5(32'hba1cdafb),
	.w6(32'h3a1468c9),
	.w7(32'h3a342112),
	.w8(32'hb982ab04),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f2d2d),
	.w1(32'h3a689bad),
	.w2(32'h38e86b78),
	.w3(32'h39340ab4),
	.w4(32'h394e87c5),
	.w5(32'hba35755c),
	.w6(32'h3986d025),
	.w7(32'h3a065f99),
	.w8(32'hb9e3b5dc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a7ac1),
	.w1(32'hba852afe),
	.w2(32'hba9b49a5),
	.w3(32'hbac1dfcf),
	.w4(32'hbacfa67c),
	.w5(32'hb92840e8),
	.w6(32'hba92ea8f),
	.w7(32'hbb006bcb),
	.w8(32'h3a594bd8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aec77),
	.w1(32'h38b1300f),
	.w2(32'hba1ce28b),
	.w3(32'hba0ae355),
	.w4(32'hba216393),
	.w5(32'h3ac38f72),
	.w6(32'h3a21d6bb),
	.w7(32'hb97d0bb2),
	.w8(32'h3a49c089),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fe598),
	.w1(32'h3a4837ef),
	.w2(32'h3a4ac5fb),
	.w3(32'h3afc7713),
	.w4(32'h3ab7ea8d),
	.w5(32'h3a1549c9),
	.w6(32'h3b02eda7),
	.w7(32'h3b0932f0),
	.w8(32'h39ec3bde),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02fa62),
	.w1(32'h3a547c0e),
	.w2(32'h390142e6),
	.w3(32'h3a640ec8),
	.w4(32'h3a906319),
	.w5(32'h3a15c0ea),
	.w6(32'h39abdb27),
	.w7(32'h3a6a4e18),
	.w8(32'h38e0ce8e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a32887),
	.w1(32'h3a3763e9),
	.w2(32'h3a817fdb),
	.w3(32'h3a29a147),
	.w4(32'h39854d0f),
	.w5(32'h3a59011a),
	.w6(32'h39eb3aa7),
	.w7(32'h3a15512d),
	.w8(32'h3af1b2f8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1fffc),
	.w1(32'h3a9d06e1),
	.w2(32'hb92e78de),
	.w3(32'h3aa034c0),
	.w4(32'h3a961172),
	.w5(32'h38f6389f),
	.w6(32'h3a6fc038),
	.w7(32'h3a7db4f0),
	.w8(32'hb9f0800f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2721b3),
	.w1(32'hba5325a2),
	.w2(32'hba065e32),
	.w3(32'hb98382a6),
	.w4(32'hba0793a1),
	.w5(32'h39c2a61d),
	.w6(32'hba7dc057),
	.w7(32'hb9ef99a8),
	.w8(32'h39c61305),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41b649),
	.w1(32'hba33c7cc),
	.w2(32'hba802050),
	.w3(32'h39d8d08e),
	.w4(32'hb92e6f96),
	.w5(32'hba0e03a3),
	.w6(32'hba41c6db),
	.w7(32'hba8f3ef0),
	.w8(32'hb9d5159a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943b242),
	.w1(32'h38d6e4f6),
	.w2(32'hb90ae0b6),
	.w3(32'hba06496c),
	.w4(32'hba1ebf07),
	.w5(32'h393ba498),
	.w6(32'hba7f44b2),
	.w7(32'hb9619f46),
	.w8(32'h36db5ab2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5721f),
	.w1(32'h390e6e5e),
	.w2(32'h3a06eca3),
	.w3(32'hb9d4d9d3),
	.w4(32'hba351d03),
	.w5(32'hb999a2f4),
	.w6(32'h38a4fe0b),
	.w7(32'hb916d0e6),
	.w8(32'hbab6300a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba329dad),
	.w1(32'hb9ca754b),
	.w2(32'hb9e5acd4),
	.w3(32'h399434cd),
	.w4(32'hb9418ff9),
	.w5(32'hba5c9115),
	.w6(32'hb9019689),
	.w7(32'hba07783c),
	.w8(32'hb9a26bd1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bb6b0),
	.w1(32'hb91d8e4f),
	.w2(32'hba1d9fef),
	.w3(32'hba500eb2),
	.w4(32'hba4dcd8c),
	.w5(32'h3a4823bf),
	.w6(32'h39cd0035),
	.w7(32'hba8abe25),
	.w8(32'hb9d8c88c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba633489),
	.w1(32'h399fd987),
	.w2(32'h39ae9307),
	.w3(32'h399aa0f5),
	.w4(32'h3a1ab4f2),
	.w5(32'h39c62a6a),
	.w6(32'h3a88983c),
	.w7(32'h39c2b575),
	.w8(32'h3a54cbcb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3f8a4),
	.w1(32'hb8f44f65),
	.w2(32'h38fdebc9),
	.w3(32'h36f6d725),
	.w4(32'hba0e78b3),
	.w5(32'h3a43aee9),
	.w6(32'h3a636a5f),
	.w7(32'hb8b4e716),
	.w8(32'hb795d92b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9c26e),
	.w1(32'h395c1074),
	.w2(32'h3a2a8066),
	.w3(32'h3a2c299b),
	.w4(32'h3a9278cf),
	.w5(32'h393da13b),
	.w6(32'h39e28f9e),
	.w7(32'h3a601501),
	.w8(32'h3a49b1d0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f29dc6),
	.w1(32'h3a5f4411),
	.w2(32'h3a116c19),
	.w3(32'hb91d4c20),
	.w4(32'hb82b108d),
	.w5(32'hb893c995),
	.w6(32'h3a27e477),
	.w7(32'h399f2128),
	.w8(32'hb83ac8ef),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983c70c),
	.w1(32'hb9db67f6),
	.w2(32'hb863ff0b),
	.w3(32'hb99d1658),
	.w4(32'h3a3b531a),
	.w5(32'hba7c7c24),
	.w6(32'hb99baaa4),
	.w7(32'hb7acad57),
	.w8(32'hba4e3338),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5be95e),
	.w1(32'hba619354),
	.w2(32'hba2c946c),
	.w3(32'hba91a481),
	.w4(32'hba6ed70e),
	.w5(32'hb9badb15),
	.w6(32'hba7d9cdf),
	.w7(32'hbaa1a964),
	.w8(32'hb9b7673b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930cbce),
	.w1(32'h38af0142),
	.w2(32'h3a5974fb),
	.w3(32'hb9718f1c),
	.w4(32'h391b5f36),
	.w5(32'h3994f21e),
	.w6(32'hba78b697),
	.w7(32'h3a380cad),
	.w8(32'h394d861f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a6d29),
	.w1(32'h379722af),
	.w2(32'h39c1444c),
	.w3(32'h39f2c7c0),
	.w4(32'h39bb2a5e),
	.w5(32'h3b37fe0d),
	.w6(32'h3a3109c5),
	.w7(32'h3a4396b1),
	.w8(32'h3a2ac679),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd0191),
	.w1(32'h3ada2ee5),
	.w2(32'h3b065596),
	.w3(32'h3b2bf296),
	.w4(32'h3b3aaec8),
	.w5(32'h3a56d6af),
	.w6(32'h3aa6bd89),
	.w7(32'h3ac1e0d6),
	.w8(32'h39edcd5b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a65ed7),
	.w1(32'h39138f88),
	.w2(32'h39e79826),
	.w3(32'h3a2b2d56),
	.w4(32'h3a6114bc),
	.w5(32'h39a87075),
	.w6(32'h3a072771),
	.w7(32'h3a3a20b6),
	.w8(32'h399f6db4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c85c6),
	.w1(32'h3a9ec9b0),
	.w2(32'h3aa0d045),
	.w3(32'hb81ce12b),
	.w4(32'h3a2980bd),
	.w5(32'hba3690a2),
	.w6(32'h39d3e7ba),
	.w7(32'h3a2931d2),
	.w8(32'hbaa85ba6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e446),
	.w1(32'hbb15c745),
	.w2(32'hba734aae),
	.w3(32'hba50e95a),
	.w4(32'hbad58d32),
	.w5(32'hbaa1c755),
	.w6(32'hbb06578c),
	.w7(32'hba9eafe6),
	.w8(32'hbaad3aa9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab54493),
	.w1(32'hbaa7a4fa),
	.w2(32'hba8fbe23),
	.w3(32'hba9a106c),
	.w4(32'hba8ce0e0),
	.w5(32'h3a93891a),
	.w6(32'hbaa8ee04),
	.w7(32'hba965615),
	.w8(32'h3a083036),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a36b7f),
	.w1(32'h39d30fdb),
	.w2(32'h3a375412),
	.w3(32'hb85457a3),
	.w4(32'h3a0dc472),
	.w5(32'h3a4594af),
	.w6(32'hb951d16e),
	.w7(32'h3a350e10),
	.w8(32'h3997258f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae597f),
	.w1(32'h3964aa52),
	.w2(32'h3997158c),
	.w3(32'h3a613f47),
	.w4(32'h3a579dc4),
	.w5(32'h38a05a29),
	.w6(32'h3a045c61),
	.w7(32'h3a16fe38),
	.w8(32'h3a0ec3d8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cbe2),
	.w1(32'h3a60a027),
	.w2(32'h3a745964),
	.w3(32'h36b4c651),
	.w4(32'hb96e5e7b),
	.w5(32'hba9adb88),
	.w6(32'hb9f78688),
	.w7(32'h3a3d3bdc),
	.w8(32'hbab6a6fb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d9e9b),
	.w1(32'hba29e198),
	.w2(32'hb9e60fa3),
	.w3(32'hba52975c),
	.w4(32'hba974a03),
	.w5(32'hb98a2563),
	.w6(32'hba8a28b6),
	.w7(32'hbab18343),
	.w8(32'hba4123ff),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7441bee),
	.w1(32'hb9d5b46e),
	.w2(32'h390d6323),
	.w3(32'hba105baa),
	.w4(32'hba877ea2),
	.w5(32'h395c0897),
	.w6(32'hb9f733d0),
	.w7(32'hb9dc7fa7),
	.w8(32'h39df7524),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a00fa5),
	.w1(32'h3a0c04eb),
	.w2(32'h39d9e0b3),
	.w3(32'h396f6cb5),
	.w4(32'h38a88d0d),
	.w5(32'h39a04f2b),
	.w6(32'h3a3da1b9),
	.w7(32'h39ddc59b),
	.w8(32'h3a0fcdad),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dbd7a),
	.w1(32'h39937a06),
	.w2(32'h3922b92d),
	.w3(32'h392e4990),
	.w4(32'h39dd9f84),
	.w5(32'hba437149),
	.w6(32'h3a4212cb),
	.w7(32'h39f368fa),
	.w8(32'hb9e23dc3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9010ef1),
	.w1(32'hba37f00e),
	.w2(32'hba15a39e),
	.w3(32'hb9f14730),
	.w4(32'h399d8bb3),
	.w5(32'hba2ea5f4),
	.w6(32'hb840b94f),
	.w7(32'h39a69977),
	.w8(32'hba2678d4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abdd7b),
	.w1(32'h3985192d),
	.w2(32'h39b274b0),
	.w3(32'h396e1a7e),
	.w4(32'hb928b48c),
	.w5(32'hba61512c),
	.w6(32'h39fa00af),
	.w7(32'h398efb6a),
	.w8(32'hba8ce379),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89f1a6),
	.w1(32'hbae2088d),
	.w2(32'hba98fda9),
	.w3(32'hba583d89),
	.w4(32'hba2035b6),
	.w5(32'hb990e2bb),
	.w6(32'hba931c05),
	.w7(32'hba6fe56f),
	.w8(32'h38a9a6ea),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6d0fb),
	.w1(32'h38809f0c),
	.w2(32'h3876b450),
	.w3(32'hb98e0067),
	.w4(32'hb9a3402e),
	.w5(32'h38bdd4eb),
	.w6(32'h3a80907d),
	.w7(32'h3817dd7f),
	.w8(32'h392d47fa),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec0e9c),
	.w1(32'hba62e349),
	.w2(32'h399f8cff),
	.w3(32'hb9ae2fcb),
	.w4(32'hb8109b9e),
	.w5(32'h3ade722f),
	.w6(32'h3a4df315),
	.w7(32'h3a1e29a6),
	.w8(32'h3ac63e54),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadf243),
	.w1(32'h3abeedbb),
	.w2(32'h3ae44cc6),
	.w3(32'h3ab92345),
	.w4(32'h3a9082d3),
	.w5(32'hb9d31341),
	.w6(32'h3ac66c61),
	.w7(32'h3ad43a76),
	.w8(32'h3985799e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f2edf),
	.w1(32'hb925d9f6),
	.w2(32'hb9ee4755),
	.w3(32'hba247cda),
	.w4(32'h377ebaff),
	.w5(32'hba1c5cfb),
	.w6(32'hb935ea5e),
	.w7(32'h385de23b),
	.w8(32'hb98ce991),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2ab3d),
	.w1(32'hb9b93e47),
	.w2(32'hb9cde256),
	.w3(32'hba2b423b),
	.w4(32'hba6bfbd2),
	.w5(32'hb917fd93),
	.w6(32'hba25c6ef),
	.w7(32'hb9dd191e),
	.w8(32'h39b35afa),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974d18b),
	.w1(32'hb86b6ff0),
	.w2(32'hb986b503),
	.w3(32'h3a1045f2),
	.w4(32'h3937886c),
	.w5(32'h3a21cdc0),
	.w6(32'h3a3420ad),
	.w7(32'hb8b95965),
	.w8(32'h3a93115d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7319e3),
	.w1(32'h3a0c43ca),
	.w2(32'hb936985a),
	.w3(32'h3a6f522f),
	.w4(32'h3a6c7eee),
	.w5(32'h3aea4a96),
	.w6(32'h3ab3022b),
	.w7(32'h3a75c36a),
	.w8(32'h3ae3b3c6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd449a),
	.w1(32'h3a3a648e),
	.w2(32'h3a6b3bc2),
	.w3(32'h3ac6a383),
	.w4(32'h3aa27c34),
	.w5(32'h3a280fe4),
	.w6(32'h3a8abf82),
	.w7(32'h3ab60784),
	.w8(32'h39180308),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f28c54),
	.w1(32'hba5a24f2),
	.w2(32'hb9dc14a7),
	.w3(32'h384b85e7),
	.w4(32'h39a42364),
	.w5(32'hb7e39b58),
	.w6(32'hba12b304),
	.w7(32'hb91f6c4f),
	.w8(32'hb98cacd9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d2cfa),
	.w1(32'hba6e98b2),
	.w2(32'hba4f628c),
	.w3(32'hb9aa16be),
	.w4(32'hba1b1e40),
	.w5(32'h39a329ce),
	.w6(32'h396df2d6),
	.w7(32'hba5b2877),
	.w8(32'h38ca660d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f61e27),
	.w1(32'h3952c4ac),
	.w2(32'hba223870),
	.w3(32'h39b82893),
	.w4(32'hb9fc158d),
	.w5(32'h3a6ef86f),
	.w6(32'h38ad0ed1),
	.w7(32'hba12ed20),
	.w8(32'h38b2bb43),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c93db9),
	.w1(32'h39b3604c),
	.w2(32'hb8fc1a2a),
	.w3(32'h38851842),
	.w4(32'h3988332c),
	.w5(32'h3a750d20),
	.w6(32'h394c9873),
	.w7(32'h39fe1e6e),
	.w8(32'h39ea71c1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53c957),
	.w1(32'h3a205d64),
	.w2(32'h3a02402d),
	.w3(32'h3a217117),
	.w4(32'h3a199f30),
	.w5(32'h3a6207e5),
	.w6(32'h3a73dab4),
	.w7(32'h3a335091),
	.w8(32'h3b0bfac4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c5924),
	.w1(32'h38919885),
	.w2(32'hb99ac8fb),
	.w3(32'h3aca0773),
	.w4(32'h3a9d1159),
	.w5(32'hbad7d5cc),
	.w6(32'h3a5c2cd4),
	.w7(32'h39dcdc89),
	.w8(32'hbaaf3c65),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ecab8),
	.w1(32'h38d5575f),
	.w2(32'hb7c410a3),
	.w3(32'hb9c5a12c),
	.w4(32'hba0fbf5d),
	.w5(32'h3a42cc9d),
	.w6(32'hb9bdeb61),
	.w7(32'hb9e60950),
	.w8(32'h39d6c95a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ce6c8),
	.w1(32'hb9faf641),
	.w2(32'hb8c97edd),
	.w3(32'h3a0e6c31),
	.w4(32'h38452ca9),
	.w5(32'hb887ca56),
	.w6(32'h3a21c5e0),
	.w7(32'hb91fcfcd),
	.w8(32'hb9d2ef74),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39487246),
	.w1(32'h39427665),
	.w2(32'h3a38fdcb),
	.w3(32'h3a2e4443),
	.w4(32'h3a94d9f7),
	.w5(32'h3a0a6293),
	.w6(32'hb6c28c83),
	.w7(32'h3a502905),
	.w8(32'h3aece4dd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22e120),
	.w1(32'h3a9178c7),
	.w2(32'h3a0b690b),
	.w3(32'h3aa5fc15),
	.w4(32'h3a982c2d),
	.w5(32'h3ab3bcb9),
	.w6(32'h3a9554bb),
	.w7(32'h3a121d78),
	.w8(32'h3a8430ea),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a572be4),
	.w1(32'h3a4fb781),
	.w2(32'h39a4f2b9),
	.w3(32'h3ac125a5),
	.w4(32'h3ac01059),
	.w5(32'hba53ce1c),
	.w6(32'h3a927cce),
	.w7(32'h3a8e8019),
	.w8(32'hb9b96b79),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17d293),
	.w1(32'hb973f711),
	.w2(32'h39006193),
	.w3(32'hba724955),
	.w4(32'hb9c138bf),
	.w5(32'hb9ba5840),
	.w6(32'h3a299d6c),
	.w7(32'hba31c40c),
	.w8(32'h3a492a57),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935b7a8),
	.w1(32'h3942f208),
	.w2(32'h3ac20e77),
	.w3(32'hba017e05),
	.w4(32'h3a116701),
	.w5(32'hb9a128be),
	.w6(32'hb8e56ddf),
	.w7(32'h3ace520d),
	.w8(32'hb74c4eb0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73ad83a),
	.w1(32'hb9cb1003),
	.w2(32'hb98bdcd4),
	.w3(32'hba20420c),
	.w4(32'hba2a7721),
	.w5(32'h3a292b9b),
	.w6(32'hb9939078),
	.w7(32'hb9d50892),
	.w8(32'h3a4276f3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23f0e3),
	.w1(32'h3a358fb1),
	.w2(32'h3a68f67b),
	.w3(32'h3a3a112b),
	.w4(32'h3a8fde01),
	.w5(32'h3a18b171),
	.w6(32'h3a54c07c),
	.w7(32'h3aceb54d),
	.w8(32'h39cb6951),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921e6a6),
	.w1(32'h39046991),
	.w2(32'hb987dae1),
	.w3(32'h3a1c48e4),
	.w4(32'h39a531cd),
	.w5(32'hb9744f86),
	.w6(32'h3a82e8a7),
	.w7(32'h3a44ba7f),
	.w8(32'hba34cc7d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a193bc),
	.w1(32'hba820f0b),
	.w2(32'hbaae9fac),
	.w3(32'hb9853e5b),
	.w4(32'hb8449363),
	.w5(32'hbb0090a5),
	.w6(32'hb8c3dde9),
	.w7(32'hb95d7c0d),
	.w8(32'hbaf5ceb7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22b6d0),
	.w1(32'hbb4a12e3),
	.w2(32'hbb13b182),
	.w3(32'hbb155a8b),
	.w4(32'hbae6c0fc),
	.w5(32'h3a61748c),
	.w6(32'hbb584d3c),
	.w7(32'hbb0e283e),
	.w8(32'h3a4d0587),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1686),
	.w1(32'h3a81556c),
	.w2(32'h3a57e592),
	.w3(32'h3a97d998),
	.w4(32'h3ae66328),
	.w5(32'h3a0f5962),
	.w6(32'h3a632412),
	.w7(32'h3b02feb4),
	.w8(32'h39c8625f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb0a64),
	.w1(32'h39fe648c),
	.w2(32'h3a2cf8ec),
	.w3(32'h3a05e8a9),
	.w4(32'h3a5d77a0),
	.w5(32'h39738e1b),
	.w6(32'hb9f827c9),
	.w7(32'h3a5fd1e0),
	.w8(32'h398e10ca),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930ca1d),
	.w1(32'h39a7f8ae),
	.w2(32'h397050d2),
	.w3(32'hb8bc88b6),
	.w4(32'hb9c5df28),
	.w5(32'hbaab0558),
	.w6(32'h39cced50),
	.w7(32'hb9ab82bf),
	.w8(32'hbad0c996),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf06c4),
	.w1(32'hbaa87f86),
	.w2(32'hbaaf12d0),
	.w3(32'hbac4b10f),
	.w4(32'hbac69fc6),
	.w5(32'h3af9fc84),
	.w6(32'hbab4d3b1),
	.w7(32'hbacd7af4),
	.w8(32'h3aca3543),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadcb98),
	.w1(32'h3ae2c62a),
	.w2(32'h3b0feb3a),
	.w3(32'h3aeb733d),
	.w4(32'h3acc9bd0),
	.w5(32'h3b29f0d8),
	.w6(32'h3af96170),
	.w7(32'h3b001ab9),
	.w8(32'h3a906276),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b039ddc),
	.w1(32'h3a9af93b),
	.w2(32'hb9d29f34),
	.w3(32'h3a977735),
	.w4(32'h3a267905),
	.w5(32'h3a95df97),
	.w6(32'h39859632),
	.w7(32'h38d68e86),
	.w8(32'h3aa59ad4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abecab5),
	.w1(32'h3a2a47d3),
	.w2(32'h3a13cab4),
	.w3(32'h3add1206),
	.w4(32'h3acb62f2),
	.w5(32'hb9e1c567),
	.w6(32'h3a994a51),
	.w7(32'h3aed3eba),
	.w8(32'hba7eee49),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388bb526),
	.w1(32'h39bb657e),
	.w2(32'h38c6a0ba),
	.w3(32'hb9430549),
	.w4(32'hb9dd862f),
	.w5(32'hba0d77b0),
	.w6(32'hba3f12b5),
	.w7(32'hb70939db),
	.w8(32'h3a4a6950),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33f015),
	.w1(32'h3a3d60d7),
	.w2(32'h38bf4060),
	.w3(32'hba00a126),
	.w4(32'h39d900fc),
	.w5(32'hba1d4794),
	.w6(32'hb80b3fee),
	.w7(32'h3967463c),
	.w8(32'hba40f589),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fe5ee),
	.w1(32'hba2504b8),
	.w2(32'hb99c1c30),
	.w3(32'hb9b44ee6),
	.w4(32'h395ec9b9),
	.w5(32'h3a8380a9),
	.w6(32'h394117d6),
	.w7(32'hb90c8091),
	.w8(32'h39cb69a4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fe3f3),
	.w1(32'hba76912d),
	.w2(32'hba48cfd7),
	.w3(32'h39c74bf0),
	.w4(32'hb89da063),
	.w5(32'hba1c855a),
	.w6(32'h3a06e599),
	.w7(32'hb965464f),
	.w8(32'hb9bca0b7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396716f8),
	.w1(32'hba228733),
	.w2(32'hba5d8777),
	.w3(32'hba5f745f),
	.w4(32'hba5b43cc),
	.w5(32'h3907058b),
	.w6(32'hba037ce7),
	.w7(32'hba623a68),
	.w8(32'h39c68768),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396775c4),
	.w1(32'h3a49bcb0),
	.w2(32'h3a177ecf),
	.w3(32'h390103a1),
	.w4(32'hb84ce0be),
	.w5(32'h3a98d749),
	.w6(32'h399c6f19),
	.w7(32'hb9a4ba4f),
	.w8(32'h3aa2f83a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab188f9),
	.w1(32'h3ad9c15e),
	.w2(32'h3b054ab7),
	.w3(32'h3abdf4d2),
	.w4(32'h3aa73f81),
	.w5(32'h3aea5fdf),
	.w6(32'h3aeaf19a),
	.w7(32'h3aed363e),
	.w8(32'h3a0b80b7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ce33c),
	.w1(32'hb5a6ffa4),
	.w2(32'hb9bdd9ba),
	.w3(32'h3a0a2344),
	.w4(32'h37d5e1c1),
	.w5(32'h39bc49bd),
	.w6(32'hba4a4c77),
	.w7(32'hba03e221),
	.w8(32'h38bd35e1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92878e6),
	.w1(32'h38d0e241),
	.w2(32'h39e2be1c),
	.w3(32'h39defe6e),
	.w4(32'h396d394e),
	.w5(32'h38c6a676),
	.w6(32'h3ab7882c),
	.w7(32'h39895f01),
	.w8(32'hb92314eb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3d177),
	.w1(32'h3a0f31b9),
	.w2(32'h39f74a2c),
	.w3(32'h3a1edc16),
	.w4(32'h3a88f642),
	.w5(32'h3a7e87e7),
	.w6(32'h39298412),
	.w7(32'h3a318d92),
	.w8(32'hb8919573),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37554586),
	.w1(32'hb965b754),
	.w2(32'h3a0192cb),
	.w3(32'h3a6ded28),
	.w4(32'h3aace873),
	.w5(32'h3a0109d1),
	.w6(32'h391b46a4),
	.w7(32'h3969c6c7),
	.w8(32'h38f6685c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c528cb),
	.w1(32'hb9c5afc1),
	.w2(32'hb9f90a95),
	.w3(32'hb872526f),
	.w4(32'hb92bd8b4),
	.w5(32'h39dbc80b),
	.w6(32'hb8d02ca3),
	.w7(32'hba5912cb),
	.w8(32'h381a5219),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f400e7),
	.w1(32'hb9e9ccfb),
	.w2(32'hba234479),
	.w3(32'hb86941e7),
	.w4(32'hba01136f),
	.w5(32'h39bc0fb3),
	.w6(32'h398835d1),
	.w7(32'hba5de723),
	.w8(32'hb9f288be),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1da8b1),
	.w1(32'hba8d2d54),
	.w2(32'hba4b9238),
	.w3(32'hb99b0904),
	.w4(32'hb98378b4),
	.w5(32'hb964602d),
	.w6(32'hb9a79749),
	.w7(32'hba2a2551),
	.w8(32'hb92a4330),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3df136),
	.w1(32'hb9a39bcb),
	.w2(32'h393f1f6b),
	.w3(32'hba1f1d76),
	.w4(32'hba1ed6f7),
	.w5(32'hbad719d8),
	.w6(32'hb9b6d36b),
	.w7(32'hb9260b84),
	.w8(32'hbaf9a523),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacb3f6),
	.w1(32'hbafcfa59),
	.w2(32'hbb345e77),
	.w3(32'hbb1fc981),
	.w4(32'hbb2d6203),
	.w5(32'h3a385f40),
	.w6(32'hbb0bc0c6),
	.w7(32'hbb4a6497),
	.w8(32'h3ac4af32),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79b74c),
	.w1(32'h38f6f041),
	.w2(32'hba0f39f8),
	.w3(32'h39b2b787),
	.w4(32'hb97581a0),
	.w5(32'h3a589957),
	.w6(32'h3a22e453),
	.w7(32'hb9cd5618),
	.w8(32'h38ae287e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd299),
	.w1(32'h3a9af0c5),
	.w2(32'h3a50635d),
	.w3(32'h3ab5b244),
	.w4(32'h3a986caa),
	.w5(32'h3a37db2b),
	.w6(32'h3a6d0699),
	.w7(32'h3aa4d8c8),
	.w8(32'h3a43ea57),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4432d),
	.w1(32'hb9020b4c),
	.w2(32'hb9423b3e),
	.w3(32'h3a4b5aa5),
	.w4(32'h39f9f626),
	.w5(32'hba8256ab),
	.w6(32'h39ebd612),
	.w7(32'h39184714),
	.w8(32'hba026c49),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bfd3a),
	.w1(32'hb9b6636c),
	.w2(32'hba127d72),
	.w3(32'hba4eac34),
	.w4(32'h3814dd6d),
	.w5(32'hba17dc4a),
	.w6(32'hb927e175),
	.w7(32'hb9c0cdd8),
	.w8(32'hba1b4548),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd6fc7),
	.w1(32'h38f204b2),
	.w2(32'hba508c56),
	.w3(32'h38656544),
	.w4(32'hb8831490),
	.w5(32'hb9f0551f),
	.w6(32'hba0dc9f0),
	.w7(32'hb98eb39d),
	.w8(32'hb9001097),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b55d1),
	.w1(32'h3a28ca3f),
	.w2(32'h38a06cfe),
	.w3(32'hb9ccea35),
	.w4(32'hba3e9914),
	.w5(32'hb8e167c1),
	.w6(32'h39433954),
	.w7(32'hba24c4d9),
	.w8(32'h3a01e8c6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecef28),
	.w1(32'h381d661c),
	.w2(32'h38b676bc),
	.w3(32'hb9791f3f),
	.w4(32'h38ae65e4),
	.w5(32'hbab6c8a2),
	.w6(32'h399278be),
	.w7(32'hb9675801),
	.w8(32'hbaa7e4ed),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857458),
	.w1(32'hba09990c),
	.w2(32'hba4deb64),
	.w3(32'hba75e033),
	.w4(32'hbad39575),
	.w5(32'hb9ed26da),
	.w6(32'hba531dbd),
	.w7(32'hbaba366c),
	.w8(32'hb9bd52d1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c72301),
	.w1(32'hba67fe54),
	.w2(32'hba97ac72),
	.w3(32'hba75705a),
	.w4(32'hba4dbf7a),
	.w5(32'hb7c84c3a),
	.w6(32'hbaa07150),
	.w7(32'hba8c2600),
	.w8(32'hb8a600e6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a576693),
	.w1(32'h38b0c306),
	.w2(32'h39882680),
	.w3(32'h39ce513c),
	.w4(32'h39b95c4b),
	.w5(32'h38c81c21),
	.w6(32'hba0a6a36),
	.w7(32'h3a15c4d7),
	.w8(32'h3969b1b8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7453e8),
	.w1(32'hb9c71751),
	.w2(32'hb9895a34),
	.w3(32'hb883f18d),
	.w4(32'hba3170f8),
	.w5(32'hba8301e0),
	.w6(32'hb9c10c3e),
	.w7(32'h39a889d2),
	.w8(32'hba786b69),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a8df),
	.w1(32'hbaaa3dfd),
	.w2(32'hbaae9f43),
	.w3(32'hbaa4164e),
	.w4(32'hba4b17fa),
	.w5(32'hbaf9fa74),
	.w6(32'hba97b4e9),
	.w7(32'hbaaa9c3f),
	.w8(32'hbb09f0a5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8a07),
	.w1(32'hbb0498b6),
	.w2(32'hbaf60019),
	.w3(32'hbb4775b9),
	.w4(32'hbb631fe7),
	.w5(32'hb99f2b15),
	.w6(32'hbb347203),
	.w7(32'hbb33f45e),
	.w8(32'hb9fe3483),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd4d3c),
	.w1(32'hb904032c),
	.w2(32'hb9cf34d3),
	.w3(32'h38b15677),
	.w4(32'h3839253f),
	.w5(32'hba2862d1),
	.w6(32'hb919756a),
	.w7(32'hb91b80f8),
	.w8(32'hb99fdcdb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf5972),
	.w1(32'hb9b80c43),
	.w2(32'hba57cc48),
	.w3(32'hba2bfd97),
	.w4(32'hb9e6d33d),
	.w5(32'h3a149ec7),
	.w6(32'hba2e7061),
	.w7(32'hb9e34a09),
	.w8(32'h39c572ed),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab9e76),
	.w1(32'hb9356cc3),
	.w2(32'hba0971ea),
	.w3(32'h39af71a8),
	.w4(32'hb6c94696),
	.w5(32'hba0a83aa),
	.w6(32'h39887a83),
	.w7(32'hb8bc9f03),
	.w8(32'h37883bf8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386dcedb),
	.w1(32'hb7f1c042),
	.w2(32'hb80b1799),
	.w3(32'hba63fe32),
	.w4(32'hba15912a),
	.w5(32'h3a877433),
	.w6(32'hb9839d17),
	.w7(32'h380c3651),
	.w8(32'h39b2ebb9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94deac4),
	.w1(32'hba2de875),
	.w2(32'hba4210ee),
	.w3(32'h39fc9a14),
	.w4(32'h3a62d44a),
	.w5(32'h395acb06),
	.w6(32'h39db3866),
	.w7(32'h3a20671e),
	.w8(32'h39ba17bf),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a277761),
	.w1(32'h3a977f3e),
	.w2(32'h3a859402),
	.w3(32'hb8a9bf41),
	.w4(32'h3a7419a6),
	.w5(32'hb93061e5),
	.w6(32'hb9e3f9d3),
	.w7(32'h3a9623e1),
	.w8(32'hb8c8dfec),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895b6d6),
	.w1(32'hba1a1aac),
	.w2(32'hb9f56b14),
	.w3(32'hb9ba762e),
	.w4(32'hba3025a8),
	.w5(32'hb769f8d3),
	.w6(32'hb785e22a),
	.w7(32'hba339419),
	.w8(32'hb93f7a56),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373495c0),
	.w1(32'hb8978e53),
	.w2(32'h39109fd5),
	.w3(32'hb911af2f),
	.w4(32'h38999a38),
	.w5(32'hb9d73eca),
	.w6(32'hb83ba095),
	.w7(32'h36d1b8f2),
	.w8(32'hb9c5bcba),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddbe2d),
	.w1(32'hba0723f8),
	.w2(32'hb89458a6),
	.w3(32'hbabfb30d),
	.w4(32'hba6e5c55),
	.w5(32'h39653596),
	.w6(32'hbaa0c9cd),
	.w7(32'hb9940c8c),
	.w8(32'hb991cca7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55d37f),
	.w1(32'h3a8675e6),
	.w2(32'h3a96f5a4),
	.w3(32'hb98995f2),
	.w4(32'h392478f7),
	.w5(32'h3a16c382),
	.w6(32'h3a8520a2),
	.w7(32'h3a1503f4),
	.w8(32'h39422c8a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f03ae),
	.w1(32'h3a42fb6c),
	.w2(32'hb9e77972),
	.w3(32'h3a1bd45c),
	.w4(32'hba4f0952),
	.w5(32'h3a86d905),
	.w6(32'h3a2269f3),
	.w7(32'hba4b37bd),
	.w8(32'h3a1447d3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a011f9a),
	.w1(32'h39a78370),
	.w2(32'h3a868e2c),
	.w3(32'h3ad399b5),
	.w4(32'h3aa98105),
	.w5(32'h3a00cbf1),
	.w6(32'h3b00f261),
	.w7(32'h3aeddac4),
	.w8(32'h3a25b92e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399749ef),
	.w1(32'h3a1cea22),
	.w2(32'h3a0025ed),
	.w3(32'h3a209ff4),
	.w4(32'hba023d2c),
	.w5(32'h3a2839a4),
	.w6(32'h39f23425),
	.w7(32'h391a2c17),
	.w8(32'h3993034a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989ab1a),
	.w1(32'h3872b3b1),
	.w2(32'hb46b6857),
	.w3(32'h39aedf3c),
	.w4(32'h3a38c2e3),
	.w5(32'h3a546666),
	.w6(32'hb910726b),
	.w7(32'h38700226),
	.w8(32'h3a920bca),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef272f),
	.w1(32'h3a92b695),
	.w2(32'h3a692f87),
	.w3(32'h3ac702c0),
	.w4(32'h3aaa65dd),
	.w5(32'h39c48820),
	.w6(32'h3afb94dd),
	.w7(32'h3ab2ce66),
	.w8(32'h3990b94b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8782f9),
	.w1(32'h39b854a6),
	.w2(32'h397cf4ac),
	.w3(32'h34459f14),
	.w4(32'hb9e4cef7),
	.w5(32'h3a9a328b),
	.w6(32'h393e5d67),
	.w7(32'h37d33c4e),
	.w8(32'h3a8c2b07),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76c4d9),
	.w1(32'hba1a2438),
	.w2(32'hba5184bc),
	.w3(32'h3a14a36d),
	.w4(32'hb98a1381),
	.w5(32'h3b58395d),
	.w6(32'h397be5fc),
	.w7(32'hba858f07),
	.w8(32'h3adc8124),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80995e),
	.w1(32'h3a82af6f),
	.w2(32'h3a91fd3b),
	.w3(32'h3b46beea),
	.w4(32'h3b2f0d0b),
	.w5(32'h399564d3),
	.w6(32'h3aefe0a8),
	.w7(32'h3a8df9ec),
	.w8(32'hba901aab),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4528c),
	.w1(32'h3af669a5),
	.w2(32'h3a852652),
	.w3(32'h3a82b8f9),
	.w4(32'h3b2f6f83),
	.w5(32'hbb500f89),
	.w6(32'h3914bd55),
	.w7(32'hbabac704),
	.w8(32'hb9acf553),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403e71),
	.w1(32'hba233521),
	.w2(32'hbb99da62),
	.w3(32'hbac17866),
	.w4(32'hbb09fcf6),
	.w5(32'h3b886e5a),
	.w6(32'h3b8c6927),
	.w7(32'hb91be04c),
	.w8(32'hbb0df6e2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c9dd),
	.w1(32'hbbb98ed7),
	.w2(32'hbbbe2338),
	.w3(32'h3ba881d7),
	.w4(32'h3b4959b7),
	.w5(32'hba4b10f5),
	.w6(32'hbb29c427),
	.w7(32'hbb4caecf),
	.w8(32'hba95f729),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39cba0),
	.w1(32'h3c13a2fa),
	.w2(32'h3c52bf26),
	.w3(32'h3ad76e51),
	.w4(32'h3c13a234),
	.w5(32'hbb6a9919),
	.w6(32'h3b354576),
	.w7(32'h3c418a55),
	.w8(32'hbbd6ec8a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c11a),
	.w1(32'hbb784204),
	.w2(32'h3a7820e8),
	.w3(32'hbb909e82),
	.w4(32'hb945e28b),
	.w5(32'h3b8271fd),
	.w6(32'hbbe2d822),
	.w7(32'hbad4edb0),
	.w8(32'h3b717ce8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921af7a),
	.w1(32'h3ab526fb),
	.w2(32'h38c8ffd1),
	.w3(32'hb950a12c),
	.w4(32'hb98ca038),
	.w5(32'h3a84f2ef),
	.w6(32'hb627b60a),
	.w7(32'hba0a4115),
	.w8(32'hb92d3bfa),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c28df0),
	.w1(32'h3a66d948),
	.w2(32'h3ade2224),
	.w3(32'h3ad9dbc8),
	.w4(32'h3b167865),
	.w5(32'h3b93aa25),
	.w6(32'h3af6ab14),
	.w7(32'h39125024),
	.w8(32'hba526f5e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fea21),
	.w1(32'hbb6cee3f),
	.w2(32'hbb90862d),
	.w3(32'h3b17d95b),
	.w4(32'h3aecc234),
	.w5(32'h3a210aa6),
	.w6(32'hbb20fe4a),
	.w7(32'hbaeec4fd),
	.w8(32'hba81a4fc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bba437),
	.w1(32'h3b30d71d),
	.w2(32'h3b352b25),
	.w3(32'h3b3a5e7a),
	.w4(32'h3b53d6c1),
	.w5(32'h3c18baef),
	.w6(32'h3afaaa69),
	.w7(32'h3b88c740),
	.w8(32'h3c111cc6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be88ee9),
	.w1(32'h3c08e514),
	.w2(32'h3c2b1778),
	.w3(32'h3c2dcfd1),
	.w4(32'h3c3c2338),
	.w5(32'hb9ad0b3a),
	.w6(32'h3c2c8251),
	.w7(32'h3c3462f2),
	.w8(32'hbb2fec5d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36c728),
	.w1(32'hbb3c549c),
	.w2(32'hbb345a18),
	.w3(32'hb971cec7),
	.w4(32'hb80d7b8a),
	.w5(32'hbb96c6d1),
	.w6(32'hbb2efa9a),
	.w7(32'hbb2defe7),
	.w8(32'hbb4e7395),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b59ce),
	.w1(32'hbb833aa0),
	.w2(32'hbb5b4947),
	.w3(32'hbacdc525),
	.w4(32'hb99a6ec8),
	.w5(32'h3b4e60be),
	.w6(32'hbaf20a2f),
	.w7(32'hbb352836),
	.w8(32'h3b7046e1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4ab68),
	.w1(32'hbb95e7d4),
	.w2(32'hbb919d31),
	.w3(32'hbab48620),
	.w4(32'hbb569a07),
	.w5(32'h3b7edd96),
	.w6(32'hbb6ce9c7),
	.w7(32'hbb94e9ff),
	.w8(32'h3b1ec053),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5731df),
	.w1(32'h3aaa146a),
	.w2(32'h3a1dc2bf),
	.w3(32'h3aa24bbe),
	.w4(32'h3990dd80),
	.w5(32'hbb5767ef),
	.w6(32'hb91aaefa),
	.w7(32'hba2ed1b5),
	.w8(32'hbaf34fd2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac3a0d),
	.w1(32'h3bc4b8e1),
	.w2(32'h3b8c6282),
	.w3(32'hbb7a7e37),
	.w4(32'hbae075c9),
	.w5(32'hba9c53ed),
	.w6(32'hbb358b11),
	.w7(32'hbaf76c50),
	.w8(32'hbad1375f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c07b7d),
	.w1(32'h3a125ddc),
	.w2(32'h3a9f2dd1),
	.w3(32'hba8401cc),
	.w4(32'h3938c743),
	.w5(32'hba9e7a37),
	.w6(32'hba025343),
	.w7(32'h37f3d5d5),
	.w8(32'hb97c7c94),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7abb60),
	.w1(32'hbc057a87),
	.w2(32'hbc141bfb),
	.w3(32'hbb418484),
	.w4(32'hbba4529c),
	.w5(32'h3b8314fa),
	.w6(32'hbb9f3f28),
	.w7(32'hbbf504cb),
	.w8(32'h3bb14f9b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8ba44),
	.w1(32'h3bd3076c),
	.w2(32'h3b8691e9),
	.w3(32'h3ba67d21),
	.w4(32'h3b4033aa),
	.w5(32'hba927ce6),
	.w6(32'h3c04d167),
	.w7(32'h3bb7242e),
	.w8(32'hb6b23432),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab3a24),
	.w1(32'h3b10c420),
	.w2(32'h3ac08ea8),
	.w3(32'hbb4a1375),
	.w4(32'hbb434fac),
	.w5(32'hbaa1a2f4),
	.w6(32'hbb76c3ba),
	.w7(32'hbb267328),
	.w8(32'hbb3eab5b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad107be),
	.w1(32'hbaf4adf2),
	.w2(32'hbb4787be),
	.w3(32'hbb17f9ee),
	.w4(32'hbb0853f8),
	.w5(32'h3b0204d1),
	.w6(32'hbb869e79),
	.w7(32'hbb62e931),
	.w8(32'hbb31518e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1840a),
	.w1(32'hbb3c170a),
	.w2(32'hbae001d0),
	.w3(32'hbaa64dd0),
	.w4(32'hba26a7bc),
	.w5(32'h3b166a1f),
	.w6(32'hbb7c32a4),
	.w7(32'hbb46cfc3),
	.w8(32'h3b4b67c8),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb45439),
	.w1(32'hbbb5db05),
	.w2(32'hbb74465d),
	.w3(32'h3adf761a),
	.w4(32'hbae4e534),
	.w5(32'hbb37a43a),
	.w6(32'h3a567c01),
	.w7(32'hba876dbf),
	.w8(32'hbb47fa90),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e59ad),
	.w1(32'hbba24c55),
	.w2(32'h3a6b39ce),
	.w3(32'hbbbb6be6),
	.w4(32'h39a3c795),
	.w5(32'hbbbbb946),
	.w6(32'hbbe15870),
	.w7(32'hba353d70),
	.w8(32'hba633025),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48cfd3),
	.w1(32'h3b6aba81),
	.w2(32'h3bd424f5),
	.w3(32'hbba96950),
	.w4(32'hbb459adf),
	.w5(32'hbac09f1b),
	.w6(32'hbaf3bb8d),
	.w7(32'hb64d7dc2),
	.w8(32'hbade9497),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5592b5),
	.w1(32'hbb49744d),
	.w2(32'hbacf2a2f),
	.w3(32'h393e71f8),
	.w4(32'h3a6b1b1c),
	.w5(32'hbba66ad1),
	.w6(32'hb9712198),
	.w7(32'h3a17f3fb),
	.w8(32'hbb9d995c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba192288),
	.w1(32'hbaed2520),
	.w2(32'hb9becded),
	.w3(32'hbb8b428e),
	.w4(32'hbb780ffc),
	.w5(32'h3a139a82),
	.w6(32'hbbb62c30),
	.w7(32'hbb9ee1b5),
	.w8(32'hba5efb7b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b691181),
	.w1(32'h3b979751),
	.w2(32'h3b9ee4f5),
	.w3(32'h3ace5942),
	.w4(32'h3be31581),
	.w5(32'hba373143),
	.w6(32'hbadd6b18),
	.w7(32'h3adb5724),
	.w8(32'hba94e023),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38954cb3),
	.w1(32'hba59e2cd),
	.w2(32'hba8af68c),
	.w3(32'hba9367cd),
	.w4(32'hba8357bc),
	.w5(32'hba6d885d),
	.w6(32'hbaffe95c),
	.w7(32'hba91687f),
	.w8(32'hbaac9176),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86cfe7),
	.w1(32'hbacfbec7),
	.w2(32'hbaa8fb5e),
	.w3(32'hbb10bbcc),
	.w4(32'hba06b791),
	.w5(32'h39bf0177),
	.w6(32'hbaed0448),
	.w7(32'hbaf51646),
	.w8(32'hba5f39a5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule