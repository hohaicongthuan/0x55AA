module top(data_in, data_out, Clk, Rst, En);
    input Clk, Rst, En;
    input [7:0] data_in;
    output [31:0] data_out;

    layer_0_top layer_0_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_1_top layer_1_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_2_top layer_2_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_3_top layer_3_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_4_top layer_4_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_5_top layer_5_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_6_top layer_6_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_7_top layer_7_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_8_top layer_8_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_9_top layer_9_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_10_top layer_10_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_11_top layer_11_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_12_top layer_12_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_13_top layer_13_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_14_top layer_14_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
    layer_15_top layer_15_top_Inst0(
        .Clk(Clk), .Rst(Rst),
        .data_in(), .data_out(),
        .valid_in(), .valid_out()
    );
endmodule