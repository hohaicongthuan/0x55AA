module layer_10_featuremap_163(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94334fa),
	.w1(32'hbc66abf1),
	.w2(32'hbc0d31ab),
	.w3(32'hbaaf7add),
	.w4(32'hba9685ef),
	.w5(32'h3c7f281d),
	.w6(32'h3c0ec11b),
	.w7(32'h3c67715c),
	.w8(32'h3c034a2e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009f38),
	.w1(32'h3ad5a40f),
	.w2(32'h3b5bf739),
	.w3(32'h3b5bc660),
	.w4(32'hbb16bfb9),
	.w5(32'hba81e3da),
	.w6(32'h3a17765f),
	.w7(32'h3a46b6b2),
	.w8(32'h3902a901),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d1dbe),
	.w1(32'h3b826ef8),
	.w2(32'hbaed757d),
	.w3(32'hb8b51248),
	.w4(32'h3aa2d4b2),
	.w5(32'h398fe880),
	.w6(32'h3b055fab),
	.w7(32'hbb1fee8c),
	.w8(32'hbafacfaa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb60c5),
	.w1(32'hbb41b379),
	.w2(32'hb92c6ff2),
	.w3(32'hbac0f2ab),
	.w4(32'h3c0de588),
	.w5(32'hbc182f80),
	.w6(32'hbc063ba6),
	.w7(32'hbb0a462c),
	.w8(32'hbac91b81),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb342320),
	.w1(32'hbc214017),
	.w2(32'hbc0d5123),
	.w3(32'hbb45a660),
	.w4(32'hbb9f448c),
	.w5(32'hbbbc2701),
	.w6(32'h39fb4586),
	.w7(32'hbc0a66ec),
	.w8(32'hba71460e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f3e78),
	.w1(32'hbbf2db45),
	.w2(32'hbaeee214),
	.w3(32'h3bb11965),
	.w4(32'hbb870094),
	.w5(32'h3ab05537),
	.w6(32'hbb82e213),
	.w7(32'hba73f597),
	.w8(32'h3b71265f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f74c8),
	.w1(32'h3b4da741),
	.w2(32'h3aa098f7),
	.w3(32'h3919db54),
	.w4(32'hba8e4556),
	.w5(32'h3b4940e5),
	.w6(32'h3b2763bc),
	.w7(32'h3afbbe0a),
	.w8(32'h3baa5645),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71e504),
	.w1(32'h3ad838d4),
	.w2(32'hbbd2a4ee),
	.w3(32'h3ae21ffc),
	.w4(32'h3ae3f65a),
	.w5(32'hbb437470),
	.w6(32'h3b20bcb2),
	.w7(32'h3b91a4be),
	.w8(32'h3b538f3d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c912f),
	.w1(32'hbbb30cca),
	.w2(32'h3affe7ef),
	.w3(32'hbabafb30),
	.w4(32'hbb06bac3),
	.w5(32'hba382470),
	.w6(32'hbaea951f),
	.w7(32'h3b4dddcb),
	.w8(32'hb9b65327),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7c2e),
	.w1(32'hbaebe6bc),
	.w2(32'h3be883ad),
	.w3(32'h3b3163db),
	.w4(32'h3a952715),
	.w5(32'h3bcd0e63),
	.w6(32'h3bdaaa30),
	.w7(32'h3c03ddfc),
	.w8(32'h3c12e967),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33fe95),
	.w1(32'hbbe9d2ec),
	.w2(32'hbc279351),
	.w3(32'h38a74a1e),
	.w4(32'h3a689919),
	.w5(32'h379bab0c),
	.w6(32'hbbafe184),
	.w7(32'hbc3cbc2f),
	.w8(32'hbbcdc633),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b9dab),
	.w1(32'hbb1a85d5),
	.w2(32'h3bd5afb1),
	.w3(32'h3af57157),
	.w4(32'h3c1cbcdb),
	.w5(32'hbb5a6ec0),
	.w6(32'h3b4a6265),
	.w7(32'h3bb5b3d5),
	.w8(32'h3bc46611),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b633),
	.w1(32'h39cc8856),
	.w2(32'hba328cfd),
	.w3(32'h3be91edd),
	.w4(32'h3893e214),
	.w5(32'h3b3ba298),
	.w6(32'h3be3c45d),
	.w7(32'h3b06c5f3),
	.w8(32'h3b723f4b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12acd3),
	.w1(32'h3c0555b5),
	.w2(32'hbb799fca),
	.w3(32'hb91fd74a),
	.w4(32'h3bed6796),
	.w5(32'hbb95bf64),
	.w6(32'h3ba100c0),
	.w7(32'h3af0a6bc),
	.w8(32'h3b424463),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fae9b),
	.w1(32'hbb060ccc),
	.w2(32'hbbe6a52f),
	.w3(32'hb992995c),
	.w4(32'h3c37bca7),
	.w5(32'hbc80866b),
	.w6(32'h3addbe97),
	.w7(32'h3b143495),
	.w8(32'h3b70618d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64976e),
	.w1(32'hbb60e585),
	.w2(32'h3bb0f074),
	.w3(32'h3c034822),
	.w4(32'hbabff175),
	.w5(32'hb9b9db99),
	.w6(32'h3b583e22),
	.w7(32'h3bb5a850),
	.w8(32'h3b1e0bf7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb24805),
	.w1(32'h3b2287cb),
	.w2(32'hb9dfea48),
	.w3(32'hbb8014f3),
	.w4(32'hbb160264),
	.w5(32'hba592e5d),
	.w6(32'h3bba3453),
	.w7(32'hb9dbeb1b),
	.w8(32'h39f77bf7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bb863),
	.w1(32'h3b090669),
	.w2(32'h3b9b57ac),
	.w3(32'h3b2ee5a2),
	.w4(32'hbb21f254),
	.w5(32'h3b6f9432),
	.w6(32'h3beadd07),
	.w7(32'h3b5734f4),
	.w8(32'h3bcf5f7c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be59d3a),
	.w1(32'h3af32b09),
	.w2(32'h3a3c0a1b),
	.w3(32'h3a70a9a1),
	.w4(32'h3b13583a),
	.w5(32'h3a595d5a),
	.w6(32'h3b151543),
	.w7(32'hba9ad4a8),
	.w8(32'h3b152b46),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98a8ac),
	.w1(32'hbb604d2d),
	.w2(32'h3aac2085),
	.w3(32'hbb728b35),
	.w4(32'hbb135e8b),
	.w5(32'hbb0f3c24),
	.w6(32'hbab13d5e),
	.w7(32'hb8b920b4),
	.w8(32'h3a86090a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0def5c),
	.w1(32'h3b1ca78e),
	.w2(32'hba9e7f03),
	.w3(32'hbab8c196),
	.w4(32'h3aa921e4),
	.w5(32'hbaa6196f),
	.w6(32'h3b2141a8),
	.w7(32'h3b3041a2),
	.w8(32'h3ad91436),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add5e21),
	.w1(32'h3b0b5f2f),
	.w2(32'hbc7a99c8),
	.w3(32'h3a159536),
	.w4(32'hba1b685b),
	.w5(32'h3c3fea3f),
	.w6(32'h3b351df3),
	.w7(32'hbb60f44b),
	.w8(32'h3b39e7e9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01bdf5),
	.w1(32'h3a2f2344),
	.w2(32'hb9a07621),
	.w3(32'h3c863e6a),
	.w4(32'h3a735538),
	.w5(32'h39e16464),
	.w6(32'h3c1a4d14),
	.w7(32'h3b4dd753),
	.w8(32'h3bb9ecc9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e846),
	.w1(32'h3b6d7ae0),
	.w2(32'h3b119130),
	.w3(32'h3bfe144b),
	.w4(32'h3b6d3966),
	.w5(32'hb9f49ee3),
	.w6(32'h3c282de9),
	.w7(32'h3bc23c49),
	.w8(32'h3b9f06d4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc8fd),
	.w1(32'hb9f293aa),
	.w2(32'h3c3b35d0),
	.w3(32'h3bc10633),
	.w4(32'h38bf408b),
	.w5(32'hbb57d50a),
	.w6(32'h3be514a7),
	.w7(32'h3bb7b446),
	.w8(32'hba956dd7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3095),
	.w1(32'hbb544db4),
	.w2(32'h3af1f693),
	.w3(32'hba7a0b2a),
	.w4(32'hbb61f395),
	.w5(32'hbb8eeffc),
	.w6(32'hba67fd0c),
	.w7(32'hbb6a8010),
	.w8(32'hbb960050),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f660d4),
	.w1(32'hbaf2cae0),
	.w2(32'hbafc03c9),
	.w3(32'h3abfb087),
	.w4(32'hbb17eb99),
	.w5(32'hbb294af2),
	.w6(32'h39ce2c92),
	.w7(32'hb9f453ba),
	.w8(32'h3b09566a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933e80a),
	.w1(32'hbc1e3f6e),
	.w2(32'h3c3eb6e0),
	.w3(32'h3b72d428),
	.w4(32'h3be50457),
	.w5(32'h3b00c0c0),
	.w6(32'hbb9d6e37),
	.w7(32'hba0cd61a),
	.w8(32'h3a8d0262),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ee7ad),
	.w1(32'h3b486c37),
	.w2(32'hbb66a6e0),
	.w3(32'h3b5e08cd),
	.w4(32'h3bb8faa5),
	.w5(32'hbba31725),
	.w6(32'h3c1c86e9),
	.w7(32'h3aba1002),
	.w8(32'h3aaa8082),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a394a),
	.w1(32'h3b79021c),
	.w2(32'h3c11306f),
	.w3(32'h3ba0e925),
	.w4(32'h3b7f2825),
	.w5(32'h3ab19493),
	.w6(32'h3c15fc10),
	.w7(32'h3c3decb2),
	.w8(32'h3a381326),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea824c),
	.w1(32'h39f1c7bf),
	.w2(32'hbaf6cc6e),
	.w3(32'hba9db8f9),
	.w4(32'h3a72080d),
	.w5(32'hb9c82e4c),
	.w6(32'h3ab33097),
	.w7(32'h3a1fa43d),
	.w8(32'h3a3ff604),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afd9e2),
	.w1(32'h389fc319),
	.w2(32'hbb081b5c),
	.w3(32'h3aa8370e),
	.w4(32'hb9c1ff32),
	.w5(32'hba2dd9d1),
	.w6(32'h3ae0672a),
	.w7(32'h3a472e2e),
	.w8(32'h3aa44801),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bfce6),
	.w1(32'hbbcfeba1),
	.w2(32'hbb5a87f4),
	.w3(32'h38dae993),
	.w4(32'hbb0118dd),
	.w5(32'hbc243bdd),
	.w6(32'h3a58be33),
	.w7(32'hbbc92a52),
	.w8(32'h3b2a061e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8443d8),
	.w1(32'hbb85cc3d),
	.w2(32'h3acc62d5),
	.w3(32'hba9364b0),
	.w4(32'hbba75bde),
	.w5(32'hba5d768f),
	.w6(32'hbb8a4f1d),
	.w7(32'hbbe22d14),
	.w8(32'hbb73d309),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f084),
	.w1(32'hbbcd935b),
	.w2(32'h3b93a188),
	.w3(32'h3a8ccf40),
	.w4(32'hbb22828a),
	.w5(32'h3b5cd62c),
	.w6(32'hbb18b0ef),
	.w7(32'h3af42058),
	.w8(32'h3b8e6828),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c184b),
	.w1(32'hbb5c290b),
	.w2(32'hbada9be5),
	.w3(32'h3b8f94e4),
	.w4(32'hba259d50),
	.w5(32'hba4e0164),
	.w6(32'hbb356e99),
	.w7(32'hbb4c17cc),
	.w8(32'hb9860e51),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d7eb0),
	.w1(32'hbc450da5),
	.w2(32'hbbc7edb6),
	.w3(32'h3bddbe75),
	.w4(32'hbbd07640),
	.w5(32'hb9ad92d4),
	.w6(32'h3b16358d),
	.w7(32'hbb6a8998),
	.w8(32'hbb3b6f82),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aa98b),
	.w1(32'hba571b25),
	.w2(32'hbc378121),
	.w3(32'h3c200f91),
	.w4(32'hbbd5fec1),
	.w5(32'hbc54e291),
	.w6(32'h3c6f06a6),
	.w7(32'h3aaac76c),
	.w8(32'hbb579095),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cf1b9),
	.w1(32'hbaf233ec),
	.w2(32'hbc25ce5a),
	.w3(32'h3c06d3af),
	.w4(32'hbaa28ce2),
	.w5(32'hbc33618b),
	.w6(32'h3c5adc42),
	.w7(32'h3b460ebd),
	.w8(32'hbb4587f9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a299e63),
	.w1(32'h3a235a2e),
	.w2(32'hba6dfcbc),
	.w3(32'h39a417bf),
	.w4(32'hbac2d5ee),
	.w5(32'hbb3121cf),
	.w6(32'h3ac57892),
	.w7(32'hbb35bc12),
	.w8(32'hbadc3801),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44643a),
	.w1(32'hbad1f2ce),
	.w2(32'h3b408b17),
	.w3(32'hba42024f),
	.w4(32'hbaa3d6d4),
	.w5(32'hbac0b455),
	.w6(32'hba1f0a1b),
	.w7(32'h3b0ab725),
	.w8(32'hbab9725b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba623fe1),
	.w1(32'hbb7bdfc7),
	.w2(32'h3bb9e43c),
	.w3(32'hb9f5f6ad),
	.w4(32'hbac1b069),
	.w5(32'hbb999c32),
	.w6(32'hbb80abb2),
	.w7(32'hbc0594e6),
	.w8(32'hbaba1204),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981c0c3),
	.w1(32'h3afe2029),
	.w2(32'hba0c345f),
	.w3(32'h38a82026),
	.w4(32'hb9729adb),
	.w5(32'h3a3d36ea),
	.w6(32'h3adb2c1e),
	.w7(32'h3936352f),
	.w8(32'h3ac217c5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43b6e2),
	.w1(32'hbb215099),
	.w2(32'h3be3a64e),
	.w3(32'h3b9e4786),
	.w4(32'hbb41fa59),
	.w5(32'h3bb99ba6),
	.w6(32'h3c32f719),
	.w7(32'h3bf800fa),
	.w8(32'h3c230f16),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde1fb8),
	.w1(32'h3c7af947),
	.w2(32'hbc4aa2ab),
	.w3(32'h3b97a781),
	.w4(32'h3bf8b42a),
	.w5(32'hb928c229),
	.w6(32'h3ca8a364),
	.w7(32'h3abee9ce),
	.w8(32'hba198d40),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5dee0),
	.w1(32'h3be56456),
	.w2(32'hbb419266),
	.w3(32'hbafc815e),
	.w4(32'hbb4a2f8d),
	.w5(32'hbae2e26e),
	.w6(32'h3bb98bde),
	.w7(32'hbb3d4c08),
	.w8(32'h3af57a85),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6f32),
	.w1(32'h3bca5397),
	.w2(32'h3bdf1f3f),
	.w3(32'h3b34caac),
	.w4(32'h3c7401b3),
	.w5(32'hbb57042d),
	.w6(32'h3b8ffa28),
	.w7(32'h3ba714d7),
	.w8(32'h3c1e46e7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe57f6e),
	.w1(32'hbb80a6be),
	.w2(32'hbb6273c7),
	.w3(32'h3acf937e),
	.w4(32'h3b01ce19),
	.w5(32'h3aa05d9b),
	.w6(32'h3b2713a2),
	.w7(32'h3aae5233),
	.w8(32'hb997aa65),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dec9b),
	.w1(32'h3997121e),
	.w2(32'h3a4e8c54),
	.w3(32'hbb2b0301),
	.w4(32'hb9c9e45f),
	.w5(32'h3a5bfd6b),
	.w6(32'h39bed6f0),
	.w7(32'hb937381c),
	.w8(32'h3b2ea747),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4e9fd),
	.w1(32'h3b6fab5d),
	.w2(32'hbb7ffe15),
	.w3(32'h3972e389),
	.w4(32'h3b022ab4),
	.w5(32'hbbad2db8),
	.w6(32'h3aeab4fb),
	.w7(32'hba904360),
	.w8(32'hbb2c6858),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab0f4),
	.w1(32'h3b55fe4f),
	.w2(32'hbc25af2d),
	.w3(32'hbad93265),
	.w4(32'hb9e31a01),
	.w5(32'hbc336515),
	.w6(32'h3b836572),
	.w7(32'hbb024606),
	.w8(32'hbb1342bb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144dca),
	.w1(32'h3b9b0e3a),
	.w2(32'h3d829b27),
	.w3(32'hbb804b8e),
	.w4(32'h3c862935),
	.w5(32'h3c37f4d4),
	.w6(32'hbb78d0d0),
	.w7(32'h3cdccaf6),
	.w8(32'h3bd2ff99),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f690c),
	.w1(32'hbbd802d0),
	.w2(32'h3a9d882b),
	.w3(32'hbbcfd8ef),
	.w4(32'hbba28dd2),
	.w5(32'hb9bfe15d),
	.w6(32'hbb8648ca),
	.w7(32'hb9e984c3),
	.w8(32'h3a22e4e2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404904),
	.w1(32'hbc07ae7c),
	.w2(32'hbafb7191),
	.w3(32'hbb11a7cf),
	.w4(32'hbbc8f045),
	.w5(32'h3b9aca49),
	.w6(32'hba6d1df4),
	.w7(32'hbba75aad),
	.w8(32'h3bb913b4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be61625),
	.w1(32'hbb138cd4),
	.w2(32'h3830a375),
	.w3(32'h3bb94eb2),
	.w4(32'hbb5c4698),
	.w5(32'h3a1177ab),
	.w6(32'hba7b00b3),
	.w7(32'hbb3a9d8b),
	.w8(32'h39ed75ff),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394553c4),
	.w1(32'hbadacf97),
	.w2(32'hbb46a335),
	.w3(32'hba821f39),
	.w4(32'hba6edd98),
	.w5(32'hbb6968dd),
	.w6(32'hb9804b6c),
	.w7(32'hb88185cb),
	.w8(32'hbaff21c2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f5c9),
	.w1(32'h3bfbe832),
	.w2(32'hb9b62114),
	.w3(32'h3a222c47),
	.w4(32'h3be638ad),
	.w5(32'h3ac4f79b),
	.w6(32'h3b835973),
	.w7(32'h3b789d0f),
	.w8(32'h3b9bc5cf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40fdc8),
	.w1(32'hbb92ad26),
	.w2(32'hbba0c99a),
	.w3(32'h3afe2f02),
	.w4(32'h39210594),
	.w5(32'hbb9fe76a),
	.w6(32'h3b9191f7),
	.w7(32'hbba16ff4),
	.w8(32'h38f8fe1a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c6912),
	.w1(32'h398f779e),
	.w2(32'h3b88b1a6),
	.w3(32'h3b1c41cc),
	.w4(32'hba4e6b53),
	.w5(32'hbaec0437),
	.w6(32'h39e3058e),
	.w7(32'h3b34aebb),
	.w8(32'hba9064ab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae41bc),
	.w1(32'h3a9a003c),
	.w2(32'hba2630bd),
	.w3(32'hbbb3e799),
	.w4(32'h3b0744b9),
	.w5(32'hba0825f4),
	.w6(32'h3abf13ec),
	.w7(32'h3b0cbf79),
	.w8(32'h3ab7d4d1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8189fe),
	.w1(32'h3a2a12ab),
	.w2(32'h3b8200b7),
	.w3(32'h3ae6faac),
	.w4(32'h3b42b29e),
	.w5(32'h3b12414a),
	.w6(32'h3b18b32c),
	.w7(32'hb9ea3a70),
	.w8(32'h3a3650d8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f85592),
	.w1(32'h3ada2076),
	.w2(32'hbb925cc8),
	.w3(32'hbac65511),
	.w4(32'h3b011a13),
	.w5(32'h3a472915),
	.w6(32'h3bb134f0),
	.w7(32'h3b1f935c),
	.w8(32'h3bd68d26),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac23d9c),
	.w1(32'hbbe9d763),
	.w2(32'hbc016b96),
	.w3(32'hba574196),
	.w4(32'hbc200364),
	.w5(32'hbc3d52f1),
	.w6(32'hb95d0a7e),
	.w7(32'hbbc0d878),
	.w8(32'hbb6a88af),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc962563),
	.w1(32'hbb7d31c8),
	.w2(32'h3abc2330),
	.w3(32'hbbb72f8f),
	.w4(32'hbb8da051),
	.w5(32'h39c796d2),
	.w6(32'hba9364b5),
	.w7(32'hb9594056),
	.w8(32'h3add5cb5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2986c),
	.w1(32'h3b13fd72),
	.w2(32'h3ac515e5),
	.w3(32'h38fa69c0),
	.w4(32'h3a80eb9c),
	.w5(32'hb8ff4c60),
	.w6(32'h3a8e180e),
	.w7(32'h3a844481),
	.w8(32'h3ac92519),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f5048),
	.w1(32'h3afe135d),
	.w2(32'h3a818322),
	.w3(32'hbb54cba5),
	.w4(32'h3b0f734d),
	.w5(32'hbb33d7e6),
	.w6(32'hba4abf3d),
	.w7(32'hbb731479),
	.w8(32'hbb69bc9c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2ea5),
	.w1(32'hbc0d0aa1),
	.w2(32'hb9b97349),
	.w3(32'hbaef5ee8),
	.w4(32'hbb87b2b2),
	.w5(32'hba2e19d1),
	.w6(32'h3af33201),
	.w7(32'h3b4e02e0),
	.w8(32'h3b059081),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badb3b1),
	.w1(32'h3bfc2148),
	.w2(32'h3bac8ef4),
	.w3(32'hbb34b052),
	.w4(32'hb89f7534),
	.w5(32'h3951f03e),
	.w6(32'h3bc4f4ed),
	.w7(32'h3bc86630),
	.w8(32'h3ba05fdd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5928),
	.w1(32'hbb33094f),
	.w2(32'h3acf7f61),
	.w3(32'h3ac324a7),
	.w4(32'hbb7554ab),
	.w5(32'hbb8b33f6),
	.w6(32'h3b8fefa8),
	.w7(32'h3a22cfdf),
	.w8(32'h39fc354c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8fd3e),
	.w1(32'h3b6c3f88),
	.w2(32'hbca955e3),
	.w3(32'h3bc814d3),
	.w4(32'hbb50e063),
	.w5(32'hbcdef4cd),
	.w6(32'h3c8af9fd),
	.w7(32'hba730afb),
	.w8(32'hbb390d4a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e7ac),
	.w1(32'h3a8e0ac4),
	.w2(32'h3b5d3615),
	.w3(32'hba6e6209),
	.w4(32'hbb00a19c),
	.w5(32'hb95bdc5d),
	.w6(32'hb9ba4f50),
	.w7(32'h39a33b07),
	.w8(32'h3a549024),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b324a2b),
	.w1(32'hbac2d8ba),
	.w2(32'hbb0c5cf0),
	.w3(32'h37b871bb),
	.w4(32'hb7b9d9fd),
	.w5(32'hbac6f468),
	.w6(32'h39ba6597),
	.w7(32'hba77a938),
	.w8(32'h39c814c2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be3a44),
	.w1(32'hb7059806),
	.w2(32'h39ba2270),
	.w3(32'h3801213d),
	.w4(32'h3ac6f328),
	.w5(32'hba5cf23a),
	.w6(32'h3a4a5ccb),
	.w7(32'h3afdcaac),
	.w8(32'h3a2c4e94),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef53fc),
	.w1(32'hbb1cba37),
	.w2(32'hbaf45efa),
	.w3(32'hbac24689),
	.w4(32'hba5b91b6),
	.w5(32'hb9deef64),
	.w6(32'h39f1ba13),
	.w7(32'h3a13808d),
	.w8(32'h3a60c501),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2e200),
	.w1(32'hbae7c4d9),
	.w2(32'h3c4780fe),
	.w3(32'hb9dfc94f),
	.w4(32'hb9b30ea1),
	.w5(32'h3b044380),
	.w6(32'hbb4bc29c),
	.w7(32'h3ab415d9),
	.w8(32'hba962894),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7514f1),
	.w1(32'hbbeb3074),
	.w2(32'h3cd7e10e),
	.w3(32'hbb9641c5),
	.w4(32'h3b22e07c),
	.w5(32'hbc965ee9),
	.w6(32'hbb9cfe81),
	.w7(32'hb8943def),
	.w8(32'hba9d84fe),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00bd53),
	.w1(32'h3b7278ce),
	.w2(32'hbbbb65ba),
	.w3(32'h3a7aa47e),
	.w4(32'h3a726ce5),
	.w5(32'hbb5aca75),
	.w6(32'h3c0bd110),
	.w7(32'h3b99ca47),
	.w8(32'h3b2bdb3f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2d299),
	.w1(32'h3b9eb62a),
	.w2(32'h3b895465),
	.w3(32'h3bab1cae),
	.w4(32'h3b18c931),
	.w5(32'hbb8f129e),
	.w6(32'h3bbd42de),
	.w7(32'hba0b1d06),
	.w8(32'hbafd5dbf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012ba0),
	.w1(32'hbb5d4ef1),
	.w2(32'h3b86e51b),
	.w3(32'hbba1a7af),
	.w4(32'hbbaf3505),
	.w5(32'hbaaeb92b),
	.w6(32'h3b5a90f3),
	.w7(32'hbb3a2d61),
	.w8(32'h3b6c5584),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5765fb),
	.w1(32'hbab7aeb1),
	.w2(32'hbb702dec),
	.w3(32'h3ab93421),
	.w4(32'h3aac6be0),
	.w5(32'h38a6c08e),
	.w6(32'h3bb41af2),
	.w7(32'h3b277130),
	.w8(32'h3b556c71),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b358e99),
	.w1(32'hba173dc0),
	.w2(32'hbae4266a),
	.w3(32'h3b5a1fdb),
	.w4(32'h39eb1745),
	.w5(32'hbafbf29a),
	.w6(32'h3b5a51ca),
	.w7(32'h3b2767d1),
	.w8(32'hb9d297d8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fe993),
	.w1(32'h3ada2018),
	.w2(32'h3b50e1e2),
	.w3(32'hbae2de47),
	.w4(32'h39fd1aea),
	.w5(32'h3b5103a7),
	.w6(32'h3b90cee6),
	.w7(32'h3b04afe8),
	.w8(32'h3a85f056),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f08a),
	.w1(32'hbbae0dc2),
	.w2(32'h390bdabe),
	.w3(32'hbb1eeea0),
	.w4(32'hbb278d7d),
	.w5(32'hbb48a216),
	.w6(32'hbb3f5f36),
	.w7(32'hbb1a668f),
	.w8(32'hba250c16),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04ab44),
	.w1(32'hba82279e),
	.w2(32'h37ad25ea),
	.w3(32'hb8b8816e),
	.w4(32'hba8616ce),
	.w5(32'h3b50a22b),
	.w6(32'h3a19bda2),
	.w7(32'h3a8bb77c),
	.w8(32'hba84ff33),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b699b),
	.w1(32'h38d039cf),
	.w2(32'hbba553e5),
	.w3(32'hbb1e159f),
	.w4(32'hba5422e9),
	.w5(32'h3a00910e),
	.w6(32'h3a94a6df),
	.w7(32'hbb5f9ab9),
	.w8(32'hbbf44ad5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a41d5),
	.w1(32'h3b93de09),
	.w2(32'h39e86df8),
	.w3(32'hbb4fec47),
	.w4(32'h3a6979e3),
	.w5(32'hba44e39e),
	.w6(32'h3b2f85b7),
	.w7(32'h3abb4e5f),
	.w8(32'h37379b8e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fd5af),
	.w1(32'hb9fce48c),
	.w2(32'hbaa75697),
	.w3(32'h3ae0cd21),
	.w4(32'h3a486279),
	.w5(32'hbc1ebc18),
	.w6(32'h3b7a79b6),
	.w7(32'hbba6ee72),
	.w8(32'hbaaf77f3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91891b),
	.w1(32'hb883756b),
	.w2(32'hba6ea9dc),
	.w3(32'hbb71d0c3),
	.w4(32'h38f7ca99),
	.w5(32'hba7a3aaa),
	.w6(32'h3ab13adc),
	.w7(32'h3ab44bf6),
	.w8(32'h39e3d5ff),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075877),
	.w1(32'h38022a8f),
	.w2(32'h3af9a87c),
	.w3(32'h3a62b63c),
	.w4(32'hbb44e559),
	.w5(32'hb90b98ac),
	.w6(32'h3a51b0ab),
	.w7(32'hba64915b),
	.w8(32'h3aadc078),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e2ea3),
	.w1(32'hb9cf1e37),
	.w2(32'hbb46d6d6),
	.w3(32'h3b10f5e1),
	.w4(32'hba67e6a2),
	.w5(32'hbb349090),
	.w6(32'h3bd955dd),
	.w7(32'h3b57d7c0),
	.w8(32'h3b4820f8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b647310),
	.w1(32'h38c8977c),
	.w2(32'hbb9809d8),
	.w3(32'h3b86a30a),
	.w4(32'hb9612ab4),
	.w5(32'hbacfec69),
	.w6(32'h3bc102ad),
	.w7(32'h3abd1844),
	.w8(32'hbaa9e496),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc039bbe),
	.w1(32'hbbf5ec0c),
	.w2(32'hbc4a457e),
	.w3(32'h3a2f0736),
	.w4(32'hbb4a8498),
	.w5(32'hbbb96548),
	.w6(32'h3b994e1a),
	.w7(32'h3a4a2ec3),
	.w8(32'h39cb09ed),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bf4a7),
	.w1(32'hbbfdbbdb),
	.w2(32'hbb115b66),
	.w3(32'hba95a5b1),
	.w4(32'hbbf10339),
	.w5(32'hbb007925),
	.w6(32'hb9a150e9),
	.w7(32'h38565a1b),
	.w8(32'hbb8ba12f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb250b22),
	.w1(32'hbae943fe),
	.w2(32'h3a0e4eab),
	.w3(32'hbac8b09f),
	.w4(32'hbaa12c47),
	.w5(32'hbb1f4d21),
	.w6(32'h3bcfb111),
	.w7(32'h3b37631a),
	.w8(32'h3b122850),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86847d),
	.w1(32'h3a8b8a2e),
	.w2(32'h375acd0a),
	.w3(32'hb94f4d23),
	.w4(32'h3abd4ce6),
	.w5(32'hba05eaee),
	.w6(32'h3ab423bd),
	.w7(32'hbac9b037),
	.w8(32'hbb370438),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba21b9e),
	.w1(32'hbb734984),
	.w2(32'hbc1bdafc),
	.w3(32'h3b33a7de),
	.w4(32'hbc1e202d),
	.w5(32'h3a149c21),
	.w6(32'h3bf2b5e1),
	.w7(32'hbaeb1018),
	.w8(32'h3b9c2b14),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc520d0),
	.w1(32'h3b150706),
	.w2(32'h3991a39c),
	.w3(32'h3bbf787e),
	.w4(32'hb9de63d4),
	.w5(32'h3ad325e6),
	.w6(32'hbb30aca0),
	.w7(32'h3b2757cc),
	.w8(32'h38ca242f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba9c22),
	.w1(32'hbbc41a7a),
	.w2(32'h3c7ec293),
	.w3(32'h3b98ad85),
	.w4(32'hbb6a544b),
	.w5(32'hba930fc7),
	.w6(32'h3af9f73f),
	.w7(32'h3ba0d56e),
	.w8(32'h3bbafea4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c4b64),
	.w1(32'hbbaef737),
	.w2(32'hbbf0f685),
	.w3(32'hbb6fdc88),
	.w4(32'hbbcebace),
	.w5(32'hbb64a019),
	.w6(32'h3b5dc248),
	.w7(32'hbbaf974f),
	.w8(32'hbb7331e1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdadb6e),
	.w1(32'hbb84e1c8),
	.w2(32'h3bd4b5df),
	.w3(32'hbb4076c8),
	.w4(32'hbbcf0bd2),
	.w5(32'hbb15daba),
	.w6(32'hba97c5a1),
	.w7(32'h3adc5068),
	.w8(32'hbbe2a7d6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a55b2),
	.w1(32'h3a328987),
	.w2(32'hbc0a9e28),
	.w3(32'h3b7b110c),
	.w4(32'h3b5eccd0),
	.w5(32'hbc08c1c2),
	.w6(32'h3c97665f),
	.w7(32'hbb154b73),
	.w8(32'h3a883663),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca00a12),
	.w1(32'h3c1bb431),
	.w2(32'h3b6623ad),
	.w3(32'h3c0bee1e),
	.w4(32'hbb0e32d3),
	.w5(32'h3adc371f),
	.w6(32'h3bf95023),
	.w7(32'hbae241ac),
	.w8(32'hbaafd5e2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e7f7),
	.w1(32'hbb33405c),
	.w2(32'hbc6ab946),
	.w3(32'h3bc7caf8),
	.w4(32'h39cfd4a0),
	.w5(32'hbb82bf67),
	.w6(32'h3c07854e),
	.w7(32'h3a1a3f9f),
	.w8(32'h3ade2109),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5623b),
	.w1(32'h3b2e412e),
	.w2(32'hba46ec70),
	.w3(32'h3ace61fa),
	.w4(32'h3ada9aad),
	.w5(32'hbb08b5a9),
	.w6(32'h3b02a7bd),
	.w7(32'hba0c05e6),
	.w8(32'h3a404b2b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00e6c),
	.w1(32'h3b3459d1),
	.w2(32'hbb8a247c),
	.w3(32'h3b2cf553),
	.w4(32'h3b3ba4b9),
	.w5(32'hbb2ffd7f),
	.w6(32'h3ba02ece),
	.w7(32'h3b56d8e0),
	.w8(32'hbabb4470),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a308479),
	.w1(32'hbb70dc2f),
	.w2(32'hbac25a27),
	.w3(32'h3ae257c4),
	.w4(32'h3a731571),
	.w5(32'hba822c78),
	.w6(32'h3a0f1483),
	.w7(32'h3a4b4885),
	.w8(32'h3b2b5eeb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4e61),
	.w1(32'h3b0a12a2),
	.w2(32'hbb5194b0),
	.w3(32'hba0bdf41),
	.w4(32'h3af1a2f1),
	.w5(32'hba0859d5),
	.w6(32'h3af38690),
	.w7(32'hbb0ea9a1),
	.w8(32'hbb901e68),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb492ac5),
	.w1(32'h3a70ea80),
	.w2(32'hb9dd01da),
	.w3(32'hbb0292b5),
	.w4(32'hb82c6a30),
	.w5(32'hb92f8a48),
	.w6(32'h3b0916d9),
	.w7(32'h3b23d1b9),
	.w8(32'h3a849895),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ace64),
	.w1(32'h3bc76ad1),
	.w2(32'hb9a8df17),
	.w3(32'h3ba78e46),
	.w4(32'h3b943adb),
	.w5(32'h3a712f53),
	.w6(32'h3c16dc0a),
	.w7(32'h3ba95549),
	.w8(32'h3bc58471),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be867e1),
	.w1(32'h3c8bb28c),
	.w2(32'hba5b9754),
	.w3(32'h3bc94691),
	.w4(32'h3c2aa480),
	.w5(32'hbb8d4014),
	.w6(32'h3c32a809),
	.w7(32'h3b8d44a1),
	.w8(32'h3a7b462e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf6730),
	.w1(32'hbb139ef2),
	.w2(32'h3c177c6b),
	.w3(32'hbbb889a0),
	.w4(32'h3b5af633),
	.w5(32'h3b1cc613),
	.w6(32'hba33b69b),
	.w7(32'h3bf1e452),
	.w8(32'h3b279a1a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882a398),
	.w1(32'h3c097adc),
	.w2(32'h3c88eccd),
	.w3(32'h3b1bd238),
	.w4(32'h3c8aee14),
	.w5(32'h3c0dd67e),
	.w6(32'h3c53b4cd),
	.w7(32'h3c879da4),
	.w8(32'h3b8ea03b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f5440),
	.w1(32'hbb0dc431),
	.w2(32'h3bd8f5e4),
	.w3(32'hbbdf7f76),
	.w4(32'h39578f99),
	.w5(32'h3a6f3002),
	.w6(32'hba894e6f),
	.w7(32'h3bb6e905),
	.w8(32'h3b296621),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfa4c),
	.w1(32'hbb3dcf44),
	.w2(32'h3bbba86f),
	.w3(32'hbacdfada),
	.w4(32'hba47a082),
	.w5(32'hbb522e83),
	.w6(32'hbad30e92),
	.w7(32'hbb229d25),
	.w8(32'hb8aa281b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b09132),
	.w1(32'h3b8d4890),
	.w2(32'hbb7d4b6c),
	.w3(32'h39b63868),
	.w4(32'h3b8362d4),
	.w5(32'hbb7deddb),
	.w6(32'h3bd78628),
	.w7(32'h3ada5b92),
	.w8(32'h3b0066b0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc52663),
	.w1(32'h3b3c985d),
	.w2(32'hbbcd1aaa),
	.w3(32'hbb228f54),
	.w4(32'h3b186bd4),
	.w5(32'hbb4b33ae),
	.w6(32'h3b96a1b8),
	.w7(32'h3a9718dc),
	.w8(32'h3b089f07),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bf07c),
	.w1(32'h39d15256),
	.w2(32'hbaf02695),
	.w3(32'h3723b9a8),
	.w4(32'h3a300b96),
	.w5(32'hbaaa41d1),
	.w6(32'h3ae16948),
	.w7(32'h3a35ca79),
	.w8(32'h3a29d455),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836a43),
	.w1(32'hb98b2bb5),
	.w2(32'hbae0e565),
	.w3(32'h399a8bf7),
	.w4(32'h3a1af0aa),
	.w5(32'h39141259),
	.w6(32'h3b00ff19),
	.w7(32'h3a15b780),
	.w8(32'h3a1ddfd7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ac336),
	.w1(32'h3b923875),
	.w2(32'hbc8d668f),
	.w3(32'h39b8ff99),
	.w4(32'h3b7241d3),
	.w5(32'h3c01cb9f),
	.w6(32'h3c1cd326),
	.w7(32'hbb973ffc),
	.w8(32'h3b0e0740),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53afc0),
	.w1(32'h3c1b2d72),
	.w2(32'h3b106f27),
	.w3(32'h3c1822dc),
	.w4(32'h3bf3fcde),
	.w5(32'hba91e372),
	.w6(32'h3c3396e8),
	.w7(32'h3b482e09),
	.w8(32'h3bb2530e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e4620),
	.w1(32'hbb5b0b0b),
	.w2(32'hbbc604cf),
	.w3(32'hbb7d1687),
	.w4(32'hb92286a3),
	.w5(32'hbb10e8d7),
	.w6(32'hbb035b37),
	.w7(32'hbb7e96ab),
	.w8(32'hba25f647),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaced82b),
	.w1(32'hbbbb6109),
	.w2(32'hba444f08),
	.w3(32'h3a75f8e8),
	.w4(32'hbaab7c60),
	.w5(32'hbac85737),
	.w6(32'hbaf13c22),
	.w7(32'h3af77f57),
	.w8(32'h3a5d2108),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e3f0c),
	.w1(32'h3baace10),
	.w2(32'hbb236787),
	.w3(32'h3a316cbb),
	.w4(32'h3ad5d4f0),
	.w5(32'hbbb09f5a),
	.w6(32'h3bf4dd1d),
	.w7(32'h3b56af5a),
	.w8(32'h3a8f4693),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8adaa),
	.w1(32'h3af69019),
	.w2(32'hbc970597),
	.w3(32'hba816304),
	.w4(32'h3aefcf49),
	.w5(32'h3c6043d5),
	.w6(32'h3c41d6d4),
	.w7(32'h3a22ada7),
	.w8(32'h3bb57be5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5157db),
	.w1(32'hbc39952f),
	.w2(32'hbb8ea60a),
	.w3(32'h3c05ec32),
	.w4(32'hbc20cab4),
	.w5(32'hb9f3d7bc),
	.w6(32'hbba673c3),
	.w7(32'hbb561cc9),
	.w8(32'hb9c9c3de),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5b8a),
	.w1(32'hbae22e7a),
	.w2(32'hba91125d),
	.w3(32'hbb9d3087),
	.w4(32'hba4f137b),
	.w5(32'hb9c0204a),
	.w6(32'h39e50015),
	.w7(32'h3a989abb),
	.w8(32'hb9d7face),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba984a17),
	.w1(32'h3a1ceaaa),
	.w2(32'h3a2e1526),
	.w3(32'h3721292a),
	.w4(32'h39e3b561),
	.w5(32'h3a088823),
	.w6(32'h39eac601),
	.w7(32'h3a04ae18),
	.w8(32'h3a410f98),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0b7fb),
	.w1(32'h3bac1913),
	.w2(32'h3bb15f81),
	.w3(32'hbb3625fe),
	.w4(32'hba1e3da8),
	.w5(32'h3a12595a),
	.w6(32'h39d1016e),
	.w7(32'h3b91cb9c),
	.w8(32'h3b976d2d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3850b3a0),
	.w1(32'hbae3633c),
	.w2(32'h3b2391b2),
	.w3(32'h3aa0cf02),
	.w4(32'h39773e19),
	.w5(32'h3b8fe59a),
	.w6(32'h3b4db163),
	.w7(32'h3b0852f6),
	.w8(32'h3b9a0aa7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6bc60),
	.w1(32'hb8e8af41),
	.w2(32'hb91dba84),
	.w3(32'hb8cda80b),
	.w4(32'h37c9db68),
	.w5(32'hb9180a21),
	.w6(32'h38f0bfdd),
	.w7(32'h380bd621),
	.w8(32'hb7c9ad40),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae03c41),
	.w1(32'h3a9b28bb),
	.w2(32'h39fdf0ab),
	.w3(32'h3a7c45de),
	.w4(32'h39618372),
	.w5(32'h39db52c1),
	.w6(32'h3a880b5f),
	.w7(32'h3aa7de89),
	.w8(32'h3ab4702f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a997954),
	.w1(32'h3a2097a7),
	.w2(32'h3a0aebe3),
	.w3(32'h3a7e2a26),
	.w4(32'h39575e91),
	.w5(32'hb923582c),
	.w6(32'h3ac5965c),
	.w7(32'h3a3ddb4e),
	.w8(32'h39ffaa14),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6149f),
	.w1(32'h39c85ade),
	.w2(32'h39e7f704),
	.w3(32'h3a885685),
	.w4(32'hb7b75ec8),
	.w5(32'h386440b9),
	.w6(32'h3b0c564d),
	.w7(32'h3a94977f),
	.w8(32'h3a9e2c72),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110e20),
	.w1(32'h3b06fa54),
	.w2(32'h3b0d78df),
	.w3(32'h39b6a437),
	.w4(32'hba59f18a),
	.w5(32'hbac95102),
	.w6(32'h3b05f085),
	.w7(32'h3a471afd),
	.w8(32'hb9277624),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005791),
	.w1(32'hbb5c828a),
	.w2(32'h3a049293),
	.w3(32'h3a76ac90),
	.w4(32'hba55225b),
	.w5(32'h3b357898),
	.w6(32'h3b7b6316),
	.w7(32'h3b1a5994),
	.w8(32'h3b7944c9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61c5a5),
	.w1(32'h3adc5b61),
	.w2(32'h39218f4b),
	.w3(32'h3b1b8a0e),
	.w4(32'hb9c72a00),
	.w5(32'hbacf8828),
	.w6(32'h3b8acc67),
	.w7(32'h3adb4656),
	.w8(32'h38fcb01e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b35b28),
	.w1(32'hba83e641),
	.w2(32'h3820ee42),
	.w3(32'hb9d0e066),
	.w4(32'hbaaad9e1),
	.w5(32'hb9820412),
	.w6(32'h3a6947d7),
	.w7(32'hba87b36e),
	.w8(32'h3a625055),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946eff6),
	.w1(32'hbb55e595),
	.w2(32'hba98e4e3),
	.w3(32'h3a3ceb79),
	.w4(32'hbac909c0),
	.w5(32'h3983b334),
	.w6(32'h3aef180c),
	.w7(32'hba7be812),
	.w8(32'hb72b24b9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dafe9),
	.w1(32'h37a2fde1),
	.w2(32'hbaa90c26),
	.w3(32'h3a0282b5),
	.w4(32'hbb0cdca5),
	.w5(32'hbb62d46a),
	.w6(32'h3b456a58),
	.w7(32'h396795e4),
	.w8(32'hbab13601),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac25c27),
	.w1(32'hba24e44d),
	.w2(32'h3b0feaa4),
	.w3(32'h3aa86c87),
	.w4(32'h3a6fa540),
	.w5(32'h3b31a724),
	.w6(32'h3b276c03),
	.w7(32'h3b1c15ac),
	.w8(32'h3b3f8874),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c348e),
	.w1(32'h3a0c9321),
	.w2(32'h3a0fc31c),
	.w3(32'h3a4fbf3e),
	.w4(32'h38ba08ac),
	.w5(32'h38d98151),
	.w6(32'h3ae5b593),
	.w7(32'h3a6f0397),
	.w8(32'h3a141ed9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd69b51),
	.w1(32'h3abdbb16),
	.w2(32'hbb9c4f4d),
	.w3(32'h3bb72e6f),
	.w4(32'hba5ceac7),
	.w5(32'hbb90115a),
	.w6(32'h3bfa9058),
	.w7(32'h3acc002a),
	.w8(32'hbae69875),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addd746),
	.w1(32'h3a58fb49),
	.w2(32'h39a9dfaa),
	.w3(32'h3aecb302),
	.w4(32'hb90e13ef),
	.w5(32'hba0430c1),
	.w6(32'h3b11b660),
	.w7(32'h3a74159f),
	.w8(32'h3a2faec4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38928d44),
	.w1(32'h383d84f6),
	.w2(32'h38e48b7e),
	.w3(32'hb90a20d0),
	.w4(32'hb8b2b8bf),
	.w5(32'hb79a0cec),
	.w6(32'hb84a918c),
	.w7(32'hb914975c),
	.w8(32'h370e1713),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb819d092),
	.w1(32'hb82f576c),
	.w2(32'h3916eefe),
	.w3(32'h38789162),
	.w4(32'h38a91e5c),
	.w5(32'h392eaf31),
	.w6(32'hb89cf6da),
	.w7(32'hb8d1bdc2),
	.w8(32'hb8f48cf4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d0e0e),
	.w1(32'hb7fa47d7),
	.w2(32'hb9ddbfd1),
	.w3(32'h3a6e88cc),
	.w4(32'h3a09416d),
	.w5(32'hb9fb2904),
	.w6(32'h3a86239b),
	.w7(32'h3a646f56),
	.w8(32'hb98ac8f2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b450047),
	.w1(32'h3ab4e3a7),
	.w2(32'h395013a5),
	.w3(32'h3b1e9b6d),
	.w4(32'hba1b991d),
	.w5(32'hb9b88510),
	.w6(32'h3b6f5e4f),
	.w7(32'h3aa38314),
	.w8(32'h39a001d2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7829af),
	.w1(32'h3a8d9d0a),
	.w2(32'h3aeab7b8),
	.w3(32'h3b84cc91),
	.w4(32'h3a04579b),
	.w5(32'h3a43cc11),
	.w6(32'h3bca5c96),
	.w7(32'h3b5e4e0c),
	.w8(32'h3b45f496),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898113e),
	.w1(32'hb89d8573),
	.w2(32'hb89ca0b8),
	.w3(32'hb8e87a7b),
	.w4(32'h3896512a),
	.w5(32'h381a5fa5),
	.w6(32'h36f15741),
	.w7(32'hb8887de4),
	.w8(32'hb83c2ac5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a505ef0),
	.w1(32'hb9378401),
	.w2(32'h3b0a27e9),
	.w3(32'h3b412791),
	.w4(32'h3ab022b3),
	.w5(32'h3b2cc7e9),
	.w6(32'h3ba0e80e),
	.w7(32'h3b748d59),
	.w8(32'h3b516e4b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87426d),
	.w1(32'h3b62aa7c),
	.w2(32'h3ab789be),
	.w3(32'h3b8c4cab),
	.w4(32'h3af64299),
	.w5(32'h3a77d141),
	.w6(32'h3b713c05),
	.w7(32'h3affce07),
	.w8(32'h3aa6aa1b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ddb70),
	.w1(32'hbb3d6712),
	.w2(32'hba946cac),
	.w3(32'h3a8ccec1),
	.w4(32'h3aaad341),
	.w5(32'h3b17cc72),
	.w6(32'h3b351e71),
	.w7(32'h3a4b121d),
	.w8(32'h3a8a9f1a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c1ff),
	.w1(32'hba4eb430),
	.w2(32'hba9a899e),
	.w3(32'h3b831a4c),
	.w4(32'hb8c538e8),
	.w5(32'h3990608a),
	.w6(32'h3bd32fc9),
	.w7(32'h3b14575e),
	.w8(32'h3a840e07),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae16846),
	.w1(32'h3adc5736),
	.w2(32'h3a988da2),
	.w3(32'h3a021971),
	.w4(32'hba4cce22),
	.w5(32'hbb000d26),
	.w6(32'h3abd19d1),
	.w7(32'hb9307cd2),
	.w8(32'hb999a94e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59ea7c),
	.w1(32'h3b21889c),
	.w2(32'h3b032260),
	.w3(32'h3b470cde),
	.w4(32'h3ae0b582),
	.w5(32'h3a8d0c2e),
	.w6(32'h3b12f576),
	.w7(32'h3a851df6),
	.w8(32'h3a5aee4d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b109c),
	.w1(32'hb994afa8),
	.w2(32'h39c45fbe),
	.w3(32'h3a18dac9),
	.w4(32'hba8803b9),
	.w5(32'hba71025c),
	.w6(32'h3b677bbf),
	.w7(32'h3a8f2a1f),
	.w8(32'hb894cfc8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b112949),
	.w1(32'hba6f865f),
	.w2(32'hbabd7ea1),
	.w3(32'h3a6bbc10),
	.w4(32'hbb53eda2),
	.w5(32'hbb1e18d5),
	.w6(32'h3b1c673c),
	.w7(32'hbb132b2e),
	.w8(32'hba476378),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41f9aa),
	.w1(32'h39e1ed6c),
	.w2(32'hbabcfc55),
	.w3(32'h3b2523c1),
	.w4(32'hb9f5460f),
	.w5(32'hbb0ffff9),
	.w6(32'h3b35bd45),
	.w7(32'h38a176bb),
	.w8(32'hba5b5514),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7707758),
	.w1(32'hba593d5c),
	.w2(32'hba83c875),
	.w3(32'h37edd9bf),
	.w4(32'h38f8a7ea),
	.w5(32'h384f5295),
	.w6(32'h398fe5d7),
	.w7(32'hb837775d),
	.w8(32'hb8ed5ed0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7d9ac),
	.w1(32'h399699e0),
	.w2(32'h399d997d),
	.w3(32'h395bd766),
	.w4(32'h39476be5),
	.w5(32'h391348ff),
	.w6(32'h38a74673),
	.w7(32'h3900b468),
	.w8(32'h39821c39),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bfe33),
	.w1(32'h3a13790d),
	.w2(32'h3b0393a5),
	.w3(32'h3ab6afaf),
	.w4(32'h3a832866),
	.w5(32'h3b0f25d4),
	.w6(32'h3b502eea),
	.w7(32'h3b09425a),
	.w8(32'h3b1dacb2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba850f96),
	.w1(32'hbaa7c38a),
	.w2(32'hb9cd521d),
	.w3(32'h37603334),
	.w4(32'hb9ba3dc9),
	.w5(32'h38d584ab),
	.w6(32'hb91258e1),
	.w7(32'hb9047bd3),
	.w8(32'hb98384ac),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b266ff0),
	.w1(32'h3b03d0ea),
	.w2(32'h3af0ade3),
	.w3(32'h3af5e551),
	.w4(32'h3a9efe14),
	.w5(32'h3a16961e),
	.w6(32'h3b7a33d5),
	.w7(32'h3b076d86),
	.w8(32'h3ad1dd83),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928d0d4),
	.w1(32'hb9cb24c9),
	.w2(32'hb9df42f0),
	.w3(32'hb94b623b),
	.w4(32'hb99dbff8),
	.w5(32'hb8d534a2),
	.w6(32'hb99a56d4),
	.w7(32'hb900cf62),
	.w8(32'h397539f0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d8b33),
	.w1(32'hb99d1639),
	.w2(32'h37715abc),
	.w3(32'h3b22af5c),
	.w4(32'hb8ac700b),
	.w5(32'hb80a5c92),
	.w6(32'h3af913fb),
	.w7(32'h39bca094),
	.w8(32'h3a97499e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bbe46),
	.w1(32'h38be0522),
	.w2(32'h39d25b8f),
	.w3(32'h3942c620),
	.w4(32'h39ebccb7),
	.w5(32'h3a14b2b1),
	.w6(32'h393c1132),
	.w7(32'h399522f2),
	.w8(32'h39c8d2f5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c65403),
	.w1(32'hb8b6f725),
	.w2(32'hba14619d),
	.w3(32'hb96adcf2),
	.w4(32'hb979b3a4),
	.w5(32'hba0a0ea5),
	.w6(32'hb892fe4f),
	.w7(32'hb8b3cf32),
	.w8(32'hb9446c69),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fc501),
	.w1(32'h3a5250df),
	.w2(32'h3b1786a1),
	.w3(32'h3a92619c),
	.w4(32'h3a72ecb0),
	.w5(32'h3b11725a),
	.w6(32'h3b34597d),
	.w7(32'h3b106b05),
	.w8(32'h3b1547ff),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba93ce1),
	.w1(32'h3b00d37c),
	.w2(32'h3a27f70a),
	.w3(32'h3b810c62),
	.w4(32'h3ac84d06),
	.w5(32'h3b17f432),
	.w6(32'h3bc7e77c),
	.w7(32'h3b90d97b),
	.w8(32'h3b48985f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2057dd),
	.w1(32'hb99af3bc),
	.w2(32'hbb019f47),
	.w3(32'h3af3a8bc),
	.w4(32'hb84e4ad6),
	.w5(32'hbaf506de),
	.w6(32'h3b20f34d),
	.w7(32'h39472430),
	.w8(32'hba1f469e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b248502),
	.w1(32'h3a89bf65),
	.w2(32'hb9f359da),
	.w3(32'h3aa5a045),
	.w4(32'hbaa5f038),
	.w5(32'hbaa80f77),
	.w6(32'h3b859559),
	.w7(32'h3ad1dd3d),
	.w8(32'h38f2b4db),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69f6e1),
	.w1(32'hba8ac3c0),
	.w2(32'hb9e6fd39),
	.w3(32'h3aa6b5d8),
	.w4(32'h3a463cf9),
	.w5(32'h3a269aa2),
	.w6(32'h3a843392),
	.w7(32'h3a3ef693),
	.w8(32'h38b60dc8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2159b),
	.w1(32'h39d692da),
	.w2(32'h3b96f5c1),
	.w3(32'h3bd6368d),
	.w4(32'h3aee2a52),
	.w5(32'h3b789c60),
	.w6(32'h3c0b8950),
	.w7(32'h3b95cb62),
	.w8(32'h3bfce44a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b5019),
	.w1(32'hbb0f2364),
	.w2(32'hbac8e4db),
	.w3(32'h38dbcabc),
	.w4(32'hbb33d19d),
	.w5(32'hbb2af8f6),
	.w6(32'h3b436b2b),
	.w7(32'h39a1b342),
	.w8(32'hb9e7f0b7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296f92),
	.w1(32'h3b2ff6bc),
	.w2(32'h3babfda0),
	.w3(32'h3b4b3ff1),
	.w4(32'h3b2f192b),
	.w5(32'h3b85ae4d),
	.w6(32'h3b96b8b3),
	.w7(32'h3b8277f9),
	.w8(32'h3b6e38f1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38153ee1),
	.w1(32'h3881a705),
	.w2(32'h3a67cb40),
	.w3(32'h3a0ecdac),
	.w4(32'h39fd3a62),
	.w5(32'h3a6bddcd),
	.w6(32'h395fde88),
	.w7(32'h39b53a08),
	.w8(32'h3a42fed3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933dcc),
	.w1(32'hba8f4605),
	.w2(32'h3a481c16),
	.w3(32'hba6b9a1b),
	.w4(32'hba6f5a68),
	.w5(32'h3a5f563d),
	.w6(32'h3a355cbb),
	.w7(32'h3a00f623),
	.w8(32'h3a1bf43e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8920144),
	.w1(32'h398c93c8),
	.w2(32'h397f65d0),
	.w3(32'hb90d537f),
	.w4(32'h3988dafb),
	.w5(32'h397b8d34),
	.w6(32'h393d6583),
	.w7(32'h394b6475),
	.w8(32'h39a9b5d0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a844a28),
	.w1(32'hb91f88a2),
	.w2(32'hb98f3868),
	.w3(32'h3a9c9f1b),
	.w4(32'h3862d122),
	.w5(32'hb964a844),
	.w6(32'h3a7e2f4c),
	.w7(32'h3a05c130),
	.w8(32'h3a2f89a7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a227bc2),
	.w1(32'h39cf77c8),
	.w2(32'hb98d805a),
	.w3(32'h39cd30cc),
	.w4(32'hb9ecb50d),
	.w5(32'hba7ae446),
	.w6(32'h3a411854),
	.w7(32'h37d9a93d),
	.w8(32'h396dff86),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a325635),
	.w1(32'hba0bfaba),
	.w2(32'h3aec177a),
	.w3(32'h3aea0f33),
	.w4(32'hb985211f),
	.w5(32'h39882371),
	.w6(32'h3b4755c7),
	.w7(32'h3ac03ac6),
	.w8(32'h3b281c06),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7951512),
	.w1(32'hb920ca68),
	.w2(32'hb9072644),
	.w3(32'hb83eb850),
	.w4(32'hb853670b),
	.w5(32'h38c9cd98),
	.w6(32'hb8a84118),
	.w7(32'hb7c42127),
	.w8(32'hb92ea980),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80cbc4b),
	.w1(32'h39a6a857),
	.w2(32'h393f83b7),
	.w3(32'h37f923a5),
	.w4(32'h38512430),
	.w5(32'hb84f3040),
	.w6(32'h372bfb31),
	.w7(32'h38b15cef),
	.w8(32'hb8c85fce),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac616a5),
	.w1(32'h3a131d73),
	.w2(32'hb94f8e0c),
	.w3(32'h3a1b6961),
	.w4(32'hb9fb2be4),
	.w5(32'hbaa876ff),
	.w6(32'h3af673e7),
	.w7(32'h3a00276c),
	.w8(32'h3960185f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391deade),
	.w1(32'h397491d4),
	.w2(32'hba01e2dc),
	.w3(32'h3a0fcad2),
	.w4(32'hba0f2171),
	.w5(32'hbae0236b),
	.w6(32'h3aee483f),
	.w7(32'h3990b71f),
	.w8(32'h398c8d34),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48b662),
	.w1(32'hbb1761c6),
	.w2(32'hbb724f16),
	.w3(32'h3b6be6da),
	.w4(32'hba222323),
	.w5(32'hbac5362f),
	.w6(32'h3aba4f9d),
	.w7(32'hb99443ec),
	.w8(32'hbb05bd70),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b5907),
	.w1(32'hba80c301),
	.w2(32'hbac4d16c),
	.w3(32'hb9f2fc1f),
	.w4(32'hba4ad54b),
	.w5(32'hba9c3c72),
	.w6(32'hb990db25),
	.w7(32'hba4e6097),
	.w8(32'hba226414),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcecc1c),
	.w1(32'h3b957453),
	.w2(32'h3c264bb7),
	.w3(32'h3bcc0e60),
	.w4(32'h3bafb307),
	.w5(32'h3bcfce22),
	.w6(32'h3be92303),
	.w7(32'h3bd280a7),
	.w8(32'h3bd186e2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9381d71),
	.w1(32'hbb8a2089),
	.w2(32'hbb413276),
	.w3(32'h3b513c43),
	.w4(32'hbae9902e),
	.w5(32'hba73ff7a),
	.w6(32'h3be424b9),
	.w7(32'h3a09d2c3),
	.w8(32'h3a7ba383),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1f970),
	.w1(32'hba995ae6),
	.w2(32'hbae197a1),
	.w3(32'h382ff499),
	.w4(32'h39690180),
	.w5(32'h3a49ea0e),
	.w6(32'h39d0b3cf),
	.w7(32'h3ab8868c),
	.w8(32'h3a76959d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38822644),
	.w1(32'hb9693593),
	.w2(32'hb9d4b93b),
	.w3(32'h3903371b),
	.w4(32'hb9a82937),
	.w5(32'hb9b4bc18),
	.w6(32'hb9fe1aaf),
	.w7(32'hb9fe5441),
	.w8(32'hb8d57b0d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fccda7),
	.w1(32'h39c02f35),
	.w2(32'h391aaceb),
	.w3(32'h394a8771),
	.w4(32'hb867f28b),
	.w5(32'hb98bc6eb),
	.w6(32'hb7edf5a8),
	.w7(32'hb995bb16),
	.w8(32'hb9ceef4d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a254fd),
	.w1(32'h388415f4),
	.w2(32'h38b015a2),
	.w3(32'hb89cb9ed),
	.w4(32'hb85bbd99),
	.w5(32'hb86be5e4),
	.w6(32'hb8d45920),
	.w7(32'hb7b58818),
	.w8(32'h38784b87),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa11acf),
	.w1(32'hba7e5dab),
	.w2(32'hb9f14970),
	.w3(32'hb9bf91a6),
	.w4(32'hb9e1b548),
	.w5(32'h3a284dcf),
	.w6(32'hb992261b),
	.w7(32'h3a8de272),
	.w8(32'h3ab0691a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad8759),
	.w1(32'hb9b83e88),
	.w2(32'hba014d4e),
	.w3(32'hbab3758a),
	.w4(32'hbaf1a11c),
	.w5(32'hba473c01),
	.w6(32'h3a9a009f),
	.w7(32'h396a1206),
	.w8(32'h3a704df4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfba26b),
	.w1(32'h3b98a2f3),
	.w2(32'h3b7ac904),
	.w3(32'h3ba92e4e),
	.w4(32'h3af7d29b),
	.w5(32'h39cdfe89),
	.w6(32'h3be01b6a),
	.w7(32'h3b977449),
	.w8(32'h3b0c6e53),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979ff94),
	.w1(32'hba101a1d),
	.w2(32'hba42749f),
	.w3(32'h39ce6ff3),
	.w4(32'hba0c1f27),
	.w5(32'hba787aad),
	.w6(32'h3a864574),
	.w7(32'hb8f3ee53),
	.w8(32'hb963ebdc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92e4b7),
	.w1(32'hb9fe56d6),
	.w2(32'h37c88cd7),
	.w3(32'h3b1a8ff8),
	.w4(32'hb908d55c),
	.w5(32'hb9805f74),
	.w6(32'h3ba800d3),
	.w7(32'h3b40407c),
	.w8(32'h3b4fb2f2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac166e0),
	.w1(32'h39986192),
	.w2(32'hb93c413a),
	.w3(32'h3951ff18),
	.w4(32'h3a817017),
	.w5(32'h3a1496fa),
	.w6(32'h3a710747),
	.w7(32'h3ad3f964),
	.w8(32'h3a072e77),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9013bdb),
	.w1(32'h38201df9),
	.w2(32'h37bf1de2),
	.w3(32'hb88b246f),
	.w4(32'h390b4dd2),
	.w5(32'h38a4e5ea),
	.w6(32'h36ed1f91),
	.w7(32'hb5bd395a),
	.w8(32'h38f4347e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9932a34),
	.w1(32'h3a1908bc),
	.w2(32'h3a4ae1c2),
	.w3(32'h3a342895),
	.w4(32'h38c35a40),
	.w5(32'h3894b630),
	.w6(32'h39d91a1f),
	.w7(32'h39e8471f),
	.w8(32'hb9a1269d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3626cad4),
	.w1(32'hb8b53fca),
	.w2(32'h37af7342),
	.w3(32'h38536f5d),
	.w4(32'hb72ba02f),
	.w5(32'h3895a1ba),
	.w6(32'hb9a50e5a),
	.w7(32'hb98afebc),
	.w8(32'hb90e7db7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269249),
	.w1(32'hba14e6b7),
	.w2(32'h3995f4c8),
	.w3(32'h3b0380b0),
	.w4(32'hba3bbb53),
	.w5(32'hba1d5e19),
	.w6(32'h3b8a5a94),
	.w7(32'h3aecb2f2),
	.w8(32'h3aee2403),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1d10d),
	.w1(32'h3ad4a2ed),
	.w2(32'hba803a3e),
	.w3(32'h3b525ad1),
	.w4(32'hbaf615ae),
	.w5(32'hbb6c9308),
	.w6(32'h3bbcda04),
	.w7(32'h3a1d6e64),
	.w8(32'hba33cc13),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cc222),
	.w1(32'h3a8ef2da),
	.w2(32'h382e9c42),
	.w3(32'h3b3e560e),
	.w4(32'h3997a8fa),
	.w5(32'hba7ffd3f),
	.w6(32'h3bad21e5),
	.w7(32'h3b39392b),
	.w8(32'h3ac26d14),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39643151),
	.w1(32'hba8a4873),
	.w2(32'hbab7e798),
	.w3(32'h39c3e405),
	.w4(32'hba86d27b),
	.w5(32'hbae1688c),
	.w6(32'h39c403b2),
	.w7(32'hba1b49e2),
	.w8(32'hba4c7fa7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e46c4),
	.w1(32'h3b5cb999),
	.w2(32'h3b286a8b),
	.w3(32'h3b41b99c),
	.w4(32'hb8f5b83a),
	.w5(32'hba213121),
	.w6(32'h3bbb3d47),
	.w7(32'h3b3ff0c8),
	.w8(32'h3afdb939),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac01fa),
	.w1(32'h3aa8b673),
	.w2(32'h3af3efac),
	.w3(32'h3aceb577),
	.w4(32'h39c88307),
	.w5(32'h3a29adc5),
	.w6(32'h3b53089d),
	.w7(32'h3b1965c3),
	.w8(32'h3acaa956),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc4627),
	.w1(32'h3b01bebd),
	.w2(32'h3b044e2c),
	.w3(32'h3bdc54ea),
	.w4(32'h3b439f51),
	.w5(32'h3afd90ad),
	.w6(32'h3c0311f7),
	.w7(32'h3bbf20e1),
	.w8(32'h3ba1d5a6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cc802),
	.w1(32'h39522a20),
	.w2(32'h395e7c25),
	.w3(32'hb8db80fa),
	.w4(32'h3968710f),
	.w5(32'h39817666),
	.w6(32'h39508c4c),
	.w7(32'h397287b2),
	.w8(32'h3991d745),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947aacf),
	.w1(32'hb9440198),
	.w2(32'hb9888751),
	.w3(32'h3996fc35),
	.w4(32'h381f993d),
	.w5(32'h3617a48b),
	.w6(32'hb8c6e670),
	.w7(32'hb993f973),
	.w8(32'hb9184d23),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd79903),
	.w1(32'h3b8ffc6a),
	.w2(32'h3937db9e),
	.w3(32'hb9b0ae74),
	.w4(32'hba43b65e),
	.w5(32'hbad8b6ad),
	.w6(32'h3b4d4387),
	.w7(32'h3b453a2b),
	.w8(32'h3b1a3160),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c3fd),
	.w1(32'h3b5d9924),
	.w2(32'h3b43ac94),
	.w3(32'h3b6b068a),
	.w4(32'h3acf114a),
	.w5(32'h3b1001ef),
	.w6(32'h3bd1b297),
	.w7(32'h3b609550),
	.w8(32'h3b804f5a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d0bd),
	.w1(32'h3b24bb22),
	.w2(32'h3ae78ae8),
	.w3(32'h3b2b615b),
	.w4(32'hb9f9a539),
	.w5(32'hbaa325f3),
	.w6(32'h3ba68527),
	.w7(32'h3b224b22),
	.w8(32'h3ab9ce08),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00df65),
	.w1(32'hbc038b10),
	.w2(32'hbb8cb446),
	.w3(32'hba47864c),
	.w4(32'hba1477a8),
	.w5(32'h3ace7fed),
	.w6(32'h3ad75bdc),
	.w7(32'h3a8b8109),
	.w8(32'h3ad2060b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9337a63),
	.w1(32'hb918cc85),
	.w2(32'h394e1b0c),
	.w3(32'hb9bca765),
	.w4(32'hb8b59468),
	.w5(32'hb923f8ba),
	.w6(32'hb856ea15),
	.w7(32'h3736d9d5),
	.w8(32'h37cebd81),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fca33d),
	.w1(32'hb8937640),
	.w2(32'h3a18b8c5),
	.w3(32'h3929304f),
	.w4(32'hb7f3c13c),
	.w5(32'h3a009e57),
	.w6(32'hb82a0e00),
	.w7(32'h3a15939b),
	.w8(32'h39cc9210),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b605608),
	.w1(32'hbaf45275),
	.w2(32'hbad2644c),
	.w3(32'hb934e09b),
	.w4(32'hbb184bb1),
	.w5(32'h3a5ca59d),
	.w6(32'hb8f1d06d),
	.w7(32'hba407ea1),
	.w8(32'hba8607c3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cbc80),
	.w1(32'h3aaf025d),
	.w2(32'h3b764ee1),
	.w3(32'h3b337f69),
	.w4(32'h3adf9d6e),
	.w5(32'h3b38be15),
	.w6(32'h3b9f905d),
	.w7(32'h3b8fbcea),
	.w8(32'h3bab433f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f12e0),
	.w1(32'h3a878096),
	.w2(32'hba913664),
	.w3(32'hb9af74e4),
	.w4(32'h3acd9290),
	.w5(32'h3a4b8463),
	.w6(32'h39f16ce0),
	.w7(32'h3a8c82d5),
	.w8(32'hb95e2837),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b5bde),
	.w1(32'hba3e453b),
	.w2(32'hbb111065),
	.w3(32'h3b23ac36),
	.w4(32'hbb11c25c),
	.w5(32'hbb8434ba),
	.w6(32'h3b7f87e8),
	.w7(32'h397f69bb),
	.w8(32'hbab54aa4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e214),
	.w1(32'h3b569b0a),
	.w2(32'h39d61395),
	.w3(32'h3b950a3d),
	.w4(32'h3a9a521c),
	.w5(32'hbb06b877),
	.w6(32'h3bc98029),
	.w7(32'h3b3c8a7e),
	.w8(32'h39bf4a6c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ca30a),
	.w1(32'h38a2612d),
	.w2(32'h38af3bd6),
	.w3(32'hb94cac41),
	.w4(32'h37452369),
	.w5(32'h37acfb78),
	.w6(32'h37e2b42c),
	.w7(32'h38175185),
	.w8(32'h390293d3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cc5320),
	.w1(32'hb8a114c2),
	.w2(32'h37fb04c7),
	.w3(32'hb7a6da7f),
	.w4(32'h3702b297),
	.w5(32'h3895f902),
	.w6(32'h394a6ed9),
	.w7(32'h38f75b23),
	.w8(32'h3872a594),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f539),
	.w1(32'hba85fcaa),
	.w2(32'hb9818e86),
	.w3(32'hbb065a26),
	.w4(32'hb9f7130b),
	.w5(32'h389d75b2),
	.w6(32'hba339c95),
	.w7(32'h39cdc8a3),
	.w8(32'h3aabdeae),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897809b),
	.w1(32'hb88f6d32),
	.w2(32'hb9bc5eef),
	.w3(32'hb9073816),
	.w4(32'hb8c4122f),
	.w5(32'hb9842acf),
	.w6(32'hb8185a5e),
	.w7(32'hb97614c9),
	.w8(32'h38934d3f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78a5e4),
	.w1(32'h3aa9b23c),
	.w2(32'h3a438e0d),
	.w3(32'hbaa16cd8),
	.w4(32'h3a28e049),
	.w5(32'h3a9a51c3),
	.w6(32'hba0e7caf),
	.w7(32'h3ab36dd5),
	.w8(32'h3abb8a24),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b459091),
	.w1(32'h3b00f103),
	.w2(32'h3b348a08),
	.w3(32'h3a9a7606),
	.w4(32'hb968584b),
	.w5(32'h3950e3b0),
	.w6(32'h3b5bf2b0),
	.w7(32'h3abcc144),
	.w8(32'h3b4d3486),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad83653),
	.w1(32'h3a075fc8),
	.w2(32'hb955ffb3),
	.w3(32'h3b12121f),
	.w4(32'h3a0bedb0),
	.w5(32'h3a17b678),
	.w6(32'h3b3f3f36),
	.w7(32'h3ad9a8a6),
	.w8(32'h3ad6c03e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96dccb1),
	.w1(32'hb8a9f5dd),
	.w2(32'h39c39942),
	.w3(32'hb98bb584),
	.w4(32'hb976e4d5),
	.w5(32'h39653dfd),
	.w6(32'h37f5d7ce),
	.w7(32'h38fab502),
	.w8(32'hb9179379),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91df58),
	.w1(32'hba3ab89f),
	.w2(32'hbb322c45),
	.w3(32'h3a445559),
	.w4(32'h3a8fd312),
	.w5(32'h39ebf53a),
	.w6(32'h3b584d40),
	.w7(32'h3b361b57),
	.w8(32'h3a78b41e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad71608),
	.w1(32'h3891e491),
	.w2(32'h3a41f891),
	.w3(32'h3ac71157),
	.w4(32'h39b96943),
	.w5(32'h39c3eb9b),
	.w6(32'h3ae5776f),
	.w7(32'h3aa04dfa),
	.w8(32'h3aa7ab89),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386ff214),
	.w1(32'h395df02c),
	.w2(32'h3938bb8b),
	.w3(32'h38d8d74d),
	.w4(32'h3995169b),
	.w5(32'h399c91a5),
	.w6(32'h392be07c),
	.w7(32'h393531ae),
	.w8(32'h39a862fb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285ae7),
	.w1(32'hbb5ab3c3),
	.w2(32'hbaf5f4c6),
	.w3(32'hb9fab350),
	.w4(32'hbacb549c),
	.w5(32'hba084c32),
	.w6(32'h3a324b45),
	.w7(32'hb7467563),
	.w8(32'hb84a7b90),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8b55b),
	.w1(32'h39b52f1f),
	.w2(32'h39c99733),
	.w3(32'h399aa438),
	.w4(32'h3987e7bb),
	.w5(32'h38e3ccc7),
	.w6(32'h39a9c1f3),
	.w7(32'h3986783f),
	.w8(32'h3938b61c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39628e26),
	.w1(32'h39a7a5be),
	.w2(32'h39e06430),
	.w3(32'h39a1b5e3),
	.w4(32'h3a19beb2),
	.w5(32'h3a3517ab),
	.w6(32'h39ee6edb),
	.w7(32'h3a10013b),
	.w8(32'h39cd442f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916b457),
	.w1(32'h3954feec),
	.w2(32'h390d5cdd),
	.w3(32'h37d8e441),
	.w4(32'h3968a3c2),
	.w5(32'h392fbf6f),
	.w6(32'h392e2ff5),
	.w7(32'h3917d804),
	.w8(32'h396f3641),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe2e5d),
	.w1(32'hb8afbb30),
	.w2(32'hb8d38492),
	.w3(32'h39628a67),
	.w4(32'hb892f2a3),
	.w5(32'hb93a1e37),
	.w6(32'hb8eb6817),
	.w7(32'hb89c3e26),
	.w8(32'h394fb2f8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc3a9),
	.w1(32'hb997c200),
	.w2(32'hba99c9cf),
	.w3(32'h3a1f661f),
	.w4(32'hba374557),
	.w5(32'hbae15f52),
	.w6(32'h3ac5b37e),
	.w7(32'h396b92a4),
	.w8(32'hb88c4599),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118646),
	.w1(32'hbb73ed88),
	.w2(32'h3a54b99a),
	.w3(32'h3b30a52f),
	.w4(32'h3a01ce09),
	.w5(32'h3b412081),
	.w6(32'h3bb4e903),
	.w7(32'h3b40928b),
	.w8(32'h3b68cfdd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dd12c),
	.w1(32'hbaaf0427),
	.w2(32'h3aa10e42),
	.w3(32'h3a3ec640),
	.w4(32'hb9ff36ea),
	.w5(32'h3ae47f2a),
	.w6(32'h3b1bba4c),
	.w7(32'h3aa037a6),
	.w8(32'h3aa6c117),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c34672),
	.w1(32'hba03a467),
	.w2(32'h3b7103a1),
	.w3(32'h3b03a6ad),
	.w4(32'h3b1edc8c),
	.w5(32'h3bb5e31f),
	.w6(32'h3b9262b0),
	.w7(32'h3b80054a),
	.w8(32'h3bbdddc2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5a598),
	.w1(32'hb86cce23),
	.w2(32'hb991429d),
	.w3(32'h3983b5b3),
	.w4(32'hb9074f79),
	.w5(32'hb98b332b),
	.w6(32'h37c97597),
	.w7(32'h38a060a9),
	.w8(32'h3984062c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e473c7),
	.w1(32'h384ff7b2),
	.w2(32'h3a0f482a),
	.w3(32'hb984e8a1),
	.w4(32'h3905052e),
	.w5(32'h39877fd9),
	.w6(32'hb88548df),
	.w7(32'h39524cc5),
	.w8(32'h3a08c64b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988e0ee),
	.w1(32'h396454b0),
	.w2(32'h396e521a),
	.w3(32'h39b35b1f),
	.w4(32'h3980aedf),
	.w5(32'h3968ca37),
	.w6(32'h393c6e07),
	.w7(32'h392a7b7f),
	.w8(32'h3959cace),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938da4b),
	.w1(32'h3958f4a4),
	.w2(32'h395caa8f),
	.w3(32'h399445c5),
	.w4(32'h3981c89f),
	.w5(32'h39615bc9),
	.w6(32'h3977b6de),
	.w7(32'h393050d5),
	.w8(32'h394614eb),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41527),
	.w1(32'h3890972c),
	.w2(32'h3b596580),
	.w3(32'hb96446c5),
	.w4(32'hba88ed05),
	.w5(32'h3aa4e070),
	.w6(32'h3a82e649),
	.w7(32'h3a0ef8b8),
	.w8(32'h3b22ea75),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25d591),
	.w1(32'h377b3add),
	.w2(32'h398604ef),
	.w3(32'hb9e7f873),
	.w4(32'hb9b305c4),
	.w5(32'hb92e1716),
	.w6(32'hb9cc195a),
	.w7(32'hb9b4f422),
	.w8(32'hb9589e73),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80ed21),
	.w1(32'hba2c5779),
	.w2(32'hbb09b8a5),
	.w3(32'h3a47b8f8),
	.w4(32'hb99b2a4d),
	.w5(32'hbb0329c2),
	.w6(32'h3a2ceb9d),
	.w7(32'hb945e587),
	.w8(32'hbab4228b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976dfcf),
	.w1(32'h38327ae1),
	.w2(32'hba482ed5),
	.w3(32'h38a2930a),
	.w4(32'hba0cf9d2),
	.w5(32'hba435c70),
	.w6(32'hb8f2b740),
	.w7(32'hb9f4f051),
	.w8(32'hba0f60fd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992acf5),
	.w1(32'h39a08e45),
	.w2(32'h3996d39f),
	.w3(32'hb996be5a),
	.w4(32'h39993243),
	.w5(32'h3981b2cd),
	.w6(32'h39523958),
	.w7(32'h393d24c0),
	.w8(32'h398513a9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a747088),
	.w1(32'hb90a98ab),
	.w2(32'h3a8cc1ad),
	.w3(32'h3a7b6e7c),
	.w4(32'h38d46c8d),
	.w5(32'h3a58d07e),
	.w6(32'h3a701720),
	.w7(32'h3a63e2ba),
	.w8(32'h3abbf112),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949d4f),
	.w1(32'h391cb25a),
	.w2(32'h39acccc9),
	.w3(32'hb9504590),
	.w4(32'h397dab2d),
	.w5(32'h396e4721),
	.w6(32'h38b19c81),
	.w7(32'h36cac83b),
	.w8(32'h396bd3c5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850eeb),
	.w1(32'hbba8b4a7),
	.w2(32'h3a45da35),
	.w3(32'hbac69677),
	.w4(32'hba659611),
	.w5(32'h3aed1e9b),
	.w6(32'h3b390927),
	.w7(32'h39353994),
	.w8(32'h3b1c8cd9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ea837),
	.w1(32'hba46334c),
	.w2(32'h3a1f584f),
	.w3(32'hb92a4710),
	.w4(32'hbb8ea684),
	.w5(32'hba38cb47),
	.w6(32'hba180937),
	.w7(32'h3bc6c018),
	.w8(32'h3ad3b0c4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa8606),
	.w1(32'h3b22824d),
	.w2(32'h3a87f1e7),
	.w3(32'h3bbc5a5e),
	.w4(32'hbaea22cb),
	.w5(32'hbac0f8b5),
	.w6(32'h3b41ed31),
	.w7(32'hb9e905f2),
	.w8(32'hbb8fb335),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule