module layer_10_featuremap_393(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2e25c),
	.w1(32'hbb9f7171),
	.w2(32'hbb3a428b),
	.w3(32'h3b1a3e7e),
	.w4(32'hbb923dca),
	.w5(32'h3b0ca28e),
	.w6(32'h3af99c94),
	.w7(32'hbb6cd646),
	.w8(32'hbb6bad7c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a36d),
	.w1(32'hbb984d25),
	.w2(32'hbb133a63),
	.w3(32'hbbc8ac9f),
	.w4(32'hbb3c4e07),
	.w5(32'hbac0ddf3),
	.w6(32'hbb998e78),
	.w7(32'hbac51df5),
	.w8(32'hba31a1d1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b45d1),
	.w1(32'hbb2ce074),
	.w2(32'hb99c0d66),
	.w3(32'hbaa9984d),
	.w4(32'h3b541667),
	.w5(32'h3bf1e278),
	.w6(32'hbb4aa9ca),
	.w7(32'h3ba441d6),
	.w8(32'h3be8f155),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca87e7),
	.w1(32'h3b032e32),
	.w2(32'hb9a5375f),
	.w3(32'h3be935ca),
	.w4(32'h3b70ecc1),
	.w5(32'hbc162c45),
	.w6(32'h3bd6fcff),
	.w7(32'h3b12df63),
	.w8(32'hbb00135c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbab3c8),
	.w1(32'h3bc0c7be),
	.w2(32'h3b9ae1f9),
	.w3(32'hbb8eaf14),
	.w4(32'h3b872fb8),
	.w5(32'h3bf84242),
	.w6(32'hbb276474),
	.w7(32'hbaf6a0ba),
	.w8(32'h3a4460f0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34c89),
	.w1(32'h3c18d3ff),
	.w2(32'h3c805424),
	.w3(32'h3bb1979b),
	.w4(32'hb98b8de1),
	.w5(32'h3c0a9648),
	.w6(32'h3b86681e),
	.w7(32'hbb0a4e95),
	.w8(32'hbb400f6e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16da9a),
	.w1(32'hbac7ad4a),
	.w2(32'h3b335200),
	.w3(32'h3c88fc55),
	.w4(32'h3a1f6439),
	.w5(32'hbb89296f),
	.w6(32'h3bd86c93),
	.w7(32'hba12dfbc),
	.w8(32'hbbb45a15),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef575b),
	.w1(32'hbb27973e),
	.w2(32'h3af87c29),
	.w3(32'h3a92c1e0),
	.w4(32'h38762b5c),
	.w5(32'h3b8f4735),
	.w6(32'h3b334541),
	.w7(32'h3a953a61),
	.w8(32'h3b21997f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f49ee5),
	.w1(32'h3b61741e),
	.w2(32'hbb13e59d),
	.w3(32'h3b57b84e),
	.w4(32'h3b7f1eeb),
	.w5(32'hbb562dc7),
	.w6(32'hb9584e5f),
	.w7(32'h3b3f4ce9),
	.w8(32'h3ae43c8f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a304874),
	.w1(32'h3b331c37),
	.w2(32'h3b4591b7),
	.w3(32'hbb85aaca),
	.w4(32'hbaceb688),
	.w5(32'hbbc34393),
	.w6(32'hb8487ccb),
	.w7(32'hbb2a0542),
	.w8(32'hbb82d70c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b577),
	.w1(32'h39b6fe39),
	.w2(32'hbb238043),
	.w3(32'hbb051328),
	.w4(32'h39ef58e5),
	.w5(32'h3abc07c3),
	.w6(32'h3aff5bb2),
	.w7(32'hba2aa858),
	.w8(32'hbb05525e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de46b4),
	.w1(32'h3bb867d2),
	.w2(32'h3a2352ce),
	.w3(32'hba985529),
	.w4(32'h3bd20dd8),
	.w5(32'h3aacf2fa),
	.w6(32'hbb5b56e3),
	.w7(32'h3be7cf1a),
	.w8(32'h3c251da3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8f024),
	.w1(32'hb930a0ec),
	.w2(32'hba3d73c8),
	.w3(32'hbbc6331c),
	.w4(32'h3b2b086c),
	.w5(32'hbc187501),
	.w6(32'h3a49116d),
	.w7(32'h3bc639d0),
	.w8(32'h3b9bb821),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3df991),
	.w1(32'hbb23dc65),
	.w2(32'hba45a825),
	.w3(32'h3a5d4ec8),
	.w4(32'h3b767b82),
	.w5(32'h3b749d19),
	.w6(32'h3ac90446),
	.w7(32'hbb21c77f),
	.w8(32'hba96ab4b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba912fa8),
	.w1(32'h3b5933c1),
	.w2(32'h3bd9251d),
	.w3(32'h3a95b404),
	.w4(32'h3bc35172),
	.w5(32'h3bde7f2b),
	.w6(32'hbad54e80),
	.w7(32'h3b24cdfd),
	.w8(32'h3bec2751),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc9a5c),
	.w1(32'h3b6681f8),
	.w2(32'h3b918b51),
	.w3(32'h3be7a1cc),
	.w4(32'h3c557317),
	.w5(32'hb9c9d578),
	.w6(32'h3bca3666),
	.w7(32'h3c2158d0),
	.w8(32'h3c0b12c9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60895c),
	.w1(32'hbaa008ff),
	.w2(32'hba866ab6),
	.w3(32'h3aba8791),
	.w4(32'h390d61da),
	.w5(32'hbb99656c),
	.w6(32'hba192ee3),
	.w7(32'h3b303b83),
	.w8(32'h3a8e90cd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349470),
	.w1(32'h3bf52f92),
	.w2(32'h3bbd5e0b),
	.w3(32'h3bc5bbac),
	.w4(32'h3c0d6342),
	.w5(32'h3bf2bf0c),
	.w6(32'h3bb33ddc),
	.w7(32'h3bcd1071),
	.w8(32'h3b03bc90),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b129c5a),
	.w1(32'h3c4b95b7),
	.w2(32'h3b609411),
	.w3(32'hbafae3da),
	.w4(32'h3c52a224),
	.w5(32'h3ba463e1),
	.w6(32'hbb03be9e),
	.w7(32'h3c34f6a4),
	.w8(32'h3c2f2753),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c20c0),
	.w1(32'hbb90f3cf),
	.w2(32'h3a0b45df),
	.w3(32'h3a3e10b7),
	.w4(32'hbc208681),
	.w5(32'h3aa2f703),
	.w6(32'h39eb51e8),
	.w7(32'hbc06c18f),
	.w8(32'hbbfc8e06),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e3bac),
	.w1(32'h3b7acc52),
	.w2(32'h3b80f83a),
	.w3(32'h3c76e04b),
	.w4(32'hbb03e09d),
	.w5(32'h3b35b88a),
	.w6(32'hbb2d1b69),
	.w7(32'hbb085b1e),
	.w8(32'h3b961efe),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e1b4a),
	.w1(32'hbb065c93),
	.w2(32'hbacc673d),
	.w3(32'h3b6eeafc),
	.w4(32'hbbae4802),
	.w5(32'hbb5c4f81),
	.w6(32'h3b235c11),
	.w7(32'hbb1de4b0),
	.w8(32'hbb3342f1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64e2ee),
	.w1(32'h3c75d6b9),
	.w2(32'h3c973213),
	.w3(32'h3cccc6c6),
	.w4(32'h3c0638a9),
	.w5(32'h3bdf4cf7),
	.w6(32'h3c8e0f6f),
	.w7(32'h3b993cbe),
	.w8(32'h3bde3867),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e1ad),
	.w1(32'hbae6c43a),
	.w2(32'hbb3fb178),
	.w3(32'h3a3ca2e0),
	.w4(32'h39273031),
	.w5(32'h3aa3fcb9),
	.w6(32'hbb3f339d),
	.w7(32'hb9e26d06),
	.w8(32'h3b1273c2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23918e),
	.w1(32'hbb27d5ef),
	.w2(32'h39d450a4),
	.w3(32'hbb6caa57),
	.w4(32'hbb5f443f),
	.w5(32'hbbd1dbf8),
	.w6(32'hbb3db5a5),
	.w7(32'h3bba535a),
	.w8(32'h3b689def),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c320c24),
	.w1(32'hbb890c87),
	.w2(32'h3c2c60a3),
	.w3(32'h3bcbdd94),
	.w4(32'hbbf024b8),
	.w5(32'h3c0ebc0a),
	.w6(32'hba17d4c6),
	.w7(32'hbbe3361b),
	.w8(32'hbb785fa6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba5b0a),
	.w1(32'h39f07544),
	.w2(32'h3b8f432f),
	.w3(32'h3b6edd59),
	.w4(32'h3a893e57),
	.w5(32'h3b5af220),
	.w6(32'h3b3af234),
	.w7(32'hba550e2b),
	.w8(32'h3b83a5eb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9796a8),
	.w1(32'hb95e763c),
	.w2(32'hba585e24),
	.w3(32'h39a8cc0d),
	.w4(32'hb941175b),
	.w5(32'hbad7c025),
	.w6(32'hbb16c0b3),
	.w7(32'h39ac61d1),
	.w8(32'hbb7599c4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b7888),
	.w1(32'h3af65054),
	.w2(32'hbac689df),
	.w3(32'hbb2528fa),
	.w4(32'hbb1165f8),
	.w5(32'hbbc61c3c),
	.w6(32'hbb8da2a9),
	.w7(32'hbab2a291),
	.w8(32'h39291589),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981367),
	.w1(32'h3b2a72eb),
	.w2(32'h3bc6e0ae),
	.w3(32'hbb30e635),
	.w4(32'hba61f0a1),
	.w5(32'h3b9f3ce8),
	.w6(32'hbb45d65f),
	.w7(32'hb9ffa9c0),
	.w8(32'h3b8148aa),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3288),
	.w1(32'h3a8019c2),
	.w2(32'h39364c4e),
	.w3(32'h39fc0744),
	.w4(32'h3b9a36b9),
	.w5(32'h3b93a2c2),
	.w6(32'hb935db85),
	.w7(32'hba92e137),
	.w8(32'hb9e57d66),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3990f),
	.w1(32'hbb13f234),
	.w2(32'h3b796858),
	.w3(32'hbb7a8bd4),
	.w4(32'h3b8d6813),
	.w5(32'h3b53355d),
	.w6(32'hbb09770d),
	.w7(32'h3b7f26f4),
	.w8(32'h3b1d67e7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35b613),
	.w1(32'hbbf6fea5),
	.w2(32'hbb8b6dce),
	.w3(32'h3b4abe8a),
	.w4(32'hbbaf1aa1),
	.w5(32'hbc229cf0),
	.w6(32'h3bea4853),
	.w7(32'hbb2578c9),
	.w8(32'hbbd0dad0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42017),
	.w1(32'hbb87d8f1),
	.w2(32'h3b8feb1d),
	.w3(32'hbb96c2b9),
	.w4(32'hbaf06a87),
	.w5(32'hbb2bc723),
	.w6(32'hbb1cb664),
	.w7(32'hbb4cc33a),
	.w8(32'hbba1285a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83f196),
	.w1(32'hbabccb0f),
	.w2(32'h3b76d4e3),
	.w3(32'h3928dd39),
	.w4(32'h397aa65b),
	.w5(32'h3b894022),
	.w6(32'hbb477722),
	.w7(32'hba8f2169),
	.w8(32'hb9dba3fc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b030ff3),
	.w1(32'hbaf0f0d7),
	.w2(32'hbb478b19),
	.w3(32'h3b627cc3),
	.w4(32'hbb175c61),
	.w5(32'hbc180daa),
	.w6(32'h3b3080b0),
	.w7(32'hba50c0a4),
	.w8(32'hbb8263f5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10a178),
	.w1(32'h3ab76b41),
	.w2(32'h39c3a38d),
	.w3(32'hbb159a4c),
	.w4(32'h3a4fd7e9),
	.w5(32'hbb247fb5),
	.w6(32'h3aa64c28),
	.w7(32'h3b931bfd),
	.w8(32'hbb95a730),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fa090),
	.w1(32'hbbe3caa5),
	.w2(32'h3ae3c4fa),
	.w3(32'hbc65b178),
	.w4(32'hbc196e94),
	.w5(32'hbb2fba60),
	.w6(32'hbbae0aef),
	.w7(32'hbbb3edf2),
	.w8(32'hb9218d69),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8750bd),
	.w1(32'hbbc5fe93),
	.w2(32'hbbb5c870),
	.w3(32'hbba3077e),
	.w4(32'hbb030fb1),
	.w5(32'h3be73530),
	.w6(32'hbb5fedd1),
	.w7(32'hbbd4579c),
	.w8(32'hbb364035),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed1e3c),
	.w1(32'hbc190911),
	.w2(32'hbbe063ac),
	.w3(32'hbadbbea5),
	.w4(32'hbbe1b77d),
	.w5(32'hbb62b184),
	.w6(32'hbbbd2fc0),
	.w7(32'hbbd4071d),
	.w8(32'hbba1e1f2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1434aa),
	.w1(32'h3a35120c),
	.w2(32'h3a5a61c0),
	.w3(32'hbae52780),
	.w4(32'h3b2b1759),
	.w5(32'hbbc296ea),
	.w6(32'hbb10d6fb),
	.w7(32'h39dba46b),
	.w8(32'hbb9b440b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d5f9),
	.w1(32'hba20a99b),
	.w2(32'hba7c4af5),
	.w3(32'hbbbf575e),
	.w4(32'hbb86ef59),
	.w5(32'hbaeae709),
	.w6(32'hbbad1b4b),
	.w7(32'hbb2ca971),
	.w8(32'hbb425ecc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2d18a),
	.w1(32'hbba51b68),
	.w2(32'h3923f798),
	.w3(32'hbb49c8fb),
	.w4(32'hbae585ae),
	.w5(32'hbc050858),
	.w6(32'hba8079a6),
	.w7(32'hbaee9a5e),
	.w8(32'hbae6312c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bec33),
	.w1(32'h3bc5c700),
	.w2(32'h3b6dc481),
	.w3(32'hb942bcd2),
	.w4(32'h3bf1fc26),
	.w5(32'h3c1d61e5),
	.w6(32'hbb3a3d89),
	.w7(32'h3b3c51d7),
	.w8(32'h3ace6f86),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37ce90),
	.w1(32'h3b336305),
	.w2(32'hbb66daa1),
	.w3(32'h3a8a0ad8),
	.w4(32'h3aa3d267),
	.w5(32'hbbd54c63),
	.w6(32'h3b02be1f),
	.w7(32'h3a9bb5d3),
	.w8(32'h3a1bec3b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fda3),
	.w1(32'h3b782fb0),
	.w2(32'h383602de),
	.w3(32'hbb1973c3),
	.w4(32'h3c172701),
	.w5(32'hbb523525),
	.w6(32'h3ac47ad5),
	.w7(32'h3c17d66c),
	.w8(32'h3bc8c124),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b580d42),
	.w1(32'h3a03e1f4),
	.w2(32'hba41685f),
	.w3(32'h3ad04e34),
	.w4(32'h3bb29a45),
	.w5(32'hbbb04663),
	.w6(32'h3b1465ad),
	.w7(32'hba9ba5d3),
	.w8(32'h3b05f365),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0546b),
	.w1(32'h3c5d76cd),
	.w2(32'h3bd67182),
	.w3(32'h3baaab4e),
	.w4(32'h3c19f900),
	.w5(32'h3a495846),
	.w6(32'h3c288ce1),
	.w7(32'h3b96a979),
	.w8(32'h3af465a9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970e17),
	.w1(32'h3b158a04),
	.w2(32'h3bb05ea4),
	.w3(32'hbb4cc19d),
	.w4(32'h3b68bbd7),
	.w5(32'h3bbfdc15),
	.w6(32'hbb99adaa),
	.w7(32'hba49217a),
	.w8(32'h3a3f04aa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbec062),
	.w1(32'h3b0f572a),
	.w2(32'h3b73f5f8),
	.w3(32'h3c240f33),
	.w4(32'h3b32029c),
	.w5(32'h3979042b),
	.w6(32'h3baf8fac),
	.w7(32'h3b418acb),
	.w8(32'h39b69009),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20082d),
	.w1(32'h3bbc074d),
	.w2(32'hba6ac3c5),
	.w3(32'hbb952a4a),
	.w4(32'h3b954a33),
	.w5(32'h3a43e6c7),
	.w6(32'hb901bbe8),
	.w7(32'h3ba464f3),
	.w8(32'h3bf03e16),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02cd59),
	.w1(32'hbb106062),
	.w2(32'hbaae712d),
	.w3(32'hb80e22ea),
	.w4(32'h3b0f96e3),
	.w5(32'hbb909e4e),
	.w6(32'h3a5ff26d),
	.w7(32'h3baf228c),
	.w8(32'hbb033bd3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c8202),
	.w1(32'h3ae83ec4),
	.w2(32'h3bd99917),
	.w3(32'h3ba556ce),
	.w4(32'h3b211193),
	.w5(32'h3bc1a42f),
	.w6(32'h39500a77),
	.w7(32'hb9838546),
	.w8(32'h3995099d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7300b),
	.w1(32'hbbac7df4),
	.w2(32'hbbd80adb),
	.w3(32'h3c22a5bc),
	.w4(32'hbaaeae1d),
	.w5(32'hbb722bd0),
	.w6(32'h3bbfffd4),
	.w7(32'hbb934935),
	.w8(32'hbb05276b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb63392),
	.w1(32'hbaf3d77d),
	.w2(32'h3a7dd177),
	.w3(32'hbba4b0fb),
	.w4(32'hb9c21400),
	.w5(32'hbb8223b6),
	.w6(32'hbb3579e0),
	.w7(32'h3b2c9da2),
	.w8(32'hbb5fc2c0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befaf47),
	.w1(32'hbb62a12e),
	.w2(32'h3b0088e3),
	.w3(32'h3b584695),
	.w4(32'hbbe72a00),
	.w5(32'h3991a970),
	.w6(32'hbab5b1cf),
	.w7(32'hbc30c50c),
	.w8(32'hbb3b3163),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919237d),
	.w1(32'h3bc82e25),
	.w2(32'h3a3baca2),
	.w3(32'hba38824a),
	.w4(32'h3bcd6498),
	.w5(32'hbb2596ec),
	.w6(32'hbb042230),
	.w7(32'h3b3552a8),
	.w8(32'h3b92a77b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64dd9a),
	.w1(32'hbbc7c0d9),
	.w2(32'h3b172605),
	.w3(32'h3b97c75b),
	.w4(32'hbbf8aba8),
	.w5(32'h3a44fbed),
	.w6(32'h3affa857),
	.w7(32'hbba17c8e),
	.w8(32'hbc3a95bb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef9ac),
	.w1(32'hbacc0b1e),
	.w2(32'h3bc2530b),
	.w3(32'h3b50fc2f),
	.w4(32'hbba7cc8b),
	.w5(32'h3b14ffce),
	.w6(32'h3b2a4f83),
	.w7(32'hb9c36561),
	.w8(32'hb9ddeb1d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd46faa),
	.w1(32'hbaa2d337),
	.w2(32'hbbb081ce),
	.w3(32'h3b9c147e),
	.w4(32'h3b053f9b),
	.w5(32'hbb6132e9),
	.w6(32'h3b163fc4),
	.w7(32'h37c443b6),
	.w8(32'h3b8d7b2c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2958ce),
	.w1(32'hbb951b1f),
	.w2(32'hba389524),
	.w3(32'hbbc2e219),
	.w4(32'hbb3ec7d8),
	.w5(32'hbb88d06a),
	.w6(32'h3b261110),
	.w7(32'hbbfe1082),
	.w8(32'hbb397e68),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b959acf),
	.w1(32'h3bf48331),
	.w2(32'h3c212598),
	.w3(32'hb98f43a4),
	.w4(32'h3c4e7f3d),
	.w5(32'h3ca3e20c),
	.w6(32'h3b0d73e6),
	.w7(32'h3b8cdcf6),
	.w8(32'h3bf8cdd1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bef2e),
	.w1(32'hbb160261),
	.w2(32'hba2bc69a),
	.w3(32'h3c359336),
	.w4(32'h3b9e272e),
	.w5(32'h3a202495),
	.w6(32'h3c30fb1a),
	.w7(32'h3ba807df),
	.w8(32'h3b548905),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2554f9),
	.w1(32'h3b720822),
	.w2(32'hbbcee1a7),
	.w3(32'hba9caa4b),
	.w4(32'h3baf6fbb),
	.w5(32'h38adf7ee),
	.w6(32'h3af34cc8),
	.w7(32'h397e0cec),
	.w8(32'h3b05bc79),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76de67),
	.w1(32'h3bbae2e2),
	.w2(32'h3b9e9b14),
	.w3(32'hbba39e23),
	.w4(32'h3b4cb47d),
	.w5(32'h3b45eadc),
	.w6(32'hbb1078ab),
	.w7(32'h3ac3032b),
	.w8(32'h3b7ae136),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6f42),
	.w1(32'hbac0bb3b),
	.w2(32'h3a969fe3),
	.w3(32'hb9a6e14d),
	.w4(32'hbaa420b3),
	.w5(32'h3c1f3bdf),
	.w6(32'h3b954fe9),
	.w7(32'hbaee79b1),
	.w8(32'hba19933d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14cab0),
	.w1(32'hbb1dab9f),
	.w2(32'hbb18a12e),
	.w3(32'h3b4c2800),
	.w4(32'h3b4b17ee),
	.w5(32'hbbebf439),
	.w6(32'h3ab9d04c),
	.w7(32'h3b24a18f),
	.w8(32'hbb562859),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af33a99),
	.w1(32'h3a2190a8),
	.w2(32'hbb89b239),
	.w3(32'hbb6973b3),
	.w4(32'h3b9e494d),
	.w5(32'hb9cda0c8),
	.w6(32'hbbe57b71),
	.w7(32'h3bca6b86),
	.w8(32'hbabba4f4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b1250),
	.w1(32'h3bd7bb34),
	.w2(32'h390b68a9),
	.w3(32'h3c0d3661),
	.w4(32'h3b8e23a1),
	.w5(32'h3a5cae05),
	.w6(32'h3b64d080),
	.w7(32'h3b42ed6c),
	.w8(32'h3b08f4f7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70f6c8),
	.w1(32'hbbe0320f),
	.w2(32'hbb916878),
	.w3(32'hbb1d89d0),
	.w4(32'hbb96dcaa),
	.w5(32'h39cf2941),
	.w6(32'h3abe67e0),
	.w7(32'h39fbd437),
	.w8(32'h3afc6c62),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e76b6c),
	.w1(32'hbaa44c8a),
	.w2(32'hbb1cfa3a),
	.w3(32'h3a916fa9),
	.w4(32'h3a24b193),
	.w5(32'hbaaa948d),
	.w6(32'hb93a5608),
	.w7(32'hba17bb60),
	.w8(32'hb9b75ae2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba750ea6),
	.w1(32'h38f7fc9f),
	.w2(32'hb9a0771e),
	.w3(32'h39a0e003),
	.w4(32'hb93b878e),
	.w5(32'h37c75a49),
	.w6(32'hb911683d),
	.w7(32'hb88a2303),
	.w8(32'h38be5bb1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62713b),
	.w1(32'hba8b5b5a),
	.w2(32'hbaa27fea),
	.w3(32'h3ac74ad9),
	.w4(32'h38840924),
	.w5(32'hb9aa179d),
	.w6(32'h3b053cf8),
	.w7(32'hb9ec9feb),
	.w8(32'h39916357),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cf523),
	.w1(32'h3ab708ef),
	.w2(32'h3b1861c2),
	.w3(32'hb9c591b8),
	.w4(32'h393b28ce),
	.w5(32'h3af687e8),
	.w6(32'h39e52962),
	.w7(32'h3ad9a96e),
	.w8(32'h3b1b0f48),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a383227),
	.w1(32'h39795f28),
	.w2(32'h3a727d76),
	.w3(32'h37b3cad9),
	.w4(32'h3ab2558e),
	.w5(32'h3a7a1630),
	.w6(32'h39aba027),
	.w7(32'h3a0e6d7f),
	.w8(32'h3ac7878c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b790ad1),
	.w1(32'h3bc44ad8),
	.w2(32'h3b840d70),
	.w3(32'h3bc26462),
	.w4(32'h3bb99a07),
	.w5(32'h3b1b1574),
	.w6(32'h3bd5308e),
	.w7(32'h3b78a97e),
	.w8(32'h3b1eab26),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba45df7),
	.w1(32'h3bab7cf9),
	.w2(32'h3bcac995),
	.w3(32'h3bebcdf9),
	.w4(32'h3bffa626),
	.w5(32'h3b91cace),
	.w6(32'h3c2e3d4a),
	.w7(32'h3bac9a9b),
	.w8(32'h3b931304),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39eda8),
	.w1(32'hbb7bc5c4),
	.w2(32'hba6c99fb),
	.w3(32'hbb994184),
	.w4(32'hbb9cae60),
	.w5(32'hbb142f9e),
	.w6(32'hbb2bd639),
	.w7(32'hbaa81bf8),
	.w8(32'hbae808a7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a45c),
	.w1(32'h3af76883),
	.w2(32'h3a0c67e8),
	.w3(32'h3b1dcf0e),
	.w4(32'h3ac27c60),
	.w5(32'hba60440c),
	.w6(32'h3b3fa70e),
	.w7(32'h3a988085),
	.w8(32'h38d77086),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083e9d),
	.w1(32'hba891fb4),
	.w2(32'hbaf5d00c),
	.w3(32'hbb044df9),
	.w4(32'hba87f9d7),
	.w5(32'hba0c47e4),
	.w6(32'hb81eeb74),
	.w7(32'hba387f78),
	.w8(32'h381a9587),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaed41d),
	.w1(32'h3aefcd78),
	.w2(32'h3b3fad21),
	.w3(32'hbb01128c),
	.w4(32'h3af159c6),
	.w5(32'h3a9e71eb),
	.w6(32'hba69aaaf),
	.w7(32'h3b2c1fbd),
	.w8(32'h3b4a37b8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2990e),
	.w1(32'h3bcdc136),
	.w2(32'h3b933b11),
	.w3(32'h3bb89121),
	.w4(32'h3ba582d1),
	.w5(32'h3b2ba513),
	.w6(32'h3bdc2da6),
	.w7(32'h3b7f8c3d),
	.w8(32'h3ad7ff99),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8446455),
	.w1(32'h380991ed),
	.w2(32'h3a8ff072),
	.w3(32'hb90bc7d8),
	.w4(32'hb9b5d218),
	.w5(32'hb9c58db3),
	.w6(32'hba56dbb8),
	.w7(32'hba968ca6),
	.w8(32'hb90f3c6a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa27651),
	.w1(32'h3a335baf),
	.w2(32'h393030f5),
	.w3(32'h392f219d),
	.w4(32'h3ae239c0),
	.w5(32'h398aa1fd),
	.w6(32'h3ab270f9),
	.w7(32'h3abfc28f),
	.w8(32'h3a32380e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f206f),
	.w1(32'h39d4fb0d),
	.w2(32'hb96ee14a),
	.w3(32'h3a00b207),
	.w4(32'h3a90a1eb),
	.w5(32'hbab96a8f),
	.w6(32'hbaa24ae9),
	.w7(32'h3a3a1d21),
	.w8(32'h3a9eedfa),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc22c1),
	.w1(32'hbb1e8558),
	.w2(32'hba00517d),
	.w3(32'h3aed32c3),
	.w4(32'hba3fc24b),
	.w5(32'hb807d972),
	.w6(32'h3a6f261d),
	.w7(32'hba6eea40),
	.w8(32'hbac37343),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15a385),
	.w1(32'hba64433e),
	.w2(32'hbb51e3ad),
	.w3(32'hbb9b03f4),
	.w4(32'hb9b09951),
	.w5(32'hba823130),
	.w6(32'hbb191d4c),
	.w7(32'h3b38a4e0),
	.w8(32'h3a8b0350),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e7e3b),
	.w1(32'h39c3991d),
	.w2(32'h3998b4fe),
	.w3(32'h3a74e414),
	.w4(32'h39375844),
	.w5(32'h3af1fc52),
	.w6(32'h3a8f5b54),
	.w7(32'h3a86eaa3),
	.w8(32'hb9bf4874),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3653b),
	.w1(32'hba894bf0),
	.w2(32'hbaed54d6),
	.w3(32'h3a79364d),
	.w4(32'h38548f9c),
	.w5(32'hb9e77010),
	.w6(32'h3b67abb4),
	.w7(32'h3a26fd43),
	.w8(32'hba9f5542),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf12654),
	.w1(32'h3c19e03a),
	.w2(32'h3c103be7),
	.w3(32'h3c248dbc),
	.w4(32'h3bd339d5),
	.w5(32'h3bcde30b),
	.w6(32'h3c3ba8b7),
	.w7(32'h3bfa356a),
	.w8(32'h3bd12d35),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf500a5),
	.w1(32'hbb04defc),
	.w2(32'hbb0c6644),
	.w3(32'hbb4f0836),
	.w4(32'hbb1909af),
	.w5(32'hbae14f43),
	.w6(32'hbac831bb),
	.w7(32'hba0cc49e),
	.w8(32'hba7488e7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21210c),
	.w1(32'hba742d37),
	.w2(32'hbb49d7f0),
	.w3(32'h3b618902),
	.w4(32'hbadc29a7),
	.w5(32'hbb4751e3),
	.w6(32'h3b2007ab),
	.w7(32'hb9e0b1fc),
	.w8(32'hba90eb18),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27dd86),
	.w1(32'hbaa7930a),
	.w2(32'hba7791b6),
	.w3(32'hbb7fe248),
	.w4(32'hba60694c),
	.w5(32'h39e93848),
	.w6(32'hbb5adc9d),
	.w7(32'hbaf1197b),
	.w8(32'hb95ae67b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3cc9e),
	.w1(32'h3aa43ebc),
	.w2(32'h3aa660c5),
	.w3(32'h3a26a1d0),
	.w4(32'h388c20b0),
	.w5(32'hb91e8b1c),
	.w6(32'h3aa1c2f6),
	.w7(32'h3aeed032),
	.w8(32'h3b502b29),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855632),
	.w1(32'hbafd77bf),
	.w2(32'hbb3a930a),
	.w3(32'h38234251),
	.w4(32'hbb15bb81),
	.w5(32'hbb33c85e),
	.w6(32'h39a7c965),
	.w7(32'hbaf2ee25),
	.w8(32'hba1411da),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf1218),
	.w1(32'hba9ebffd),
	.w2(32'h3a7906e9),
	.w3(32'hbb7dc1e9),
	.w4(32'hbb1905e5),
	.w5(32'hbad7e6d4),
	.w6(32'hbb089853),
	.w7(32'h39dbe832),
	.w8(32'h3b09d1db),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39777ca4),
	.w1(32'h3a45f2dc),
	.w2(32'h3a0364c8),
	.w3(32'hbab6aecb),
	.w4(32'hb9ede059),
	.w5(32'hbb24adb1),
	.w6(32'hbafdbfb6),
	.w7(32'hba021a8c),
	.w8(32'hbac1f85f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02cf45),
	.w1(32'hbb0af4e0),
	.w2(32'hba913559),
	.w3(32'h3ab3edef),
	.w4(32'hbaaf837b),
	.w5(32'hba99b0d1),
	.w6(32'h3ac97b7d),
	.w7(32'hba89f8cc),
	.w8(32'h3a05f59c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c60d1d),
	.w1(32'hbb2114fc),
	.w2(32'hbb2b8e63),
	.w3(32'hbadfb1b2),
	.w4(32'hba50ef1f),
	.w5(32'hb95a8977),
	.w6(32'hba9cf2d5),
	.w7(32'hb89a0229),
	.w8(32'hba42bff1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b263b58),
	.w1(32'h3c1a2939),
	.w2(32'h3be4cf50),
	.w3(32'h3c0e57dc),
	.w4(32'h3be2aa56),
	.w5(32'h3b05a7a4),
	.w6(32'h3c107f48),
	.w7(32'h3bbcdd7b),
	.w8(32'hbabf9615),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85c3b7),
	.w1(32'hbb65f366),
	.w2(32'hbb2275ce),
	.w3(32'hbbb85f6d),
	.w4(32'hbb26c8f2),
	.w5(32'hb9c3e67c),
	.w6(32'hbb765214),
	.w7(32'hbb10d79b),
	.w8(32'hbab21c64),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43e3c1),
	.w1(32'hbb1f832f),
	.w2(32'hbb362a7b),
	.w3(32'hbb6a5b1f),
	.w4(32'hbaa6cc4c),
	.w5(32'hbb65c973),
	.w6(32'hbb187977),
	.w7(32'h3aa1f9a1),
	.w8(32'h3af5448e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d35a1),
	.w1(32'h3b454a8e),
	.w2(32'h3a4d0ae0),
	.w3(32'h3b4725fa),
	.w4(32'h3a147309),
	.w5(32'hb9fa0edd),
	.w6(32'h3b9142dc),
	.w7(32'h39e77c83),
	.w8(32'hbae77ae8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dd2f9),
	.w1(32'hba27aa52),
	.w2(32'hb9fc12fd),
	.w3(32'h3904f22c),
	.w4(32'hba208063),
	.w5(32'hbb7d6c89),
	.w6(32'hb9b9893d),
	.w7(32'hba382c9d),
	.w8(32'hba954851),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff1de4),
	.w1(32'h3c819f2c),
	.w2(32'h3c8292f3),
	.w3(32'h3c3e8a00),
	.w4(32'h3c57636d),
	.w5(32'h3bf017b7),
	.w6(32'h3c64a801),
	.w7(32'h3c366f11),
	.w8(32'h3be829f2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a402518),
	.w1(32'hb990c7c5),
	.w2(32'hbaa4e6a0),
	.w3(32'hbace1191),
	.w4(32'h393d6296),
	.w5(32'hb77850fc),
	.w6(32'h3a16cec5),
	.w7(32'hbaa02010),
	.w8(32'hbb117f3b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90da170),
	.w1(32'hb9095f3b),
	.w2(32'h39944cd2),
	.w3(32'hb9df50cd),
	.w4(32'h3874b506),
	.w5(32'hb996d25e),
	.w6(32'hbae6f9ef),
	.w7(32'h39627cc8),
	.w8(32'h38df6aee),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34bc1),
	.w1(32'hb975305e),
	.w2(32'hb92192d9),
	.w3(32'h3a79df87),
	.w4(32'h39fcb300),
	.w5(32'hba4cb14c),
	.w6(32'h3ad394e2),
	.w7(32'h38f42ef5),
	.w8(32'hb94a5064),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8a3a),
	.w1(32'h3a0ecbdc),
	.w2(32'h3910aecb),
	.w3(32'hb94827bb),
	.w4(32'h37f1048e),
	.w5(32'hbb0a2773),
	.w6(32'hb9b2d0f2),
	.w7(32'h3b32aa75),
	.w8(32'h3b0293fe),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a660cbb),
	.w1(32'hbb642291),
	.w2(32'hbaae3c7f),
	.w3(32'hbb08665c),
	.w4(32'hbb22bd00),
	.w5(32'hbb1e7216),
	.w6(32'hb9bbda4f),
	.w7(32'hbabf3f85),
	.w8(32'h3a2fe8fd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981b6f2),
	.w1(32'hba73abc4),
	.w2(32'h3b5b1dc4),
	.w3(32'hba7a0c49),
	.w4(32'h39a960a3),
	.w5(32'h3b115b9a),
	.w6(32'h384f8134),
	.w7(32'hb97dfe03),
	.w8(32'h396ece59),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d9c81),
	.w1(32'hbadcdc59),
	.w2(32'hba84c7b9),
	.w3(32'hb9592a9d),
	.w4(32'hbaaafd73),
	.w5(32'h3a01878f),
	.w6(32'hbabe5a27),
	.w7(32'h39ef9ef9),
	.w8(32'h39d23e27),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ba8ad),
	.w1(32'hba1cc6fb),
	.w2(32'h3a01e03d),
	.w3(32'h3a88bb0e),
	.w4(32'hba71d10b),
	.w5(32'hbacf72df),
	.w6(32'h3a3bf84d),
	.w7(32'h3a17939e),
	.w8(32'h3ad12efe),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39518a),
	.w1(32'h39108796),
	.w2(32'hbb02e618),
	.w3(32'h3b8892a7),
	.w4(32'h3a3f673a),
	.w5(32'hbb5885cd),
	.w6(32'h3bad58d2),
	.w7(32'hb98623e2),
	.w8(32'h3abf68b0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7fc9f),
	.w1(32'hb9824ef8),
	.w2(32'h3913fd35),
	.w3(32'hbba5f986),
	.w4(32'hba8a94c5),
	.w5(32'hb99e4121),
	.w6(32'hbb45ef98),
	.w7(32'hba7fcc21),
	.w8(32'hba167f15),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d25fd),
	.w1(32'hba9224b8),
	.w2(32'hbad1e14b),
	.w3(32'hb9726a74),
	.w4(32'hb9a6c10c),
	.w5(32'h3992654b),
	.w6(32'h39bab0f8),
	.w7(32'hba6a9246),
	.w8(32'hba8b5161),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c60d9),
	.w1(32'h39f9e8f1),
	.w2(32'h3a7665cf),
	.w3(32'hb9dfa966),
	.w4(32'h3a841ea6),
	.w5(32'h38b576fa),
	.w6(32'hba6c1e93),
	.w7(32'h3a9ef267),
	.w8(32'h3aa795a4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87a02f),
	.w1(32'h39a45f7c),
	.w2(32'hb892986e),
	.w3(32'h3abaf078),
	.w4(32'hba8b352c),
	.w5(32'h3a61acd6),
	.w6(32'h3a361902),
	.w7(32'hba19d03e),
	.w8(32'h3999e95d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe8768),
	.w1(32'h3afe2cc5),
	.w2(32'h3b261eca),
	.w3(32'hba228479),
	.w4(32'hb8f09dba),
	.w5(32'h3a9b8c86),
	.w6(32'hb9c0a13f),
	.w7(32'h3af2b809),
	.w8(32'h3af872c9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a3203),
	.w1(32'hbb87c21d),
	.w2(32'hbb2411cb),
	.w3(32'hbb5b98a8),
	.w4(32'hbb3e3159),
	.w5(32'hbb84d8bf),
	.w6(32'hb990d6c9),
	.w7(32'hbb3cc3a0),
	.w8(32'hbb1d7a41),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5342e),
	.w1(32'h38fe759a),
	.w2(32'hb983bd5f),
	.w3(32'h3b45524e),
	.w4(32'h39becc09),
	.w5(32'h39959999),
	.w6(32'h3ae547dc),
	.w7(32'h39c1e4c9),
	.w8(32'h3a14a19d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b4eb2),
	.w1(32'h3a3a39ed),
	.w2(32'h3967607c),
	.w3(32'h3b4bed89),
	.w4(32'h3b22fc2a),
	.w5(32'hb96c6719),
	.w6(32'h3b63fc6e),
	.w7(32'h3b235ba9),
	.w8(32'h3ab672e2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cde26),
	.w1(32'hbb70a6d9),
	.w2(32'hbb845d98),
	.w3(32'hbb72b976),
	.w4(32'hbae0f076),
	.w5(32'hbb08c248),
	.w6(32'hbb3d27a1),
	.w7(32'hba99007a),
	.w8(32'hba715493),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61cc4d),
	.w1(32'hb95f88f3),
	.w2(32'hba537bf7),
	.w3(32'hba054017),
	.w4(32'hb9841111),
	.w5(32'hba639f6e),
	.w6(32'hb9bd098f),
	.w7(32'hba92ecd6),
	.w8(32'hba5f7e52),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59aa6),
	.w1(32'h3a39b37f),
	.w2(32'hb7e9a775),
	.w3(32'hbae6a37d),
	.w4(32'h391d455e),
	.w5(32'h39ff4151),
	.w6(32'hbaffa6b2),
	.w7(32'h3a255ae2),
	.w8(32'h39f28563),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cad7d3),
	.w1(32'hba0aab7d),
	.w2(32'hb99f0899),
	.w3(32'h39ab9a50),
	.w4(32'hb931406d),
	.w5(32'hba95b850),
	.w6(32'h36a80923),
	.w7(32'hb8d89d8a),
	.w8(32'hba2e1070),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251f1e),
	.w1(32'hbb008c59),
	.w2(32'hbb375fe8),
	.w3(32'hbb7bf84f),
	.w4(32'h3978f1d5),
	.w5(32'h3ab1c512),
	.w6(32'hbb2d8c04),
	.w7(32'hba5f9123),
	.w8(32'hbb1156f8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd7c79),
	.w1(32'h38b98ce5),
	.w2(32'hba29aee9),
	.w3(32'hb8f97a83),
	.w4(32'h3aae5388),
	.w5(32'h3a6514ef),
	.w6(32'h38882773),
	.w7(32'h3b12078c),
	.w8(32'h3ab6d83a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac39dcb),
	.w1(32'h399aca48),
	.w2(32'hb802105c),
	.w3(32'hb88d1411),
	.w4(32'h3ae67885),
	.w5(32'h3b1a11e4),
	.w6(32'h3a012c83),
	.w7(32'h3b036755),
	.w8(32'h3a69bd4a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992c923),
	.w1(32'h3a15a570),
	.w2(32'h3aa099ff),
	.w3(32'h3a5e71d1),
	.w4(32'h3a0abf05),
	.w5(32'h39f31dea),
	.w6(32'h3a8d7647),
	.w7(32'hba1f5251),
	.w8(32'hb7abb259),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaeb9a2),
	.w1(32'hbaf8a827),
	.w2(32'h39f40588),
	.w3(32'h3a923f2d),
	.w4(32'hbb0a79c7),
	.w5(32'hb97e83f5),
	.w6(32'h3a54fc6d),
	.w7(32'hbab5246f),
	.w8(32'hba6e723a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a406bbc),
	.w1(32'h3ae22e8b),
	.w2(32'hb94cd9b5),
	.w3(32'hba7fe513),
	.w4(32'h3aec8535),
	.w5(32'hbb75e91f),
	.w6(32'hba64a3f9),
	.w7(32'h3ab67936),
	.w8(32'hb9daaa6d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d0f58),
	.w1(32'hba368e42),
	.w2(32'h3a0204d7),
	.w3(32'hb99a0baf),
	.w4(32'hba0cdc4c),
	.w5(32'h3a27bf23),
	.w6(32'h3a507143),
	.w7(32'h398d9860),
	.w8(32'h3abaf92b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce1b87),
	.w1(32'hbb1b04f1),
	.w2(32'hbb2d946b),
	.w3(32'hba28b3f2),
	.w4(32'hbadc3d75),
	.w5(32'hba5e0a1c),
	.w6(32'h38f20201),
	.w7(32'hbaae2a86),
	.w8(32'hba07dc9a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9898d3),
	.w1(32'h3bc6257f),
	.w2(32'h3bdb584a),
	.w3(32'h3bc3e3b7),
	.w4(32'h3b66e11d),
	.w5(32'h3b3de4bd),
	.w6(32'h3be28ab9),
	.w7(32'h3b9f3dbf),
	.w8(32'h3b4b22ec),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbd93f),
	.w1(32'hba91dade),
	.w2(32'hba82a67a),
	.w3(32'hbb0b5673),
	.w4(32'h390bc36d),
	.w5(32'h3a31f917),
	.w6(32'hbacd10a9),
	.w7(32'h3a5f3cce),
	.w8(32'h3a9ae09d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a253),
	.w1(32'hb9dd6295),
	.w2(32'h39546f0a),
	.w3(32'h3b00c157),
	.w4(32'h39cff8b2),
	.w5(32'hb99c4637),
	.w6(32'h3b285c3a),
	.w7(32'h3a9ff79d),
	.w8(32'h3b1118a6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba37c57),
	.w1(32'h3ba1c891),
	.w2(32'h3b592552),
	.w3(32'h3bea64ab),
	.w4(32'h3b59bbeb),
	.w5(32'h3a217719),
	.w6(32'h3bc4320f),
	.w7(32'h3addfe74),
	.w8(32'h39957288),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820a30),
	.w1(32'hba4a28c9),
	.w2(32'hbb5107a5),
	.w3(32'hba895930),
	.w4(32'h3b1c4770),
	.w5(32'hba9547f5),
	.w6(32'h3b0a8828),
	.w7(32'h3ab1b291),
	.w8(32'h3a811a85),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfbc3b),
	.w1(32'h3a0ace27),
	.w2(32'hb964e302),
	.w3(32'h3a6e5eaf),
	.w4(32'h3a30e5e3),
	.w5(32'h395ec979),
	.w6(32'h3aaab257),
	.w7(32'h38c81a8c),
	.w8(32'hb9ba8a1d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5756ae),
	.w1(32'h3a5dbe49),
	.w2(32'h3b12e028),
	.w3(32'h3a605dff),
	.w4(32'h3a64ed85),
	.w5(32'hb7cbd572),
	.w6(32'h39f0bc3a),
	.w7(32'h3aa6e74e),
	.w8(32'h3b25b154),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994c33b),
	.w1(32'hbb173514),
	.w2(32'h39b34fce),
	.w3(32'hbb64d5af),
	.w4(32'hbb56eedc),
	.w5(32'h39faa890),
	.w6(32'hbb067823),
	.w7(32'hba3edf31),
	.w8(32'h3ad658ba),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b833ab7),
	.w1(32'h3b15907e),
	.w2(32'h3a8813fa),
	.w3(32'h3b8444e4),
	.w4(32'h3b10b704),
	.w5(32'h3a36d536),
	.w6(32'h3b6f6817),
	.w7(32'h3afd64a6),
	.w8(32'h3abfa3b1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b3059),
	.w1(32'h3ac99a48),
	.w2(32'h3a568351),
	.w3(32'h3a37d580),
	.w4(32'h3ab066de),
	.w5(32'h3b1ac71d),
	.w6(32'hba680cd2),
	.w7(32'h3ad45ce5),
	.w8(32'h3ac85021),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd2a4f),
	.w1(32'hb9e78d3a),
	.w2(32'hbaca45db),
	.w3(32'h3b1058a3),
	.w4(32'h39a211c7),
	.w5(32'hb9d5c51f),
	.w6(32'h3af85c22),
	.w7(32'hb9aad9df),
	.w8(32'hba60dc8d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62cf6),
	.w1(32'hb6bc732c),
	.w2(32'hbaa2ea15),
	.w3(32'hbb1faca7),
	.w4(32'h39900cd2),
	.w5(32'hba4993b0),
	.w6(32'hbb0e5653),
	.w7(32'h3952846c),
	.w8(32'h39b2b61b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa75af4),
	.w1(32'hba1203b1),
	.w2(32'h3a80f1f8),
	.w3(32'hbb4b893c),
	.w4(32'h3985f735),
	.w5(32'hbaa6b3fa),
	.w6(32'hba70711b),
	.w7(32'h3a973242),
	.w8(32'h3aa9d648),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa43301),
	.w1(32'hba769f66),
	.w2(32'hbb1686e4),
	.w3(32'h3a299dfd),
	.w4(32'hb9f2bbb5),
	.w5(32'hba8c150d),
	.w6(32'h39c66b69),
	.w7(32'h3927431d),
	.w8(32'h38118728),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7557a0),
	.w1(32'hb94a0a55),
	.w2(32'hb9df725a),
	.w3(32'h3b0da2ac),
	.w4(32'hb9b81cf5),
	.w5(32'hba1cb25c),
	.w6(32'h39d44e2c),
	.w7(32'hb9f999d5),
	.w8(32'hba0c67cb),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d55785),
	.w1(32'hba6e619a),
	.w2(32'hb93e034a),
	.w3(32'hb8e80104),
	.w4(32'hbb0e7357),
	.w5(32'h3903c999),
	.w6(32'h39e9fe47),
	.w7(32'hbafe534a),
	.w8(32'h3b217e2d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26463c),
	.w1(32'hbacce7b3),
	.w2(32'hbaabd1df),
	.w3(32'hbb4f0f5c),
	.w4(32'hbb0c26eb),
	.w5(32'hb9a0ee49),
	.w6(32'hba7c0d97),
	.w7(32'hb9d845a6),
	.w8(32'hb916ec81),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a92eb),
	.w1(32'h3b837174),
	.w2(32'h3bb2a9fc),
	.w3(32'h3b4236c3),
	.w4(32'h39bec87a),
	.w5(32'h3acb61f7),
	.w6(32'h3b2d67f3),
	.w7(32'h3b066e4f),
	.w8(32'h3b289299),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb116a4a),
	.w1(32'h39ceec4e),
	.w2(32'h3ac57659),
	.w3(32'hbbd72f9c),
	.w4(32'hbb001ee6),
	.w5(32'h3ae5b9d3),
	.w6(32'hbba5b719),
	.w7(32'h3af790fa),
	.w8(32'h3b1cca08),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a618a90),
	.w1(32'hbb3f1a12),
	.w2(32'hba90f7f5),
	.w3(32'hba615615),
	.w4(32'hbaedce94),
	.w5(32'h3aed84e8),
	.w6(32'hbac7a7c3),
	.w7(32'hbafc3310),
	.w8(32'hbb1336da),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c52e),
	.w1(32'hbac54d5d),
	.w2(32'hbaca4be7),
	.w3(32'hbb3236b6),
	.w4(32'hbb2340df),
	.w5(32'hbb573a4a),
	.w6(32'hbb8e19e5),
	.w7(32'hbb0bacf2),
	.w8(32'hba73aeef),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3044f1),
	.w1(32'h39318d7b),
	.w2(32'h3a25a754),
	.w3(32'h3a03af5e),
	.w4(32'h3931ead9),
	.w5(32'h3a0316bb),
	.w6(32'hb89e1309),
	.w7(32'h3ab11318),
	.w8(32'h3b1f1484),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c97b3),
	.w1(32'hbaf4a926),
	.w2(32'hbb3ca2b4),
	.w3(32'hba58600b),
	.w4(32'hbb424284),
	.w5(32'hb9f55d9f),
	.w6(32'hb9249f97),
	.w7(32'hbb01cb4e),
	.w8(32'hbb19e87b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb311768),
	.w1(32'h396836a7),
	.w2(32'h3a201fd6),
	.w3(32'hbad2a8e2),
	.w4(32'hb907cd7f),
	.w5(32'h3a2caaa2),
	.w6(32'hbb62f2c0),
	.w7(32'hb821674e),
	.w8(32'hbab7ca09),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5d684),
	.w1(32'h3a2bd5c8),
	.w2(32'h386dc851),
	.w3(32'h3ac36cfc),
	.w4(32'h39cbdbda),
	.w5(32'h3a8a15c0),
	.w6(32'h3a38fde8),
	.w7(32'h3a43439a),
	.w8(32'hb9814c2e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f80dd),
	.w1(32'hba09836b),
	.w2(32'h3a319c6d),
	.w3(32'hbaa2b9e6),
	.w4(32'h3a15c123),
	.w5(32'hb7ff7fe7),
	.w6(32'hba8c9b5b),
	.w7(32'h3820893a),
	.w8(32'h396152e4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea86f7),
	.w1(32'hba264817),
	.w2(32'hba8d5392),
	.w3(32'h3b5184b8),
	.w4(32'hba0a61d1),
	.w5(32'h3927086d),
	.w6(32'h3b74ffee),
	.w7(32'h3a55a925),
	.w8(32'h3ad6ea38),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b302a),
	.w1(32'h3a1ac415),
	.w2(32'h3a378135),
	.w3(32'h3a2a22f8),
	.w4(32'hba350220),
	.w5(32'hb616908c),
	.w6(32'h3a399751),
	.w7(32'hb8eef817),
	.w8(32'hbb12d78d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83b03c),
	.w1(32'hbb2c57e4),
	.w2(32'hbadfde60),
	.w3(32'hba9386eb),
	.w4(32'hbb02c3c6),
	.w5(32'hb9604bfe),
	.w6(32'hbacbea1a),
	.w7(32'hbaf2577f),
	.w8(32'hba738463),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2c177),
	.w1(32'h38c2ca0e),
	.w2(32'hbabcdcfe),
	.w3(32'h3913423b),
	.w4(32'h38bb583d),
	.w5(32'hbaead923),
	.w6(32'h3a1fccf4),
	.w7(32'hba18550e),
	.w8(32'hba8ca081),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6def),
	.w1(32'h3a7b8e03),
	.w2(32'hb9fac265),
	.w3(32'hbb1bd925),
	.w4(32'h3a9358cf),
	.w5(32'hb82b6b9b),
	.w6(32'hba631873),
	.w7(32'h39647ece),
	.w8(32'h3aea7efe),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9334f),
	.w1(32'h3a88df9c),
	.w2(32'h3ab554a0),
	.w3(32'h3a804bb6),
	.w4(32'h3a053cfb),
	.w5(32'hba38733e),
	.w6(32'hb99aaba1),
	.w7(32'h3abf0ac4),
	.w8(32'h3a7dd119),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09839c),
	.w1(32'hba05ff96),
	.w2(32'h3a486050),
	.w3(32'h3b1d84b7),
	.w4(32'h3957cf2e),
	.w5(32'h38f474b5),
	.w6(32'h3b2b2012),
	.w7(32'h397eda65),
	.w8(32'h3a9f8fb1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88001e),
	.w1(32'h38007d2a),
	.w2(32'hbabb7c14),
	.w3(32'hba5be4aa),
	.w4(32'h3a064607),
	.w5(32'hbb39af03),
	.w6(32'hba9c04ac),
	.w7(32'h3aa117db),
	.w8(32'hbad6e95e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5ae38),
	.w1(32'h3b0f3ed9),
	.w2(32'h3b2700a4),
	.w3(32'h3b830f8e),
	.w4(32'h3af18d6d),
	.w5(32'h3a85a053),
	.w6(32'h3bd64e46),
	.w7(32'h3ad4b07c),
	.w8(32'h38126e86),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9086e9),
	.w1(32'hb89a8f73),
	.w2(32'hba22d3f7),
	.w3(32'hb9c76f09),
	.w4(32'hb9cc9378),
	.w5(32'hbb398392),
	.w6(32'hba9c706c),
	.w7(32'hba9feb68),
	.w8(32'hbab714af),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac127ac),
	.w1(32'hbb106305),
	.w2(32'hb9d61596),
	.w3(32'hbb235da1),
	.w4(32'hbb06cc7c),
	.w5(32'hbb42ac0e),
	.w6(32'hbb310cf9),
	.w7(32'hba94b977),
	.w8(32'hb9a2df4f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf1e6b),
	.w1(32'h3a81c042),
	.w2(32'h39c8f48d),
	.w3(32'hb9df6acd),
	.w4(32'h3afc74a6),
	.w5(32'h39d01076),
	.w6(32'hb977d396),
	.w7(32'h3a47b168),
	.w8(32'hba0064bc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01f941),
	.w1(32'hb9c9d392),
	.w2(32'h3a1c7797),
	.w3(32'h3ae6f977),
	.w4(32'hb8a97ae2),
	.w5(32'hba56276a),
	.w6(32'h3a784a0c),
	.w7(32'h3a820602),
	.w8(32'h3b1e204e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a078fb3),
	.w1(32'h3ad7cad5),
	.w2(32'hb96f2c16),
	.w3(32'h3a812d13),
	.w4(32'h3ae48327),
	.w5(32'h3b2cf670),
	.w6(32'h3b1bc943),
	.w7(32'h3b101b7e),
	.w8(32'h3b0ce939),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99976f),
	.w1(32'h3b97b2d6),
	.w2(32'h3b9fca01),
	.w3(32'h3be0f76d),
	.w4(32'h3b3e8044),
	.w5(32'h3b45b7f6),
	.w6(32'h3bc4c6ef),
	.w7(32'h3acac6fe),
	.w8(32'h3a7cbb96),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f37d9),
	.w1(32'hbad5c477),
	.w2(32'hba4951d4),
	.w3(32'h39e36d66),
	.w4(32'hbaa6634c),
	.w5(32'hb9f56c3c),
	.w6(32'h39184502),
	.w7(32'hbac082cc),
	.w8(32'hbaea0619),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24725f),
	.w1(32'h3b092755),
	.w2(32'h3addf9af),
	.w3(32'h3a33a587),
	.w4(32'h3b20dcca),
	.w5(32'h3a5a2347),
	.w6(32'h3a07929d),
	.w7(32'h3aaaa32c),
	.w8(32'h3ae100ca),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957b461),
	.w1(32'h39873ccf),
	.w2(32'h3992fc79),
	.w3(32'h3921081d),
	.w4(32'hb7f7e85a),
	.w5(32'hbad0c3e9),
	.w6(32'h36a0dafb),
	.w7(32'hbac4d8f6),
	.w8(32'hbacf5e73),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a973831),
	.w1(32'hbaa11314),
	.w2(32'h39844a77),
	.w3(32'h38824d56),
	.w4(32'hbb0ab5de),
	.w5(32'h3abcc90e),
	.w6(32'h3a964770),
	.w7(32'hbb083fc0),
	.w8(32'hb9d0443e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5314fd),
	.w1(32'hbae0d58c),
	.w2(32'hba36a07d),
	.w3(32'h3a0f7cbf),
	.w4(32'hba8e233c),
	.w5(32'h39c51b46),
	.w6(32'h3a59a28c),
	.w7(32'hbab46ec0),
	.w8(32'h3b251de2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f4099),
	.w1(32'hba11ef97),
	.w2(32'hba1969df),
	.w3(32'hbae4f778),
	.w4(32'hba8ef276),
	.w5(32'hb8a58e57),
	.w6(32'h3a399d24),
	.w7(32'h3ad18d7a),
	.w8(32'h3a3a849a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef5847),
	.w1(32'hba0385e4),
	.w2(32'h383cff2e),
	.w3(32'hbaa697dd),
	.w4(32'h3a5b27a3),
	.w5(32'h3acb426f),
	.w6(32'hb9d5e795),
	.w7(32'h3a94f7eb),
	.w8(32'hb64260eb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c1081),
	.w1(32'hba0d39f3),
	.w2(32'hba8f414c),
	.w3(32'h37805d49),
	.w4(32'h394debcd),
	.w5(32'hbad44913),
	.w6(32'h396076df),
	.w7(32'h3a310245),
	.w8(32'hba185810),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15ba95),
	.w1(32'h3a7950ce),
	.w2(32'h39cb7e9b),
	.w3(32'hba97d62b),
	.w4(32'hba058121),
	.w5(32'hbb78e745),
	.w6(32'h3a097d32),
	.w7(32'h3abf2ee0),
	.w8(32'h3a07e974),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97aec1b),
	.w1(32'h3b1bbc62),
	.w2(32'h3b00e1db),
	.w3(32'hbb3f1fcb),
	.w4(32'h3b0f3c07),
	.w5(32'h3b70ce4d),
	.w6(32'hb9281467),
	.w7(32'h3b16efa6),
	.w8(32'h3af194d3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb86f),
	.w1(32'hb93cdee4),
	.w2(32'hbacbd09f),
	.w3(32'h3b1c679a),
	.w4(32'h39bd61df),
	.w5(32'hba48f6f4),
	.w6(32'h3b07bf61),
	.w7(32'hba2a9939),
	.w8(32'h3a21caee),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa752ef),
	.w1(32'hb9ff252a),
	.w2(32'h3653d8d4),
	.w3(32'h3aaebd9d),
	.w4(32'hba79658b),
	.w5(32'h3ae7ab7e),
	.w6(32'h39d4106e),
	.w7(32'hb9e68314),
	.w8(32'h3a0f3d35),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39f8f8),
	.w1(32'h3b9e2d78),
	.w2(32'h3ad68618),
	.w3(32'h3aa760e7),
	.w4(32'h3b09d324),
	.w5(32'h3aa210fa),
	.w6(32'h3b023a4c),
	.w7(32'h3b0762ba),
	.w8(32'hbaa7ec04),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf721b9),
	.w1(32'hbbeea75d),
	.w2(32'hbba1ef6a),
	.w3(32'hbb918995),
	.w4(32'hbbcad268),
	.w5(32'hbab17a2f),
	.w6(32'hbb61eb47),
	.w7(32'hbad418c3),
	.w8(32'h39df5ed0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeda68b),
	.w1(32'h3a68b9f0),
	.w2(32'h3a585501),
	.w3(32'hbafc449c),
	.w4(32'h3ae69a97),
	.w5(32'hbadb92f5),
	.w6(32'hbac8bd6c),
	.w7(32'h3aa12018),
	.w8(32'h3aa52222),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ab3d3),
	.w1(32'hb992e42e),
	.w2(32'hba136e3e),
	.w3(32'h3b585505),
	.w4(32'hbad96177),
	.w5(32'hbb1e2c93),
	.w6(32'h3af516f5),
	.w7(32'hba1d32ab),
	.w8(32'h39bfb559),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e735f9),
	.w1(32'hb9b0003a),
	.w2(32'h3aab3d74),
	.w3(32'hb9195761),
	.w4(32'h3a0914f3),
	.w5(32'h3b340cff),
	.w6(32'h3a5e7c88),
	.w7(32'h37f85fda),
	.w8(32'hb9f3be0f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a07279),
	.w1(32'h3b4b4b55),
	.w2(32'h3b424a5a),
	.w3(32'hb9e9761f),
	.w4(32'h3b1c5a07),
	.w5(32'h39ae6328),
	.w6(32'hba85e0bc),
	.w7(32'h3b2bd187),
	.w8(32'h3b120545),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d979e),
	.w1(32'h3a693846),
	.w2(32'h3ad550ba),
	.w3(32'h3ac4d3e7),
	.w4(32'h39d28224),
	.w5(32'hba532429),
	.w6(32'h3b472711),
	.w7(32'h3a3e7283),
	.w8(32'h3a5d0540),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab244f0),
	.w1(32'h3ad062b1),
	.w2(32'h3ac4de8a),
	.w3(32'h3a270f8c),
	.w4(32'h3b30efe9),
	.w5(32'h3b13dd82),
	.w6(32'h3a672514),
	.w7(32'h3b148013),
	.w8(32'h3a80298f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57ba26),
	.w1(32'h39a74dda),
	.w2(32'hbb3bd63c),
	.w3(32'hba2aefcf),
	.w4(32'h39a6975a),
	.w5(32'hbab962db),
	.w6(32'hba9136bb),
	.w7(32'h3b46052a),
	.w8(32'h3a5065f1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad159f9),
	.w1(32'hb956d764),
	.w2(32'hbaf0f827),
	.w3(32'h3b0717fa),
	.w4(32'h3aaae5fe),
	.w5(32'hb8b8bc58),
	.w6(32'h3826df11),
	.w7(32'h39e578ab),
	.w8(32'hb9d1795c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc5216),
	.w1(32'hbb0ffd01),
	.w2(32'hbc123501),
	.w3(32'hbb06b3f5),
	.w4(32'h3ae5462f),
	.w5(32'hbb95711f),
	.w6(32'h3a70e8d2),
	.w7(32'h3bef5bb1),
	.w8(32'h3a24f347),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffa9d7),
	.w1(32'hbb7ca828),
	.w2(32'hbb580569),
	.w3(32'hbb86cf90),
	.w4(32'hbbc6a3b0),
	.w5(32'hbc28364c),
	.w6(32'hb9fa1936),
	.w7(32'hbb65ecbb),
	.w8(32'h3a6e27b5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60a6fd),
	.w1(32'hbb354d62),
	.w2(32'h3af1c67a),
	.w3(32'hba1808fd),
	.w4(32'h3882b78a),
	.w5(32'hbbbcf12c),
	.w6(32'h3c02dced),
	.w7(32'hbb4eb7f6),
	.w8(32'hbb904c25),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1b0dc),
	.w1(32'h3b2e008a),
	.w2(32'hbb77dad3),
	.w3(32'hbc2dd668),
	.w4(32'h3b8a9187),
	.w5(32'hbb454d3c),
	.w6(32'hbadfc413),
	.w7(32'h3c33e128),
	.w8(32'h3b2766e0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5337a),
	.w1(32'h3a01313a),
	.w2(32'h3a818a8b),
	.w3(32'hbbbf37db),
	.w4(32'h3a358147),
	.w5(32'h3a278204),
	.w6(32'hbb1e47da),
	.w7(32'hba883539),
	.w8(32'hba9883d3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2788a1),
	.w1(32'h398c9903),
	.w2(32'h3c00bdab),
	.w3(32'h3789dfe6),
	.w4(32'h3a23f625),
	.w5(32'h3c50881b),
	.w6(32'h3bbd381a),
	.w7(32'h3a04ffd4),
	.w8(32'h3b3075be),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4efcf),
	.w1(32'hbb267f79),
	.w2(32'h3b1805a5),
	.w3(32'h3b2c526b),
	.w4(32'h3b0f3f1e),
	.w5(32'h3c117728),
	.w6(32'hbb79ba35),
	.w7(32'hb93854cb),
	.w8(32'h3b0c3e5e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea92a7),
	.w1(32'hbb58c405),
	.w2(32'hbba97c1e),
	.w3(32'hba0f3e67),
	.w4(32'h3a8d56a1),
	.w5(32'hba82f3c6),
	.w6(32'hbb0f1599),
	.w7(32'hbb175aa6),
	.w8(32'hbada08e1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318044),
	.w1(32'hba2c5c20),
	.w2(32'hb880f920),
	.w3(32'hbb23c7ef),
	.w4(32'h3acd23d3),
	.w5(32'hbba4ee64),
	.w6(32'hba3de4be),
	.w7(32'hbb9329ce),
	.w8(32'h3ba3dcbb),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0987b),
	.w1(32'hbb058989),
	.w2(32'h3bc235e2),
	.w3(32'hbbc160c5),
	.w4(32'h3b20ce56),
	.w5(32'h3b74ebb4),
	.w6(32'hbb5ca8a2),
	.w7(32'hbb48b728),
	.w8(32'h39eb08b4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b126422),
	.w1(32'hba5ed880),
	.w2(32'hbb881362),
	.w3(32'h3b2dfbf1),
	.w4(32'hbb01eac3),
	.w5(32'hbb0902c4),
	.w6(32'hbb0a924d),
	.w7(32'hb96a7f9a),
	.w8(32'h39c6318d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfcb6b),
	.w1(32'h3aabda8e),
	.w2(32'h3c3bdb0b),
	.w3(32'hbbb3eb53),
	.w4(32'h3a1a54a0),
	.w5(32'h3a244534),
	.w6(32'h3a8a3feb),
	.w7(32'hbb943df6),
	.w8(32'hbb9988fc),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b1ca7),
	.w1(32'h3bb81c48),
	.w2(32'h3b52ce65),
	.w3(32'h3b45e86f),
	.w4(32'h3a9f1fba),
	.w5(32'hb9ae7eab),
	.w6(32'hbb6c2182),
	.w7(32'hba8a1d6e),
	.w8(32'hbb2ecc1f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80cd0c),
	.w1(32'h388f9979),
	.w2(32'h3b1eaabf),
	.w3(32'h3a70f96f),
	.w4(32'h3ad78baf),
	.w5(32'h3c0a7c93),
	.w6(32'hbb1729a9),
	.w7(32'hbac47c88),
	.w8(32'h3896df09),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7abadc),
	.w1(32'h3ba769ce),
	.w2(32'hb967a46d),
	.w3(32'hbaaee3e7),
	.w4(32'h3b9540a3),
	.w5(32'h3ae49b69),
	.w6(32'h3a756bec),
	.w7(32'hba3f555e),
	.w8(32'h3c24cea7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33365f),
	.w1(32'h3b6143f1),
	.w2(32'h3ac7c71c),
	.w3(32'h3c0ede6c),
	.w4(32'hbace2d62),
	.w5(32'h39611b18),
	.w6(32'h3bfa84fe),
	.w7(32'h3b69bb17),
	.w8(32'h3ab0805d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d658e),
	.w1(32'hbbc1ddfe),
	.w2(32'hbc10cb46),
	.w3(32'hbaf17436),
	.w4(32'hbc80648e),
	.w5(32'h3d141b2d),
	.w6(32'h3b8c0633),
	.w7(32'h3c54644d),
	.w8(32'h3cdd9991),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381cacc9),
	.w1(32'hbb555f32),
	.w2(32'hba30f7b1),
	.w3(32'h3b142635),
	.w4(32'hbba60a2d),
	.w5(32'hbbed6f35),
	.w6(32'hbbeab383),
	.w7(32'h3a5f3c0d),
	.w8(32'h3bc21919),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5cff5),
	.w1(32'hbb94bb5f),
	.w2(32'hbba4616f),
	.w3(32'h3b0fd5c8),
	.w4(32'h3ba46d40),
	.w5(32'h3be2d874),
	.w6(32'h3b1c3a2c),
	.w7(32'hbb3b8849),
	.w8(32'hbabe3dd5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa72fd),
	.w1(32'h3a70d9a6),
	.w2(32'hbb18ca5b),
	.w3(32'h3ba73d36),
	.w4(32'h3bad9bd8),
	.w5(32'hbadf89bd),
	.w6(32'h3b11545b),
	.w7(32'hbbab8ae4),
	.w8(32'h3baeb431),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba565dea),
	.w1(32'h3b862bcd),
	.w2(32'h3ba6baa5),
	.w3(32'h3b75b7bc),
	.w4(32'h3b7dc95b),
	.w5(32'hbb005d1d),
	.w6(32'h3bb36936),
	.w7(32'h3c10c7d3),
	.w8(32'hba4dbecc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c076709),
	.w1(32'h3b818cc6),
	.w2(32'h3ac6110a),
	.w3(32'h3b6a8b78),
	.w4(32'h3c00dd41),
	.w5(32'hbb58f4e4),
	.w6(32'hbb053128),
	.w7(32'h3ba392d2),
	.w8(32'hbaa08f85),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b790578),
	.w1(32'h3b42fed8),
	.w2(32'h3b0a6048),
	.w3(32'h3c3c8933),
	.w4(32'h3caeb0df),
	.w5(32'h3cec1337),
	.w6(32'h3c88e0a6),
	.w7(32'h3c068839),
	.w8(32'h3bbbbc81),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2163a),
	.w1(32'h3a6dad9e),
	.w2(32'h3b721c56),
	.w3(32'h3c73a0ae),
	.w4(32'h3ae74dc5),
	.w5(32'h3c081575),
	.w6(32'hbb39c8bf),
	.w7(32'h3a8becb6),
	.w8(32'h3ba5e240),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38635e),
	.w1(32'hbae89700),
	.w2(32'hb96c9993),
	.w3(32'h39e771b3),
	.w4(32'h3ae9db30),
	.w5(32'h3a30dbe7),
	.w6(32'h3b26c7bd),
	.w7(32'h3bb8cc18),
	.w8(32'h3b99609c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8971ec),
	.w1(32'h3b45c6bf),
	.w2(32'h3a2b6b64),
	.w3(32'h3b4b1e3d),
	.w4(32'h3b0400f6),
	.w5(32'h3c05618f),
	.w6(32'h3bbbc5cc),
	.w7(32'h38b5d36e),
	.w8(32'h3c14a7ed),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e3b5b),
	.w1(32'h39bca6f7),
	.w2(32'h3aa7b9b9),
	.w3(32'hbb0bb36c),
	.w4(32'h3bb65e6c),
	.w5(32'hbb391e06),
	.w6(32'hbbaa946b),
	.w7(32'hba9bb538),
	.w8(32'hbb9c4d3e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bcfe7),
	.w1(32'hbaf45586),
	.w2(32'hbbdc9393),
	.w3(32'hbbf779f2),
	.w4(32'hbbb3c224),
	.w5(32'hb9c899ae),
	.w6(32'hb9f52b0a),
	.w7(32'h38962a79),
	.w8(32'h3a6c494f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0264e0),
	.w1(32'h3b2d1b1c),
	.w2(32'hbaafd3f8),
	.w3(32'hbb2cf75a),
	.w4(32'hba29e13b),
	.w5(32'h3a82ccbb),
	.w6(32'hbbbaccc4),
	.w7(32'h3c146728),
	.w8(32'h3ba2e3cc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7337f5),
	.w1(32'h3ba9a708),
	.w2(32'h3b2828c3),
	.w3(32'h3ae5083d),
	.w4(32'h3c43a2e1),
	.w5(32'hbab72dfd),
	.w6(32'hbb8e955d),
	.w7(32'h3c80a022),
	.w8(32'h3bb96039),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ce9b9),
	.w1(32'hbb32d886),
	.w2(32'h3bab9237),
	.w3(32'h3bff1440),
	.w4(32'hb8007a1e),
	.w5(32'hbb862e59),
	.w6(32'h3c0ca4b4),
	.w7(32'hba74fe42),
	.w8(32'hbb8d21e0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb160c45),
	.w1(32'h3b255683),
	.w2(32'h3b8b8a97),
	.w3(32'hb9142ffe),
	.w4(32'h3a467d11),
	.w5(32'h3951b7a4),
	.w6(32'hbc077dd6),
	.w7(32'hbb7e731e),
	.w8(32'hb9c64a99),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b057aaf),
	.w1(32'hbac57622),
	.w2(32'hbb326690),
	.w3(32'hbaa00213),
	.w4(32'hbae3fea4),
	.w5(32'h3a813de5),
	.w6(32'h3b07ecc4),
	.w7(32'h38ae924e),
	.w8(32'hbb8c8b79),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8187dc),
	.w1(32'h3b0271c5),
	.w2(32'h3b6022aa),
	.w3(32'h3bc0ba14),
	.w4(32'h3c480348),
	.w5(32'h3b7c1912),
	.w6(32'h3ba68a10),
	.w7(32'h3b1f8587),
	.w8(32'hbafae2ef),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7f463),
	.w1(32'h3ba58b92),
	.w2(32'h3af6ee74),
	.w3(32'h3b1af067),
	.w4(32'h3ba21fa5),
	.w5(32'h3a1cdb7f),
	.w6(32'hb95f0597),
	.w7(32'h3b4f46e1),
	.w8(32'hb844d3ce),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa00dbc),
	.w1(32'h3b6b0718),
	.w2(32'h3b53a203),
	.w3(32'hbbea5610),
	.w4(32'hbbb7b483),
	.w5(32'h3a936293),
	.w6(32'hbbd85af1),
	.w7(32'hbb583eb0),
	.w8(32'hbc04983a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4cb9),
	.w1(32'h3bb0f4af),
	.w2(32'h3baaf03a),
	.w3(32'hbbda3c18),
	.w4(32'h3a6891d5),
	.w5(32'h3af8993b),
	.w6(32'hbb666125),
	.w7(32'h3b283004),
	.w8(32'hb7a15b8b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5b416),
	.w1(32'hbb372b09),
	.w2(32'hb975a6ee),
	.w3(32'h3b09120c),
	.w4(32'hbae48132),
	.w5(32'h3a275a32),
	.w6(32'hbb9436a1),
	.w7(32'hba573b8f),
	.w8(32'h3a6976d5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ca52),
	.w1(32'h3c1cfeeb),
	.w2(32'hba73c36d),
	.w3(32'hb9582ef0),
	.w4(32'h3ae8aebc),
	.w5(32'hbbf1cc45),
	.w6(32'hbae4ab7e),
	.w7(32'h3b01a6a4),
	.w8(32'hbbb8f12d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d8c8e),
	.w1(32'hbae3d172),
	.w2(32'h3ba99e21),
	.w3(32'h3bc90be4),
	.w4(32'hba7ef510),
	.w5(32'hb9f50a5b),
	.w6(32'h3a319a47),
	.w7(32'h3a177b73),
	.w8(32'h3b811907),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2384),
	.w1(32'hba4cc734),
	.w2(32'hbb3bf510),
	.w3(32'h3ada097c),
	.w4(32'h3b914c8b),
	.w5(32'h3c035392),
	.w6(32'h3a2cdb37),
	.w7(32'hbb21a4ed),
	.w8(32'hbb5eb755),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f33d3e),
	.w1(32'hbbbc3cce),
	.w2(32'hb9b7180b),
	.w3(32'h3b291ffb),
	.w4(32'h3acdbaf9),
	.w5(32'h3b6bd71d),
	.w6(32'hba43d101),
	.w7(32'h3b9e2cb3),
	.w8(32'hbb1d0db7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87f51b),
	.w1(32'hbb099226),
	.w2(32'h3ab1f976),
	.w3(32'h3b65b9be),
	.w4(32'hbc244408),
	.w5(32'hbbe2a2f0),
	.w6(32'hbb546ebc),
	.w7(32'hb934cc48),
	.w8(32'hb9961ed6),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b6e1),
	.w1(32'h3b20d80f),
	.w2(32'h3b77b565),
	.w3(32'hba953062),
	.w4(32'hbb493821),
	.w5(32'h3b67ccfe),
	.w6(32'hbbf9ae78),
	.w7(32'h3b138420),
	.w8(32'h3b915e49),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85a6eb),
	.w1(32'h3a2b9d1f),
	.w2(32'h3b744ca8),
	.w3(32'hba949f35),
	.w4(32'h3b9a5ba8),
	.w5(32'h3c7d169a),
	.w6(32'h3aaf7db6),
	.w7(32'h39b7a07c),
	.w8(32'h3c0dbff0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9c390),
	.w1(32'h3b86a5bb),
	.w2(32'hbbb025fb),
	.w3(32'hbaaed953),
	.w4(32'h3a39b07b),
	.w5(32'h3bc33369),
	.w6(32'hbab70c4f),
	.w7(32'hbad2940e),
	.w8(32'h3bc25573),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec3441),
	.w1(32'h38e6a5c2),
	.w2(32'hbb6798ac),
	.w3(32'hbb7bc0c4),
	.w4(32'hbb784056),
	.w5(32'hbb7d760f),
	.w6(32'hbad6f0fb),
	.w7(32'hbbd9e63d),
	.w8(32'h3b011c58),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eb451),
	.w1(32'h3b13f202),
	.w2(32'hbb135ab3),
	.w3(32'h3b541fdc),
	.w4(32'h3b1ff93f),
	.w5(32'h3be878d2),
	.w6(32'h3bb95e8d),
	.w7(32'h3b250561),
	.w8(32'h3b4d9a56),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93d7d6),
	.w1(32'h3adff59d),
	.w2(32'h3b48b990),
	.w3(32'h3af82f7a),
	.w4(32'h3b118f1d),
	.w5(32'hbaf425c9),
	.w6(32'h3b67cf6a),
	.w7(32'h3b70501a),
	.w8(32'h3a8ceed8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32448a),
	.w1(32'hbad914f4),
	.w2(32'h3b9b686f),
	.w3(32'h3b70177a),
	.w4(32'h3b37b53a),
	.w5(32'hbaaf8e08),
	.w6(32'h3b927f3f),
	.w7(32'h3ae5397a),
	.w8(32'h3b9173db),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b568b2f),
	.w1(32'h3ba62612),
	.w2(32'h3b8cd6c5),
	.w3(32'hbb4c5e15),
	.w4(32'hbb2f58f6),
	.w5(32'hbabb1f08),
	.w6(32'hba90bf0b),
	.w7(32'hbb5e2814),
	.w8(32'h3b00a0f0),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0a075),
	.w1(32'hbbb98774),
	.w2(32'hbb9641f8),
	.w3(32'hbb88475c),
	.w4(32'hbbb6922c),
	.w5(32'hbab4b23f),
	.w6(32'hbb09ebe9),
	.w7(32'hbc049f7e),
	.w8(32'hbbd0791a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f399),
	.w1(32'hb928b7a0),
	.w2(32'h3b25a7f1),
	.w3(32'hbb92ce4b),
	.w4(32'h3b16deab),
	.w5(32'hbb037581),
	.w6(32'hbbe27dbf),
	.w7(32'h3b317c7d),
	.w8(32'hbacb7bca),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ebce0),
	.w1(32'hbaca81b1),
	.w2(32'hbbad3423),
	.w3(32'h3ad24c5e),
	.w4(32'hbb24d168),
	.w5(32'hba503a36),
	.w6(32'h39cdd617),
	.w7(32'hba9053d4),
	.w8(32'hbae6c262),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b0de),
	.w1(32'hbb3b035d),
	.w2(32'hbb131a4d),
	.w3(32'h3906e35d),
	.w4(32'hbb33b27f),
	.w5(32'h3bb16e64),
	.w6(32'hbaa592e1),
	.w7(32'hbbdb56a5),
	.w8(32'hbc14c0c5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eb2e5),
	.w1(32'hbb70df5b),
	.w2(32'h3bc34f2e),
	.w3(32'h3b4ef5ba),
	.w4(32'hbb444f6d),
	.w5(32'hbb473f94),
	.w6(32'hbbb5a158),
	.w7(32'h3aaaf84a),
	.w8(32'hba061126),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe421a),
	.w1(32'h3b487a96),
	.w2(32'h3a01ca0d),
	.w3(32'h3b5f6b49),
	.w4(32'h3bdd2850),
	.w5(32'h3c4d11a2),
	.w6(32'h3b550d2f),
	.w7(32'h3a5a382e),
	.w8(32'hba55b760),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71d121),
	.w1(32'hbb1da0ff),
	.w2(32'hbbdec4df),
	.w3(32'hbb4c562e),
	.w4(32'hbab0d229),
	.w5(32'hbc367cf1),
	.w6(32'hba0e1149),
	.w7(32'h38a863e2),
	.w8(32'hba9a01da),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d5614),
	.w1(32'h3ae0ed17),
	.w2(32'hbb37af1d),
	.w3(32'hb9637744),
	.w4(32'h3a310b9b),
	.w5(32'h3c34b851),
	.w6(32'hbaed16e3),
	.w7(32'h3b3cdd3e),
	.w8(32'h3c1a47d3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule