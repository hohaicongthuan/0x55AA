module layer_10_featuremap_30(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbc79d),
	.w1(32'h3be3918f),
	.w2(32'h3afb8c76),
	.w3(32'h3bae5d97),
	.w4(32'h3bce8b54),
	.w5(32'hba07d84b),
	.w6(32'hbac2a194),
	.w7(32'hba3d6a05),
	.w8(32'hbb949126),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a834304),
	.w1(32'h3b7af94c),
	.w2(32'h3b3e2a0a),
	.w3(32'h3aefa19c),
	.w4(32'hbaf59073),
	.w5(32'h3b55c075),
	.w6(32'h3af9136a),
	.w7(32'h3b9dd043),
	.w8(32'h3b0b476a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab310b),
	.w1(32'hbba5c77f),
	.w2(32'h3ba4461e),
	.w3(32'h3c012a41),
	.w4(32'hbb2bd729),
	.w5(32'hba95d2a2),
	.w6(32'h3b082346),
	.w7(32'h3af98d01),
	.w8(32'hbb397d90),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ae8e2),
	.w1(32'h3ae48c0f),
	.w2(32'h3a7eba72),
	.w3(32'hbba4a614),
	.w4(32'hbb22f63d),
	.w5(32'h3a974dc3),
	.w6(32'hbae53c51),
	.w7(32'h3af5fa42),
	.w8(32'hbb9c76f0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b128318),
	.w1(32'h3afd98a2),
	.w2(32'hbad27ce2),
	.w3(32'h3b996605),
	.w4(32'h3a3774df),
	.w5(32'hbbf6e03d),
	.w6(32'hbc091b83),
	.w7(32'h3b1c0070),
	.w8(32'hbbfd06e0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32f4c2),
	.w1(32'h3b5cddf6),
	.w2(32'hbd3bb682),
	.w3(32'hbb287ed5),
	.w4(32'h3a4337b8),
	.w5(32'hbd2b7d80),
	.w6(32'hb9607073),
	.w7(32'h3b2be45f),
	.w8(32'hbd1648d7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70853d),
	.w1(32'h3ce69a0f),
	.w2(32'hbbdd9ea3),
	.w3(32'h3d567318),
	.w4(32'h3db1f4e1),
	.w5(32'hbbea3198),
	.w6(32'h3d3bdd79),
	.w7(32'h3d7f61a2),
	.w8(32'hbb969da8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9301),
	.w1(32'hba1d7590),
	.w2(32'hbacc0d55),
	.w3(32'h37b8a70f),
	.w4(32'hbb850fe0),
	.w5(32'h39b0c0d0),
	.w6(32'h3a0e7168),
	.w7(32'hbb90d2d9),
	.w8(32'hbab97063),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc542),
	.w1(32'h3bf37629),
	.w2(32'h3bb78587),
	.w3(32'h3a3ed7e2),
	.w4(32'h3baf6614),
	.w5(32'h3b39ac84),
	.w6(32'h3a8ab519),
	.w7(32'h3aae3e83),
	.w8(32'h3bf0c587),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b679e6a),
	.w1(32'h3bc22b4f),
	.w2(32'hbc63029a),
	.w3(32'h3ba87e10),
	.w4(32'h3ad5a80a),
	.w5(32'hbc86c588),
	.w6(32'h3c0f8ccc),
	.w7(32'h3b39b054),
	.w8(32'hbc2f1f19),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb7f31),
	.w1(32'h3c33b1d9),
	.w2(32'h3c093cd6),
	.w3(32'h3c545915),
	.w4(32'h3cdf5426),
	.w5(32'h3a5ecfa8),
	.w6(32'h3c69857a),
	.w7(32'h3cd15db1),
	.w8(32'hb9c1ffde),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab32f2),
	.w1(32'h3b3fba87),
	.w2(32'h3b56e93f),
	.w3(32'hbac493e7),
	.w4(32'hbb84e90f),
	.w5(32'h3b0c4e66),
	.w6(32'hbb1ada9c),
	.w7(32'hbb0b2958),
	.w8(32'h3b0df7cc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf461cc),
	.w1(32'hbc25343b),
	.w2(32'hbb025654),
	.w3(32'hbc0f6665),
	.w4(32'hbc8aad2c),
	.w5(32'h37d01e6a),
	.w6(32'hbbaecba3),
	.w7(32'hbc826785),
	.w8(32'hbaa05855),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc183e64),
	.w1(32'hbc0b7a93),
	.w2(32'hba8776ad),
	.w3(32'hbb8e5bb4),
	.w4(32'hbbf7b468),
	.w5(32'hbbbc8f07),
	.w6(32'hbb98245d),
	.w7(32'hbba45a9b),
	.w8(32'hb9c7a062),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45fef),
	.w1(32'h3b679470),
	.w2(32'hbae01690),
	.w3(32'hbbddd012),
	.w4(32'h3abe83df),
	.w5(32'hba4037b3),
	.w6(32'hbaf99d7b),
	.w7(32'h3b56a584),
	.w8(32'hbbbbf671),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1f77b),
	.w1(32'h3986942d),
	.w2(32'hbccc3bd3),
	.w3(32'h39f3069c),
	.w4(32'h3aaa6226),
	.w5(32'hbcca665a),
	.w6(32'hb8d8cd65),
	.w7(32'hbb1fda65),
	.w8(32'hbc8d94af),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012364),
	.w1(32'h3cfba75e),
	.w2(32'h3b181b8c),
	.w3(32'h3d1dcf2c),
	.w4(32'h3d84cad1),
	.w5(32'hbabe6a2a),
	.w6(32'h3d0e8cd8),
	.w7(32'h3d5ac4c5),
	.w8(32'hbb853554),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0302b4),
	.w1(32'h3be33353),
	.w2(32'h38f28e09),
	.w3(32'h3b45df39),
	.w4(32'h3bd5df20),
	.w5(32'h399a0fb9),
	.w6(32'hb9616054),
	.w7(32'h3b13d9d5),
	.w8(32'hba8d5777),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c023f8),
	.w1(32'hba7381a5),
	.w2(32'hbb4e8570),
	.w3(32'hbb87a500),
	.w4(32'hba9eafe0),
	.w5(32'hba04f903),
	.w6(32'hbb220ad8),
	.w7(32'hbb40c159),
	.w8(32'h3bc90a04),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13778b),
	.w1(32'h3c05dac6),
	.w2(32'hbad170ee),
	.w3(32'hbbecf949),
	.w4(32'h3bc60adc),
	.w5(32'h3af878d1),
	.w6(32'h3b35833b),
	.w7(32'h3b9bc5ab),
	.w8(32'hbb360217),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821008),
	.w1(32'h3b0ec456),
	.w2(32'hba5d4755),
	.w3(32'h3b8d7c69),
	.w4(32'h3abe4b05),
	.w5(32'hb7db259d),
	.w6(32'hba959a44),
	.w7(32'h3ab2994d),
	.w8(32'h3a019b5f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941f2d),
	.w1(32'h3abdc7f1),
	.w2(32'h3b1d4968),
	.w3(32'h3adde794),
	.w4(32'h3b892503),
	.w5(32'h3a310039),
	.w6(32'hba072f7a),
	.w7(32'h3af5528c),
	.w8(32'h3b07613b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf674a),
	.w1(32'hbb50bfa1),
	.w2(32'h3ca88414),
	.w3(32'hbb3d9e24),
	.w4(32'hbbaaaa75),
	.w5(32'h3c92562a),
	.w6(32'h3b608676),
	.w7(32'h37152770),
	.w8(32'h3ccd4200),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cc441),
	.w1(32'hbc561946),
	.w2(32'h3a94ff80),
	.w3(32'hbcab8764),
	.w4(32'hbcf78445),
	.w5(32'hba3b6a74),
	.w6(32'hbbd32668),
	.w7(32'hbc6d5684),
	.w8(32'hbb620ab7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32a627),
	.w1(32'hbbb7331f),
	.w2(32'hbb611776),
	.w3(32'hbbee76c8),
	.w4(32'hbbc628cd),
	.w5(32'hbbfd38f0),
	.w6(32'h3acc1797),
	.w7(32'hbbbb7ae3),
	.w8(32'hbbcf0d6e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fb979),
	.w1(32'h3b848422),
	.w2(32'h383488ad),
	.w3(32'hbbf661e0),
	.w4(32'hbaa40f10),
	.w5(32'hbb9a3276),
	.w6(32'hbb7cbb49),
	.w7(32'hbb0a8b13),
	.w8(32'hba6d2493),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb62b40),
	.w1(32'h3ad89ea4),
	.w2(32'h394e0d21),
	.w3(32'hbb24a731),
	.w4(32'hbb9c230b),
	.w5(32'hbab88890),
	.w6(32'hbb31aa0d),
	.w7(32'hbb71accc),
	.w8(32'hb83054da),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585c5b),
	.w1(32'h3a355eb5),
	.w2(32'hbbb522ba),
	.w3(32'h3af5a3d9),
	.w4(32'hb9f83e21),
	.w5(32'hbc0d1076),
	.w6(32'hba42a330),
	.w7(32'h3a27d07a),
	.w8(32'hbbdd44b3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4b8ef),
	.w1(32'hbc07f2ca),
	.w2(32'hb9ba4500),
	.w3(32'h3c630a97),
	.w4(32'hbb687b87),
	.w5(32'h3a3968a0),
	.w6(32'h3b81276c),
	.w7(32'h3a541f34),
	.w8(32'h3af4ce5d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca33423),
	.w1(32'hbc477cb9),
	.w2(32'hbafe9bd7),
	.w3(32'hbc44c9e2),
	.w4(32'h38cb8d76),
	.w5(32'h3b01e2ab),
	.w6(32'hbc32d974),
	.w7(32'h3c866529),
	.w8(32'hba00d651),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28d166),
	.w1(32'hbaa95617),
	.w2(32'h3a8eb25f),
	.w3(32'h3b69d101),
	.w4(32'h3a66a29f),
	.w5(32'h39f50d0c),
	.w6(32'h3ae53e80),
	.w7(32'h3883ef99),
	.w8(32'hba21b589),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8155b7),
	.w1(32'hbbf1a714),
	.w2(32'hbb51dd76),
	.w3(32'h3bc897b7),
	.w4(32'hbc323ba4),
	.w5(32'hbbda6354),
	.w6(32'h3b9b2542),
	.w7(32'hba74f36b),
	.w8(32'hba9670e2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc6b23),
	.w1(32'hbb5b341f),
	.w2(32'h3a04725a),
	.w3(32'hbbdfa8b9),
	.w4(32'hbc625b77),
	.w5(32'h3a3fb4b2),
	.w6(32'hbc047d2d),
	.w7(32'hbc02782c),
	.w8(32'hba8110da),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c789c),
	.w1(32'hb9bed961),
	.w2(32'hbae77a27),
	.w3(32'h3b711e6f),
	.w4(32'hba22af55),
	.w5(32'hb954a899),
	.w6(32'h3b41682c),
	.w7(32'hbaaa3e23),
	.w8(32'h39e9c18b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf3bd5),
	.w1(32'h3bddeffe),
	.w2(32'hbb14b76e),
	.w3(32'hbb59c425),
	.w4(32'h3c854774),
	.w5(32'hbae096c8),
	.w6(32'h3b579263),
	.w7(32'h3c80166f),
	.w8(32'hbb10f8a7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf8371),
	.w1(32'hbba43b63),
	.w2(32'h3c37b822),
	.w3(32'h3b4e03eb),
	.w4(32'hbb52728e),
	.w5(32'h3b85a002),
	.w6(32'h3b2e1011),
	.w7(32'hbb581b7a),
	.w8(32'hbae2e383),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9da313),
	.w1(32'hbaeb9944),
	.w2(32'hbb924bc3),
	.w3(32'hbc6bda0c),
	.w4(32'h3b9fb088),
	.w5(32'hbae2af89),
	.w6(32'hbbec2c0a),
	.w7(32'h3cb788d1),
	.w8(32'hbb6d7c83),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500545),
	.w1(32'hbb638fce),
	.w2(32'h3ada7c62),
	.w3(32'h3b421569),
	.w4(32'h3b049eb9),
	.w5(32'hbb7a8e1c),
	.w6(32'hba09ed0c),
	.w7(32'h3b23cc93),
	.w8(32'hb9ce190f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65a25c),
	.w1(32'hbad915bd),
	.w2(32'hbc90667e),
	.w3(32'h3c56cc06),
	.w4(32'h3aa50735),
	.w5(32'hbcaf7bf4),
	.w6(32'h3c340105),
	.w7(32'hbb4a9926),
	.w8(32'hbc75184e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78c32f),
	.w1(32'hbbbb73ca),
	.w2(32'hb9a416ce),
	.w3(32'h3ce4f384),
	.w4(32'hbc07d1b5),
	.w5(32'h3c11b75d),
	.w6(32'h3c4710f2),
	.w7(32'h3ba64a4e),
	.w8(32'hbb0f5475),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e6c10),
	.w1(32'hbc181e8b),
	.w2(32'h3b025d94),
	.w3(32'h3a9b7455),
	.w4(32'hba2b1a6f),
	.w5(32'hba2b698a),
	.w6(32'h3b592629),
	.w7(32'hbb78c1cd),
	.w8(32'hbc247467),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebe4f),
	.w1(32'hb8bf3f0f),
	.w2(32'hba5e0f1d),
	.w3(32'hbaf803f8),
	.w4(32'hbaad3e23),
	.w5(32'hbab183d9),
	.w6(32'hbb8d8269),
	.w7(32'hbb341abb),
	.w8(32'hbb1cda03),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9407ac),
	.w1(32'h3a489a8f),
	.w2(32'hbaff70b8),
	.w3(32'hbc378c29),
	.w4(32'hbc22ec19),
	.w5(32'hba6c4be8),
	.w6(32'hbab19e3c),
	.w7(32'h3b0d8a79),
	.w8(32'h3ac34078),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96e966),
	.w1(32'hbb859a37),
	.w2(32'hbc25f5a8),
	.w3(32'h3bc17e7d),
	.w4(32'h39a9c447),
	.w5(32'hbbb7abeb),
	.w6(32'h3bfd64d8),
	.w7(32'h3b32722c),
	.w8(32'hbc4bd417),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c172c04),
	.w1(32'hbc38950e),
	.w2(32'h3c012158),
	.w3(32'hbb910f16),
	.w4(32'hb7af26c2),
	.w5(32'hbb3efb00),
	.w6(32'hbc504deb),
	.w7(32'h3bd7b104),
	.w8(32'h3b92b6c7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76c841),
	.w1(32'hbc5876fd),
	.w2(32'hbcb3f780),
	.w3(32'h3b9f76b6),
	.w4(32'hbbff51ec),
	.w5(32'hbbe5e574),
	.w6(32'h3b921cac),
	.w7(32'hbb9e54e9),
	.w8(32'h391d297c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc313e04),
	.w1(32'h3bb6d09c),
	.w2(32'h3c9528a8),
	.w3(32'hbce22f4b),
	.w4(32'h3ca82d69),
	.w5(32'h3ca70dc7),
	.w6(32'hbcef1d34),
	.w7(32'h3c653920),
	.w8(32'h3c2fbbb0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1292e6),
	.w1(32'h3cfeda6d),
	.w2(32'h3a83ca52),
	.w3(32'hbce63170),
	.w4(32'h3ce54fd1),
	.w5(32'hb80c1f8f),
	.w6(32'hbc440f59),
	.w7(32'h3c6e97fb),
	.w8(32'h3af04d70),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bbbd5),
	.w1(32'hbb7906e4),
	.w2(32'h3b8db352),
	.w3(32'h3ae5c2a5),
	.w4(32'hbaacd5d4),
	.w5(32'h3b5daaa1),
	.w6(32'h3b5de03a),
	.w7(32'hb84e2092),
	.w8(32'h3aee5713),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37705faa),
	.w1(32'h3bb9de9b),
	.w2(32'h3bf1cd8e),
	.w3(32'h3c6f1486),
	.w4(32'hbac1c737),
	.w5(32'hbb288b95),
	.w6(32'h3c0d07b8),
	.w7(32'hbba6eeb5),
	.w8(32'h3c0827e7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbf96c),
	.w1(32'hbbe43f13),
	.w2(32'hbbcd3e7e),
	.w3(32'h39349d1b),
	.w4(32'hbb7e1050),
	.w5(32'hbc56e60a),
	.w6(32'h3bbea1bb),
	.w7(32'h3c2c0a23),
	.w8(32'hbc864a5a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3672d3),
	.w1(32'hbc320d6f),
	.w2(32'h3b2faa64),
	.w3(32'hbbd28738),
	.w4(32'hbc27d50b),
	.w5(32'hbab7bef6),
	.w6(32'hbb11449a),
	.w7(32'hbbfd1343),
	.w8(32'h3926d18a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c2973),
	.w1(32'hbbfa5646),
	.w2(32'h3b5c8fc5),
	.w3(32'h3b25941b),
	.w4(32'hbc793212),
	.w5(32'h3ab87174),
	.w6(32'h3bf36843),
	.w7(32'hbbbddeb6),
	.w8(32'hbaa48078),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073788),
	.w1(32'h3adfe836),
	.w2(32'h3bd5efa2),
	.w3(32'h3bc7c246),
	.w4(32'hba0d6931),
	.w5(32'h3ad91011),
	.w6(32'h3b16f357),
	.w7(32'hbab4f94d),
	.w8(32'hbc11a132),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c330f22),
	.w1(32'hba9545bb),
	.w2(32'h3bdd858f),
	.w3(32'hba23b590),
	.w4(32'h3c52347b),
	.w5(32'hb987421a),
	.w6(32'h39b88ccc),
	.w7(32'h3c68c98e),
	.w8(32'hbaba2d78),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94959c),
	.w1(32'h3bbead92),
	.w2(32'hbc699f33),
	.w3(32'h3c8c20c8),
	.w4(32'hbbee257a),
	.w5(32'hbca8b8b9),
	.w6(32'h3c9a588f),
	.w7(32'hbb9dd037),
	.w8(32'hbbb77509),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d61ba),
	.w1(32'hbcbe737f),
	.w2(32'h3aecf10f),
	.w3(32'h3c76ebe4),
	.w4(32'hbc4f3b11),
	.w5(32'h3b5cc729),
	.w6(32'hbbdf3f1c),
	.w7(32'h3bbc5387),
	.w8(32'h3baf0c50),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15fdc5),
	.w1(32'hba2c16fe),
	.w2(32'hba2e7879),
	.w3(32'hbb72979b),
	.w4(32'h3b81607c),
	.w5(32'hbab88229),
	.w6(32'hba92dce1),
	.w7(32'h3b2ccf74),
	.w8(32'h3b9b6eeb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20683),
	.w1(32'hbc406b6d),
	.w2(32'hba83e79f),
	.w3(32'h3a699928),
	.w4(32'hbbf62bad),
	.w5(32'hbaa34200),
	.w6(32'h3b5d2a13),
	.w7(32'hb9ad45d6),
	.w8(32'h3acaaae1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67f89a),
	.w1(32'h3b5dd7f6),
	.w2(32'h3c6f83c2),
	.w3(32'hb9bb7836),
	.w4(32'h3acac2e9),
	.w5(32'h3bee2ebd),
	.w6(32'h3b8aae7f),
	.w7(32'h3b97a49e),
	.w8(32'h3bd02996),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea265),
	.w1(32'hba9ebb1c),
	.w2(32'hbc2ef6e5),
	.w3(32'hbb8c306b),
	.w4(32'h3a99b64c),
	.w5(32'h3c151acc),
	.w6(32'h3aa5ab9e),
	.w7(32'hbacf32d4),
	.w8(32'h3bf84b81),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52ff20),
	.w1(32'h3b9114d6),
	.w2(32'hbaec4bd5),
	.w3(32'h3ba42164),
	.w4(32'h3c08625c),
	.w5(32'h3bc1a943),
	.w6(32'hbc0dbe15),
	.w7(32'h3c176341),
	.w8(32'h3bcabecd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2059a7),
	.w1(32'h3b59611b),
	.w2(32'hba920a7e),
	.w3(32'hbc1034f1),
	.w4(32'hbb1148b3),
	.w5(32'hbb956ff2),
	.w6(32'h3a084271),
	.w7(32'hbbe7fba1),
	.w8(32'hbba2a647),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1e88d),
	.w1(32'hbbb04002),
	.w2(32'h3ba8f9bd),
	.w3(32'hba4cf707),
	.w4(32'h3a2a61c4),
	.w5(32'hbc136d43),
	.w6(32'hbb17a513),
	.w7(32'hbb7b8eae),
	.w8(32'h37cc7bbd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2332c),
	.w1(32'hbb488bd8),
	.w2(32'h3bbf1805),
	.w3(32'h3ad835d7),
	.w4(32'hbb9061ae),
	.w5(32'h3b9c2796),
	.w6(32'h3c079752),
	.w7(32'h399f75c5),
	.w8(32'h3b9b6379),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e873c),
	.w1(32'h3a52b657),
	.w2(32'hbaf956de),
	.w3(32'h3b9105bc),
	.w4(32'h3b5c6b90),
	.w5(32'hbb09fa5e),
	.w6(32'h3beb90be),
	.w7(32'h3b5460d4),
	.w8(32'hb9f2916a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e80a8),
	.w1(32'h3a46caa3),
	.w2(32'hbbc809ad),
	.w3(32'h3bb1287b),
	.w4(32'h3b1be7ca),
	.w5(32'hbb238c37),
	.w6(32'h3bb1023f),
	.w7(32'h3bccf9ea),
	.w8(32'hbac5531c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb81f84),
	.w1(32'hbb080425),
	.w2(32'h3b2b34d7),
	.w3(32'hbcaf5b52),
	.w4(32'hbc42e662),
	.w5(32'h3aa9b81d),
	.w6(32'hbcb800a8),
	.w7(32'hbb7f3b20),
	.w8(32'h3a07e8b9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e77a),
	.w1(32'h39886a56),
	.w2(32'hbb978a4d),
	.w3(32'h3bf636c8),
	.w4(32'hb97fae5a),
	.w5(32'hbb808460),
	.w6(32'h3bc6c189),
	.w7(32'hbaec4e88),
	.w8(32'hbafb955a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ecf93),
	.w1(32'hb97247dc),
	.w2(32'hbbe888a0),
	.w3(32'hbb17c510),
	.w4(32'h3a98baab),
	.w5(32'hbb600027),
	.w6(32'hbab3a7a5),
	.w7(32'h3ab9799f),
	.w8(32'hbaab49cd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c256f15),
	.w1(32'h374f5606),
	.w2(32'hbc78acc4),
	.w3(32'h3c161886),
	.w4(32'h3baeb3f1),
	.w5(32'hbc1a8573),
	.w6(32'h3adcae0c),
	.w7(32'h3bd27655),
	.w8(32'hbb5bcfe6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce0721),
	.w1(32'hbbc565e1),
	.w2(32'h3b03c8f1),
	.w3(32'hbac9549b),
	.w4(32'h3b3a5d36),
	.w5(32'h3c30143c),
	.w6(32'hbb59839b),
	.w7(32'h3baca41f),
	.w8(32'h3c4e8fff),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc302581),
	.w1(32'h3c31843d),
	.w2(32'hbba26d43),
	.w3(32'hbc488bd5),
	.w4(32'h3d066458),
	.w5(32'hbb8ac458),
	.w6(32'hbc73a96a),
	.w7(32'h3ce5413c),
	.w8(32'hbc53f27f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7983a2),
	.w1(32'hbd1adb61),
	.w2(32'hbafd6fcb),
	.w3(32'h3cdb18ef),
	.w4(32'hbd47e325),
	.w5(32'h3983aa81),
	.w6(32'h3ccac766),
	.w7(32'hbce197f7),
	.w8(32'hba55b578),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7434e3),
	.w1(32'hbbb90aee),
	.w2(32'hb890d2d9),
	.w3(32'h3bc0d13a),
	.w4(32'hbb09fd8f),
	.w5(32'hbac47e60),
	.w6(32'h3bb5527d),
	.w7(32'hba27a89a),
	.w8(32'hba882c59),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d653f),
	.w1(32'hbc3ecabc),
	.w2(32'h3a6ffc7c),
	.w3(32'h399e083f),
	.w4(32'hbbf9153d),
	.w5(32'hbb9370dc),
	.w6(32'h3a4871bd),
	.w7(32'hbc332c99),
	.w8(32'hbb51ce0c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae16feb),
	.w1(32'hbb8106e7),
	.w2(32'hba15cff5),
	.w3(32'h3c3fcfa8),
	.w4(32'hbb4d0ece),
	.w5(32'hbbcc3e50),
	.w6(32'h3c06ccf1),
	.w7(32'h3b9fbf58),
	.w8(32'hbc097ad9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac2c0f),
	.w1(32'hbb8dce04),
	.w2(32'h3b4658b8),
	.w3(32'h3c4386d0),
	.w4(32'hbc0279ca),
	.w5(32'h3a0d6524),
	.w6(32'hbb23747f),
	.w7(32'h3bb30c78),
	.w8(32'hbbdce97f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb82aeb),
	.w1(32'h3c0d82fd),
	.w2(32'hba3aebbf),
	.w3(32'hbd0d7df6),
	.w4(32'h3c858716),
	.w5(32'h3a297944),
	.w6(32'hbcc60e50),
	.w7(32'h3c6b71d1),
	.w8(32'hbae6324e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85c435),
	.w1(32'h3a8e5366),
	.w2(32'hbb39fe39),
	.w3(32'h3c1ff63d),
	.w4(32'h3ac2cdfe),
	.w5(32'hb9c38245),
	.w6(32'hba932ec0),
	.w7(32'hba2aa108),
	.w8(32'h35c71e42),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc390ddb),
	.w1(32'h3bb13a07),
	.w2(32'hbb4e418d),
	.w3(32'hbc4ada63),
	.w4(32'h3bbdfef7),
	.w5(32'hbb5b8b76),
	.w6(32'hbc2cb79c),
	.w7(32'h3b724ae7),
	.w8(32'hbb453756),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3352d),
	.w1(32'hbba2d767),
	.w2(32'h3c2c6230),
	.w3(32'hb92c1e0a),
	.w4(32'hbaff6324),
	.w5(32'h3ca7daa4),
	.w6(32'hbb1a5399),
	.w7(32'hbad31719),
	.w8(32'h3c924f47),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cb314),
	.w1(32'h3c9c3e10),
	.w2(32'hbbbd403c),
	.w3(32'hbcba8b86),
	.w4(32'h3cf12445),
	.w5(32'hbbbea4d6),
	.w6(32'hbc9532f7),
	.w7(32'h3d00e683),
	.w8(32'hbbcbe885),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfea313),
	.w1(32'hbbb3d7a1),
	.w2(32'hbafc05d5),
	.w3(32'hbcb7acec),
	.w4(32'h3c64ad67),
	.w5(32'h3a2135cd),
	.w6(32'hbc3b0901),
	.w7(32'h3b01ca44),
	.w8(32'h3bd79294),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf18a9a),
	.w1(32'h3b7016aa),
	.w2(32'hbbbb78a3),
	.w3(32'hbcc57d57),
	.w4(32'h3c9315f1),
	.w5(32'hbc58ff8a),
	.w6(32'hbce624ef),
	.w7(32'h3c348a5c),
	.w8(32'hbc1d67fc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb10b0b),
	.w1(32'hbc66465e),
	.w2(32'h3a56e438),
	.w3(32'h3cbbfca0),
	.w4(32'hbc0e3b00),
	.w5(32'h3bbb7c20),
	.w6(32'h3c28ac62),
	.w7(32'hbc2e3b15),
	.w8(32'h3be5ab92),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097c16),
	.w1(32'hbbdcb63f),
	.w2(32'hbabc238f),
	.w3(32'hbb92266a),
	.w4(32'hbb31de45),
	.w5(32'hbab4b48e),
	.w6(32'h3a4d2029),
	.w7(32'h3ada75b4),
	.w8(32'h3a695118),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919a5ef),
	.w1(32'hbb56f3a9),
	.w2(32'h3ae78ef3),
	.w3(32'h3ab1de60),
	.w4(32'hba6e2667),
	.w5(32'hba9eb7db),
	.w6(32'h3b2ac4e7),
	.w7(32'hba8b58de),
	.w8(32'hbb0295b1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c4114),
	.w1(32'hbbf6b8fa),
	.w2(32'h3ab54d3f),
	.w3(32'hbc2fec9c),
	.w4(32'hbc24b9ee),
	.w5(32'hbb86e449),
	.w6(32'hbb9a08e2),
	.w7(32'hbb212dba),
	.w8(32'hbbabf083),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb8a62),
	.w1(32'hbba1d1de),
	.w2(32'h3b16afd3),
	.w3(32'hbb4f6dfc),
	.w4(32'hbb005a0d),
	.w5(32'hbbec4e71),
	.w6(32'hbc051c52),
	.w7(32'hbb66f61c),
	.w8(32'hbb3aa88c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73f450),
	.w1(32'hbaf3d0f6),
	.w2(32'h3bcd160c),
	.w3(32'h3b92575a),
	.w4(32'hba0c4e7b),
	.w5(32'hba947a4a),
	.w6(32'h3b9d5b8d),
	.w7(32'hb9e18193),
	.w8(32'hbb7a3a43),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2cd7),
	.w1(32'h3ba49cfc),
	.w2(32'hbb6aefe8),
	.w3(32'hbb39b08d),
	.w4(32'h3c0a2b53),
	.w5(32'h3b5edaea),
	.w6(32'hb9c9a256),
	.w7(32'h3b8954c6),
	.w8(32'h3b10fcd3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb3d9),
	.w1(32'hbb0386c6),
	.w2(32'h39c673c4),
	.w3(32'h3bd81741),
	.w4(32'h3b2bc1ca),
	.w5(32'h3b2dfcb6),
	.w6(32'h3bae1dbc),
	.w7(32'hb7c8c1c1),
	.w8(32'h3b18f927),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319aac),
	.w1(32'hbb2cb574),
	.w2(32'h398887ac),
	.w3(32'h3b2b81e6),
	.w4(32'h38ca015e),
	.w5(32'hbba34487),
	.w6(32'h3b5a8233),
	.w7(32'h399ca446),
	.w8(32'h3b822b5b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34ebc3),
	.w1(32'hb98fc5dc),
	.w2(32'hbb70c929),
	.w3(32'h3c159834),
	.w4(32'hbc06ab62),
	.w5(32'h3b1e91e6),
	.w6(32'h3c0768af),
	.w7(32'hbb522a52),
	.w8(32'hbaa03e05),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b585f),
	.w1(32'h3a383558),
	.w2(32'hb9d16e63),
	.w3(32'hbabf3ded),
	.w4(32'hbadeee47),
	.w5(32'hbbd6c3fb),
	.w6(32'hbbe57ff4),
	.w7(32'hbc330047),
	.w8(32'h3b0422e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd39d),
	.w1(32'hbc2717e7),
	.w2(32'hbbacf615),
	.w3(32'hbc661f07),
	.w4(32'hbc66558f),
	.w5(32'h3b129a12),
	.w6(32'hbc4e1bb1),
	.w7(32'hb90e44ea),
	.w8(32'h3c29f172),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b369335),
	.w1(32'hbbeb8ffc),
	.w2(32'h3bab07e5),
	.w3(32'hbcdd56d1),
	.w4(32'h3ac7d4bd),
	.w5(32'hba6994c9),
	.w6(32'hbc4f85d3),
	.w7(32'h3b54075e),
	.w8(32'hbbdc8739),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01b3f),
	.w1(32'hbb2cd7f8),
	.w2(32'hbb878f67),
	.w3(32'h389fed5b),
	.w4(32'hbb698ffd),
	.w5(32'h3928dd73),
	.w6(32'h3bf8aeb3),
	.w7(32'hbb538743),
	.w8(32'h3b501cff),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb155cad),
	.w1(32'hbae667ec),
	.w2(32'h3c1c1665),
	.w3(32'h39bd14ed),
	.w4(32'h3aef6675),
	.w5(32'hb9eca787),
	.w6(32'h3abf8b1b),
	.w7(32'h3a47ffdd),
	.w8(32'hbc195bcc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7100),
	.w1(32'hbc495bfa),
	.w2(32'hba39b877),
	.w3(32'h3c425354),
	.w4(32'hbc06bc31),
	.w5(32'hbbca39e0),
	.w6(32'h3c331be6),
	.w7(32'hbb53f1af),
	.w8(32'hbc04cc00),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a972431),
	.w1(32'h3ae76bef),
	.w2(32'h39f16185),
	.w3(32'h3bf357f8),
	.w4(32'hbb7ad73f),
	.w5(32'h3ae08696),
	.w6(32'h3bd913d5),
	.w7(32'hba8069be),
	.w8(32'h3af02508),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cee0d),
	.w1(32'hbb182ffe),
	.w2(32'hbb26acfd),
	.w3(32'h3c0415a0),
	.w4(32'hbbbab8ab),
	.w5(32'hba02b193),
	.w6(32'h3b8b94f5),
	.w7(32'hbba030d6),
	.w8(32'h3ac4ae18),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b019ceb),
	.w1(32'hb99e5190),
	.w2(32'hbcc54290),
	.w3(32'h3b6476cb),
	.w4(32'hbaf385a2),
	.w5(32'hbc81ee44),
	.w6(32'hbab697f2),
	.w7(32'hbb454547),
	.w8(32'hbc60d077),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35c5cd),
	.w1(32'h3b84e179),
	.w2(32'hbc493733),
	.w3(32'hbc4678d3),
	.w4(32'h3b7612ad),
	.w5(32'hbb8961b9),
	.w6(32'hbc8b5f00),
	.w7(32'h3b967ffb),
	.w8(32'hbb180b7b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e807),
	.w1(32'h3af4bfa9),
	.w2(32'hbc00886c),
	.w3(32'hbb0bdd21),
	.w4(32'h3baa3bc8),
	.w5(32'hbb0a7896),
	.w6(32'hbbcaa114),
	.w7(32'h3bafbaf7),
	.w8(32'h3a2c73b6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdad3cd),
	.w1(32'h3bff0b69),
	.w2(32'hbba2a55a),
	.w3(32'hbbf9c473),
	.w4(32'h3c32f6d2),
	.w5(32'h3b72cd8e),
	.w6(32'hbc0d2c02),
	.w7(32'h3c4eec60),
	.w8(32'h3b2bb9d1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5880e),
	.w1(32'h3b9be347),
	.w2(32'hbcd186b6),
	.w3(32'hbc4d2f74),
	.w4(32'h3c5a065c),
	.w5(32'hbc80e7a5),
	.w6(32'hbb214d07),
	.w7(32'h3c64f0e4),
	.w8(32'hbbea0de7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b568),
	.w1(32'hbca033f5),
	.w2(32'h3bbf6f10),
	.w3(32'hbc5ca80d),
	.w4(32'hbbcaf53c),
	.w5(32'h3bb39ad0),
	.w6(32'hbcd6950a),
	.w7(32'h3c1f4c57),
	.w8(32'h3b65547e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b998b),
	.w1(32'hbb90673b),
	.w2(32'hb95b0573),
	.w3(32'h3c1edd50),
	.w4(32'hbbf4fae7),
	.w5(32'h3c1fd46d),
	.w6(32'h3c81c369),
	.w7(32'hbb01165e),
	.w8(32'h3c00f751),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fabfc),
	.w1(32'hbb91ef23),
	.w2(32'hbba97694),
	.w3(32'hbc612750),
	.w4(32'hbada96e1),
	.w5(32'hbaa5e673),
	.w6(32'hbb20f4e4),
	.w7(32'hbae49d98),
	.w8(32'h3bd46c80),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac782bb),
	.w1(32'h3c8fad25),
	.w2(32'h3b5edec2),
	.w3(32'hbbab4f4f),
	.w4(32'h3cacc90f),
	.w5(32'h3c111b52),
	.w6(32'hbbe434f9),
	.w7(32'h3cbc1376),
	.w8(32'h3b205932),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b6c18),
	.w1(32'h3b9ff59f),
	.w2(32'hbb474f44),
	.w3(32'hbc2bb9eb),
	.w4(32'h3c7425f3),
	.w5(32'h3aa9d541),
	.w6(32'hbb9837a3),
	.w7(32'h3b7cf057),
	.w8(32'hbafb2389),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18f2d0),
	.w1(32'h3aaf90f3),
	.w2(32'hbbbe94cc),
	.w3(32'hbc3b0c91),
	.w4(32'hbbe9c445),
	.w5(32'hbb8d5be0),
	.w6(32'h38e5708b),
	.w7(32'h3b0a8ff7),
	.w8(32'hbc85ef8c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb1daf),
	.w1(32'hbbc1c769),
	.w2(32'hba0265eb),
	.w3(32'h3bac9151),
	.w4(32'hbc45224d),
	.w5(32'hb7a28e0e),
	.w6(32'hbb383e81),
	.w7(32'hbb12a8ca),
	.w8(32'h3b5a0e06),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e2f9),
	.w1(32'hbb4c64e5),
	.w2(32'h3b577c17),
	.w3(32'hbaede394),
	.w4(32'hbb1c7398),
	.w5(32'h3bacb3f5),
	.w6(32'h3b94465f),
	.w7(32'hba97ef60),
	.w8(32'h3aa663fc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7387a),
	.w1(32'hbbb09ab7),
	.w2(32'hb9711b89),
	.w3(32'h3ac954cd),
	.w4(32'h3bb4182e),
	.w5(32'h3ad574c8),
	.w6(32'hbb14daa9),
	.w7(32'h3a96b548),
	.w8(32'h39b996e6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1603),
	.w1(32'hba6a339e),
	.w2(32'h3b7ccce3),
	.w3(32'h3acbd30d),
	.w4(32'h3b7fb0ac),
	.w5(32'hbbcb123a),
	.w6(32'h3b66f2a4),
	.w7(32'h3b62a9b2),
	.w8(32'hbbd83b97),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d069f),
	.w1(32'hbb85c5cf),
	.w2(32'hba18bdab),
	.w3(32'h3bf13fec),
	.w4(32'hbc566df5),
	.w5(32'hba4acd17),
	.w6(32'h3bd3be13),
	.w7(32'hbb7baf79),
	.w8(32'hbbc4ef63),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1c66d),
	.w1(32'hb92e8ef8),
	.w2(32'h3b49bce7),
	.w3(32'h3a9dafdc),
	.w4(32'hbc089c10),
	.w5(32'h3beaf7f1),
	.w6(32'h3bd7ee12),
	.w7(32'hbaf93782),
	.w8(32'h3b3f66b3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c366826),
	.w1(32'hbba195bd),
	.w2(32'hba889c13),
	.w3(32'hbb5b536b),
	.w4(32'hbb9e0b35),
	.w5(32'h3a2c30d0),
	.w6(32'h3b36acdc),
	.w7(32'hbc0aec7b),
	.w8(32'hba5d4630),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c8f7),
	.w1(32'hbb92f694),
	.w2(32'h3ab5bb2a),
	.w3(32'h3ac87d40),
	.w4(32'hbbbf2d82),
	.w5(32'h3b117548),
	.w6(32'h3ad17c84),
	.w7(32'hbb026f48),
	.w8(32'h3a6eed0a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bc635),
	.w1(32'hbb1a7f6d),
	.w2(32'h3c4fc25a),
	.w3(32'h39c991dd),
	.w4(32'hbac1a56e),
	.w5(32'h3c38a18f),
	.w6(32'h3a27f867),
	.w7(32'hbb2a0bb9),
	.w8(32'h3be03298),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc7f7b),
	.w1(32'h3c4f4a10),
	.w2(32'h3baa986a),
	.w3(32'hbcf8985a),
	.w4(32'h3c050adb),
	.w5(32'h3b171205),
	.w6(32'hbc9bf656),
	.w7(32'hbba0a1d0),
	.w8(32'hbacc36af),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348531),
	.w1(32'h3b103d96),
	.w2(32'hbbe70a97),
	.w3(32'h3b86683c),
	.w4(32'h3b69204b),
	.w5(32'hbc2bae15),
	.w6(32'hba68940f),
	.w7(32'h3b6328b2),
	.w8(32'hbc235dd5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccae197),
	.w1(32'h3c3fdb87),
	.w2(32'h3a1fe915),
	.w3(32'hbcbebb68),
	.w4(32'h39b5bde6),
	.w5(32'h3c011af1),
	.w6(32'hbc9bde9a),
	.w7(32'h3983a49f),
	.w8(32'h3c52134e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf0504e),
	.w1(32'h3c9d1d34),
	.w2(32'h3aed1477),
	.w3(32'hbd1f16ec),
	.w4(32'h3cd03c66),
	.w5(32'h3bd72fcf),
	.w6(32'hbcd51106),
	.w7(32'h3c76e6b9),
	.w8(32'h3babf5af),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f2c2f),
	.w1(32'hbb32b3f9),
	.w2(32'hbc51d88d),
	.w3(32'hbc72e859),
	.w4(32'h3c18f467),
	.w5(32'hbc376d14),
	.w6(32'hbc68427a),
	.w7(32'h3bdd2a69),
	.w8(32'hbb1e6dd0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c299bf2),
	.w1(32'hbc43e8a4),
	.w2(32'hbb15ceaa),
	.w3(32'h3c927dfd),
	.w4(32'hbb794a9a),
	.w5(32'h3ba280a5),
	.w6(32'h3b506a8c),
	.w7(32'h3bdb8989),
	.w8(32'h3c3092a5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48ff16),
	.w1(32'h3c7bae87),
	.w2(32'hba60c874),
	.w3(32'hbc869672),
	.w4(32'h3c7cd342),
	.w5(32'hbba8ccfe),
	.w6(32'hbcf22af9),
	.w7(32'h3c30ea4b),
	.w8(32'hbc1afa4f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fdc32),
	.w1(32'hbc918ca3),
	.w2(32'h3c40e881),
	.w3(32'h3d09937d),
	.w4(32'hbcd5a007),
	.w5(32'h3bb66677),
	.w6(32'h3d000d55),
	.w7(32'hbc85d8b1),
	.w8(32'h3c543ae1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b488dc8),
	.w1(32'hbaf175b4),
	.w2(32'hbb7b8570),
	.w3(32'h3a697e6e),
	.w4(32'hbab65dcc),
	.w5(32'hbb952b0f),
	.w6(32'h3c271c63),
	.w7(32'hbb057fb4),
	.w8(32'hb9b8421b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c486d),
	.w1(32'h3b5fad34),
	.w2(32'hbb2cb70a),
	.w3(32'hbb7c1c22),
	.w4(32'hb9d565b7),
	.w5(32'hba853ae2),
	.w6(32'hbbe945be),
	.w7(32'hbbaa385e),
	.w8(32'hbb511c4d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf18d77),
	.w1(32'h3b5dc594),
	.w2(32'hbaa5463d),
	.w3(32'h3d176d77),
	.w4(32'hbaf9ee82),
	.w5(32'h3b0279ac),
	.w6(32'h3c985a8f),
	.w7(32'h3b9aff20),
	.w8(32'hb998b717),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934acc),
	.w1(32'hbbe68dd9),
	.w2(32'hbb81878f),
	.w3(32'h3ba23da5),
	.w4(32'hbb3dd8a4),
	.w5(32'h3a8e9a91),
	.w6(32'h3b083518),
	.w7(32'hb95919d6),
	.w8(32'hbb9c6564),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67dcf),
	.w1(32'h3a6bc192),
	.w2(32'hbb7b146f),
	.w3(32'h3a469b77),
	.w4(32'hba66eb8b),
	.w5(32'hbbd94a92),
	.w6(32'hbad9fdec),
	.w7(32'hba929348),
	.w8(32'h3b2dd480),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddb4c8),
	.w1(32'hbadfb48c),
	.w2(32'h3b87025b),
	.w3(32'hbc1d922b),
	.w4(32'h3bc84228),
	.w5(32'h3ab485a5),
	.w6(32'hbba24715),
	.w7(32'h3b429ca7),
	.w8(32'h3b217af8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27067f),
	.w1(32'hbb9c96e0),
	.w2(32'h3b0748b6),
	.w3(32'hbc05191b),
	.w4(32'hbb563383),
	.w5(32'h3b166539),
	.w6(32'hbbad84d5),
	.w7(32'hbbfe6d16),
	.w8(32'h3aa0b814),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac82b34),
	.w1(32'h3a1f799b),
	.w2(32'h3b9acbdb),
	.w3(32'h3b0b1a7b),
	.w4(32'h3a050152),
	.w5(32'h3c1667c5),
	.w6(32'h3a8a3cf0),
	.w7(32'h3a7b8250),
	.w8(32'h3bdfcfbb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c182d6e),
	.w1(32'hbb183323),
	.w2(32'hbad93bb6),
	.w3(32'h3af3f4f5),
	.w4(32'h3949cb17),
	.w5(32'h3b0a62bc),
	.w6(32'h3c2c8102),
	.w7(32'h3b05eb38),
	.w8(32'h3a4a973c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14e976),
	.w1(32'hba0f0e00),
	.w2(32'hbbbc26ee),
	.w3(32'h39af94de),
	.w4(32'h3b13fe2f),
	.w5(32'h3a4e802d),
	.w6(32'h3a9e2a1d),
	.w7(32'h3afb23c4),
	.w8(32'h3b8d444b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60a9f6),
	.w1(32'hbb38f14c),
	.w2(32'hbbceadd3),
	.w3(32'h3c086980),
	.w4(32'h3b7dc860),
	.w5(32'hbb38ad1c),
	.w6(32'h3aa9f79d),
	.w7(32'h3a931465),
	.w8(32'hbb8c50ae),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f4b6),
	.w1(32'h3a972405),
	.w2(32'hbad39cd9),
	.w3(32'h3ae6a30f),
	.w4(32'h3b9b0ed0),
	.w5(32'hbadb21cf),
	.w6(32'h3b89e9aa),
	.w7(32'h3babb54f),
	.w8(32'hbb86047e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ff40c8),
	.w1(32'hbacb10c7),
	.w2(32'hbb2d843f),
	.w3(32'hbb17b46d),
	.w4(32'h3ad600ce),
	.w5(32'hbb01939b),
	.w6(32'h3b7612a5),
	.w7(32'h3ad2c138),
	.w8(32'hbb522aaa),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a04b),
	.w1(32'hbb5e7123),
	.w2(32'h3b6a9f61),
	.w3(32'hbb672adf),
	.w4(32'hbb3bac89),
	.w5(32'h3ab75a43),
	.w6(32'hbb5a28ae),
	.w7(32'hbb2595bf),
	.w8(32'h395710df),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b2263),
	.w1(32'h3a21f13c),
	.w2(32'h3b479fd2),
	.w3(32'h3b91394d),
	.w4(32'hbb224f68),
	.w5(32'h3a99ad3f),
	.w6(32'h3bb7df60),
	.w7(32'h3bcb5103),
	.w8(32'h3a9196a2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe4fe),
	.w1(32'h3a8e5396),
	.w2(32'h3bc71efd),
	.w3(32'hba57325a),
	.w4(32'h3aea017f),
	.w5(32'h3c778787),
	.w6(32'h3b35a66f),
	.w7(32'h3bb2568f),
	.w8(32'h3b1ce01f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d4c82),
	.w1(32'h3a8509ea),
	.w2(32'h3b89295e),
	.w3(32'hbccf1fb6),
	.w4(32'h3c5f119b),
	.w5(32'h3b120eb3),
	.w6(32'hbbb2dac3),
	.w7(32'h3c0b100e),
	.w8(32'h3ad0e3a3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba14c70),
	.w1(32'h3a333371),
	.w2(32'h3a1169ba),
	.w3(32'h3b873bdf),
	.w4(32'hbae12487),
	.w5(32'h3c095168),
	.w6(32'h3940e049),
	.w7(32'h3b66765d),
	.w8(32'h3bd1931c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b931b7c),
	.w1(32'hbbbb8fdb),
	.w2(32'hbbf05c17),
	.w3(32'hbc64e277),
	.w4(32'h3c407f15),
	.w5(32'h3bb1d56f),
	.w6(32'hbb858b1c),
	.w7(32'h3b3a2a6b),
	.w8(32'h3b15b163),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53149),
	.w1(32'hbc41da0a),
	.w2(32'h3b5f7778),
	.w3(32'hbc434576),
	.w4(32'hbb192ebe),
	.w5(32'h3bcbf408),
	.w6(32'hbb700cf1),
	.w7(32'hbaa0bc28),
	.w8(32'h3b7272d3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5da6a),
	.w1(32'h3ad62d7c),
	.w2(32'h3b981271),
	.w3(32'h3be45af1),
	.w4(32'h3afe8346),
	.w5(32'hbb7a91de),
	.w6(32'h3bb05497),
	.w7(32'h3a5ebcbc),
	.w8(32'h3a907d4b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b139e49),
	.w1(32'h3bcdd9a3),
	.w2(32'hb9b1f5d6),
	.w3(32'h3c3f1fe2),
	.w4(32'h3b70efc1),
	.w5(32'hbbfddcff),
	.w6(32'h3bde6ae1),
	.w7(32'h39e1d219),
	.w8(32'hbbb92e38),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1b57a),
	.w1(32'h3a444612),
	.w2(32'hbaeaec54),
	.w3(32'hbc30c746),
	.w4(32'hbc50f86c),
	.w5(32'hbb774865),
	.w6(32'h39aaa904),
	.w7(32'hbc5d8e43),
	.w8(32'hbaa84713),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e7fe3),
	.w1(32'h3b6a3a7c),
	.w2(32'hba996c1e),
	.w3(32'h3c70baf6),
	.w4(32'hbb498a9e),
	.w5(32'hbab38f74),
	.w6(32'h3bf75e60),
	.w7(32'h3b4ff63a),
	.w8(32'hba5d3363),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39b33),
	.w1(32'hb9784a62),
	.w2(32'h3b8202c7),
	.w3(32'hbb240173),
	.w4(32'hb9c508da),
	.w5(32'h3b421666),
	.w6(32'hbb150ada),
	.w7(32'hb974550f),
	.w8(32'hba3a8d29),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9202),
	.w1(32'hbb528376),
	.w2(32'hbbd7e0b6),
	.w3(32'h3a6a492f),
	.w4(32'hbc095f88),
	.w5(32'hbc2aab9b),
	.w6(32'hbb933c19),
	.w7(32'hbc8231ff),
	.w8(32'h3a28ba41),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40805a),
	.w1(32'h3b0f61e9),
	.w2(32'hb930343b),
	.w3(32'hbb904d51),
	.w4(32'hbb926bf6),
	.w5(32'hbaaa1fe8),
	.w6(32'hba0f9f03),
	.w7(32'h3a5ae390),
	.w8(32'hbaf6cd00),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38445095),
	.w1(32'hbae8130c),
	.w2(32'hbbf51a1b),
	.w3(32'hba5d4dc0),
	.w4(32'hba33719c),
	.w5(32'hbc5338ce),
	.w6(32'hbae0dfcb),
	.w7(32'hbb4e4836),
	.w8(32'h39a241aa),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226bb6),
	.w1(32'hbbed234b),
	.w2(32'hbaab6305),
	.w3(32'hbc52d22d),
	.w4(32'hbc7ae6ce),
	.w5(32'hbbaac73d),
	.w6(32'hbc003199),
	.w7(32'hbbeea26d),
	.w8(32'h3ba1f245),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07ab62),
	.w1(32'h3b96409d),
	.w2(32'h3b7a08c7),
	.w3(32'hbc371331),
	.w4(32'hbb7003bf),
	.w5(32'h3acfb29c),
	.w6(32'h3bcf033b),
	.w7(32'h3b47ac2b),
	.w8(32'h39c07351),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9fdfa),
	.w1(32'hbb24c5ce),
	.w2(32'hbbc75b6e),
	.w3(32'h3a91c9b8),
	.w4(32'hbb9ada9e),
	.w5(32'hbbdac0ad),
	.w6(32'h3a48ea4f),
	.w7(32'hbb680436),
	.w8(32'hbc0fa9eb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080813),
	.w1(32'h3c192998),
	.w2(32'h3b2a48bb),
	.w3(32'hbba4a87b),
	.w4(32'h3cce8d7c),
	.w5(32'h3b762316),
	.w6(32'h3c4f13f5),
	.w7(32'h3c77985c),
	.w8(32'h3baa5ce2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b6478),
	.w1(32'h3b1e0492),
	.w2(32'h3ba077e8),
	.w3(32'h3b6dec16),
	.w4(32'h3ac5ea1e),
	.w5(32'h39807efc),
	.w6(32'h3b800314),
	.w7(32'h3b740bfe),
	.w8(32'hbbb46da7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a9af),
	.w1(32'h398ffe9c),
	.w2(32'h396b8233),
	.w3(32'hbbff27b0),
	.w4(32'hbbae76e4),
	.w5(32'hbb4d674e),
	.w6(32'hbc691efd),
	.w7(32'h3c173c7d),
	.w8(32'hbb8b9677),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa60ca5),
	.w1(32'hbb7d6a26),
	.w2(32'hbb938bac),
	.w3(32'hbbb59f12),
	.w4(32'hbb2ae23d),
	.w5(32'hbc27c2c6),
	.w6(32'hbb66e084),
	.w7(32'hbb360808),
	.w8(32'h39cf5172),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12979f),
	.w1(32'hbc088274),
	.w2(32'hbc3dae14),
	.w3(32'hbbe167dc),
	.w4(32'hbb5cf2cf),
	.w5(32'hbc020657),
	.w6(32'h3b16bedd),
	.w7(32'h3b8809c1),
	.w8(32'hb94a4948),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5514a),
	.w1(32'h3beb5710),
	.w2(32'hba982fdb),
	.w3(32'hbc198525),
	.w4(32'h3bbfefe5),
	.w5(32'hb93ca7ae),
	.w6(32'hbc4a60ce),
	.w7(32'h3c00fee2),
	.w8(32'h3b843569),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57cedf),
	.w1(32'hba9c1d20),
	.w2(32'hbb8c902a),
	.w3(32'h3c0be4fe),
	.w4(32'h393442b2),
	.w5(32'hbbd98f0b),
	.w6(32'h3bf36f74),
	.w7(32'h3b1873fb),
	.w8(32'h3ab2648d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a123180),
	.w1(32'h3bad0d77),
	.w2(32'hbba96f85),
	.w3(32'hba8fb961),
	.w4(32'h3bf0d649),
	.w5(32'hbbafb8cf),
	.w6(32'h3b9f51a2),
	.w7(32'h3c76de92),
	.w8(32'hbbead017),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e93bcf),
	.w1(32'h39bccef9),
	.w2(32'hbb5971b2),
	.w3(32'hbac38022),
	.w4(32'hbc489e9f),
	.w5(32'hbb3e7562),
	.w6(32'hba1e13ab),
	.w7(32'hbc071700),
	.w8(32'hbaa061d5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e6e61),
	.w1(32'hba9634a0),
	.w2(32'hbc208fa0),
	.w3(32'hbb71b284),
	.w4(32'hbad27aa7),
	.w5(32'hbbc75349),
	.w6(32'hbab511af),
	.w7(32'h3a51af41),
	.w8(32'hbb9104a5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befcd4a),
	.w1(32'h3c74c0cf),
	.w2(32'hbb9233e4),
	.w3(32'h3c99fb5d),
	.w4(32'h3ccfb888),
	.w5(32'hbbb6b9c5),
	.w6(32'h3c58af71),
	.w7(32'h3c437a46),
	.w8(32'h3b9d4f1e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bdd845),
	.w1(32'h3bdd4ca1),
	.w2(32'hbc367c2a),
	.w3(32'hbb196feb),
	.w4(32'h3bd5c107),
	.w5(32'hbb8fce6c),
	.w6(32'h3c07b78e),
	.w7(32'h3a39e0e3),
	.w8(32'hbc250d44),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13b40c),
	.w1(32'hbb3b4033),
	.w2(32'hbb40f0bd),
	.w3(32'hbbbabe55),
	.w4(32'hbb124680),
	.w5(32'h39cd34cc),
	.w6(32'hbbf3c124),
	.w7(32'hbb5b9ce8),
	.w8(32'h3b836ea8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16f173),
	.w1(32'h3c51b121),
	.w2(32'hb9d6afb3),
	.w3(32'h3bea8591),
	.w4(32'h3c885626),
	.w5(32'h39d31458),
	.w6(32'h3bc1a563),
	.w7(32'h3aed3ca8),
	.w8(32'h3b36d12a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24a93d),
	.w1(32'h3ba5ecb2),
	.w2(32'hbc1ad524),
	.w3(32'h3a892e26),
	.w4(32'h3b8d2783),
	.w5(32'hbc6f0a68),
	.w6(32'h3b455e09),
	.w7(32'h3bcbe301),
	.w8(32'hbbb830cf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99d2c5),
	.w1(32'hbac790f7),
	.w2(32'hbbbd7806),
	.w3(32'hbc2e81ab),
	.w4(32'hbb3f343a),
	.w5(32'hbbf3befd),
	.w6(32'h3a334314),
	.w7(32'hbb553a8b),
	.w8(32'hbc265dcb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ecbd),
	.w1(32'hbb613adf),
	.w2(32'hbc13d246),
	.w3(32'hbc4b446d),
	.w4(32'hbbbd2f81),
	.w5(32'hbc0152a2),
	.w6(32'hba8ca133),
	.w7(32'hb9886255),
	.w8(32'hbc703e18),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc608b59),
	.w1(32'hbb975e90),
	.w2(32'h3ae9c165),
	.w3(32'hbc4036df),
	.w4(32'hbbd03f76),
	.w5(32'h3b319e14),
	.w6(32'hbbdad88f),
	.w7(32'h3a8fc3c7),
	.w8(32'hbab4cb6d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af76986),
	.w1(32'hba0c82fa),
	.w2(32'h3ba79547),
	.w3(32'hbb751f0d),
	.w4(32'h3aff7896),
	.w5(32'h3b910d36),
	.w6(32'hbb593a7f),
	.w7(32'hbb741e34),
	.w8(32'h3b6e9b4e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb23b27),
	.w1(32'h3b2788be),
	.w2(32'hbbe281ec),
	.w3(32'h3b972009),
	.w4(32'h3c16c632),
	.w5(32'hbc6dcf85),
	.w6(32'h3ba18521),
	.w7(32'h3c0acdce),
	.w8(32'hbc14b66e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7f1ab),
	.w1(32'hbc2ee0fe),
	.w2(32'hbc0397ed),
	.w3(32'hbc3a3935),
	.w4(32'hba429a33),
	.w5(32'hbc3e13ed),
	.w6(32'hbc2fad86),
	.w7(32'h3be149ce),
	.w8(32'h3b9b9f42),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04c6a8),
	.w1(32'hbac5a739),
	.w2(32'hbc4c33db),
	.w3(32'hbc04db26),
	.w4(32'h3b89fd7a),
	.w5(32'hbc07ef77),
	.w6(32'h3bc1e3e0),
	.w7(32'h3c2ed619),
	.w8(32'hbbdcd41f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4365f0),
	.w1(32'hba50e243),
	.w2(32'h3b2451b2),
	.w3(32'hbbc62df8),
	.w4(32'hbb808047),
	.w5(32'h3bb6d7be),
	.w6(32'hbb0c68ae),
	.w7(32'h3ba4b053),
	.w8(32'h3ae3f1c0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac51f5c),
	.w1(32'h3bc17f06),
	.w2(32'h3b0b00d6),
	.w3(32'hba4936b5),
	.w4(32'h3c06ddc9),
	.w5(32'h3a65b881),
	.w6(32'hb9f4c2d1),
	.w7(32'h3b01a2d1),
	.w8(32'h3b21021c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac60aba),
	.w1(32'hbbe5e026),
	.w2(32'hbb5c0e6f),
	.w3(32'hbb530382),
	.w4(32'hbc03b24b),
	.w5(32'h3a8021b3),
	.w6(32'hbada9ce3),
	.w7(32'hbbb70e0e),
	.w8(32'hb95b452f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8f47),
	.w1(32'hbb4985df),
	.w2(32'h3b998857),
	.w3(32'hb8e29926),
	.w4(32'hba6841d4),
	.w5(32'h3c23f56a),
	.w6(32'h3b160ad7),
	.w7(32'hbb135685),
	.w8(32'h3c3101ea),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd14a8c),
	.w1(32'h3bb4358a),
	.w2(32'hbbfc1453),
	.w3(32'h3bf4dece),
	.w4(32'h3bdb0cd2),
	.w5(32'hbc8c805f),
	.w6(32'h3b8d15f0),
	.w7(32'h3a8b9bc0),
	.w8(32'hbc184b34),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb5019),
	.w1(32'hbae321dc),
	.w2(32'h3a64246c),
	.w3(32'hbbaa71d6),
	.w4(32'hbb07c929),
	.w5(32'h3bbb59dc),
	.w6(32'hbafc8507),
	.w7(32'hb9e22f9b),
	.w8(32'hba150bbd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14db34),
	.w1(32'h39efaef7),
	.w2(32'h3a12ef99),
	.w3(32'h3b709d9d),
	.w4(32'h3bbd92a2),
	.w5(32'h39e79b7c),
	.w6(32'h3b71948a),
	.w7(32'hbb734ffb),
	.w8(32'hba86b043),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eca23),
	.w1(32'h3ba08ead),
	.w2(32'hba6b63b9),
	.w3(32'hbb8bbe12),
	.w4(32'h3b686669),
	.w5(32'hbb2bcf78),
	.w6(32'hbb526c15),
	.w7(32'h3b937a9b),
	.w8(32'h3b3a7941),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfbc74),
	.w1(32'h3b2d18f4),
	.w2(32'h3a44f5f1),
	.w3(32'h3ba6bdc9),
	.w4(32'hbb2e1df0),
	.w5(32'hba222538),
	.w6(32'hbb86a659),
	.w7(32'hbaf2611f),
	.w8(32'hbab83bc6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931c33e),
	.w1(32'hba8151ab),
	.w2(32'h3ba58534),
	.w3(32'h392174d4),
	.w4(32'h3b3b3db3),
	.w5(32'h3b8b3772),
	.w6(32'h3a2bc225),
	.w7(32'h3ba1b76d),
	.w8(32'h3b904bc0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab5b87),
	.w1(32'h3b89bfa3),
	.w2(32'h39c9c285),
	.w3(32'h3b8f09e1),
	.w4(32'h3b50e891),
	.w5(32'h39caf76f),
	.w6(32'h3b9c0ec5),
	.w7(32'h3b5c6990),
	.w8(32'h399aef9c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26c1e1),
	.w1(32'hbbf679f7),
	.w2(32'h3baf3ab7),
	.w3(32'hba8ff9b5),
	.w4(32'hbba94511),
	.w5(32'h3bdbfb36),
	.w6(32'hbbb4df47),
	.w7(32'hbb9aec10),
	.w8(32'h3c43d6f0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baed594),
	.w1(32'h3b977abe),
	.w2(32'hba3b1a94),
	.w3(32'h3bb413e8),
	.w4(32'hba572b04),
	.w5(32'h3a3daac6),
	.w6(32'h3b88aff0),
	.w7(32'hba135c4d),
	.w8(32'h3a90e330),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842afb7),
	.w1(32'h3af8f63e),
	.w2(32'h3bc6d541),
	.w3(32'h38f1c37c),
	.w4(32'h3b04fad7),
	.w5(32'h3bb02c88),
	.w6(32'h3ac03c57),
	.w7(32'h3afeb642),
	.w8(32'h3be4495f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0eba9),
	.w1(32'h3b1b24d2),
	.w2(32'hba168ba3),
	.w3(32'h3bc63bb3),
	.w4(32'h3aba8d00),
	.w5(32'hbb665224),
	.w6(32'h3bb77446),
	.w7(32'h3b09c58b),
	.w8(32'hbb1b09b2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894097),
	.w1(32'hba8b8125),
	.w2(32'hbbb0752b),
	.w3(32'h3adf7d5a),
	.w4(32'h37a69ec8),
	.w5(32'hba69c33c),
	.w6(32'hbb082926),
	.w7(32'h3a90de66),
	.w8(32'hbb8fd97b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3da3c2),
	.w1(32'h397bade4),
	.w2(32'h396abf5d),
	.w3(32'h3b6923e1),
	.w4(32'hbb5040dc),
	.w5(32'hbbf24f5a),
	.w6(32'hbb59b59a),
	.w7(32'hbb8fbd06),
	.w8(32'hbbe39a94),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abee4f9),
	.w1(32'hbc05d410),
	.w2(32'hbbf22875),
	.w3(32'h399c0475),
	.w4(32'h3aa04f5e),
	.w5(32'hbbe83b93),
	.w6(32'hb92ae34f),
	.w7(32'h3b4be567),
	.w8(32'hbb73d120),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb109d),
	.w1(32'h398cdf5e),
	.w2(32'h3c01768b),
	.w3(32'hbbe7ed36),
	.w4(32'hba16c111),
	.w5(32'h3c0e98dd),
	.w6(32'hbb520168),
	.w7(32'h3b463f9c),
	.w8(32'h3b8ec463),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6579a),
	.w1(32'h3b4c1cfd),
	.w2(32'h3b8a9003),
	.w3(32'h3c02f4d5),
	.w4(32'hbb44c249),
	.w5(32'hbaa6f403),
	.w6(32'h3b8fc597),
	.w7(32'hbafbb221),
	.w8(32'hbb0088bd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6185e3),
	.w1(32'h3c08ce87),
	.w2(32'hbbd70548),
	.w3(32'h3b61d256),
	.w4(32'h3ae7add5),
	.w5(32'h3a066846),
	.w6(32'h3bc20ca2),
	.w7(32'h3b16d164),
	.w8(32'hbc1ba0cc),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddc753),
	.w1(32'hba86376c),
	.w2(32'hbc0c5740),
	.w3(32'hbc34e65b),
	.w4(32'hbb4ade40),
	.w5(32'hbc1ef133),
	.w6(32'hbb8d9078),
	.w7(32'h3ba43012),
	.w8(32'h3918360d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2574f),
	.w1(32'h3b60a67b),
	.w2(32'hb9ae2635),
	.w3(32'hbb8fd8f8),
	.w4(32'h3bb610ee),
	.w5(32'hb99e644d),
	.w6(32'hbc36ecc2),
	.w7(32'h3b82dd07),
	.w8(32'hb90f2919),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c20525),
	.w1(32'h39feb7dc),
	.w2(32'h3bbcd096),
	.w3(32'hbb05c291),
	.w4(32'hb938c5eb),
	.w5(32'h3b73e071),
	.w6(32'hba404b91),
	.w7(32'hba7baade),
	.w8(32'h3b813147),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061f73),
	.w1(32'h3ae9a4c2),
	.w2(32'hb987dacb),
	.w3(32'hb9a52d83),
	.w4(32'h37ae7e11),
	.w5(32'hba73d503),
	.w6(32'h3b656bf1),
	.w7(32'h3b0105b4),
	.w8(32'hba9160de),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65c65a),
	.w1(32'hbb078579),
	.w2(32'h3c44313b),
	.w3(32'hbaf022b2),
	.w4(32'hbb0dc4f6),
	.w5(32'h3b980b9e),
	.w6(32'hbafaab62),
	.w7(32'hbaac72f7),
	.w8(32'h3ac3bfd2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd16849),
	.w1(32'h3c68d5a2),
	.w2(32'hbc216ae4),
	.w3(32'h3b96aa31),
	.w4(32'h3c597a6c),
	.w5(32'hbc9bc178),
	.w6(32'hbb7b8978),
	.w7(32'h3c6560d9),
	.w8(32'hbc0e80af),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbbfb3),
	.w1(32'h3b652d49),
	.w2(32'hbbaa5d84),
	.w3(32'hbb7e7d98),
	.w4(32'h3b702d0a),
	.w5(32'hbc07932c),
	.w6(32'hbb9d6e67),
	.w7(32'h3ac723c1),
	.w8(32'h3a0f1da9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a235a47),
	.w1(32'hbb8f74fc),
	.w2(32'hbbf8dfa5),
	.w3(32'h3ac40b77),
	.w4(32'hbbe3fad5),
	.w5(32'hbc6b1389),
	.w6(32'h3b548a55),
	.w7(32'h3b1834f4),
	.w8(32'hbc04a556),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dff3c),
	.w1(32'h3b629f1f),
	.w2(32'h3b3c9d7a),
	.w3(32'h3a4d3677),
	.w4(32'hbb092384),
	.w5(32'h3b2d95c5),
	.w6(32'h3b235023),
	.w7(32'h3ae74b7e),
	.w8(32'h3b956ecb),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b93ae),
	.w1(32'h3b54d628),
	.w2(32'h3b78e4be),
	.w3(32'h3b1e9258),
	.w4(32'h3b4b3b37),
	.w5(32'h3bb36618),
	.w6(32'h3b05d670),
	.w7(32'h3b93ee3d),
	.w8(32'h3bb4a8ff),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a893ea3),
	.w1(32'h3b146f1a),
	.w2(32'hbb141428),
	.w3(32'h3b6a8304),
	.w4(32'h3b40dedc),
	.w5(32'hbbd00cf7),
	.w6(32'h3b92ff64),
	.w7(32'h3b0492ec),
	.w8(32'hbb5d7372),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc143f29),
	.w1(32'hbba0c473),
	.w2(32'hbc1f5841),
	.w3(32'hbb931e1d),
	.w4(32'hbb6656f7),
	.w5(32'hbc076451),
	.w6(32'hbbad5a3d),
	.w7(32'hbb97efd9),
	.w8(32'hbad53887),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf77fcd),
	.w1(32'hbaf231c0),
	.w2(32'h3bd7d694),
	.w3(32'h36d90ab9),
	.w4(32'h3b9892b5),
	.w5(32'h3c0f011b),
	.w6(32'h378773e8),
	.w7(32'h3bc43a60),
	.w8(32'h3bc835f9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd703),
	.w1(32'h3ad072ff),
	.w2(32'h3c1cdc67),
	.w3(32'h3b5b7b6d),
	.w4(32'h3bcc3622),
	.w5(32'h3c0d5cfd),
	.w6(32'h3b2c4d52),
	.w7(32'h3be74a20),
	.w8(32'h3c253b57),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c029c0a),
	.w1(32'h3c16d3ec),
	.w2(32'h3b1780b4),
	.w3(32'h3bf4508a),
	.w4(32'h3c7007cb),
	.w5(32'h39ab7da6),
	.w6(32'h3bd8a709),
	.w7(32'h3c0f430d),
	.w8(32'h3ab294ca),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea8c4b),
	.w1(32'hb8980bc8),
	.w2(32'h3b27323b),
	.w3(32'h3b0e5f46),
	.w4(32'hb9268aca),
	.w5(32'h3b4cdbe4),
	.w6(32'h3b25a036),
	.w7(32'hbb1b141f),
	.w8(32'h3b91614d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e6338c),
	.w1(32'h3a701755),
	.w2(32'h3afda6d1),
	.w3(32'h3a55b6f9),
	.w4(32'h3b3563b5),
	.w5(32'h3bdf537d),
	.w6(32'h3adf952d),
	.w7(32'h3b00f944),
	.w8(32'h3bf6c4f7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51a591),
	.w1(32'h3bbde67d),
	.w2(32'hbc2cfa05),
	.w3(32'h3c20ecd1),
	.w4(32'h3bf1e408),
	.w5(32'hbac2c432),
	.w6(32'h3c0e6381),
	.w7(32'h3bbfe059),
	.w8(32'h3c2cad05),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c585d),
	.w1(32'h3bf7aa7d),
	.w2(32'h3b7ba2df),
	.w3(32'h3c64f7da),
	.w4(32'h3cbbe882),
	.w5(32'hbae444eb),
	.w6(32'h3cda3eab),
	.w7(32'h3c933494),
	.w8(32'h3b797ce6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c00f),
	.w1(32'h395fcbb9),
	.w2(32'hbb700e8d),
	.w3(32'hbbe62fc6),
	.w4(32'hbbb40121),
	.w5(32'hbaea1edf),
	.w6(32'hba23830d),
	.w7(32'h3ba88796),
	.w8(32'h3b0c7664),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2054a),
	.w1(32'hbb964642),
	.w2(32'hbb91cb24),
	.w3(32'h3bbc4908),
	.w4(32'hbafe6525),
	.w5(32'hbc48ed96),
	.w6(32'h39f5d797),
	.w7(32'h3a8d95c1),
	.w8(32'hbbd871a5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2adf3a),
	.w1(32'hbb311c21),
	.w2(32'h3bc86e99),
	.w3(32'hbc6bede1),
	.w4(32'hbc10ee6b),
	.w5(32'h3bc00cfb),
	.w6(32'hbc174d76),
	.w7(32'hba431dcb),
	.w8(32'h3c09296a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6bdc6),
	.w1(32'h3bd1f9af),
	.w2(32'h3bbc5250),
	.w3(32'h3b4d38c5),
	.w4(32'h3bc62ead),
	.w5(32'h3bfb2aaf),
	.w6(32'h3bb80c95),
	.w7(32'h3bf2d94e),
	.w8(32'h39ecbcc8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eee9e),
	.w1(32'h3b294b77),
	.w2(32'hbb206b03),
	.w3(32'h3bbca8ca),
	.w4(32'hbb81aac8),
	.w5(32'h3b1ca297),
	.w6(32'hbbe30af9),
	.w7(32'hbba037e5),
	.w8(32'h3b9534d1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7704e),
	.w1(32'hbac122bc),
	.w2(32'hbbba0ab0),
	.w3(32'h3bd04e29),
	.w4(32'h3a83e657),
	.w5(32'hbb36ace9),
	.w6(32'h3a8374de),
	.w7(32'h3aba04a4),
	.w8(32'hbc04f69a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94da3bb),
	.w1(32'hbb9be812),
	.w2(32'hbaa821af),
	.w3(32'hba6aea70),
	.w4(32'hbbcc089c),
	.w5(32'h3bbd299f),
	.w6(32'hbaa220f2),
	.w7(32'hbb2bc985),
	.w8(32'h3bca9d52),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97de7d),
	.w1(32'h3bb4e227),
	.w2(32'hbb748109),
	.w3(32'h3bba6eb9),
	.w4(32'h3c2eb18b),
	.w5(32'hbb250da1),
	.w6(32'h3c00eb6d),
	.w7(32'h3c64d0c1),
	.w8(32'h3aa94167),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b0603),
	.w1(32'hbb5af288),
	.w2(32'hba1cf4a9),
	.w3(32'hbc3169c0),
	.w4(32'hbbcbaf02),
	.w5(32'hbb2db63f),
	.w6(32'hbc22d0f3),
	.w7(32'hbb7e98bf),
	.w8(32'hbb3fd1d4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ece9c),
	.w1(32'hbac47ba0),
	.w2(32'h3a14a839),
	.w3(32'hbaabbe99),
	.w4(32'h39332e98),
	.w5(32'h3a0013bf),
	.w6(32'h3a3d681f),
	.w7(32'h3b9126b1),
	.w8(32'h39549e24),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2217d9),
	.w1(32'hb901a925),
	.w2(32'hb8cfcb9c),
	.w3(32'hba34abc3),
	.w4(32'h3a6c60fc),
	.w5(32'h3a2ee821),
	.w6(32'hbaf1bc58),
	.w7(32'h3aebb649),
	.w8(32'hbadaa257),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e850d),
	.w1(32'hbb319874),
	.w2(32'hbb4b1ee1),
	.w3(32'hba18f097),
	.w4(32'hbb63ec16),
	.w5(32'h3a72a45b),
	.w6(32'hbabe4145),
	.w7(32'hbb342585),
	.w8(32'hb94b3ec3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb487dad),
	.w1(32'h38b28f4d),
	.w2(32'hbc1f4fb8),
	.w3(32'hbc00fab7),
	.w4(32'hbb89be32),
	.w5(32'hbc261529),
	.w6(32'hbb9942f9),
	.w7(32'hbbec3219),
	.w8(32'hbc22db10),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc572c9c),
	.w1(32'hbbffab64),
	.w2(32'h3a88a82c),
	.w3(32'hbc28452b),
	.w4(32'hbc7077ef),
	.w5(32'h3bfdb224),
	.w6(32'hbb940e9d),
	.w7(32'hbbb04f05),
	.w8(32'h3a498a77),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab01dc),
	.w1(32'hb9b9b7ea),
	.w2(32'hbb6f5033),
	.w3(32'h3b36ab40),
	.w4(32'h3b9b67fe),
	.w5(32'hbbf77069),
	.w6(32'h3b43e916),
	.w7(32'hbab5600f),
	.w8(32'hbbb47321),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1598d4),
	.w1(32'hbbe81eef),
	.w2(32'h3b83f736),
	.w3(32'hbc1e8cb7),
	.w4(32'hba88dabf),
	.w5(32'h3a16f94a),
	.w6(32'hbbea49f6),
	.w7(32'hbb67e05f),
	.w8(32'h3ac88340),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a203d24),
	.w1(32'h3bab852e),
	.w2(32'hbc81c0e4),
	.w3(32'hbabdb32e),
	.w4(32'h3c11c461),
	.w5(32'hbc3044d6),
	.w6(32'h3c01a3c9),
	.w7(32'h3c749542),
	.w8(32'hbc0d0d7d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009fbc),
	.w1(32'hbc0c8948),
	.w2(32'hbb8a2f02),
	.w3(32'hbc333f2a),
	.w4(32'hbc255a15),
	.w5(32'h3b171e02),
	.w6(32'hbc165354),
	.w7(32'hbc689971),
	.w8(32'h3c2028b3),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0c7d),
	.w1(32'h3bfd3b65),
	.w2(32'h39edb4ec),
	.w3(32'h3c24043d),
	.w4(32'h3c3194f7),
	.w5(32'h3b4ffdba),
	.w6(32'h3c58e126),
	.w7(32'h3c6793be),
	.w8(32'h3bc29ec6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a4fee),
	.w1(32'h3b30c2d3),
	.w2(32'h3bb22a04),
	.w3(32'h3a9e9acc),
	.w4(32'h3b78debc),
	.w5(32'h3b8828c8),
	.w6(32'h3b990242),
	.w7(32'h3b2ba14f),
	.w8(32'hba58f092),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3704273e),
	.w1(32'hbaec07ae),
	.w2(32'h3aeeec4b),
	.w3(32'hbb271c50),
	.w4(32'h3a78fe89),
	.w5(32'h3bc3251a),
	.w6(32'hbb7c44c7),
	.w7(32'hba3335fd),
	.w8(32'h3bc44935),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b0e47),
	.w1(32'h3baa3e25),
	.w2(32'hbbe8a697),
	.w3(32'h3b8be25d),
	.w4(32'h3bbf6b67),
	.w5(32'hbc6b132a),
	.w6(32'h3bc9cfb4),
	.w7(32'h3b574e60),
	.w8(32'hbc04ce96),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc582c94),
	.w1(32'hbbd585d4),
	.w2(32'h3ab76118),
	.w3(32'hbc78bf7a),
	.w4(32'hbc878a43),
	.w5(32'h3b922d9c),
	.w6(32'hbc13b103),
	.w7(32'hbb998dcb),
	.w8(32'hba26f7ac),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829ffa),
	.w1(32'h3bc93ac3),
	.w2(32'h3c609081),
	.w3(32'h3b85a395),
	.w4(32'hbbc5e098),
	.w5(32'h3c61692f),
	.w6(32'h3b4f5708),
	.w7(32'hbc03af43),
	.w8(32'h3bcf4a36),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b991f51),
	.w1(32'h3b8098fb),
	.w2(32'h3a587c31),
	.w3(32'h3b9744b1),
	.w4(32'hba30f8ab),
	.w5(32'h3b41c0d2),
	.w6(32'h3c013e03),
	.w7(32'h3a916d0e),
	.w8(32'h3b14d850),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b1a75),
	.w1(32'h3ab8618d),
	.w2(32'h3a2e9cc1),
	.w3(32'h3b9869ba),
	.w4(32'h3b833f26),
	.w5(32'h3b32a40b),
	.w6(32'h3ba091f9),
	.w7(32'h394e6ea6),
	.w8(32'h3ad0b951),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b188ada),
	.w1(32'h3b4b78a0),
	.w2(32'h3bb7ff68),
	.w3(32'h3b8faa17),
	.w4(32'h3abfdf8a),
	.w5(32'hbbbbb22e),
	.w6(32'h3b167623),
	.w7(32'h3a13c913),
	.w8(32'h3ba31c4d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c795e8c),
	.w1(32'h3c8d905f),
	.w2(32'hbae64d4e),
	.w3(32'h3b8a3296),
	.w4(32'h3c9b0ac4),
	.w5(32'hba40959b),
	.w6(32'h3be1b4d1),
	.w7(32'h3c279fc8),
	.w8(32'h38a7d4c9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb8a5d),
	.w1(32'h3af9e67d),
	.w2(32'hbb8f5a16),
	.w3(32'h3ab5fcdc),
	.w4(32'h3ad398bf),
	.w5(32'hbc093459),
	.w6(32'h3afc4a72),
	.w7(32'hb959a721),
	.w8(32'hbc40ff97),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c9168),
	.w1(32'hbc131810),
	.w2(32'hbaf0ea72),
	.w3(32'hbc605ba5),
	.w4(32'hbc3b3257),
	.w5(32'hbb3fcc91),
	.w6(32'hbbf9aa6e),
	.w7(32'hbb9bf914),
	.w8(32'hbbea37b3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2176b6),
	.w1(32'h3a05ba53),
	.w2(32'hb97e2e9e),
	.w3(32'h3bd8132a),
	.w4(32'hba47467a),
	.w5(32'h3b7e534a),
	.w6(32'h3961a8d1),
	.w7(32'hba4e7ba8),
	.w8(32'h3aa622f9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c591b),
	.w1(32'hbb21392b),
	.w2(32'hbc0f4b1b),
	.w3(32'h3bcc2ddb),
	.w4(32'h3a00e3ce),
	.w5(32'hbbb5fc58),
	.w6(32'h3ad17a7a),
	.w7(32'hba2f4bed),
	.w8(32'hba4c6964),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule