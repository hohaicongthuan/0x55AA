module layer_8_featuremap_224(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0a98e),
	.w1(32'hbbec1331),
	.w2(32'hbc733ec5),
	.w3(32'hbc6a4b27),
	.w4(32'h3be78b39),
	.w5(32'h3c62468c),
	.w6(32'hbc2ec877),
	.w7(32'hbc5c05a8),
	.w8(32'hbc0e0ab3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe8f10),
	.w1(32'hbb0006d9),
	.w2(32'hbace74c3),
	.w3(32'hbb228efa),
	.w4(32'h3b5113ac),
	.w5(32'h3b2ad62a),
	.w6(32'hbbb45d73),
	.w7(32'hbbcdd26c),
	.w8(32'hbbc8999c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ca988),
	.w1(32'hbb3d833b),
	.w2(32'h3bb79bd4),
	.w3(32'h3b50ee80),
	.w4(32'h3c488438),
	.w5(32'h3c6c353c),
	.w6(32'hbae9a8bf),
	.w7(32'hbaa87c23),
	.w8(32'h3a08cfed),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d5cd),
	.w1(32'hbc8da386),
	.w2(32'hbc97c599),
	.w3(32'h3a931cff),
	.w4(32'h3b22e8f5),
	.w5(32'h3afe9a10),
	.w6(32'hbc46d0ea),
	.w7(32'hbcb154ed),
	.w8(32'hbcac5787),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc995389),
	.w1(32'hba138fb8),
	.w2(32'hbba3fa4e),
	.w3(32'hbba7d596),
	.w4(32'h3a1a7850),
	.w5(32'hbbbee052),
	.w6(32'hbb2d6269),
	.w7(32'hbbc1382b),
	.w8(32'hbb828e67),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12bd61),
	.w1(32'h3b03eb6a),
	.w2(32'h3bea94d5),
	.w3(32'hbb23cad2),
	.w4(32'h3c215891),
	.w5(32'h3cea9aff),
	.w6(32'h3bd34731),
	.w7(32'h3a977056),
	.w8(32'hba07a5ca),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26c945),
	.w1(32'hbb4709c3),
	.w2(32'hbb90e3ca),
	.w3(32'h3c8e6f8a),
	.w4(32'hbb74a366),
	.w5(32'hbbc45dc4),
	.w6(32'h3a7989ca),
	.w7(32'hbaf67c18),
	.w8(32'hb93680cc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7222b3),
	.w1(32'h3b2fdb9c),
	.w2(32'hbb78d699),
	.w3(32'hbb00819a),
	.w4(32'h3b1601d2),
	.w5(32'hbba04af9),
	.w6(32'h3bca7e11),
	.w7(32'h3b8f3f80),
	.w8(32'h3bde5432),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3881c),
	.w1(32'hbbb74279),
	.w2(32'hbc1dae38),
	.w3(32'hbc19f240),
	.w4(32'hbc29bfd0),
	.w5(32'hbc61508e),
	.w6(32'hba4c84bd),
	.w7(32'hba229837),
	.w8(32'h3b0d5eed),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361172),
	.w1(32'h3c93efad),
	.w2(32'h3caa9f28),
	.w3(32'h3a191fe3),
	.w4(32'h3c21d545),
	.w5(32'h3c9d51b8),
	.w6(32'hbbd010e7),
	.w7(32'hbad8dec0),
	.w8(32'hbc08b46c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab30c8),
	.w1(32'h3a894eca),
	.w2(32'hbbd15a97),
	.w3(32'hbb82f6a5),
	.w4(32'h3c0b029e),
	.w5(32'h3bb35ae3),
	.w6(32'h3b714629),
	.w7(32'hbb5d5b28),
	.w8(32'hbbab9ce8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3bf8f),
	.w1(32'hbc16fcea),
	.w2(32'hbc3cd182),
	.w3(32'h3b9fff4c),
	.w4(32'h3be0b4d8),
	.w5(32'h3c1dfa3c),
	.w6(32'hbb569233),
	.w7(32'hbbce692f),
	.w8(32'hbb92068a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1fce3),
	.w1(32'hbbbb9118),
	.w2(32'hbaceb149),
	.w3(32'hbafdb858),
	.w4(32'h3c2eff41),
	.w5(32'h3c9e92ee),
	.w6(32'hbc0475af),
	.w7(32'hbc608783),
	.w8(32'hbc3745de),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc067ae3),
	.w1(32'h3bbc88fe),
	.w2(32'h3bf5a68a),
	.w3(32'h3bb1b745),
	.w4(32'h3bc792bc),
	.w5(32'h3c89de9f),
	.w6(32'hbae1e578),
	.w7(32'hbb7dbdc4),
	.w8(32'hbb052456),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf78f4),
	.w1(32'hbb79bce2),
	.w2(32'hbb13a01d),
	.w3(32'h3a6d0d4b),
	.w4(32'hbc0bd050),
	.w5(32'hbbb3b5c2),
	.w6(32'h3b13c6e4),
	.w7(32'h3b7d09ab),
	.w8(32'h3bb206d8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba106e22),
	.w1(32'hbc2dc387),
	.w2(32'h3bf11b91),
	.w3(32'hbb85bfe3),
	.w4(32'hbba0fa08),
	.w5(32'h3c69bfc4),
	.w6(32'hbc27923b),
	.w7(32'h3bdf860f),
	.w8(32'h3c4965c4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c806960),
	.w1(32'hbba8e899),
	.w2(32'hbb1b1639),
	.w3(32'h3c8e5d41),
	.w4(32'h3a8246ce),
	.w5(32'hbbb2cee6),
	.w6(32'hbb0041ca),
	.w7(32'h39a62b3c),
	.w8(32'h3a2cdccb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa6363),
	.w1(32'h3ba2407a),
	.w2(32'h3b726162),
	.w3(32'h3af3d4de),
	.w4(32'h3aaf98a4),
	.w5(32'h3adca9ea),
	.w6(32'h3c300037),
	.w7(32'h3b99b660),
	.w8(32'h3c02cee3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2989b),
	.w1(32'hbc8d772b),
	.w2(32'hbc4a51bb),
	.w3(32'h3c9ab5d3),
	.w4(32'h3af32f6e),
	.w5(32'h3cfe4e1f),
	.w6(32'h3b12c6bb),
	.w7(32'hbbf372a7),
	.w8(32'hba0ec2fc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391faabe),
	.w1(32'hbb6f1b34),
	.w2(32'h3a43db04),
	.w3(32'h3c40c613),
	.w4(32'hbb936c99),
	.w5(32'h3a90d4e5),
	.w6(32'h3b06cbc6),
	.w7(32'h3b986544),
	.w8(32'h3ba95a07),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97626),
	.w1(32'h3bbce20c),
	.w2(32'h3cb61ed6),
	.w3(32'h3b212716),
	.w4(32'h3c72edb9),
	.w5(32'h3c84d31a),
	.w6(32'h3b99dd43),
	.w7(32'hbbc67d6b),
	.w8(32'hbbbfebeb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf96627),
	.w1(32'h3b3bc5c2),
	.w2(32'h3b959bf3),
	.w3(32'h3bf31791),
	.w4(32'h3bf83c2f),
	.w5(32'h3c1ea26b),
	.w6(32'hbbca398c),
	.w7(32'hbacf8f90),
	.w8(32'hba98bf9a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb8543),
	.w1(32'hbc0621f2),
	.w2(32'hbb3dd3fd),
	.w3(32'h3c22c8e3),
	.w4(32'h3c005d76),
	.w5(32'h3cceff6d),
	.w6(32'hba386a85),
	.w7(32'hb6144550),
	.w8(32'hbc6e8742),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d48520),
	.w1(32'h3b11f45d),
	.w2(32'h3ba2de60),
	.w3(32'h3b460bdf),
	.w4(32'hbb1a2219),
	.w5(32'h3a9d7e9e),
	.w6(32'h3b6e7e96),
	.w7(32'h39c4c582),
	.w8(32'h3a2800cf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a631e),
	.w1(32'h3ab69427),
	.w2(32'hbbc0d14a),
	.w3(32'h3b6f8be1),
	.w4(32'h3c140c7c),
	.w5(32'h3c27c675),
	.w6(32'hbc525ca0),
	.w7(32'hbc7d1574),
	.w8(32'hbc7cd995),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68e2d5),
	.w1(32'hb86c13f5),
	.w2(32'h3b97eb19),
	.w3(32'h3c0e8769),
	.w4(32'h394c0548),
	.w5(32'hba33ee3a),
	.w6(32'hbbb2108e),
	.w7(32'h3aca1f13),
	.w8(32'hba3584c3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac095c6),
	.w1(32'hbc4b4ab7),
	.w2(32'hbc225943),
	.w3(32'h3b230297),
	.w4(32'hbaa228df),
	.w5(32'h3b86001b),
	.w6(32'hbc45da22),
	.w7(32'hbcbcdf3c),
	.w8(32'hbca26c54),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc628f5e),
	.w1(32'h3bc18b9f),
	.w2(32'hbc4cc44b),
	.w3(32'h3cd06df1),
	.w4(32'h3c92078b),
	.w5(32'h3b8b0390),
	.w6(32'h3c8d716c),
	.w7(32'h3b87a60d),
	.w8(32'h3c10356c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e89c2),
	.w1(32'hbc0c44da),
	.w2(32'hbb1babfd),
	.w3(32'hba81d003),
	.w4(32'hba3660d1),
	.w5(32'h3bba60f2),
	.w6(32'h3b625aba),
	.w7(32'h3b4beda7),
	.w8(32'hbb361447),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3fde7),
	.w1(32'hbb22cd48),
	.w2(32'hbbea4035),
	.w3(32'h3b869e3b),
	.w4(32'hbb905f25),
	.w5(32'hbb977623),
	.w6(32'hba9cbf36),
	.w7(32'hbb2ea04f),
	.w8(32'hbba4a0bf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9cf9e),
	.w1(32'hbb69d7c7),
	.w2(32'hbbf92524),
	.w3(32'hbaec650b),
	.w4(32'h3aef088d),
	.w5(32'hbabf360e),
	.w6(32'hbc10091a),
	.w7(32'hbc0bbb57),
	.w8(32'hbc3a89b4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fc9f1),
	.w1(32'h390148cb),
	.w2(32'h3c3255b2),
	.w3(32'hbc25af56),
	.w4(32'hbb80f982),
	.w5(32'hbbdd4833),
	.w6(32'h3baa10a3),
	.w7(32'h3c9d82f1),
	.w8(32'h3c914d27),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2ca0d),
	.w1(32'h3be3950e),
	.w2(32'h3b1d73ff),
	.w3(32'hbb433cbf),
	.w4(32'h3c0265a9),
	.w5(32'h3c7f453c),
	.w6(32'hbb1db660),
	.w7(32'hbc00cdb2),
	.w8(32'hbc23ed51),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d590),
	.w1(32'hbb3a58c5),
	.w2(32'hb913d589),
	.w3(32'h3af09ed0),
	.w4(32'hbbc4a3dd),
	.w5(32'hbc059745),
	.w6(32'h39908d0e),
	.w7(32'h3947fd87),
	.w8(32'h3be5361b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1bc81),
	.w1(32'h3a22fe51),
	.w2(32'h3bd7172e),
	.w3(32'hbbafc905),
	.w4(32'hbabc5ca8),
	.w5(32'hb7e7071a),
	.w6(32'hbb4900bd),
	.w7(32'hba82eca9),
	.w8(32'hbb759998),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9321a8),
	.w1(32'hbb56bdf5),
	.w2(32'hbb97a346),
	.w3(32'h3b7200cc),
	.w4(32'hbb287fa8),
	.w5(32'hbb57ce51),
	.w6(32'h3adc3cd2),
	.w7(32'h3bc3044c),
	.w8(32'h3bf7df9f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77b887),
	.w1(32'hbc0bf61c),
	.w2(32'hbc509e2d),
	.w3(32'hbaa91e5b),
	.w4(32'hbaef96b2),
	.w5(32'hbbad8423),
	.w6(32'hbbfd4732),
	.w7(32'hbc0e7d0b),
	.w8(32'hbc1e2ad0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43a5d1),
	.w1(32'hba83df0a),
	.w2(32'hbb4254e7),
	.w3(32'hbba33b96),
	.w4(32'hbbb2c54a),
	.w5(32'hbc34499c),
	.w6(32'h3b93b865),
	.w7(32'h3bc22e96),
	.w8(32'h3bdd23eb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86b3bc),
	.w1(32'hbb7a1f65),
	.w2(32'hbb4d6717),
	.w3(32'hbbc3cdd3),
	.w4(32'hbbf98115),
	.w5(32'h3b4fd69d),
	.w6(32'hbbc8dbf9),
	.w7(32'hbadedce3),
	.w8(32'hbb274fb9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac24e36),
	.w1(32'hbacf50cf),
	.w2(32'hbb0aa4fb),
	.w3(32'hba9d20fc),
	.w4(32'hbb736bb5),
	.w5(32'hbc109c80),
	.w6(32'h389ff174),
	.w7(32'h3b1035c5),
	.w8(32'hbb87bc31),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ec77b),
	.w1(32'hbbd661cb),
	.w2(32'hbb42b040),
	.w3(32'h3b5bfd83),
	.w4(32'h3b5bf9aa),
	.w5(32'h3c0ffdd5),
	.w6(32'h3be39e8b),
	.w7(32'h3c0477fa),
	.w8(32'h3b906382),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2388b),
	.w1(32'hbc0ee204),
	.w2(32'h3a996123),
	.w3(32'hbb2cad5c),
	.w4(32'hbb261269),
	.w5(32'h3c34d675),
	.w6(32'hbc035781),
	.w7(32'hbb45e49f),
	.w8(32'h3a969928),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac04ee),
	.w1(32'hbb984742),
	.w2(32'hbbdaf28c),
	.w3(32'hbab1c653),
	.w4(32'hba014953),
	.w5(32'hbb3fc048),
	.w6(32'hba4c9ab6),
	.w7(32'hbb7d1ab6),
	.w8(32'hbba57517),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30af8),
	.w1(32'h39df6f22),
	.w2(32'h3b2c6851),
	.w3(32'h39bd3c3b),
	.w4(32'hbbdf11c6),
	.w5(32'h3be567ea),
	.w6(32'h3b75c072),
	.w7(32'hba0702c0),
	.w8(32'h3ac4c05e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d3fce),
	.w1(32'h3bd72338),
	.w2(32'h3ba4ca06),
	.w3(32'h3becc4aa),
	.w4(32'h3c01cc8b),
	.w5(32'h3cab6b03),
	.w6(32'h3c307ace),
	.w7(32'h3c1363d0),
	.w8(32'h3b749418),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb322431),
	.w1(32'hbbc7ae08),
	.w2(32'hbbb56217),
	.w3(32'h3c0859fd),
	.w4(32'hbb677815),
	.w5(32'hbb5edce0),
	.w6(32'h3a8e547b),
	.w7(32'hbb6f7a7c),
	.w8(32'h3818757c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0398fa),
	.w1(32'h381ce7b7),
	.w2(32'h3b041bf9),
	.w3(32'hbae74416),
	.w4(32'h3b92661b),
	.w5(32'h3c5a7b21),
	.w6(32'hbb9f7b7a),
	.w7(32'hbc0013ad),
	.w8(32'hbc19342d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27aa82),
	.w1(32'hbc2d79b2),
	.w2(32'h3b144f89),
	.w3(32'h3c214b38),
	.w4(32'h3b4dfc0a),
	.w5(32'h3b15d202),
	.w6(32'h3947117d),
	.w7(32'h3ba8b8c3),
	.w8(32'hbb8d49fb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e51e1),
	.w1(32'hba84cd3e),
	.w2(32'hbac3beb7),
	.w3(32'h3aab2cb0),
	.w4(32'h3c292478),
	.w5(32'h3ca275ba),
	.w6(32'hba958eda),
	.w7(32'hbbc92fda),
	.w8(32'hbb7430ac),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a22d2),
	.w1(32'hbc142b25),
	.w2(32'h3ba0eccd),
	.w3(32'h3bd6c8ef),
	.w4(32'hba95fbc3),
	.w5(32'h3b847ebf),
	.w6(32'h3bb1c5e8),
	.w7(32'h3bcc1cb2),
	.w8(32'hb989cb72),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c295167),
	.w1(32'hbbd8f51c),
	.w2(32'hbc49d7f4),
	.w3(32'hbaece1d7),
	.w4(32'h3b7c04b4),
	.w5(32'h3b90113d),
	.w6(32'h3b0cfca8),
	.w7(32'h3b80343c),
	.w8(32'h3ae62881),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c7978),
	.w1(32'hbc2a1a5e),
	.w2(32'hbba5abe4),
	.w3(32'h3bc5cafc),
	.w4(32'hbb296f92),
	.w5(32'h3c37fdcd),
	.w6(32'h3b8ea78e),
	.w7(32'hbb4b4923),
	.w8(32'hba928640),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61871e),
	.w1(32'hba6d30d0),
	.w2(32'hbbc67250),
	.w3(32'h3bffbcea),
	.w4(32'h3b09fe91),
	.w5(32'hbba236a9),
	.w6(32'h3b0ee0c8),
	.w7(32'h3aa35b74),
	.w8(32'h3a951a8e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919cc6),
	.w1(32'h3ba348fb),
	.w2(32'hbb0b69cc),
	.w3(32'hba3c9b6a),
	.w4(32'h3c080d03),
	.w5(32'h3bdcb8d3),
	.w6(32'h3bc73a49),
	.w7(32'h3bf6b9a6),
	.w8(32'h3b8d2625),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb7090),
	.w1(32'hbb3df36e),
	.w2(32'h3b7e519d),
	.w3(32'h3ab152f8),
	.w4(32'hbc419905),
	.w5(32'h3b308b8f),
	.w6(32'h3afbe268),
	.w7(32'hbbc95703),
	.w8(32'hbb9a5987),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6cbe3),
	.w1(32'hbb450d85),
	.w2(32'hb94f2a42),
	.w3(32'h3c8b9796),
	.w4(32'h3afffcdc),
	.w5(32'h3c585193),
	.w6(32'h3bc8fb09),
	.w7(32'h3ab5991f),
	.w8(32'hbba7d800),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea480),
	.w1(32'hba3dbd35),
	.w2(32'h3ac6fe68),
	.w3(32'h3993ebb9),
	.w4(32'h3c84e450),
	.w5(32'h3bb70f7c),
	.w6(32'hbbce8283),
	.w7(32'hbbb1fad8),
	.w8(32'h3b0ef95f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93c8d3),
	.w1(32'hbb7de1d0),
	.w2(32'hbc282fa4),
	.w3(32'hbb6daec7),
	.w4(32'h3b257231),
	.w5(32'hbb99d10b),
	.w6(32'h3b3702f6),
	.w7(32'hbb84b235),
	.w8(32'hba2fbd28),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa62f8),
	.w1(32'h39d7c004),
	.w2(32'h3a57eaec),
	.w3(32'hb8ec6665),
	.w4(32'h3b57b79c),
	.w5(32'h3b3f66e8),
	.w6(32'hb9c6698a),
	.w7(32'hbb02e08a),
	.w8(32'hbb4d206a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada453b),
	.w1(32'hbaac1e62),
	.w2(32'hbb9228fb),
	.w3(32'h3b3cc7f3),
	.w4(32'hbb87f596),
	.w5(32'h3b3de021),
	.w6(32'h3b0569fc),
	.w7(32'hbb938b59),
	.w8(32'hbbcb75f0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031db0),
	.w1(32'hbb186c81),
	.w2(32'hbb747319),
	.w3(32'h3aba41c9),
	.w4(32'h3c9fe375),
	.w5(32'h3cd9c97b),
	.w6(32'hbba9ac06),
	.w7(32'hbc873c00),
	.w8(32'hbc1609c0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc42f96),
	.w1(32'hbca5d0f9),
	.w2(32'hbce66be7),
	.w3(32'h3c2194f0),
	.w4(32'hbc7d02f5),
	.w5(32'hbc8743f2),
	.w6(32'hbc3c0c6d),
	.w7(32'hbc4c1094),
	.w8(32'hbb79b9e3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb59a6c),
	.w1(32'hbc0e2912),
	.w2(32'hbc5276ca),
	.w3(32'hbb82c0a0),
	.w4(32'hbc459283),
	.w5(32'hbcc1f2be),
	.w6(32'h3c3fc6f8),
	.w7(32'h3cbd35f1),
	.w8(32'h3c9995ae),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb663952),
	.w1(32'hbb229de2),
	.w2(32'h3b051372),
	.w3(32'hbc92e41c),
	.w4(32'h3af01ca5),
	.w5(32'h3c00ecc7),
	.w6(32'hbbc19437),
	.w7(32'hbb2aa475),
	.w8(32'hbb39223e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba281d68),
	.w1(32'hb8e03764),
	.w2(32'h3aa5b19c),
	.w3(32'h3b21e6f3),
	.w4(32'h3b287e2f),
	.w5(32'h3bb4760f),
	.w6(32'h3aae555f),
	.w7(32'h3b6a6358),
	.w8(32'h3b21f61b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392107f3),
	.w1(32'h3994b7ef),
	.w2(32'hbb5af438),
	.w3(32'h3b738fb2),
	.w4(32'hbb3c259d),
	.w5(32'hbadbd77f),
	.w6(32'h3b74e002),
	.w7(32'h3b9bd05e),
	.w8(32'h3b707172),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7b7d0),
	.w1(32'hbc034af2),
	.w2(32'hbc8b7ec4),
	.w3(32'hbb13e8a5),
	.w4(32'h3bad71c0),
	.w5(32'h3c6362b9),
	.w6(32'hbc172277),
	.w7(32'hbc8f405c),
	.w8(32'hbc52d998),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b864),
	.w1(32'hbb03c19d),
	.w2(32'h3ad6ad94),
	.w3(32'h3c900e56),
	.w4(32'h3be8c993),
	.w5(32'h3c84930c),
	.w6(32'hbb0b7af0),
	.w7(32'hbb6b9fad),
	.w8(32'hbbae158b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8ea9f),
	.w1(32'hbaa8bab6),
	.w2(32'h398ab756),
	.w3(32'h3b8bba3d),
	.w4(32'h3b2a2b98),
	.w5(32'h3b908099),
	.w6(32'hbb8df0dd),
	.w7(32'hbaa6333f),
	.w8(32'hbbc22b30),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bf452),
	.w1(32'h3acfcd41),
	.w2(32'h3b972afd),
	.w3(32'h3c32c4c7),
	.w4(32'h3c9a8b53),
	.w5(32'h3c9a0835),
	.w6(32'h3c04187f),
	.w7(32'h3b8997eb),
	.w8(32'hbb0b5feb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9fd9),
	.w1(32'hbbfe530a),
	.w2(32'hbb213838),
	.w3(32'h3c9604ca),
	.w4(32'hbc92209d),
	.w5(32'hbbc44ed1),
	.w6(32'h3c1256f4),
	.w7(32'h3b9e9649),
	.w8(32'h3bec7318),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc19682),
	.w1(32'hbb2280d6),
	.w2(32'hbab8717a),
	.w3(32'h3c114969),
	.w4(32'h3c0e79e2),
	.w5(32'h3c6f6a84),
	.w6(32'hbb951b60),
	.w7(32'hbb3312c1),
	.w8(32'hbbd3da15),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca811),
	.w1(32'hbb77bb33),
	.w2(32'hbb8fd3f0),
	.w3(32'h3bac5a01),
	.w4(32'h39adda56),
	.w5(32'h3c7de4d9),
	.w6(32'hbc34a1f0),
	.w7(32'hbb5fdbc6),
	.w8(32'hb943cd79),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a498db5),
	.w1(32'h3abff9df),
	.w2(32'hbb8e5d8d),
	.w3(32'h3bd16ce9),
	.w4(32'h3a6d4a6f),
	.w5(32'hbaf2023b),
	.w6(32'hbaf61b9d),
	.w7(32'hbbd226b4),
	.w8(32'hbbc1d82f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967b08),
	.w1(32'hbc5568c6),
	.w2(32'hbc8a90a2),
	.w3(32'hbae8992b),
	.w4(32'hbc0a6134),
	.w5(32'hbaf00f30),
	.w6(32'hbc64b84f),
	.w7(32'hbca2d9f4),
	.w8(32'hbc56512f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f11c4),
	.w1(32'hbac456ce),
	.w2(32'h3b040309),
	.w3(32'h3b8c370c),
	.w4(32'hbb48a5f3),
	.w5(32'hbb4bf4c1),
	.w6(32'h3b2ce0f0),
	.w7(32'h3be99f0f),
	.w8(32'h3bf5b7ea),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892b78d),
	.w1(32'hb973f3dd),
	.w2(32'hbb34a9ff),
	.w3(32'hbaab0d9d),
	.w4(32'h3b7758c0),
	.w5(32'h3bb4f600),
	.w6(32'hbbc759af),
	.w7(32'hbbebb300),
	.w8(32'hbbaeb93c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c47cf),
	.w1(32'hbb56fe19),
	.w2(32'hbbd5e333),
	.w3(32'h3ad0d8b4),
	.w4(32'h3c45e486),
	.w5(32'h3c1bd3d6),
	.w6(32'hbc087060),
	.w7(32'hbc0b6db2),
	.w8(32'hbc338afd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff2bb),
	.w1(32'h385c0c60),
	.w2(32'h3c3591f8),
	.w3(32'hbaf8ebe3),
	.w4(32'h3c31a1ea),
	.w5(32'h3cb22ffc),
	.w6(32'hb95a57c8),
	.w7(32'hbbb82eef),
	.w8(32'hbc3dbd98),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac02a3c),
	.w1(32'h3b2101f3),
	.w2(32'hba380114),
	.w3(32'h3bc250ad),
	.w4(32'hba789f5e),
	.w5(32'h3b464f91),
	.w6(32'h3bb628f0),
	.w7(32'h3a0e72d6),
	.w8(32'hbbcdcdaa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be335ca),
	.w1(32'h3b85ef69),
	.w2(32'h3c1f5d5b),
	.w3(32'hbad11027),
	.w4(32'h3c1e8125),
	.w5(32'h3cc50ad0),
	.w6(32'hbc22b2b5),
	.w7(32'hba952825),
	.w8(32'hbb811316),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5c811),
	.w1(32'h3b865007),
	.w2(32'hbad388ab),
	.w3(32'h3c3b3bce),
	.w4(32'hbae47af3),
	.w5(32'h39c5499b),
	.w6(32'hba1e429f),
	.w7(32'h3b07bc9e),
	.w8(32'h3bb5cd73),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6ff08),
	.w1(32'hbc1218e5),
	.w2(32'h3b2013a3),
	.w3(32'hb9b47d55),
	.w4(32'h39283876),
	.w5(32'h3c4f3e5d),
	.w6(32'h3bc19ff1),
	.w7(32'h3bfa6dc7),
	.w8(32'h3c607270),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54255e),
	.w1(32'hbc98890a),
	.w2(32'hbcb0a33d),
	.w3(32'hbb1cd1e7),
	.w4(32'hbc850ab9),
	.w5(32'hbb67e2fb),
	.w6(32'hbb2192bc),
	.w7(32'hbc3e41d6),
	.w8(32'hbc72324a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20ab3b),
	.w1(32'h3b252890),
	.w2(32'h3abc8b53),
	.w3(32'h3c3930c3),
	.w4(32'h3c518f12),
	.w5(32'h3ca72e6f),
	.w6(32'h3b0d35c8),
	.w7(32'hbb46c620),
	.w8(32'h3a8eba3a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bf082),
	.w1(32'hbbf5a959),
	.w2(32'h3bd079d6),
	.w3(32'h3c3806db),
	.w4(32'h3a939c7f),
	.w5(32'h3c123403),
	.w6(32'hbb81b255),
	.w7(32'hbc46b42d),
	.w8(32'hbbcae616),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11181c),
	.w1(32'h3c3fd13c),
	.w2(32'h3c670774),
	.w3(32'h3bba4eb5),
	.w4(32'hbac0696c),
	.w5(32'hba86cb1c),
	.w6(32'h3c1ecf4f),
	.w7(32'h3c68366b),
	.w8(32'h3c0f6024),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39d032),
	.w1(32'h3b5d65de),
	.w2(32'h3bd9868e),
	.w3(32'hbbdf43ce),
	.w4(32'hba338b2e),
	.w5(32'h3ba3e82b),
	.w6(32'hbba1c6f5),
	.w7(32'hbb67e0de),
	.w8(32'hbae1cb00),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3da4a),
	.w1(32'hbb6a776e),
	.w2(32'h39cb17a9),
	.w3(32'h3b9cc319),
	.w4(32'h3b77e1d4),
	.w5(32'h3b979416),
	.w6(32'hbb64624f),
	.w7(32'hba227c5f),
	.w8(32'hbb75911c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3c92),
	.w1(32'h3ac75889),
	.w2(32'h3c24df6b),
	.w3(32'hbb6acb6c),
	.w4(32'h3c7fa58c),
	.w5(32'h3c798ef1),
	.w6(32'hbc180007),
	.w7(32'hbba3ca3c),
	.w8(32'hbbe95b1e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26333),
	.w1(32'hbb675dbf),
	.w2(32'h3bb3bbc4),
	.w3(32'h3b379dd4),
	.w4(32'h3b1921db),
	.w5(32'h3aadcf5e),
	.w6(32'hbbdd8733),
	.w7(32'h3ad0c883),
	.w8(32'hbad7fd48),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70cac2),
	.w1(32'hbbcbac18),
	.w2(32'hbafaee45),
	.w3(32'hba98ffe4),
	.w4(32'hbbd2ff9d),
	.w5(32'hbc11ed5a),
	.w6(32'hba9d9e45),
	.w7(32'hba421bca),
	.w8(32'h3b2b11e7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90bc3f),
	.w1(32'hbb0c1073),
	.w2(32'hbb0e5b08),
	.w3(32'hba58d60c),
	.w4(32'hbb0bd040),
	.w5(32'hbb7966a4),
	.w6(32'hbb057e01),
	.w7(32'hbb7a76f7),
	.w8(32'hbb7ffcf8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3838),
	.w1(32'hb9fcfe71),
	.w2(32'h3afb76d9),
	.w3(32'hbb4aa154),
	.w4(32'h3bc6ab9c),
	.w5(32'h3c351740),
	.w6(32'hba9abddd),
	.w7(32'hbb918d99),
	.w8(32'hbb64742e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab10386),
	.w1(32'hbafe7c3f),
	.w2(32'hbb2e9c3e),
	.w3(32'h3bfb089c),
	.w4(32'hbbcd3a2f),
	.w5(32'h3b015064),
	.w6(32'h3b0addb1),
	.w7(32'h3b4e74a1),
	.w8(32'h38f1f41a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ba3cc),
	.w1(32'h3b7648d6),
	.w2(32'h3aea84ea),
	.w3(32'h3bb98ef2),
	.w4(32'h3ab4c041),
	.w5(32'hba318527),
	.w6(32'h3bd8aef0),
	.w7(32'h3ba4e64d),
	.w8(32'h3af6a8f3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc3c1),
	.w1(32'h3a0dfc46),
	.w2(32'h3a8f17e5),
	.w3(32'hbbdbadbd),
	.w4(32'h3b0fc835),
	.w5(32'h3bfa5e31),
	.w6(32'hb80b5fa9),
	.w7(32'h3c00d997),
	.w8(32'h3bb5e556),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba262ffb),
	.w1(32'hbb64c188),
	.w2(32'h3a0959cc),
	.w3(32'h3c10cc83),
	.w4(32'hbb2ddcab),
	.w5(32'h3b5849ac),
	.w6(32'hbab4d085),
	.w7(32'h3acd967b),
	.w8(32'h3bc8da4a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3785cce1),
	.w1(32'hbbbf603a),
	.w2(32'hb9afc29c),
	.w3(32'h3a8e5aa9),
	.w4(32'hbaa3d5c5),
	.w5(32'h3c0b5b17),
	.w6(32'hbb4764c1),
	.w7(32'hbae1de6f),
	.w8(32'hbac84d1f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57371f),
	.w1(32'h398cf4a0),
	.w2(32'hbbcdfa3d),
	.w3(32'h3aaef1ff),
	.w4(32'h3c439503),
	.w5(32'h3b914bd9),
	.w6(32'hbb33bbda),
	.w7(32'hbc37e0b1),
	.w8(32'hbca4348f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafccbb),
	.w1(32'h3c2ec35c),
	.w2(32'h3bcf0e2f),
	.w3(32'h3b92da1a),
	.w4(32'h3c224a7b),
	.w5(32'h3c3a1cd9),
	.w6(32'h3c33c2ff),
	.w7(32'hbb900bb3),
	.w8(32'hbc868ece),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39088cab),
	.w1(32'h39ee84b9),
	.w2(32'hbc127166),
	.w3(32'h3b38d253),
	.w4(32'h3b8cf02c),
	.w5(32'h3933322e),
	.w6(32'hbb2c7421),
	.w7(32'hbc0aa064),
	.w8(32'hbc5ed391),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51d5f1),
	.w1(32'h3b05c6f2),
	.w2(32'h3ab8fb52),
	.w3(32'h3a16d25a),
	.w4(32'h3b1efe75),
	.w5(32'h3c2bddfa),
	.w6(32'h3a4ddb96),
	.w7(32'h3b099ec1),
	.w8(32'h3c068b3a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a7fb5),
	.w1(32'h3c58ad7f),
	.w2(32'h3c118f7e),
	.w3(32'h3c0c6429),
	.w4(32'h3c2e7ca4),
	.w5(32'h3a85068b),
	.w6(32'hba3a1dc9),
	.w7(32'hbb3e35d3),
	.w8(32'hbba8a9ef),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e0a81),
	.w1(32'hbbdeca18),
	.w2(32'hbc4b25ac),
	.w3(32'hbc4815a9),
	.w4(32'h3b195a69),
	.w5(32'h3b290ccb),
	.w6(32'hbbc4d754),
	.w7(32'hbb620e76),
	.w8(32'h3ba681e7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc6b5),
	.w1(32'hbbe148e0),
	.w2(32'hbc02d307),
	.w3(32'h3c76a75f),
	.w4(32'hbbd17146),
	.w5(32'hbc16e1b1),
	.w6(32'h3bcb0364),
	.w7(32'h3aeca841),
	.w8(32'h3b4e756d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacc475),
	.w1(32'h3c04bf08),
	.w2(32'h3c9cc8d2),
	.w3(32'hbbd02508),
	.w4(32'h3c1c1ca7),
	.w5(32'h3c7a77ca),
	.w6(32'hbc008bb0),
	.w7(32'hbbb8bf8f),
	.w8(32'hbbd55490),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e707a),
	.w1(32'hbc46ee8d),
	.w2(32'hbc86d18f),
	.w3(32'h3b95d04e),
	.w4(32'hbbc904bf),
	.w5(32'hbbd2e113),
	.w6(32'hbc4845d2),
	.w7(32'hbc530e3d),
	.w8(32'hbc8a3b25),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e906f),
	.w1(32'hbb7fe0fd),
	.w2(32'hbc78326e),
	.w3(32'h39de9287),
	.w4(32'hbc7d40b9),
	.w5(32'hbcda5a5a),
	.w6(32'h3be8cbad),
	.w7(32'h3c03a914),
	.w8(32'h3b9aee48),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0869),
	.w1(32'h3a9724f2),
	.w2(32'h3a06a8f4),
	.w3(32'hbc7f67c2),
	.w4(32'h3b1c6675),
	.w5(32'hba5a2692),
	.w6(32'h3abae373),
	.w7(32'h3b46bc8e),
	.w8(32'h3aebeee9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a794e6e),
	.w1(32'hbb8b230a),
	.w2(32'h3b4dc63c),
	.w3(32'h3b2353c0),
	.w4(32'h392f9d54),
	.w5(32'h3bcc94cf),
	.w6(32'hbb0f7338),
	.w7(32'h3b58a6c6),
	.w8(32'hb82dc61a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6df17),
	.w1(32'hbb5ceff6),
	.w2(32'hbaaad10e),
	.w3(32'h3b36b9aa),
	.w4(32'h3b83e9d8),
	.w5(32'h3c3abed8),
	.w6(32'hbb84d0c8),
	.w7(32'hbb83ed53),
	.w8(32'hbb70be8d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245db6),
	.w1(32'hbae6eec0),
	.w2(32'h3b021d41),
	.w3(32'h3b8cbd96),
	.w4(32'h3bb36098),
	.w5(32'h3b4a97f0),
	.w6(32'hbb77b296),
	.w7(32'hb9a54a32),
	.w8(32'h3af0b92d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e3492),
	.w1(32'h3ba6e9c5),
	.w2(32'h3b0ee482),
	.w3(32'hbb1ab61a),
	.w4(32'h3b01ea5b),
	.w5(32'h3c264385),
	.w6(32'hbba8d5a1),
	.w7(32'hbc1e3a18),
	.w8(32'hbc4643a0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3931f6f4),
	.w1(32'hbbd71cc8),
	.w2(32'hbb9e8476),
	.w3(32'h3b26e4a0),
	.w4(32'hbb3460f3),
	.w5(32'h3b3dea3c),
	.w6(32'hbb9958f7),
	.w7(32'hbb8e5dc4),
	.w8(32'hbb871ebd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2e55c),
	.w1(32'h3af89506),
	.w2(32'h3b193f63),
	.w3(32'hbb89ac5e),
	.w4(32'h3b7d7ee9),
	.w5(32'h3b29458f),
	.w6(32'h3ae6feb6),
	.w7(32'h3b8bf8a7),
	.w8(32'h3ac7e433),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96d0da),
	.w1(32'h3b0b1886),
	.w2(32'h39ebe056),
	.w3(32'h39f2b872),
	.w4(32'hbb7e5fce),
	.w5(32'h3b234e30),
	.w6(32'h3b9ffafe),
	.w7(32'h3abbe7bd),
	.w8(32'h3b5bb9bb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95216aa),
	.w1(32'h3a22a3a4),
	.w2(32'hbb46dc55),
	.w3(32'h3c197a8f),
	.w4(32'h3a0f2173),
	.w5(32'h3aee4302),
	.w6(32'h3b384d4b),
	.w7(32'h3ba58b7f),
	.w8(32'hbaa25ee0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e848d0),
	.w1(32'h3bf7ef4e),
	.w2(32'hbba5092a),
	.w3(32'h3b9c1af1),
	.w4(32'h3c79e13e),
	.w5(32'h3cad3771),
	.w6(32'hbb47eb7c),
	.w7(32'hbc1730bc),
	.w8(32'hbc0b3ad3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d87f7),
	.w1(32'hba1285fc),
	.w2(32'hbb47cd1a),
	.w3(32'hbb34b972),
	.w4(32'hba19d3a6),
	.w5(32'hb995ed4b),
	.w6(32'hbafbe3e6),
	.w7(32'hba0604e6),
	.w8(32'hb7b44cff),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb14866),
	.w1(32'h3aa321c4),
	.w2(32'h3b24502e),
	.w3(32'h3b4018e1),
	.w4(32'hbc221d6b),
	.w5(32'hbafda952),
	.w6(32'h3bc54a83),
	.w7(32'hbb6a0167),
	.w8(32'hbb7c8003),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8de0af),
	.w1(32'h3bb86230),
	.w2(32'h3c4469df),
	.w3(32'hbb64f064),
	.w4(32'h3c05cd02),
	.w5(32'h3c9af341),
	.w6(32'hba5e2daa),
	.w7(32'hbb089657),
	.w8(32'hbb186474),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2245c1),
	.w1(32'h3b64e9b4),
	.w2(32'h3a652ba0),
	.w3(32'h3c0ee371),
	.w4(32'h3b9cbf08),
	.w5(32'h3bb22dbf),
	.w6(32'hba518c2a),
	.w7(32'hbb0046e8),
	.w8(32'hbb14a2d8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf1982),
	.w1(32'h3aa836de),
	.w2(32'h3b935c84),
	.w3(32'h3b75803d),
	.w4(32'h3a86b91d),
	.w5(32'h3c0235de),
	.w6(32'h3a433905),
	.w7(32'h3a8ce9a1),
	.w8(32'hba889dda),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11bdf1),
	.w1(32'hba7ee45d),
	.w2(32'hbbb4baba),
	.w3(32'h3b104d61),
	.w4(32'hbc015492),
	.w5(32'hbbab0bf3),
	.w6(32'h3adfb746),
	.w7(32'h3995a41f),
	.w8(32'h39ac0c30),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17776a),
	.w1(32'h38ec61d5),
	.w2(32'h3b78239e),
	.w3(32'hbbacedbc),
	.w4(32'hbb0a793d),
	.w5(32'hbb0580ad),
	.w6(32'h39133940),
	.w7(32'h3821b56d),
	.w8(32'hbb78bb56),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74aed6),
	.w1(32'hbac3b03e),
	.w2(32'hbb2ad4f6),
	.w3(32'hbae2ca34),
	.w4(32'h3a235b7e),
	.w5(32'hb98b3a95),
	.w6(32'h3a0928da),
	.w7(32'h3a0552ad),
	.w8(32'h3a4bad92),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5300),
	.w1(32'h37a1e652),
	.w2(32'hb95624c9),
	.w3(32'h3b556e60),
	.w4(32'h3b8a9ec0),
	.w5(32'h3b17bf5d),
	.w6(32'h3a5b5ddc),
	.w7(32'hb9e881e5),
	.w8(32'hbb0af32b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule