module layer_10_featuremap_156(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363cf6f7),
	.w1(32'h3677cac7),
	.w2(32'h36d96566),
	.w3(32'h36798ad3),
	.w4(32'h365ed848),
	.w5(32'h36886a7f),
	.w6(32'h35f288b3),
	.w7(32'h369683b6),
	.w8(32'h3681fef9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a200677),
	.w1(32'h3a1440d7),
	.w2(32'h39e0ceac),
	.w3(32'h3a184228),
	.w4(32'h3a0d3cc6),
	.w5(32'h39b810c6),
	.w6(32'h39924898),
	.w7(32'h39cd9efd),
	.w8(32'h3943b007),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64c3b66),
	.w1(32'hb4104f45),
	.w2(32'hb42492b7),
	.w3(32'hb65b5874),
	.w4(32'hb5d039e7),
	.w5(32'h3534c4db),
	.w6(32'hb6077367),
	.w7(32'hb5607985),
	.w8(32'hb507e773),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8719e),
	.w1(32'hb9df163c),
	.w2(32'hb9e7ff05),
	.w3(32'hb9918a99),
	.w4(32'hb9e24f9f),
	.w5(32'hb99207e8),
	.w6(32'hb95fbc08),
	.w7(32'hb98a5266),
	.w8(32'hb9643366),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f77682),
	.w1(32'hb7ce61ef),
	.w2(32'hb78d1cd0),
	.w3(32'hb7d6bee5),
	.w4(32'hb7de91d7),
	.w5(32'hb793364b),
	.w6(32'hb7bee1bd),
	.w7(32'hb79801a6),
	.w8(32'hb79e4a29),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b2e0e1),
	.w1(32'hb6ac98e2),
	.w2(32'hb6ae470b),
	.w3(32'hb7176c6c),
	.w4(32'hb7010c1b),
	.w5(32'hb6e3121f),
	.w6(32'hb669aafe),
	.w7(32'hb6425692),
	.w8(32'hb62d7c2e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bedd58),
	.w1(32'hb76bf776),
	.w2(32'hb82619ae),
	.w3(32'hb7f4a850),
	.w4(32'hb79c6c00),
	.w5(32'hb780ea7f),
	.w6(32'hb78a83b9),
	.w7(32'hb7193a0b),
	.w8(32'hb71b9a22),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c0aab),
	.w1(32'hb9948f13),
	.w2(32'h38081852),
	.w3(32'h39211d96),
	.w4(32'h38ea375a),
	.w5(32'h3772cf9f),
	.w6(32'h3992859a),
	.w7(32'h37a57dbd),
	.w8(32'hb9073e04),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396259ba),
	.w1(32'h398b95e8),
	.w2(32'h3943d586),
	.w3(32'h39900189),
	.w4(32'h39dd1d3e),
	.w5(32'h395367d8),
	.w6(32'h39195f54),
	.w7(32'h3934e933),
	.w8(32'h391ea26b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1def),
	.w1(32'hbbb23406),
	.w2(32'hbbbe15d4),
	.w3(32'hbb884e50),
	.w4(32'hbb9609ab),
	.w5(32'hbb801baa),
	.w6(32'hbb3cd593),
	.w7(32'hbb35219b),
	.w8(32'hbb165908),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b14f16),
	.w1(32'hb92a9988),
	.w2(32'hb9804515),
	.w3(32'hb76851b6),
	.w4(32'h37861847),
	.w5(32'hb8dc70da),
	.w6(32'h38cb6367),
	.w7(32'h3718a48c),
	.w8(32'hb86a1df9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d73b),
	.w1(32'h3a82f3f8),
	.w2(32'h3a73af9d),
	.w3(32'h3a4cd0ca),
	.w4(32'h3a1e989f),
	.w5(32'h3a0e1e25),
	.w6(32'h3a016193),
	.w7(32'h3a175d19),
	.w8(32'h39e7b52a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866101),
	.w1(32'hbb854a58),
	.w2(32'hbb804490),
	.w3(32'hbb719a72),
	.w4(32'hbb9303bc),
	.w5(32'hbb5c0a22),
	.w6(32'hbb38b0e6),
	.w7(32'hbb43d701),
	.w8(32'hbb02207c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c092),
	.w1(32'hbac01f6f),
	.w2(32'hbaccd928),
	.w3(32'hba9fba6b),
	.w4(32'hba966746),
	.w5(32'hba9f97c8),
	.w6(32'hba919995),
	.w7(32'hba92e76c),
	.w8(32'hba88b7b0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983e1fc),
	.w1(32'hb9c05750),
	.w2(32'hba31094d),
	.w3(32'hb99d6c9c),
	.w4(32'hb985e5b6),
	.w5(32'hb9478ecb),
	.w6(32'hb8230fb1),
	.w7(32'h39c6772c),
	.w8(32'h39c88002),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2443c4),
	.w1(32'hbb2f934b),
	.w2(32'hbb370de0),
	.w3(32'hbb05880f),
	.w4(32'hbb20263e),
	.w5(32'hbb117550),
	.w6(32'hbab7eb48),
	.w7(32'hba95cb76),
	.w8(32'hbaa652f8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39667721),
	.w1(32'hb83e0a92),
	.w2(32'hb9fb2c48),
	.w3(32'h38a1fbf2),
	.w4(32'hb9335050),
	.w5(32'hb9cb96e0),
	.w6(32'h378899c6),
	.w7(32'hb9b79368),
	.w8(32'hb9ee9710),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a3a3),
	.w1(32'hbae3b271),
	.w2(32'hbb0c7aa3),
	.w3(32'hbadb5cd7),
	.w4(32'hbacad51a),
	.w5(32'hbabd2d00),
	.w6(32'hba80c6c9),
	.w7(32'hba70012c),
	.w8(32'hbaa3b8ed),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bbd39),
	.w1(32'hbb128251),
	.w2(32'hbb1382d0),
	.w3(32'hbaf52f39),
	.w4(32'hbaf8220c),
	.w5(32'hbade7411),
	.w6(32'hba75a1e6),
	.w7(32'hba56a98c),
	.w8(32'hba731aa6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e1369b),
	.w1(32'h372171cc),
	.w2(32'h3706d756),
	.w3(32'h36c9e992),
	.w4(32'h3761a221),
	.w5(32'h372f9c89),
	.w6(32'h3692d911),
	.w7(32'h372b0da1),
	.w8(32'h37156a2b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5dbfe80),
	.w1(32'h3634c93e),
	.w2(32'h36923a4e),
	.w3(32'hb556ab4d),
	.w4(32'h35473c5d),
	.w5(32'h364edbf2),
	.w6(32'h35e2edf5),
	.w7(32'h36a48744),
	.w8(32'h36dab042),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b3c35),
	.w1(32'h3a0218e1),
	.w2(32'h3a0371e0),
	.w3(32'h3990c8ed),
	.w4(32'h3988afdf),
	.w5(32'h39731bd4),
	.w6(32'h38d74de7),
	.w7(32'h39666257),
	.w8(32'h394d2054),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa58af6),
	.w1(32'hbb09f430),
	.w2(32'hbb00be03),
	.w3(32'hbb07cfd9),
	.w4(32'hbb21d534),
	.w5(32'hbaf13848),
	.w6(32'hba925c8d),
	.w7(32'hbac88728),
	.w8(32'hbac0e73c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dc97d),
	.w1(32'hbb3ae413),
	.w2(32'hbb404b9e),
	.w3(32'hbafb77d2),
	.w4(32'hbb0f6e7a),
	.w5(32'hbb017e9a),
	.w6(32'hbac69ec3),
	.w7(32'hbad3c418),
	.w8(32'hbabfea7b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887412d),
	.w1(32'h398e82a5),
	.w2(32'h383ed449),
	.w3(32'h3989e4df),
	.w4(32'h39d15397),
	.w5(32'h38aa5606),
	.w6(32'h38fcfa43),
	.w7(32'h3985aedb),
	.w8(32'h39395f73),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba417a6f),
	.w1(32'hbaaddd0f),
	.w2(32'hba969eb6),
	.w3(32'hba07d540),
	.w4(32'hba9c5802),
	.w5(32'hba308069),
	.w6(32'hb9b060a9),
	.w7(32'hba0931fd),
	.w8(32'hb941531b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383b035c),
	.w1(32'h38917e86),
	.w2(32'h38a2dade),
	.w3(32'h37f00493),
	.w4(32'h38599b6d),
	.w5(32'h38873292),
	.w6(32'h37ea81e7),
	.w7(32'h385678cd),
	.w8(32'h3883f121),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7891644),
	.w1(32'h3949944f),
	.w2(32'h3916b14d),
	.w3(32'hb8e156b4),
	.w4(32'h3942248b),
	.w5(32'h38a8e61c),
	.w6(32'h37394181),
	.w7(32'h397c1e5e),
	.w8(32'h394964b2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a084bc8),
	.w1(32'h3a18ac3e),
	.w2(32'h3a30b4ba),
	.w3(32'h39a05d3b),
	.w4(32'h395ec20a),
	.w5(32'h3994ba29),
	.w6(32'hb8d92dc5),
	.w7(32'h38dbed4a),
	.w8(32'h393fad7f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68e010),
	.w1(32'hbb8bfedc),
	.w2(32'hbb901a5f),
	.w3(32'hbb42c8d9),
	.w4(32'hbb6f3758),
	.w5(32'hbb4621b3),
	.w6(32'hbb17fc8d),
	.w7(32'hbb213c20),
	.w8(32'hbb011123),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34226ccb),
	.w1(32'hb65c7a07),
	.w2(32'hb7a0ea64),
	.w3(32'h36824c7c),
	.w4(32'h33391546),
	.w5(32'hb7813e92),
	.w6(32'h3559d212),
	.w7(32'hb6d70924),
	.w8(32'hb7895d3e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388dd28b),
	.w1(32'h38200c49),
	.w2(32'hb76bb6d4),
	.w3(32'h38790916),
	.w4(32'h3858eab9),
	.w5(32'h378ee4f3),
	.w6(32'h37fbe543),
	.w7(32'h37f2e018),
	.w8(32'hb7df25cc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c1245),
	.w1(32'hbab51890),
	.w2(32'hbab1caa7),
	.w3(32'hba48a578),
	.w4(32'hba81991f),
	.w5(32'hba768b64),
	.w6(32'hba00067e),
	.w7(32'hba4ae6d5),
	.w8(32'hba4aa8d6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cabe6a),
	.w1(32'h38ab6ba1),
	.w2(32'h380bfc15),
	.w3(32'h397146e7),
	.w4(32'h39646190),
	.w5(32'h3871c63c),
	.w6(32'h3970d224),
	.w7(32'h3973cf77),
	.w8(32'h38955738),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d23bd),
	.w1(32'h3880d2a8),
	.w2(32'h385923ea),
	.w3(32'h38985d8c),
	.w4(32'h38a2027d),
	.w5(32'h38a1b333),
	.w6(32'h383ae2e8),
	.w7(32'h38843a6d),
	.w8(32'h3829a06b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8483842),
	.w1(32'hb8214c06),
	.w2(32'hb810dd6c),
	.w3(32'hb71a45bb),
	.w4(32'hb7b45850),
	.w5(32'hb7aae684),
	.w6(32'h3786ad7a),
	.w7(32'hb766ec21),
	.w8(32'hb7ba3e37),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0e30d),
	.w1(32'hbaa259b9),
	.w2(32'hbabf701e),
	.w3(32'hb91d90ab),
	.w4(32'hba60a9be),
	.w5(32'hba047be7),
	.w6(32'hb8a1ff73),
	.w7(32'hb96f8ac8),
	.w8(32'hb9f57869),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897ab0),
	.w1(32'h3b856c1e),
	.w2(32'h3b561828),
	.w3(32'h3b5d0983),
	.w4(32'h3b64486a),
	.w5(32'h3b0a6f4d),
	.w6(32'h3ae4aa98),
	.w7(32'h3aeddb90),
	.w8(32'h3a6db893),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39680b),
	.w1(32'h3b769668),
	.w2(32'h3b4f132a),
	.w3(32'h3b091a16),
	.w4(32'h3b2f94c4),
	.w5(32'h3af8a603),
	.w6(32'h3aa15750),
	.w7(32'h3ae38dbe),
	.w8(32'h3aa5b0df),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37531daf),
	.w1(32'h36c87746),
	.w2(32'hb8b4788d),
	.w3(32'h37db4ad5),
	.w4(32'h36f653fb),
	.w5(32'hb8bc153f),
	.w6(32'hb7f93789),
	.w7(32'h37958a6e),
	.w8(32'hb8278404),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce0f28),
	.w1(32'h37958d37),
	.w2(32'h3852df2d),
	.w3(32'h385002c7),
	.w4(32'h39162880),
	.w5(32'h3878d6af),
	.w6(32'h3813257f),
	.w7(32'h38fa5715),
	.w8(32'h38811e71),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3800e6a3),
	.w1(32'h38f94311),
	.w2(32'h390a5fe6),
	.w3(32'h37d0aee2),
	.w4(32'h38bbf638),
	.w5(32'h385eaa75),
	.w6(32'h3711e64a),
	.w7(32'h384199bc),
	.w8(32'h3882b3bd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398466c5),
	.w1(32'hb7b377ea),
	.w2(32'h3982d8d3),
	.w3(32'h38e94353),
	.w4(32'hb8f8aa72),
	.w5(32'h38a1e8b5),
	.w6(32'hb801cd62),
	.w7(32'hb9595d85),
	.w8(32'h38f30acf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd49777),
	.w1(32'hbbd73106),
	.w2(32'hbbb89008),
	.w3(32'hbbc6ec98),
	.w4(32'hbb9ee911),
	.w5(32'hbb861f11),
	.w6(32'hbb7dc0c8),
	.w7(32'hbb436362),
	.w8(32'hbb255e79),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada5053),
	.w1(32'hbb1c1f7c),
	.w2(32'hbb22411b),
	.w3(32'hbaad2eb4),
	.w4(32'hbaf7885c),
	.w5(32'hbadac0b7),
	.w6(32'hba866abd),
	.w7(32'hbaa4605e),
	.w8(32'hba83406c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481f43),
	.w1(32'hbb6139fb),
	.w2(32'hbb62741f),
	.w3(32'hbb20d1c1),
	.w4(32'hbb31f595),
	.w5(32'hbb1f7d47),
	.w6(32'hbaf73b6b),
	.w7(32'hbafd74ea),
	.w8(32'hbad85c3b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd904c),
	.w1(32'h39422a8d),
	.w2(32'h37288d12),
	.w3(32'h3a14aa01),
	.w4(32'h3a400fac),
	.w5(32'h39fbb71a),
	.w6(32'h39fd94e9),
	.w7(32'h3a0f49fb),
	.w8(32'h393a3870),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643969),
	.w1(32'hbb82d028),
	.w2(32'hbb780fc6),
	.w3(32'hbb4cf6b8),
	.w4(32'hbb803123),
	.w5(32'hbb62c966),
	.w6(32'hbac0826b),
	.w7(32'hbb098d6f),
	.w8(32'hbb0f0ad7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2572c),
	.w1(32'hb89f1b84),
	.w2(32'h39985e4e),
	.w3(32'hb995a59f),
	.w4(32'h388aa8da),
	.w5(32'h39984bfd),
	.w6(32'hb8f60232),
	.w7(32'h386a332f),
	.w8(32'h3985fe68),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60a1f8),
	.w1(32'hb9e68b5a),
	.w2(32'hb8fbca26),
	.w3(32'hba24d8d8),
	.w4(32'hb9854efe),
	.w5(32'hb90a350f),
	.w6(32'hb9958e36),
	.w7(32'hb89a73c2),
	.w8(32'hb921d83d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b898b),
	.w1(32'hb9692474),
	.w2(32'h383db1fb),
	.w3(32'hb980b66e),
	.w4(32'hb96d09f8),
	.w5(32'hb8ff969d),
	.w6(32'hb9bc3767),
	.w7(32'hb954bf00),
	.w8(32'hb952c9ae),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab03171),
	.w1(32'hbb258955),
	.w2(32'hbb177866),
	.w3(32'hbaa82c19),
	.w4(32'hbb0abb3e),
	.w5(32'hbaf811ba),
	.w6(32'hba470730),
	.w7(32'hbac2c3ef),
	.w8(32'hba978edc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c29e1e),
	.w1(32'hb79cfa82),
	.w2(32'h38cc9fa6),
	.w3(32'h3809d388),
	.w4(32'h390130b3),
	.w5(32'h390b1654),
	.w6(32'h38b4b24e),
	.w7(32'h38ec4e80),
	.w8(32'h38cee2ca),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913013),
	.w1(32'hbb8694ec),
	.w2(32'hbb86d84a),
	.w3(32'hbb733f92),
	.w4(32'hbb568ab1),
	.w5(32'hbb2c2498),
	.w6(32'hbb13be9e),
	.w7(32'hbaf0252f),
	.w8(32'hbae62771),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993967c),
	.w1(32'h39c427fb),
	.w2(32'h39cba4d4),
	.w3(32'h3976d4cc),
	.w4(32'h39b6c086),
	.w5(32'h39a34204),
	.w6(32'h395957f9),
	.w7(32'h397920df),
	.w8(32'h392c0bc0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999896c),
	.w1(32'hb9a39b45),
	.w2(32'hb9b20d05),
	.w3(32'hb98fcd2a),
	.w4(32'hb9af9992),
	.w5(32'hb98d0e03),
	.w6(32'hb934f173),
	.w7(32'hb93fb6b2),
	.w8(32'hb91b57ee),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a90f9e),
	.w1(32'h36197931),
	.w2(32'hb6121ed5),
	.w3(32'hb403548e),
	.w4(32'h3624226a),
	.w5(32'hb570ab72),
	.w6(32'h35c94c77),
	.w7(32'h36a24bb6),
	.w8(32'h3620bd5b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66eae8b),
	.w1(32'h366003a5),
	.w2(32'hb627a186),
	.w3(32'hb6ec0292),
	.w4(32'hb6359cfd),
	.w5(32'hb70e51bb),
	.w6(32'hb710bd99),
	.w7(32'hb6d2649f),
	.w8(32'hb640883e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397debb1),
	.w1(32'h38e8b6d7),
	.w2(32'h39024ef7),
	.w3(32'h395eae6c),
	.w4(32'h38cd254e),
	.w5(32'h3842b207),
	.w6(32'h38fcc31e),
	.w7(32'h37cd3448),
	.w8(32'hb8511afe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38548e0c),
	.w1(32'hb9800ad2),
	.w2(32'hb95be417),
	.w3(32'h38b9c4f6),
	.w4(32'hb907233c),
	.w5(32'hb8f0eb5e),
	.w6(32'h390f6d5f),
	.w7(32'hb90b965e),
	.w8(32'hb7902b27),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65a7e7),
	.w1(32'hba50b782),
	.w2(32'hba52a64d),
	.w3(32'hba6130fe),
	.w4(32'hb9f0e59a),
	.w5(32'hb9e5f455),
	.w6(32'hb9de5627),
	.w7(32'hb8eeaa6c),
	.w8(32'hb9c24447),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3056e),
	.w1(32'hba85a172),
	.w2(32'hba54bfe5),
	.w3(32'hb9bdb447),
	.w4(32'hba419679),
	.w5(32'hba270ced),
	.w6(32'hb9060ec1),
	.w7(32'hba0a0655),
	.w8(32'hb9c1363d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84f731d),
	.w1(32'hb7532bf2),
	.w2(32'hb6430bfa),
	.w3(32'hb7e50ce5),
	.w4(32'hb684e3d6),
	.w5(32'hb677a88e),
	.w6(32'hb6a0f14a),
	.w7(32'hb5903861),
	.w8(32'hb70d91b2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ab5c74),
	.w1(32'hb78ddd5b),
	.w2(32'hb74d1094),
	.w3(32'hb7959b15),
	.w4(32'hb742b3ec),
	.w5(32'hb65a7e11),
	.w6(32'hb71fcb23),
	.w7(32'hb6b68613),
	.w8(32'h36a4057e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5f174),
	.w1(32'h3827e665),
	.w2(32'h37f05f1b),
	.w3(32'h36d3e129),
	.w4(32'hb7101ea9),
	.w5(32'hb7bbfc12),
	.w6(32'hb805b3f1),
	.w7(32'hb7ed1cf3),
	.w8(32'hb86189bb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37db05d9),
	.w1(32'h37f6b0dd),
	.w2(32'h37d15a4f),
	.w3(32'h37951f54),
	.w4(32'h3790abce),
	.w5(32'h37a39099),
	.w6(32'h37bc932a),
	.w7(32'h37ad065c),
	.w8(32'h3794d6e4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d7c87),
	.w1(32'hb641be70),
	.w2(32'hb86d2b97),
	.w3(32'hb70a9148),
	.w4(32'h3804c9c9),
	.w5(32'hb77d6f6f),
	.w6(32'h38c62560),
	.w7(32'h386d3684),
	.w8(32'hb87c9065),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0a686),
	.w1(32'h3908630a),
	.w2(32'hb91b110e),
	.w3(32'h39f59433),
	.w4(32'h3998e5f9),
	.w5(32'hb8b98bef),
	.w6(32'h395077f1),
	.w7(32'h3944a4ca),
	.w8(32'hb9176470),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa111ad),
	.w1(32'h3ac189f9),
	.w2(32'h3abd30a4),
	.w3(32'h3a87e8dc),
	.w4(32'h3ac00a44),
	.w5(32'h3a7cb356),
	.w6(32'h3a383dec),
	.w7(32'h3a37e562),
	.w8(32'h39d0eaf3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a40e8a),
	.w1(32'h39a18063),
	.w2(32'hb9a2191d),
	.w3(32'h3a0ebdd9),
	.w4(32'h3a014cbd),
	.w5(32'hb7e9daa6),
	.w6(32'h38e9cf8d),
	.w7(32'h399df1bc),
	.w8(32'hb8e601db),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7648ff7),
	.w1(32'hb7a4b9fd),
	.w2(32'hb78565e1),
	.w3(32'hb786f9aa),
	.w4(32'hb7a0064b),
	.w5(32'hb771deb9),
	.w6(32'hb6666b5e),
	.w7(32'hb6dd64d6),
	.w8(32'h34148e25),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6894a03),
	.w1(32'h36ba83a5),
	.w2(32'h376bdb05),
	.w3(32'hb620933b),
	.w4(32'h36f2a616),
	.w5(32'h375a643f),
	.w6(32'h36a41d50),
	.w7(32'h375e3994),
	.w8(32'h37a2ce3a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8588562),
	.w1(32'hb807744d),
	.w2(32'hb7e781af),
	.w3(32'hb841646b),
	.w4(32'hb7d85785),
	.w5(32'hb7dcd4ed),
	.w6(32'hb8253046),
	.w7(32'hb76ba3ab),
	.w8(32'hb7aa64ad),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e0bb9),
	.w1(32'h389d5c7c),
	.w2(32'hb8f539f1),
	.w3(32'h38a0136a),
	.w4(32'hb6e55414),
	.w5(32'hb8fb45f2),
	.w6(32'h38825521),
	.w7(32'h388d1da9),
	.w8(32'hb80ab852),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86b440d),
	.w1(32'h3715497e),
	.w2(32'h3751d1d4),
	.w3(32'hb8389315),
	.w4(32'h3651609e),
	.w5(32'h375985e2),
	.w6(32'hb7ca3066),
	.w7(32'hb6aebffa),
	.w8(32'h3714869c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac0f86),
	.w1(32'hb8d50548),
	.w2(32'hb884f9a4),
	.w3(32'hb90848ab),
	.w4(32'hb90167bb),
	.w5(32'hb7cde471),
	.w6(32'h38b70aca),
	.w7(32'h38d292d4),
	.w8(32'hb8ff93c1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19cdd9),
	.w1(32'hbaa2181e),
	.w2(32'hbabc2156),
	.w3(32'h37be9cc9),
	.w4(32'h3a0aca2d),
	.w5(32'hb99b0e20),
	.w6(32'hb9558474),
	.w7(32'h3a2ab4a4),
	.w8(32'h3976ecc8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba7fa4),
	.w1(32'hbae53b90),
	.w2(32'hbaf8332a),
	.w3(32'hba94859d),
	.w4(32'hbac65fac),
	.w5(32'hbab77553),
	.w6(32'hba744a01),
	.w7(32'hba805391),
	.w8(32'hba78aa15),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855946),
	.w1(32'hba8431a6),
	.w2(32'hba81c775),
	.w3(32'hba58ad19),
	.w4(32'hba3f6e9a),
	.w5(32'hba30a9f9),
	.w6(32'hb9dbe7a3),
	.w7(32'hb9e75d41),
	.w8(32'hb9fec253),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995675b),
	.w1(32'hb9d09a80),
	.w2(32'hb9dd3eb9),
	.w3(32'hb90fff39),
	.w4(32'hb98135b9),
	.w5(32'hb9885f03),
	.w6(32'hb88ab426),
	.w7(32'hb93d0d39),
	.w8(32'hb8f46df2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6b42b),
	.w1(32'hbaecec35),
	.w2(32'hbaf57092),
	.w3(32'hbaaceb0e),
	.w4(32'hbac0292e),
	.w5(32'hba9f87cb),
	.w6(32'hba860e03),
	.w7(32'hba810fc6),
	.w8(32'hba49a9ab),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba807375),
	.w1(32'hbab1741a),
	.w2(32'hba9b2eaa),
	.w3(32'hba6f873e),
	.w4(32'hbaa7e361),
	.w5(32'hba81752e),
	.w6(32'hba01721e),
	.w7(32'hba42ce13),
	.w8(32'hba3bc7b6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67e7bc1),
	.w1(32'h3707c6e8),
	.w2(32'h378e43f8),
	.w3(32'hb628f85a),
	.w4(32'h373c7741),
	.w5(32'h37ab6840),
	.w6(32'h358022b3),
	.w7(32'h37080569),
	.w8(32'h37875440),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb633f753),
	.w1(32'hb5fa77ec),
	.w2(32'h359df88a),
	.w3(32'h3679bc37),
	.w4(32'h36d47de3),
	.w5(32'h36b497bb),
	.w6(32'hb590a329),
	.w7(32'h36cfa17c),
	.w8(32'h36e7c60b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36382439),
	.w1(32'h37779810),
	.w2(32'hb786d987),
	.w3(32'hb644ee33),
	.w4(32'h37594b4c),
	.w5(32'hb780428d),
	.w6(32'hb624e787),
	.w7(32'hb6f73f98),
	.w8(32'hb67cd31a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36689c66),
	.w1(32'h36cc6729),
	.w2(32'h36c9818f),
	.w3(32'h3611ae8b),
	.w4(32'h36d14f0c),
	.w5(32'h36bbf292),
	.w6(32'h362b1474),
	.w7(32'h368bc806),
	.w8(32'h36a9723c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5a09e),
	.w1(32'h3a9215cc),
	.w2(32'h3a73f114),
	.w3(32'h3ab60054),
	.w4(32'h3aa9e13b),
	.w5(32'h39996f36),
	.w6(32'h3a86d53b),
	.w7(32'h3a42e67e),
	.w8(32'h38fa25a8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3aec9),
	.w1(32'h39a7329c),
	.w2(32'h39a99b27),
	.w3(32'h39949d6b),
	.w4(32'h39637a4b),
	.w5(32'h39a37ebf),
	.w6(32'h395f8132),
	.w7(32'h39327ef1),
	.w8(32'h394808e3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a1495),
	.w1(32'hbb0cf55f),
	.w2(32'hbb0bcec0),
	.w3(32'hbaec65cb),
	.w4(32'hbb007411),
	.w5(32'hbac36ba7),
	.w6(32'hbaa8dfa0),
	.w7(32'hba9e5c72),
	.w8(32'hba89e113),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1465),
	.w1(32'hbaac07e5),
	.w2(32'hba51c8d1),
	.w3(32'hba4355b6),
	.w4(32'hbab1b2fb),
	.w5(32'hba85c5fc),
	.w6(32'hb90f3bc4),
	.w7(32'hba279169),
	.w8(32'hba85b07e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7a9cb),
	.w1(32'h3ad1c4dd),
	.w2(32'h3ab12f7d),
	.w3(32'h3aac1fca),
	.w4(32'h3a9a45c8),
	.w5(32'h3a8ae18e),
	.w6(32'h3a529cfd),
	.w7(32'h3a5fa57f),
	.w8(32'h3a3764c8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e00b6),
	.w1(32'hbafbbf42),
	.w2(32'hbad55043),
	.w3(32'hb9bcebb7),
	.w4(32'hbac662ce),
	.w5(32'hba7d2f6c),
	.w6(32'hb9d505cd),
	.w7(32'hba636691),
	.w8(32'hba0e4b81),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b0aa9),
	.w1(32'h39f88b96),
	.w2(32'h3a1a8341),
	.w3(32'h3a35727d),
	.w4(32'h3a5f5740),
	.w5(32'h39ce9371),
	.w6(32'h3a11558e),
	.w7(32'h39dea66f),
	.w8(32'hb8b165c6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dee90),
	.w1(32'hbaf7d58b),
	.w2(32'hbadd4fc8),
	.w3(32'hbae44c03),
	.w4(32'hbaab9477),
	.w5(32'hba776ba9),
	.w6(32'hba39bb00),
	.w7(32'hb9cf1541),
	.w8(32'hb948aad4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50d8a5),
	.w1(32'hb9b4cfac),
	.w2(32'hb9f829bf),
	.w3(32'hb9e05bdc),
	.w4(32'hb92cef59),
	.w5(32'hb9af13c4),
	.w6(32'hb9da1f93),
	.w7(32'h38bc8cff),
	.w8(32'hb8c6ac6b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d492f),
	.w1(32'hba07ee0c),
	.w2(32'hba27eab1),
	.w3(32'hb7989b6e),
	.w4(32'hb9ba61ba),
	.w5(32'hb9b7b45c),
	.w6(32'hb90d9716),
	.w7(32'hb856b240),
	.w8(32'hb917fdf6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f25dd3),
	.w1(32'h392269c8),
	.w2(32'h39b26647),
	.w3(32'hb8cb9d09),
	.w4(32'h39a2b057),
	.w5(32'hb69f76fa),
	.w6(32'hb96a670f),
	.w7(32'hb96df122),
	.w8(32'hb9636e28),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5a60),
	.w1(32'hbb212d15),
	.w2(32'hbab7e724),
	.w3(32'hbb1586bc),
	.w4(32'hbad83dc9),
	.w5(32'hba785767),
	.w6(32'hbad8c8c4),
	.w7(32'hbaa93989),
	.w8(32'hba139628),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a124882),
	.w1(32'h3a1ab80a),
	.w2(32'h3a42f5ab),
	.w3(32'h3a451429),
	.w4(32'h3a20d78f),
	.w5(32'h3a481ab9),
	.w6(32'h39eb4988),
	.w7(32'h39fbc5f8),
	.w8(32'h3a0a90c7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b42a0),
	.w1(32'h3a59d5bc),
	.w2(32'h3a3aab81),
	.w3(32'h3a4a0eeb),
	.w4(32'h3a322969),
	.w5(32'h3a2d6263),
	.w6(32'h3a65fa86),
	.w7(32'h3a118f10),
	.w8(32'hb72a7651),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b728ea5),
	.w1(32'h3b45b351),
	.w2(32'h3b6e74ce),
	.w3(32'h3b8a64c8),
	.w4(32'h3b65057d),
	.w5(32'h3b35c507),
	.w6(32'h3b529d49),
	.w7(32'h3b387ca7),
	.w8(32'h3b0f0cf4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c504),
	.w1(32'hbb8a1139),
	.w2(32'hbb79dae9),
	.w3(32'hbb811e94),
	.w4(32'hbb663ea0),
	.w5(32'hbb244f98),
	.w6(32'hbb4e0742),
	.w7(32'hbb178c63),
	.w8(32'hbad90492),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ec043),
	.w1(32'hbab354a8),
	.w2(32'hba9bdca8),
	.w3(32'hba578e63),
	.w4(32'hbaa199ea),
	.w5(32'hba264239),
	.w6(32'hb8dbb4f3),
	.w7(32'hba072452),
	.w8(32'hb9916baf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cff2e),
	.w1(32'hb9bc5f6f),
	.w2(32'h3958bf9a),
	.w3(32'hb9c189dd),
	.w4(32'h370bd45d),
	.w5(32'h3a269b03),
	.w6(32'hba374c27),
	.w7(32'hba4b840b),
	.w8(32'hb944725e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eba9f),
	.w1(32'h3a43c13d),
	.w2(32'h3a3baf40),
	.w3(32'h3a482766),
	.w4(32'h3a88dc0c),
	.w5(32'h3a8c2dba),
	.w6(32'h3a99d131),
	.w7(32'h3a7cd093),
	.w8(32'h3a2a2810),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a0a43),
	.w1(32'h39309947),
	.w2(32'h38636ac4),
	.w3(32'h3a202329),
	.w4(32'h3913cef0),
	.w5(32'hb8c79db2),
	.w6(32'h3a2733f1),
	.w7(32'h39982954),
	.w8(32'hb8308aca),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3785f07e),
	.w1(32'hb80929ff),
	.w2(32'hb804ced4),
	.w3(32'h38b412a9),
	.w4(32'h369a678b),
	.w5(32'hb7284db0),
	.w6(32'h37d72c2d),
	.w7(32'h36448c6f),
	.w8(32'h3688b233),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e9ab55),
	.w1(32'h382ca852),
	.w2(32'h380ca5aa),
	.w3(32'h38592144),
	.w4(32'h38821bab),
	.w5(32'h37e12c1c),
	.w6(32'h382d55af),
	.w7(32'h384651b7),
	.w8(32'h381897e5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9944a8),
	.w1(32'hbb9b4eeb),
	.w2(32'hbb8a8964),
	.w3(32'hbb92fb81),
	.w4(32'hbb81a9e0),
	.w5(32'hbb46aa09),
	.w6(32'hbb3fa734),
	.w7(32'hbb08cce9),
	.w8(32'hbad19784),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308be5),
	.w1(32'hbb206c78),
	.w2(32'hbb02b05b),
	.w3(32'hbb0b230f),
	.w4(32'hbae6481d),
	.w5(32'hbad2e127),
	.w6(32'hbaae55e7),
	.w7(32'hba9781ba),
	.w8(32'hba811620),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8083ec),
	.w1(32'h3a4c76d5),
	.w2(32'h3a5ef049),
	.w3(32'h3a6ef11a),
	.w4(32'h3a31d971),
	.w5(32'h3a4e54eb),
	.w6(32'h39e6be54),
	.w7(32'h39ff4af2),
	.w8(32'h3a355e12),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e28313),
	.w1(32'hba66dd16),
	.w2(32'hba455dc4),
	.w3(32'hb982113b),
	.w4(32'hba218dd5),
	.w5(32'hba14cfd9),
	.w6(32'hb9d1b69a),
	.w7(32'hba1f357e),
	.w8(32'hba279ce1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dbd25),
	.w1(32'h3a25c21d),
	.w2(32'h3a0bf1da),
	.w3(32'h3a2440b3),
	.w4(32'h3a1f2d48),
	.w5(32'h39c5cf18),
	.w6(32'h39e8144f),
	.w7(32'h39897a78),
	.w8(32'h384b53d5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0256),
	.w1(32'hbb1ba368),
	.w2(32'hbb1f0875),
	.w3(32'hbab45f13),
	.w4(32'hbaf35a91),
	.w5(32'hbacedb63),
	.w6(32'hba8bb41a),
	.w7(32'hbab21ec6),
	.w8(32'hba8f1edf),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06873f),
	.w1(32'hbb1699b2),
	.w2(32'hbb16d03e),
	.w3(32'hbae1564f),
	.w4(32'hbb026bba),
	.w5(32'hbad99e3b),
	.w6(32'hba9d1b51),
	.w7(32'hbab0821e),
	.w8(32'hba91eb87),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361c3fa4),
	.w1(32'hb6cba80c),
	.w2(32'h36f98b72),
	.w3(32'h37dccd1b),
	.w4(32'h37e2cb98),
	.w5(32'h3732d96a),
	.w6(32'hb75027f1),
	.w7(32'hb7c97249),
	.w8(32'hb6a60997),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6db71a5),
	.w1(32'hb6d8b5d3),
	.w2(32'hb70a4c1b),
	.w3(32'hb6e89080),
	.w4(32'hb6c0dcf6),
	.w5(32'hb6b2bb0c),
	.w6(32'hb6cd7193),
	.w7(32'hb6809cb8),
	.w8(32'hb68cd7f8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d6135a),
	.w1(32'h36023d97),
	.w2(32'h361bcd74),
	.w3(32'h35d04035),
	.w4(32'h35a770f1),
	.w5(32'h348687f5),
	.w6(32'h365fdf6f),
	.w7(32'h36122873),
	.w8(32'h353df41f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863d239),
	.w1(32'hb6db26f0),
	.w2(32'h382a9036),
	.w3(32'hb7460fa3),
	.w4(32'h384c9453),
	.w5(32'h36f89155),
	.w6(32'hb32eaf3e),
	.w7(32'hb78c5978),
	.w8(32'hb7ed070c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7f26c),
	.w1(32'hbb0e5ea8),
	.w2(32'hbb0f67af),
	.w3(32'hbac08daa),
	.w4(32'hbae7f140),
	.w5(32'hbab1c39a),
	.w6(32'hbab70853),
	.w7(32'hbaaceaeb),
	.w8(32'hba5dba8d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d373a0),
	.w1(32'hb8916d1d),
	.w2(32'hb91bbffa),
	.w3(32'hb6363cff),
	.w4(32'h3716da18),
	.w5(32'hb8b81338),
	.w6(32'hb806bf32),
	.w7(32'hb8765abf),
	.w8(32'hb8ad7442),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998d502),
	.w1(32'hb97d456d),
	.w2(32'hb93ffc0c),
	.w3(32'hb9864210),
	.w4(32'hb9545812),
	.w5(32'hb8de0805),
	.w6(32'hb896d02d),
	.w7(32'h374d33b3),
	.w8(32'hb76de21b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65ffa3),
	.w1(32'h3a20f2b0),
	.w2(32'h3959e64f),
	.w3(32'h3a4bec2d),
	.w4(32'h39f90d02),
	.w5(32'h3916ff3d),
	.w6(32'h39791841),
	.w7(32'h3946fba5),
	.w8(32'hb5a505af),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a8d11b),
	.w1(32'hb6c22699),
	.w2(32'hb601bc02),
	.w3(32'hb696ac9a),
	.w4(32'hb70aad6c),
	.w5(32'hb601ae0a),
	.w6(32'h36412fe4),
	.w7(32'h367ec71f),
	.w8(32'h35344c92),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ec1cc),
	.w1(32'h395ef3d4),
	.w2(32'h394b9689),
	.w3(32'h393b425c),
	.w4(32'h392fb97d),
	.w5(32'h391b4c47),
	.w6(32'h391ba178),
	.w7(32'h392521e5),
	.w8(32'h38bc9529),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d537ea),
	.w1(32'h37493536),
	.w2(32'h36450b7b),
	.w3(32'hb70f8f16),
	.w4(32'hb6bf9ed6),
	.w5(32'hb6a11a75),
	.w6(32'hb77e0189),
	.w7(32'h371b65b7),
	.w8(32'h378545fa),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392797bf),
	.w1(32'h38f34dc8),
	.w2(32'h3a295c86),
	.w3(32'h38ecbf86),
	.w4(32'h3a95644f),
	.w5(32'h3a0f6231),
	.w6(32'h3a9e1c26),
	.w7(32'h39f263bf),
	.w8(32'h3af26b5c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad9b57),
	.w1(32'hbb4646f0),
	.w2(32'hbb5834d2),
	.w3(32'h3a99ea8b),
	.w4(32'hbb276131),
	.w5(32'hbb5429bf),
	.w6(32'hbb0bb4ef),
	.w7(32'hbb1df55b),
	.w8(32'hbafa9e05),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb658ee5),
	.w1(32'hba5a2196),
	.w2(32'hba59a188),
	.w3(32'hbb0fffe0),
	.w4(32'h39bac0df),
	.w5(32'hba1e53d1),
	.w6(32'hbb0eb048),
	.w7(32'hbb17181b),
	.w8(32'hbaddce2b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb023225),
	.w1(32'h3a42e249),
	.w2(32'h3ad69dfc),
	.w3(32'hb9c20a42),
	.w4(32'h3ab61ae1),
	.w5(32'h3b184392),
	.w6(32'h3a0ef4cb),
	.w7(32'h3acc7a06),
	.w8(32'h3a8024ae),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af47dc9),
	.w1(32'hbafde4fc),
	.w2(32'hb9b2e596),
	.w3(32'h3b05c67b),
	.w4(32'hba9ce9c5),
	.w5(32'h39bc5682),
	.w6(32'h39c6b101),
	.w7(32'h3a2d0ca9),
	.w8(32'h3a730a42),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a016624),
	.w1(32'hba97ec66),
	.w2(32'h3b2b4ab5),
	.w3(32'h3a8a5720),
	.w4(32'h39b2e817),
	.w5(32'h3af7c806),
	.w6(32'hba9a6d8e),
	.w7(32'hba970ae9),
	.w8(32'h3a160327),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0adbb),
	.w1(32'h391cd45f),
	.w2(32'hb9bc9d1a),
	.w3(32'h3971e698),
	.w4(32'h3941008e),
	.w5(32'h394c3fd9),
	.w6(32'hb9ea19c1),
	.w7(32'hb9087cb1),
	.w8(32'h3a4e43bc),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eb131),
	.w1(32'hba36663d),
	.w2(32'hbadcfca8),
	.w3(32'h3abcabef),
	.w4(32'h37cd11fe),
	.w5(32'hbafbf651),
	.w6(32'hba20e0c0),
	.w7(32'hbab6ca99),
	.w8(32'hbaf30f23),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb760d70),
	.w1(32'hbb47aaa8),
	.w2(32'hbae9b9f3),
	.w3(32'hbb3792e9),
	.w4(32'hbb0d71c8),
	.w5(32'hb8407010),
	.w6(32'hbb1e1292),
	.w7(32'hba99c1f3),
	.w8(32'hbadd0b8e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a239),
	.w1(32'hbaa3bf9c),
	.w2(32'hba8325dd),
	.w3(32'hb9a0265e),
	.w4(32'hba900830),
	.w5(32'hba7017f3),
	.w6(32'hba49d64a),
	.w7(32'hb91610ff),
	.w8(32'h3795a312),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34c661),
	.w1(32'hba95c596),
	.w2(32'hba933dea),
	.w3(32'h3a007a74),
	.w4(32'hba0c16fa),
	.w5(32'hbafa92fd),
	.w6(32'hb8c17093),
	.w7(32'hba3be587),
	.w8(32'hb993ff2e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7300a8),
	.w1(32'hbaad5081),
	.w2(32'hba9b1da6),
	.w3(32'hb96bec24),
	.w4(32'hba213ba0),
	.w5(32'hbacf00ca),
	.w6(32'hb8f5b7f2),
	.w7(32'hb94dfd3a),
	.w8(32'hbab395f6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd39da),
	.w1(32'hbb3e694a),
	.w2(32'hbb18523d),
	.w3(32'hbb09054b),
	.w4(32'hbba6f64f),
	.w5(32'hbb8588c2),
	.w6(32'h3a6d4380),
	.w7(32'h3b19735e),
	.w8(32'h3a62d553),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79361d),
	.w1(32'hbbbc9939),
	.w2(32'hbb8bb138),
	.w3(32'hbb81bbe3),
	.w4(32'hbb8f6698),
	.w5(32'hbb58ab05),
	.w6(32'hbb8d48e2),
	.w7(32'hbb7a225c),
	.w8(32'hbb4bfc96),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb363f76),
	.w1(32'hba7c8ac6),
	.w2(32'h394260a5),
	.w3(32'hbb0fdd31),
	.w4(32'hba69f97a),
	.w5(32'hb9336365),
	.w6(32'hba484679),
	.w7(32'hb9a6413d),
	.w8(32'hb9c531d4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a8c91),
	.w1(32'hbac8f25d),
	.w2(32'hb97e0467),
	.w3(32'h3a4fb170),
	.w4(32'hbaebb970),
	.w5(32'hba444505),
	.w6(32'h39e733dd),
	.w7(32'h3ad3d465),
	.w8(32'h3a0ba2f4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30c278),
	.w1(32'hbaf93b83),
	.w2(32'hb9a3787a),
	.w3(32'h3a55b7a1),
	.w4(32'h3a43ca07),
	.w5(32'h3a8df422),
	.w6(32'hbaa4478f),
	.w7(32'hba94a937),
	.w8(32'hba529d1d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7e292),
	.w1(32'hb9acdeb7),
	.w2(32'hba7bd584),
	.w3(32'h390fc1af),
	.w4(32'h3a2967d7),
	.w5(32'hba1313a3),
	.w6(32'hb96960be),
	.w7(32'hba6292c9),
	.w8(32'hb9f76a4d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38413dce),
	.w1(32'hbab21ccc),
	.w2(32'hbb29f7bc),
	.w3(32'h3a4a52c4),
	.w4(32'h3b1a6315),
	.w5(32'h398e6a36),
	.w6(32'hbb2c4cd4),
	.w7(32'hbb6ff7d8),
	.w8(32'hba6160e6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab46d0a),
	.w1(32'h3794f676),
	.w2(32'h3a6ce38d),
	.w3(32'h3b07e2a3),
	.w4(32'h3aa5a0c3),
	.w5(32'h3ac9b6f5),
	.w6(32'hb8f26f91),
	.w7(32'h3a750e57),
	.w8(32'h37d2146b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af185a6),
	.w1(32'h38aa1bb4),
	.w2(32'hba21da07),
	.w3(32'h3b05b57d),
	.w4(32'h3a78efb2),
	.w5(32'hb9b8edfd),
	.w6(32'h3a382247),
	.w7(32'h3a2bc600),
	.w8(32'h3a8be275),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21358c),
	.w1(32'hbb95a570),
	.w2(32'hbbb731ae),
	.w3(32'hbb2128bd),
	.w4(32'hbb4a8ae2),
	.w5(32'hbb9ce84c),
	.w6(32'hbb4e41e2),
	.w7(32'hbb6a203e),
	.w8(32'hbb3586be),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ec85d),
	.w1(32'h3ac38538),
	.w2(32'h3acae066),
	.w3(32'hb88b647f),
	.w4(32'h3b49639d),
	.w5(32'h3b0fd3c6),
	.w6(32'h3b83c6af),
	.w7(32'h3b13c15d),
	.w8(32'h3a854559),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fde29),
	.w1(32'hbb98ea93),
	.w2(32'hbad677a4),
	.w3(32'hba1b9232),
	.w4(32'hbbb69d06),
	.w5(32'hba882056),
	.w6(32'hbb3db4ce),
	.w7(32'hbb2824b7),
	.w8(32'hbb4df2f2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a584bc),
	.w1(32'hbb8b5600),
	.w2(32'hbbac1fb7),
	.w3(32'h36e11e01),
	.w4(32'hbb05c68c),
	.w5(32'hbb906c45),
	.w6(32'hbb6f02b9),
	.w7(32'hbbf803ae),
	.w8(32'hbb0f25a2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39924fe8),
	.w1(32'hbb3a5bf6),
	.w2(32'hbb0c380e),
	.w3(32'h3b6a0ecc),
	.w4(32'hbb0c690c),
	.w5(32'hbab79f51),
	.w6(32'hbae0a419),
	.w7(32'hbaa9a52a),
	.w8(32'hba3d4b14),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9082133),
	.w1(32'hb90dd9e1),
	.w2(32'hbab3618a),
	.w3(32'h3a5478e7),
	.w4(32'h3ab5c9f0),
	.w5(32'hba6276ed),
	.w6(32'h3aedb629),
	.w7(32'h3b1838d8),
	.w8(32'h3b14fa63),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88756a2),
	.w1(32'hbb73a24e),
	.w2(32'hbb9d085b),
	.w3(32'h3a610466),
	.w4(32'h399b3fe1),
	.w5(32'hbacaf3c5),
	.w6(32'hbbcce259),
	.w7(32'hbbbf702c),
	.w8(32'hbb72c966),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1ad5b),
	.w1(32'hbb438bbe),
	.w2(32'hbb157e0a),
	.w3(32'hbaf786db),
	.w4(32'hbab18aaa),
	.w5(32'hbac4ffd0),
	.w6(32'hbb6e3f8a),
	.w7(32'hbb46ba5e),
	.w8(32'hbacc9522),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51e26b),
	.w1(32'hba94f69e),
	.w2(32'hbb007fa9),
	.w3(32'hbac2f551),
	.w4(32'hb907fd63),
	.w5(32'hbaae6f40),
	.w6(32'hba4356fc),
	.w7(32'hba6192c5),
	.w8(32'hba45e620),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adeda22),
	.w1(32'h3bc83845),
	.w2(32'hba03dc75),
	.w3(32'h3b0fd7ed),
	.w4(32'h3c15483b),
	.w5(32'h3a4511ba),
	.w6(32'h3c516ff4),
	.w7(32'h3be3ed43),
	.w8(32'h3bb4cb41),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb119213),
	.w1(32'h3c8013e6),
	.w2(32'h3c35ad96),
	.w3(32'h3af56a76),
	.w4(32'h3c804967),
	.w5(32'h3c2ec5dd),
	.w6(32'h3c84ac7f),
	.w7(32'h3c2d31ad),
	.w8(32'h3bcfc6f0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd58a2),
	.w1(32'hb9807807),
	.w2(32'hb88ffd22),
	.w3(32'h3b206a64),
	.w4(32'h39b7b2f3),
	.w5(32'h3970f809),
	.w6(32'h3a812e2d),
	.w7(32'h3a46f0f3),
	.w8(32'h396f405a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991595e),
	.w1(32'hbacc4134),
	.w2(32'hb9a68967),
	.w3(32'h39907893),
	.w4(32'hb9c63eb4),
	.w5(32'hb96a5865),
	.w6(32'hba7a5eac),
	.w7(32'hba14393d),
	.w8(32'h3717f0de),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16f099),
	.w1(32'hbb0ec5ba),
	.w2(32'hbb3f94d7),
	.w3(32'h39a95daf),
	.w4(32'hbabcc4ac),
	.w5(32'hbb3287e7),
	.w6(32'hbb30577d),
	.w7(32'hbb5b2236),
	.w8(32'hba8186df),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a390ec5),
	.w1(32'hbb0e1d6c),
	.w2(32'hbbd692da),
	.w3(32'h3a660e86),
	.w4(32'hb948ca79),
	.w5(32'hbbabd185),
	.w6(32'hbad56020),
	.w7(32'hbbe08f85),
	.w8(32'hbbae7e41),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03bcdc),
	.w1(32'hbb4faaca),
	.w2(32'hbb79bac0),
	.w3(32'hbbf0457e),
	.w4(32'hbadf0103),
	.w5(32'hbb58bd09),
	.w6(32'hbabcd9ff),
	.w7(32'hbb3b61c2),
	.w8(32'hbb56719b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489052),
	.w1(32'hbaec4f45),
	.w2(32'hb9f53fa2),
	.w3(32'hbb4ab644),
	.w4(32'hba20eb7d),
	.w5(32'hb8bbb54f),
	.w6(32'hb8de3448),
	.w7(32'h3a5b1439),
	.w8(32'h3a99f091),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc4594),
	.w1(32'h3a27cbc0),
	.w2(32'h3a5bb659),
	.w3(32'h3a6e8ca0),
	.w4(32'h3ab471a1),
	.w5(32'h3a62e8ce),
	.w6(32'hba340d6e),
	.w7(32'h38fcb08a),
	.w8(32'h388313ef),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e83be),
	.w1(32'h3959d027),
	.w2(32'h3aa39edd),
	.w3(32'h3936c3a5),
	.w4(32'h3a8b8739),
	.w5(32'h3b09245b),
	.w6(32'hb933343d),
	.w7(32'h3a8c19ac),
	.w8(32'h39b95b22),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2f218),
	.w1(32'hba83bb0a),
	.w2(32'hba804a2b),
	.w3(32'h3a8a9c13),
	.w4(32'hba48b212),
	.w5(32'hba813b09),
	.w6(32'hbab29b21),
	.w7(32'hbaabf888),
	.w8(32'hba4cf616),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9add8a),
	.w1(32'hbadd988f),
	.w2(32'hb9f6f9d7),
	.w3(32'hb94fcede),
	.w4(32'hba322bfc),
	.w5(32'h3a37fdea),
	.w6(32'hbaa3832d),
	.w7(32'h3950e5fa),
	.w8(32'h39d1cf10),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e87c),
	.w1(32'h3a7c1d48),
	.w2(32'h3b2dac89),
	.w3(32'hbb32764c),
	.w4(32'h3ba6a8f2),
	.w5(32'h3bdcde34),
	.w6(32'h3bc38821),
	.w7(32'h3baad097),
	.w8(32'hb9ced25f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7422c),
	.w1(32'hba8e1452),
	.w2(32'hbac6a3fb),
	.w3(32'hbade62fe),
	.w4(32'h36b04e7f),
	.w5(32'hba186ad7),
	.w6(32'h380e4d8a),
	.w7(32'hb9799f9c),
	.w8(32'hba321e3b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99ed7),
	.w1(32'hbbbe57cb),
	.w2(32'hbb8276ba),
	.w3(32'hbb640bf0),
	.w4(32'hbb863f4d),
	.w5(32'hbb453405),
	.w6(32'hbb3112e0),
	.w7(32'hbb6012d3),
	.w8(32'hbae403ff),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba262a87),
	.w1(32'h393207a6),
	.w2(32'h3a3b12db),
	.w3(32'h3a215c9d),
	.w4(32'h3a0f9951),
	.w5(32'hb92d8e75),
	.w6(32'h36786b2d),
	.w7(32'h3aa48c1a),
	.w8(32'hba9710b8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadee167),
	.w1(32'hbad3ab0b),
	.w2(32'hb8c2cdab),
	.w3(32'hbb94ec19),
	.w4(32'hb97f1641),
	.w5(32'h3aac5b7a),
	.w6(32'hba860c49),
	.w7(32'h39f68256),
	.w8(32'hba3dc6ac),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0698db),
	.w1(32'hbaf2c18f),
	.w2(32'hba95b9e4),
	.w3(32'h3ab35eee),
	.w4(32'hba8c37f5),
	.w5(32'h3990d579),
	.w6(32'hba1dc553),
	.w7(32'hb9b2cc72),
	.w8(32'hb9d4090f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb858490),
	.w1(32'hbbc14a77),
	.w2(32'hbac5d09b),
	.w3(32'hbb1eed0e),
	.w4(32'hbb33de58),
	.w5(32'hbab472e5),
	.w6(32'hbb963057),
	.w7(32'hbaff5739),
	.w8(32'hbac64d26),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a2f8),
	.w1(32'h3aba0393),
	.w2(32'hbb6c0a31),
	.w3(32'hba42be4c),
	.w4(32'h3bd6b8fc),
	.w5(32'h3a75fec6),
	.w6(32'h3c0feb99),
	.w7(32'h3b7c1045),
	.w8(32'h3ba662f4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c5e7),
	.w1(32'hbb94faed),
	.w2(32'hbb4cc7e8),
	.w3(32'h3a84b7ba),
	.w4(32'hbb3015d3),
	.w5(32'hbb215ded),
	.w6(32'hbb5b56d5),
	.w7(32'hbb11536d),
	.w8(32'hbad3b347),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c81b4),
	.w1(32'h38d4de26),
	.w2(32'h3a1ed8c6),
	.w3(32'h386dc3e8),
	.w4(32'h38db9518),
	.w5(32'h3a34d14b),
	.w6(32'hb6f2e7a2),
	.w7(32'h3a393986),
	.w8(32'h3a6bb79f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13d90a),
	.w1(32'hbaad1cf6),
	.w2(32'hba70338a),
	.w3(32'h3acb5124),
	.w4(32'hba931e55),
	.w5(32'hba16cbe2),
	.w6(32'hbacae49a),
	.w7(32'hba3c755b),
	.w8(32'hba704ef3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd4687),
	.w1(32'h3aaa74ff),
	.w2(32'hba8ae729),
	.w3(32'hba902cf2),
	.w4(32'h3b381a8f),
	.w5(32'h3a61a1d0),
	.w6(32'h3a7e163f),
	.w7(32'hba8efb2a),
	.w8(32'hb7daf7bf),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a1a29),
	.w1(32'h3aa2ce3b),
	.w2(32'h3a07a377),
	.w3(32'h3b276cd6),
	.w4(32'h3b5eed96),
	.w5(32'h3ada5977),
	.w6(32'h3ad68a3b),
	.w7(32'h3ab5b2c8),
	.w8(32'h3a89bbdc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa87471),
	.w1(32'hbb100b07),
	.w2(32'hbb38bc29),
	.w3(32'h3b026f97),
	.w4(32'hbb18d1f7),
	.w5(32'hbb384a0b),
	.w6(32'hbb25d302),
	.w7(32'hbb285b79),
	.w8(32'hbb5009cc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158f54),
	.w1(32'hba8dd1e2),
	.w2(32'h3a84f42c),
	.w3(32'hbb2d6a80),
	.w4(32'h3a6ebc4e),
	.w5(32'h3a93492d),
	.w6(32'hbab5bde3),
	.w7(32'hb84f0e8e),
	.w8(32'h3a0ed352),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c1e67),
	.w1(32'h3b4e3587),
	.w2(32'h3b8ffe19),
	.w3(32'h3abcfa49),
	.w4(32'h3b77eafc),
	.w5(32'h3b3ea347),
	.w6(32'h3bc5250d),
	.w7(32'h3be67291),
	.w8(32'h3b5912d9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22d80c),
	.w1(32'hbb0c7fc9),
	.w2(32'h3ac680f4),
	.w3(32'hba5cae92),
	.w4(32'hb92fd901),
	.w5(32'h3b2c4ed5),
	.w6(32'hb9edbec1),
	.w7(32'h3aa5a691),
	.w8(32'hba5ad074),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba574f97),
	.w1(32'h3a6b219b),
	.w2(32'hba2e5de0),
	.w3(32'hb9a07a4e),
	.w4(32'hb9c28812),
	.w5(32'hba7eb5ab),
	.w6(32'hba905bc5),
	.w7(32'hbacd89a3),
	.w8(32'h390dbbab),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10fe43),
	.w1(32'hb9d3b4e6),
	.w2(32'hb9b3e108),
	.w3(32'hb8db68db),
	.w4(32'hb9291221),
	.w5(32'hb9683959),
	.w6(32'hba2d52af),
	.w7(32'hb9f573f4),
	.w8(32'hbaa4c740),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdae76),
	.w1(32'hbbd5b37e),
	.w2(32'hbbbdebb6),
	.w3(32'hbb9a37ab),
	.w4(32'hbba43685),
	.w5(32'hbb896fd9),
	.w6(32'hbbab903e),
	.w7(32'hbb804e5e),
	.w8(32'hbb4f50c8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ada6b7),
	.w1(32'hba1dd8ac),
	.w2(32'h3964078b),
	.w3(32'h3ac289cc),
	.w4(32'h39907bac),
	.w5(32'h3a5a22e2),
	.w6(32'hb92c0ac5),
	.w7(32'h3a28bb1c),
	.w8(32'h393fc23f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39984985),
	.w1(32'h385db693),
	.w2(32'h39922684),
	.w3(32'h3988544a),
	.w4(32'h3a47272d),
	.w5(32'h3a925739),
	.w6(32'hb9fa45ab),
	.w7(32'h3a07d05e),
	.w8(32'h3a509dc4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996f3e0),
	.w1(32'hbab842e1),
	.w2(32'hb9d5a7ec),
	.w3(32'h3aa9c687),
	.w4(32'hbadb3689),
	.w5(32'hba2467a1),
	.w6(32'hbb480277),
	.w7(32'hbafa121d),
	.w8(32'h39919d6a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4a10f),
	.w1(32'h399f79c9),
	.w2(32'h3a291d28),
	.w3(32'h3b0269f9),
	.w4(32'h3a26aec1),
	.w5(32'hb91b9db7),
	.w6(32'hb88c022b),
	.w7(32'h3a22dc29),
	.w8(32'hba6ccb20),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88c985),
	.w1(32'h3926dc3f),
	.w2(32'h3957225d),
	.w3(32'hbb423e02),
	.w4(32'h386a8ef0),
	.w5(32'hb9a76562),
	.w6(32'h39d00bce),
	.w7(32'hb9c02643),
	.w8(32'hb9a284c5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9106151),
	.w1(32'h3aae3a6d),
	.w2(32'hb8f9e6a0),
	.w3(32'h39c63a61),
	.w4(32'h391170c7),
	.w5(32'hb82cddd0),
	.w6(32'h3a533c93),
	.w7(32'hba05b774),
	.w8(32'h3a7bbbf2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac99288),
	.w1(32'h3c6b7345),
	.w2(32'h3c8030f2),
	.w3(32'h3acd3d0a),
	.w4(32'h3c801b6d),
	.w5(32'h3c819cc8),
	.w6(32'h3c4a1500),
	.w7(32'h3c3bf670),
	.w8(32'h3c124dbc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48056e),
	.w1(32'hbb7d4db7),
	.w2(32'h3a5c65a1),
	.w3(32'h3bbafb5c),
	.w4(32'h3b9cb080),
	.w5(32'h3be38358),
	.w6(32'h3965465e),
	.w7(32'h3966530c),
	.w8(32'h3a3e47ec),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee0433),
	.w1(32'hbb032a6f),
	.w2(32'hbb13517b),
	.w3(32'h3bbb76eb),
	.w4(32'hba20a310),
	.w5(32'hbac5481b),
	.w6(32'hba295ebb),
	.w7(32'hbabb6eac),
	.w8(32'hbadc2877),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043f39),
	.w1(32'hbb075f6b),
	.w2(32'hbb4ba80d),
	.w3(32'hbaac4e7d),
	.w4(32'hbb43f921),
	.w5(32'hbb0c0eba),
	.w6(32'hbac5226c),
	.w7(32'hbb32b80e),
	.w8(32'hbb2d6ab2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff175c),
	.w1(32'hba511cbc),
	.w2(32'hba13bf54),
	.w3(32'hba872c65),
	.w4(32'h39fdab4e),
	.w5(32'h3974f63e),
	.w6(32'hb97fb9ba),
	.w7(32'hb8218856),
	.w8(32'hb9bce270),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987805e),
	.w1(32'hbacbfe00),
	.w2(32'hbacd6de5),
	.w3(32'h39968de1),
	.w4(32'hba8cbcb4),
	.w5(32'hba874eec),
	.w6(32'hbad866e7),
	.w7(32'hbab0b528),
	.w8(32'hba992465),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994899f),
	.w1(32'hbaa21ae7),
	.w2(32'hba9bb99a),
	.w3(32'hb7ae4e13),
	.w4(32'hba5b8a48),
	.w5(32'hba95fa09),
	.w6(32'hbab39055),
	.w7(32'hbaada074),
	.w8(32'hba27f3d2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2da86),
	.w1(32'hbb0c761a),
	.w2(32'hba3f4570),
	.w3(32'h39d60f6f),
	.w4(32'hba42d317),
	.w5(32'hb8e81907),
	.w6(32'hba2e6e2a),
	.w7(32'hb8b4a27d),
	.w8(32'h3a04a44b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf14ccc),
	.w1(32'hba517933),
	.w2(32'hba872a17),
	.w3(32'h399dfc6d),
	.w4(32'h3a090eb3),
	.w5(32'hb8b11e52),
	.w6(32'h3a47a2a9),
	.w7(32'h3a2aa9e7),
	.w8(32'hb9c2a176),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094e41),
	.w1(32'h3aee63d7),
	.w2(32'h3af1bf03),
	.w3(32'h3b29897e),
	.w4(32'h3bae91eb),
	.w5(32'h3b42f3bc),
	.w6(32'hba0e3908),
	.w7(32'h3a7e447c),
	.w8(32'h3b027cad),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f29b),
	.w1(32'hb9bf7c38),
	.w2(32'hb8dcc572),
	.w3(32'h3b374d5f),
	.w4(32'hba04f07c),
	.w5(32'hba701029),
	.w6(32'h395be682),
	.w7(32'h3a8f0b40),
	.w8(32'h3a22b8f5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372e2a34),
	.w1(32'h3a946765),
	.w2(32'hba999a62),
	.w3(32'h3914f710),
	.w4(32'h3ad7e756),
	.w5(32'hba94a19e),
	.w6(32'h39aea42f),
	.w7(32'hba8a7446),
	.w8(32'hb9811fee),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d359f),
	.w1(32'hbb966975),
	.w2(32'hbb0e30c1),
	.w3(32'hba0cbd75),
	.w4(32'hba535cdf),
	.w5(32'hb9d7436d),
	.w6(32'hbbae1700),
	.w7(32'hbb5dc16c),
	.w8(32'hba0fc6d7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba406888),
	.w1(32'hbb48071f),
	.w2(32'hbb138d7b),
	.w3(32'h3a5dd747),
	.w4(32'hbae69a0a),
	.w5(32'hbb0104a1),
	.w6(32'hb74005c3),
	.w7(32'hba1d6ff4),
	.w8(32'h38b4f89a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4763),
	.w1(32'hb78ecd48),
	.w2(32'h3a98f139),
	.w3(32'hb8c35b3e),
	.w4(32'h3bd44014),
	.w5(32'h3c00340e),
	.w6(32'h3be9d3cc),
	.w7(32'h3bcd17bb),
	.w8(32'h3b84002e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affd672),
	.w1(32'h3b0b91b4),
	.w2(32'h3aeb4027),
	.w3(32'h3ba89256),
	.w4(32'h3b007d31),
	.w5(32'h3b0373bf),
	.w6(32'h3addf9f4),
	.w7(32'h3ad1d800),
	.w8(32'hb9d2b99d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391976c7),
	.w1(32'h39929137),
	.w2(32'hba921688),
	.w3(32'hb93aa285),
	.w4(32'h3af5e907),
	.w5(32'h37af2b13),
	.w6(32'h3b939007),
	.w7(32'h3b87a978),
	.w8(32'h3b7e6841),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1567c4),
	.w1(32'h3a13d2d6),
	.w2(32'h3a38fe8c),
	.w3(32'h388788e8),
	.w4(32'h3a143179),
	.w5(32'h3a432a9a),
	.w6(32'hb81197d6),
	.w7(32'h39b392d9),
	.w8(32'hba8071da),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1920f6),
	.w1(32'hbba1bb75),
	.w2(32'hbb96ccec),
	.w3(32'hbad8dd4f),
	.w4(32'hb9e37a26),
	.w5(32'hb7956f4c),
	.w6(32'hbaac4e6e),
	.w7(32'hbb3cbb5d),
	.w8(32'hb9c8fce6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d31e),
	.w1(32'h3b862db8),
	.w2(32'h3ba15b8f),
	.w3(32'h3b18b69c),
	.w4(32'h3b9d5ab0),
	.w5(32'h3bcf2a26),
	.w6(32'h3b7117af),
	.w7(32'h3bafb80d),
	.w8(32'h3b9cca80),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd52f43),
	.w1(32'hb8aabc56),
	.w2(32'hbad3e62c),
	.w3(32'h3bab191d),
	.w4(32'hb8a3ab65),
	.w5(32'hbaf98063),
	.w6(32'hb89b8b89),
	.w7(32'hba235a22),
	.w8(32'hba9eca05),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1024),
	.w1(32'hb9c100bc),
	.w2(32'hb717fd27),
	.w3(32'hbab9fb80),
	.w4(32'h39b1bb64),
	.w5(32'h39ded798),
	.w6(32'h3a839526),
	.w7(32'h3a790d6b),
	.w8(32'h3a1c981a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b0375),
	.w1(32'hba59187c),
	.w2(32'h3a2f7304),
	.w3(32'h3999e76c),
	.w4(32'h3a438d43),
	.w5(32'h3a5ed21e),
	.w6(32'hba55267a),
	.w7(32'h39897789),
	.w8(32'hb9d0acaa),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd3aa3),
	.w1(32'hba3a49cf),
	.w2(32'h39b8ee3c),
	.w3(32'h3929a166),
	.w4(32'h3a390347),
	.w5(32'h3a4e333c),
	.w6(32'h3a3e34e6),
	.w7(32'h3a2bc1e9),
	.w8(32'h3a48414a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4c823),
	.w1(32'hba977327),
	.w2(32'hba670913),
	.w3(32'h3a3ffd12),
	.w4(32'hba34620a),
	.w5(32'hba66b58f),
	.w6(32'hb8d56644),
	.w7(32'h39d3ec4e),
	.w8(32'hb8cf6af3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e95e88),
	.w1(32'h3aba9efd),
	.w2(32'h3b3d4fa6),
	.w3(32'h398a7797),
	.w4(32'h3b344247),
	.w5(32'h3b6514d0),
	.w6(32'h3acbd1ad),
	.w7(32'h3b4261e9),
	.w8(32'h3adbd983),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69f1f4),
	.w1(32'h3b36fc43),
	.w2(32'h3b104287),
	.w3(32'h3b138b64),
	.w4(32'h3b80700c),
	.w5(32'h3b256224),
	.w6(32'h3b587527),
	.w7(32'h3b19a06b),
	.w8(32'h3a9dec23),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398673fb),
	.w1(32'h39c8b186),
	.w2(32'h3a961296),
	.w3(32'hb7074d7f),
	.w4(32'h3ba09e7e),
	.w5(32'h3b8295a7),
	.w6(32'h3bf39f73),
	.w7(32'h3bae47f4),
	.w8(32'h3b875386),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57e2cd),
	.w1(32'hbb006733),
	.w2(32'hba816be2),
	.w3(32'h3b417516),
	.w4(32'hbad7ffd6),
	.w5(32'hb92984bf),
	.w6(32'hba4de0db),
	.w7(32'hb96e7b71),
	.w8(32'hba34291d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cfdd9),
	.w1(32'hba6862fc),
	.w2(32'hbac7ac22),
	.w3(32'h38ef093f),
	.w4(32'hbace1f67),
	.w5(32'hbacf0955),
	.w6(32'hbae331a5),
	.w7(32'hbb06cc1e),
	.w8(32'hbb2df177),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9b11c),
	.w1(32'hbb382693),
	.w2(32'hbafa6bca),
	.w3(32'hba9d5082),
	.w4(32'h38958d5a),
	.w5(32'h39bd1a58),
	.w6(32'hbb937fcf),
	.w7(32'hbbd33d49),
	.w8(32'hbaa544f4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45dfcc),
	.w1(32'h3b991b1b),
	.w2(32'h3af95204),
	.w3(32'h3b64c16b),
	.w4(32'h3baf8c06),
	.w5(32'h3a2e6d4d),
	.w6(32'h3b72a367),
	.w7(32'h39b7a86b),
	.w8(32'h3948505f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a851b0a),
	.w1(32'h3a7a9c64),
	.w2(32'h3af16ab0),
	.w3(32'h3b091cc6),
	.w4(32'h3a481656),
	.w5(32'h3ad190e6),
	.w6(32'h3a894856),
	.w7(32'h3ac38b6b),
	.w8(32'h377d507e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1e229),
	.w1(32'h3b5f8046),
	.w2(32'h3a8d5d83),
	.w3(32'hba2e04c2),
	.w4(32'h3bae1fe3),
	.w5(32'h3b0bf8ef),
	.w6(32'h3bb71c5d),
	.w7(32'h3b8425fd),
	.w8(32'h3b2dc09f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a741e1c),
	.w1(32'hbb1525c1),
	.w2(32'hbaa8de97),
	.w3(32'h3ab97583),
	.w4(32'hbaf6309d),
	.w5(32'hb986b6b8),
	.w6(32'hbb2a8c0e),
	.w7(32'hbb170ee0),
	.w8(32'h3a92638c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35d264),
	.w1(32'h3aead240),
	.w2(32'h3a119dc8),
	.w3(32'h3af4048b),
	.w4(32'h3a949307),
	.w5(32'h3ab2ca45),
	.w6(32'hb9e37989),
	.w7(32'h3a0861e3),
	.w8(32'hba79af00),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7152d),
	.w1(32'hb9bbdd5b),
	.w2(32'h3a179c75),
	.w3(32'h3a5353cc),
	.w4(32'hba4e17ef),
	.w5(32'hba36da84),
	.w6(32'h3a8b7421),
	.w7(32'h3af115fe),
	.w8(32'h3ab3ec55),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93626e),
	.w1(32'hbb370efd),
	.w2(32'hbb1f00fc),
	.w3(32'hb9f3cf4e),
	.w4(32'hbaded56c),
	.w5(32'hbae148d3),
	.w6(32'hbb1319ee),
	.w7(32'hbab298b8),
	.w8(32'hba705f1a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0338e2),
	.w1(32'h3957a717),
	.w2(32'h3a1a16cc),
	.w3(32'h37e42527),
	.w4(32'h38a9d595),
	.w5(32'hb9551b46),
	.w6(32'h3a055c6a),
	.w7(32'h3a8e7f20),
	.w8(32'h3a6a1e92),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad1caf),
	.w1(32'hbb4d09cb),
	.w2(32'hbb4206cd),
	.w3(32'hba76a96d),
	.w4(32'hbaf11a26),
	.w5(32'hbb23b6a5),
	.w6(32'hbb11d8d0),
	.w7(32'hbb1d1c75),
	.w8(32'hba9ff091),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0615e9),
	.w1(32'h389b0878),
	.w2(32'h3a35a2fb),
	.w3(32'h39d2dd50),
	.w4(32'h38fc7ee5),
	.w5(32'h3a33e45b),
	.w6(32'h3a7b230d),
	.w7(32'h3a96b776),
	.w8(32'hb838cd73),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c790e),
	.w1(32'h3a0143df),
	.w2(32'h390127da),
	.w3(32'h3a8c1dd3),
	.w4(32'h3a6b74cd),
	.w5(32'h3a20d06a),
	.w6(32'h3b385d91),
	.w7(32'h3af6873d),
	.w8(32'h3a58e72b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1f43f),
	.w1(32'h3987bbc3),
	.w2(32'h3a4c8bd8),
	.w3(32'hb93ff842),
	.w4(32'hb7045fcb),
	.w5(32'hb82d7865),
	.w6(32'h39f0a4c7),
	.w7(32'h3a966863),
	.w8(32'h3a60f413),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce4e0f),
	.w1(32'hba8943c4),
	.w2(32'hba43ebc8),
	.w3(32'h384946fc),
	.w4(32'hba24bc04),
	.w5(32'hb9aba7b2),
	.w6(32'hbae3f75d),
	.w7(32'hba781fd4),
	.w8(32'hbad21bca),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a274d62),
	.w1(32'h3a4762bb),
	.w2(32'h3a47f2fb),
	.w3(32'h3aea85ee),
	.w4(32'h3ac959aa),
	.w5(32'h3a838f15),
	.w6(32'h3a516fc8),
	.w7(32'h3a736261),
	.w8(32'h3aace602),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6365b5),
	.w1(32'hbb1c1e43),
	.w2(32'hbafd25a0),
	.w3(32'hbabf15a1),
	.w4(32'hba64a79e),
	.w5(32'hba755ba3),
	.w6(32'hbb112169),
	.w7(32'hbad3ab1e),
	.w8(32'hba2204e2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83534a),
	.w1(32'hbb8ca91d),
	.w2(32'hbb8ba811),
	.w3(32'hbaeb8549),
	.w4(32'hbb347c57),
	.w5(32'hbb32d314),
	.w6(32'hbb18cd2f),
	.w7(32'hbb032b0f),
	.w8(32'hba796b44),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305a92),
	.w1(32'hbb771db0),
	.w2(32'hbb8ec2f7),
	.w3(32'hbaac067e),
	.w4(32'hbb0e76e1),
	.w5(32'hbb036a17),
	.w6(32'hbb11844d),
	.w7(32'hbb22fea4),
	.w8(32'hbb082ee8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbe149),
	.w1(32'hbb85d541),
	.w2(32'hba9016ab),
	.w3(32'hb615cb74),
	.w4(32'hbaf6bdcf),
	.w5(32'hb9bbfe69),
	.w6(32'hbb6575f5),
	.w7(32'hbac177d3),
	.w8(32'hba6411d9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1d8ef),
	.w1(32'h39ad57f5),
	.w2(32'h3a894db7),
	.w3(32'h39ec7972),
	.w4(32'h36e39d89),
	.w5(32'hb94a3821),
	.w6(32'h3a28f6cd),
	.w7(32'h3acfc9ec),
	.w8(32'h3aa5598b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908df33),
	.w1(32'hb71910f3),
	.w2(32'hb6fe5f62),
	.w3(32'h38d8f384),
	.w4(32'hb794639a),
	.w5(32'hb9540459),
	.w6(32'h3765ffc3),
	.w7(32'h3884e1e5),
	.w8(32'h39128536),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b1c8b),
	.w1(32'h39b803f5),
	.w2(32'h389aa3c8),
	.w3(32'h398680bd),
	.w4(32'h39b93771),
	.w5(32'hb9c79eab),
	.w6(32'h39d91d87),
	.w7(32'h39ca4142),
	.w8(32'h39f8834b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995598c),
	.w1(32'hba153c7c),
	.w2(32'h3a475243),
	.w3(32'h3a27b081),
	.w4(32'hb9a3c00e),
	.w5(32'h3afc3ff5),
	.w6(32'hba38219d),
	.w7(32'hba4780a1),
	.w8(32'hbacc5d80),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380cb6e5),
	.w1(32'hba9ef50a),
	.w2(32'hba7e217b),
	.w3(32'h3aa47423),
	.w4(32'hb99d9d9a),
	.w5(32'hb9f5dc0c),
	.w6(32'hba511b9d),
	.w7(32'hbad00369),
	.w8(32'h3b2de4de),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74988c),
	.w1(32'hbb037355),
	.w2(32'hbb1501f2),
	.w3(32'h3b483d1d),
	.w4(32'hba4b7283),
	.w5(32'hbade0645),
	.w6(32'hba426ba4),
	.w7(32'hba88a2db),
	.w8(32'h393fd2fe),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96666f),
	.w1(32'h388c8561),
	.w2(32'hbb28aab0),
	.w3(32'h39e375d9),
	.w4(32'h3a24e1f6),
	.w5(32'hbb10bf69),
	.w6(32'hb83212a9),
	.w7(32'hbae69af5),
	.w8(32'hbb0dbfa0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2be31d),
	.w1(32'hba86c3e2),
	.w2(32'hba100477),
	.w3(32'hba8cff02),
	.w4(32'hba365c44),
	.w5(32'hba05ccfb),
	.w6(32'hbaa365e5),
	.w7(32'hba19c164),
	.w8(32'hb8c45f38),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9682940),
	.w1(32'hbb1c5105),
	.w2(32'hbaaf9e90),
	.w3(32'h3a6b6608),
	.w4(32'hbaeb0883),
	.w5(32'h3a3a034e),
	.w6(32'hbb449b5f),
	.w7(32'hbb34b271),
	.w8(32'hbb6e4f4d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb8e05),
	.w1(32'h3b69a4b2),
	.w2(32'h3a6fc71f),
	.w3(32'hba6c2d92),
	.w4(32'h3b97ea18),
	.w5(32'h3acf0b94),
	.w6(32'h3b760139),
	.w7(32'h3aec88eb),
	.w8(32'h3a6081c9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c77e89),
	.w1(32'hba9314f3),
	.w2(32'hbac1c999),
	.w3(32'h35870329),
	.w4(32'hb9afea66),
	.w5(32'hbab15de4),
	.w6(32'h3b24f15c),
	.w7(32'h3ab8c7fc),
	.w8(32'h3a934254),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d0d9c),
	.w1(32'hb5b7e062),
	.w2(32'hb690dda3),
	.w3(32'h3a16cca4),
	.w4(32'hb7301994),
	.w5(32'h36762502),
	.w6(32'hb675e25b),
	.w7(32'hb6241b8c),
	.w8(32'h37068f79),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c79f),
	.w1(32'hbba83ed1),
	.w2(32'hbb479b2c),
	.w3(32'hbb4c6ce9),
	.w4(32'hbb55a620),
	.w5(32'hbb253fe5),
	.w6(32'h3adeb49f),
	.w7(32'h3aa7bcba),
	.w8(32'h38fa625c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule