module layer_10_featuremap_184(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be76b0),
	.w1(32'hb76ebabe),
	.w2(32'hb6802674),
	.w3(32'hb7d383cf),
	.w4(32'hb781d33a),
	.w5(32'hb72b1601),
	.w6(32'hb8657088),
	.w7(32'hb7ecfe43),
	.w8(32'hb795f6bf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3a731),
	.w1(32'hba321e10),
	.w2(32'h3a122f57),
	.w3(32'h3989cde2),
	.w4(32'hbb0b842d),
	.w5(32'h3a3f6be9),
	.w6(32'hbb717d0e),
	.w7(32'hbb94f9fc),
	.w8(32'hbb2c35b9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b9d91e),
	.w1(32'hb74c3099),
	.w2(32'hb7580520),
	.w3(32'hb65ea8e6),
	.w4(32'hb6b2c5cd),
	.w5(32'hb5f377fe),
	.w6(32'hb6c78501),
	.w7(32'hb6c262d2),
	.w8(32'hb6af31b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01800f),
	.w1(32'h39d7e6da),
	.w2(32'h3a1b4e78),
	.w3(32'hb7fe9416),
	.w4(32'h39b95872),
	.w5(32'h3a26ab5e),
	.w6(32'h3a122bc4),
	.w7(32'h38d10f37),
	.w8(32'h39ca82f1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5f5d1),
	.w1(32'hb9c59f3e),
	.w2(32'hb71c9b3e),
	.w3(32'hb9d6d5c9),
	.w4(32'hb9ff7435),
	.w5(32'hb915e675),
	.w6(32'hb9e686f2),
	.w7(32'hba0abad1),
	.w8(32'hb99e21ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b1ce20),
	.w1(32'h383a1fcf),
	.w2(32'h37aa8fe6),
	.w3(32'h3737348b),
	.w4(32'h37bfd08e),
	.w5(32'hb61cae97),
	.w6(32'hb6e60bfb),
	.w7(32'hb720f232),
	.w8(32'hb8552d5b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc445a7e),
	.w1(32'hba87dd39),
	.w2(32'hba3d83ce),
	.w3(32'hbbde1e5c),
	.w4(32'hbad28bc2),
	.w5(32'hbb83bdc9),
	.w6(32'h3bb2785e),
	.w7(32'h3bc7aa2b),
	.w8(32'h3ae35e1d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6edd5e),
	.w1(32'h3b8f1de5),
	.w2(32'hbbd5dbd9),
	.w3(32'hbbbc2bad),
	.w4(32'hbab64028),
	.w5(32'hbbbe1e5b),
	.w6(32'h3c1ce468),
	.w7(32'h3cc1c608),
	.w8(32'h3c697ec5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10fa21),
	.w1(32'h393dfcb3),
	.w2(32'h3a8db2e0),
	.w3(32'hb980c889),
	.w4(32'h39a7b006),
	.w5(32'h3a65836f),
	.w6(32'hb9f232fa),
	.w7(32'hb90ae071),
	.w8(32'h3a2aaf54),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3733e13e),
	.w1(32'hba8944b7),
	.w2(32'hbb4482a2),
	.w3(32'hbb8b8fd9),
	.w4(32'hbb302b21),
	.w5(32'hbba0375a),
	.w6(32'h3ba54984),
	.w7(32'h3bacb3be),
	.w8(32'hba41b337),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d09c9b),
	.w1(32'hba24bc60),
	.w2(32'hb8bb6ca9),
	.w3(32'hb9d9662b),
	.w4(32'hb93784b4),
	.w5(32'hb8d26789),
	.w6(32'hb9fd1e2b),
	.w7(32'hb9899b32),
	.w8(32'hb9652e8d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc353408),
	.w1(32'h3bfab004),
	.w2(32'hbb27126a),
	.w3(32'hbc2eabc7),
	.w4(32'hbac3eab6),
	.w5(32'hbc1db938),
	.w6(32'hba6e50e4),
	.w7(32'h3c0bf05e),
	.w8(32'hb99f10ea),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e558),
	.w1(32'hbac7084a),
	.w2(32'hbb8ef85e),
	.w3(32'hbb27af64),
	.w4(32'hbb0c16cc),
	.w5(32'hbb95e7ef),
	.w6(32'h3b9c4454),
	.w7(32'h3c020085),
	.w8(32'h3b4285ec),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e82b6),
	.w1(32'hbb61ff06),
	.w2(32'hbb92be80),
	.w3(32'hbbc48d16),
	.w4(32'hbc00de4b),
	.w5(32'hbc00bc4e),
	.w6(32'hbb81da2e),
	.w7(32'hbb91f420),
	.w8(32'hbb86c0b6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e87161),
	.w1(32'hba01bf2a),
	.w2(32'h3adf0c52),
	.w3(32'hb79fbfd4),
	.w4(32'hb90357c2),
	.w5(32'h3ad6d6ad),
	.w6(32'hbb0e53a3),
	.w7(32'hbb2a422f),
	.w8(32'hbb29d384),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf72899),
	.w1(32'hbb13136c),
	.w2(32'hba6f7588),
	.w3(32'hb936f648),
	.w4(32'hbbaf92ea),
	.w5(32'hbb9c1563),
	.w6(32'h3b545ea0),
	.w7(32'hbace06ff),
	.w8(32'hbb127870),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8553),
	.w1(32'hb9c93e76),
	.w2(32'hb99e0e94),
	.w3(32'hb853f954),
	.w4(32'h381179e5),
	.w5(32'hb91a3854),
	.w6(32'hb8b118e1),
	.w7(32'hb881bf02),
	.w8(32'hb9b15cc4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad266a6),
	.w1(32'h3b0b227b),
	.w2(32'hbb18760e),
	.w3(32'h3b9f64a3),
	.w4(32'h3a75d054),
	.w5(32'hbc2a29c3),
	.w6(32'h3c64c086),
	.w7(32'h3c5fc8d2),
	.w8(32'h3c04b817),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3b9c8),
	.w1(32'h39bece3a),
	.w2(32'hbb2141a4),
	.w3(32'h3b126168),
	.w4(32'h3ab36ac3),
	.w5(32'hbb881b40),
	.w6(32'h3beaac40),
	.w7(32'h3c0bd2a2),
	.w8(32'h3b8ba24e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d568b9),
	.w1(32'h38174641),
	.w2(32'hb80ea78f),
	.w3(32'hb8ee7f37),
	.w4(32'h382b62cd),
	.w5(32'hb83c5dcb),
	.w6(32'hb84feef2),
	.w7(32'hb754cb80),
	.w8(32'h37f2029e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f8bb55),
	.w1(32'h395da79c),
	.w2(32'hb9580a5b),
	.w3(32'hb8901145),
	.w4(32'h39b45b37),
	.w5(32'h37e0e41e),
	.w6(32'hb9089d9a),
	.w7(32'h38dba521),
	.w8(32'hb7d92761),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20651),
	.w1(32'hbabe8953),
	.w2(32'hba45315f),
	.w3(32'hbab8948e),
	.w4(32'hba93b571),
	.w5(32'h3938f7b5),
	.w6(32'hbb3e777f),
	.w7(32'hbb253531),
	.w8(32'hbaa39691),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b91d2),
	.w1(32'h3bbc5c28),
	.w2(32'hba3c5d15),
	.w3(32'hbab8f966),
	.w4(32'hbb347145),
	.w5(32'hb933d04a),
	.w6(32'h3c7c0470),
	.w7(32'h3c09c132),
	.w8(32'h39f0a830),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0c566),
	.w1(32'hbae02d9c),
	.w2(32'hbb2681b5),
	.w3(32'hba50428b),
	.w4(32'h3a5b8c02),
	.w5(32'hba0866b6),
	.w6(32'h3b0df945),
	.w7(32'h3b1b2ac4),
	.w8(32'hb8a8871b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60e497),
	.w1(32'hbb6bc12f),
	.w2(32'h391b66f8),
	.w3(32'h3b6fcc9c),
	.w4(32'hbb129906),
	.w5(32'h3badbe2e),
	.w6(32'hbbf312ec),
	.w7(32'hbbf8c5f4),
	.w8(32'hbb192cbc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dc7af),
	.w1(32'hba917d7f),
	.w2(32'hba5b92a0),
	.w3(32'hb954ccc9),
	.w4(32'hba07107b),
	.w5(32'hb99aa2f6),
	.w6(32'h38f49d75),
	.w7(32'hb9a454c6),
	.w8(32'hb9b6fc33),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8631da6),
	.w1(32'h37ca220e),
	.w2(32'hb8511e57),
	.w3(32'hb7895bde),
	.w4(32'h3677fc03),
	.w5(32'hb848e837),
	.w6(32'hb959433e),
	.w7(32'hb8f6a2bb),
	.w8(32'hb91ad471),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f5e5c),
	.w1(32'h3bcff622),
	.w2(32'h3bfaaafe),
	.w3(32'hb927c7ac),
	.w4(32'h3b56b0f9),
	.w5(32'h3b64b8c3),
	.w6(32'hbc40792d),
	.w7(32'hbbbd1b43),
	.w8(32'hbb827ef6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8c193),
	.w1(32'hba4f22bb),
	.w2(32'hbac1cbe7),
	.w3(32'hba3194a7),
	.w4(32'hbaa78d41),
	.w5(32'hbad6bc66),
	.w6(32'hbaa3d1cf),
	.w7(32'hbab289eb),
	.w8(32'hbac50596),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92afb1),
	.w1(32'hbb8c0861),
	.w2(32'h3b019ad9),
	.w3(32'hbb276223),
	.w4(32'hbab9208b),
	.w5(32'h3bddf001),
	.w6(32'hbc503be0),
	.w7(32'hbc10a701),
	.w8(32'hbb868b86),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8487b5b),
	.w1(32'hb7cf3803),
	.w2(32'hb86d9e18),
	.w3(32'hb803ac00),
	.w4(32'hb783d17d),
	.w5(32'hb7e78893),
	.w6(32'hb871892a),
	.w7(32'hb81c2730),
	.w8(32'hb875333e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37657168),
	.w1(32'h38342116),
	.w2(32'hb8d6ce8a),
	.w3(32'h38885ce5),
	.w4(32'h3779ef9e),
	.w5(32'hb91fd021),
	.w6(32'hb77ba06d),
	.w7(32'hb8eff0c8),
	.w8(32'hb99ea6c9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7cf70),
	.w1(32'hb9e6dfd9),
	.w2(32'hba184956),
	.w3(32'hbaa10229),
	.w4(32'hbaaf024f),
	.w5(32'hbb43f454),
	.w6(32'h3b26c908),
	.w7(32'h3b1ba7c9),
	.w8(32'h3988de56),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a45bdc),
	.w1(32'hba786085),
	.w2(32'h3a97631d),
	.w3(32'hba8f4aaa),
	.w4(32'hbb0e2ea4),
	.w5(32'h3ac4410e),
	.w6(32'hbb849416),
	.w7(32'hbb7763b0),
	.w8(32'hba48cf92),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d0f9f),
	.w1(32'h3a72e278),
	.w2(32'hb9d461d7),
	.w3(32'hb9fb2340),
	.w4(32'h39b6ed8c),
	.w5(32'hba7d8028),
	.w6(32'hba0c624a),
	.w7(32'h390e58ef),
	.w8(32'hba636e43),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0eb26),
	.w1(32'hba3fc0a2),
	.w2(32'hbb504b7b),
	.w3(32'hbb332cdf),
	.w4(32'h39d6b747),
	.w5(32'hbaf22900),
	.w6(32'h3b4262c4),
	.w7(32'h3b51157c),
	.w8(32'h3b6fcad4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5069b7),
	.w1(32'h3cbbae59),
	.w2(32'hbc3e7441),
	.w3(32'hbcbc65c4),
	.w4(32'h3c15e01c),
	.w5(32'hbbfe1595),
	.w6(32'hbc42af0b),
	.w7(32'h3c45e02b),
	.w8(32'hbc2fbcab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b271042),
	.w1(32'h39c2fdaa),
	.w2(32'hbae00499),
	.w3(32'h3bbd1b3f),
	.w4(32'h3b33b75d),
	.w5(32'h3bf97ac2),
	.w6(32'hbb265f0d),
	.w7(32'hbbd0f08a),
	.w8(32'hbb652a1c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c6bc8),
	.w1(32'hbc03a9a7),
	.w2(32'hbbc11b14),
	.w3(32'hbb82edea),
	.w4(32'hbb785c87),
	.w5(32'h3b6df7d2),
	.w6(32'hbc6d6d9d),
	.w7(32'hbc359025),
	.w8(32'hbb4d881f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4b62d),
	.w1(32'h3aac3574),
	.w2(32'h3a1aad0f),
	.w3(32'h3a716e74),
	.w4(32'h3ae4ac78),
	.w5(32'h3a556ad5),
	.w6(32'hbadc5a58),
	.w7(32'hba8a0c9f),
	.w8(32'hbac6667e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979614b),
	.w1(32'h392157f0),
	.w2(32'hb62ea32f),
	.w3(32'h398b1bca),
	.w4(32'h397104c4),
	.w5(32'h39088cfa),
	.w6(32'h391b2256),
	.w7(32'hb6f9beb2),
	.w8(32'hb6a6930f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b238b),
	.w1(32'h3978e8f9),
	.w2(32'hb7ba6ef0),
	.w3(32'hb68d9d9e),
	.w4(32'hb7de01f8),
	.w5(32'hb851dde4),
	.w6(32'hb98d4e2e),
	.w7(32'hb8b18224),
	.w8(32'hb88a74a8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bab62),
	.w1(32'hba9e0451),
	.w2(32'hbb118a8b),
	.w3(32'hba4755eb),
	.w4(32'hbae6c391),
	.w5(32'hbac158cd),
	.w6(32'h38e7ca2f),
	.w7(32'hba0b44e3),
	.w8(32'hba15d7b4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada0424),
	.w1(32'hba9dafb2),
	.w2(32'hbb8b27e1),
	.w3(32'h3b85230c),
	.w4(32'hb9be1a25),
	.w5(32'hbc297f3a),
	.w6(32'h3b966481),
	.w7(32'h3bd255d0),
	.w8(32'hbb315730),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ffad2),
	.w1(32'hbab37ae6),
	.w2(32'hbaa7c733),
	.w3(32'h3b4d8c7d),
	.w4(32'h3a587f64),
	.w5(32'h3b258896),
	.w6(32'hba706906),
	.w7(32'hbaaed90c),
	.w8(32'hba38620f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a033937),
	.w1(32'hbb135318),
	.w2(32'hbbfe3c88),
	.w3(32'h3b261cde),
	.w4(32'h3b33d7c8),
	.w5(32'h3a92d790),
	.w6(32'h3afeb377),
	.w7(32'h3bb84f25),
	.w8(32'h3a3a9374),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73a6b9),
	.w1(32'hba97d9ff),
	.w2(32'hbaa2f786),
	.w3(32'h3986e4f3),
	.w4(32'hbac9d0da),
	.w5(32'hba86303d),
	.w6(32'h3b1a44c4),
	.w7(32'h39fcc8d7),
	.w8(32'hb9c41ee2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13e72b),
	.w1(32'h3aeef281),
	.w2(32'hbb6b1256),
	.w3(32'hbb47efa4),
	.w4(32'hb7430ba2),
	.w5(32'hbc1e0878),
	.w6(32'h3c666149),
	.w7(32'h3c716014),
	.w8(32'h3c0c2215),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36929090),
	.w1(32'hb8174a26),
	.w2(32'h373a6982),
	.w3(32'hb888cdbb),
	.w4(32'hb8f551d9),
	.w5(32'hb915dcee),
	.w6(32'hb86a32af),
	.w7(32'hb97cc646),
	.w8(32'hb9849eb8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4861ab),
	.w1(32'h39f911c0),
	.w2(32'h3aa0f790),
	.w3(32'h3a658517),
	.w4(32'h3a8a3b22),
	.w5(32'h3aee57be),
	.w6(32'h3a96c5ae),
	.w7(32'h3acc1fb4),
	.w8(32'h3b1957fa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f3b81),
	.w1(32'hb9bbeb1f),
	.w2(32'h385e6a0a),
	.w3(32'hba211816),
	.w4(32'hba26986d),
	.w5(32'hb78e0809),
	.w6(32'hb9d6a00c),
	.w7(32'hb9b6c6bf),
	.w8(32'h393eff31),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06ea73),
	.w1(32'hba56745b),
	.w2(32'hbb0612dd),
	.w3(32'h3ac495ac),
	.w4(32'h3a33108a),
	.w5(32'hb992b184),
	.w6(32'h3b068405),
	.w7(32'h3b4afc13),
	.w8(32'h3a03f5f7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980179a),
	.w1(32'h3990c11e),
	.w2(32'h3a658f28),
	.w3(32'hb9e08ed7),
	.w4(32'hb9674a03),
	.w5(32'hb8b128a0),
	.w6(32'hb923a6a6),
	.w7(32'h3a4fd8d7),
	.w8(32'h3ac2fe4d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a913e2e),
	.w1(32'h3bbef9d4),
	.w2(32'h38c1c95e),
	.w3(32'h3b1575bd),
	.w4(32'hb97b35de),
	.w5(32'hbc56c593),
	.w6(32'h3c58add7),
	.w7(32'h3c6b45d6),
	.w8(32'h3b708cc7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a997aec),
	.w1(32'h3912d8c8),
	.w2(32'hbb29f703),
	.w3(32'h3a0221b7),
	.w4(32'h3a776609),
	.w5(32'hbaa606ac),
	.w6(32'hba9259e4),
	.w7(32'h3ad86d9d),
	.w8(32'h3b2b1040),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d062b),
	.w1(32'hb98d1380),
	.w2(32'hb917fc49),
	.w3(32'hb91080c6),
	.w4(32'hb9e11323),
	.w5(32'hb82eaada),
	.w6(32'hb9df1717),
	.w7(32'hba1d2c27),
	.w8(32'hb9b23976),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37110e3c),
	.w1(32'h37f5a67a),
	.w2(32'h3763cf13),
	.w3(32'hb5ff5731),
	.w4(32'h35a51dd7),
	.w5(32'h375e4d58),
	.w6(32'hb8c76875),
	.w7(32'hb887346d),
	.w8(32'hb8a33f7e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d2ff2),
	.w1(32'hb9b3e40b),
	.w2(32'h38789ba6),
	.w3(32'hb9d8967b),
	.w4(32'h3a8972a5),
	.w5(32'h3a74585c),
	.w6(32'hb9dcb52e),
	.w7(32'hb98904a3),
	.w8(32'h38a9425a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b57e80),
	.w1(32'hba0f5025),
	.w2(32'hba56a5a1),
	.w3(32'hba0026c8),
	.w4(32'hba126665),
	.w5(32'hba079276),
	.w6(32'hba7236a4),
	.w7(32'hba262e82),
	.w8(32'hba1b1e56),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba132417),
	.w1(32'hb981d52b),
	.w2(32'hb9939801),
	.w3(32'hba739404),
	.w4(32'hba28e062),
	.w5(32'hba21f6b1),
	.w6(32'h39fe4a29),
	.w7(32'h395e85bb),
	.w8(32'h399c09b0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba577ac8),
	.w1(32'h38651285),
	.w2(32'hbaca332b),
	.w3(32'hb94094b7),
	.w4(32'hb9fb6010),
	.w5(32'hbb96708d),
	.w6(32'h3b832691),
	.w7(32'h3b474a66),
	.w8(32'h3a3e33e7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a0ff4),
	.w1(32'h3a07ab2c),
	.w2(32'hbb0303b3),
	.w3(32'h3b3f50ea),
	.w4(32'hbb3b5130),
	.w5(32'hbbbbbeed),
	.w6(32'hba069363),
	.w7(32'hba9a3cf3),
	.w8(32'h39da3c75),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d8be62),
	.w1(32'h38213ce8),
	.w2(32'hb7df1042),
	.w3(32'h38711441),
	.w4(32'hb5fb80ee),
	.w5(32'hb886802f),
	.w6(32'h35885b56),
	.w7(32'hb805b7f0),
	.w8(32'hb896196d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377880b9),
	.w1(32'h37443da0),
	.w2(32'h3784f0d3),
	.w3(32'h37e935af),
	.w4(32'h37f43f29),
	.w5(32'h3811a9dc),
	.w6(32'h365eb48c),
	.w7(32'h37304c6c),
	.w8(32'hb6fc5fe3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bef158),
	.w1(32'hb839f89a),
	.w2(32'hb8f1b145),
	.w3(32'hb878d2c1),
	.w4(32'h37156de2),
	.w5(32'hb8868348),
	.w6(32'hb8c96077),
	.w7(32'hb8a6a226),
	.w8(32'hb90e52d5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b30a65),
	.w1(32'h37eaa643),
	.w2(32'hb83419da),
	.w3(32'h3729079d),
	.w4(32'h384ffeb1),
	.w5(32'hb80512db),
	.w6(32'hb8a02713),
	.w7(32'hb80f974f),
	.w8(32'hb8af4b99),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84f53d),
	.w1(32'h3c0554ba),
	.w2(32'hbb16f47f),
	.w3(32'hbb036c33),
	.w4(32'hbc1cf2ee),
	.w5(32'hbc743043),
	.w6(32'hbbc46c9f),
	.w7(32'hb98b6982),
	.w8(32'hbc1ac602),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857f95),
	.w1(32'hbbdde965),
	.w2(32'hbc6289af),
	.w3(32'h3b926250),
	.w4(32'h3a3646ec),
	.w5(32'hbaa08388),
	.w6(32'h3b6ee873),
	.w7(32'h3bc911be),
	.w8(32'h3c00cc5e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac520a6),
	.w1(32'hbb01c4c5),
	.w2(32'hbb2bec41),
	.w3(32'h3b4b2cdf),
	.w4(32'hbac173cc),
	.w5(32'hbb769275),
	.w6(32'h3b84f069),
	.w7(32'h3b271786),
	.w8(32'h3bc6cb9e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabe327),
	.w1(32'hbb6ecf3d),
	.w2(32'hba9ced1c),
	.w3(32'h3b83ab41),
	.w4(32'h39b36d85),
	.w5(32'h3bf95754),
	.w6(32'hbb8499d8),
	.w7(32'hbb81a959),
	.w8(32'h397c6715),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8020849),
	.w1(32'h37a742d4),
	.w2(32'hb85392c9),
	.w3(32'h37dcefff),
	.w4(32'h389bfeb2),
	.w5(32'h3779940a),
	.w6(32'h37a418d4),
	.w7(32'h3886d642),
	.w8(32'h37d9f344),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3631ac13),
	.w1(32'h363318bb),
	.w2(32'hb7a13c42),
	.w3(32'h378b9ae3),
	.w4(32'h381509fc),
	.w5(32'h36e8c261),
	.w6(32'hb886d975),
	.w7(32'hb80d932e),
	.w8(32'hb816c5c4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815c699),
	.w1(32'h38cb5f43),
	.w2(32'hb5d135da),
	.w3(32'h38b3b5ee),
	.w4(32'h392337c3),
	.w5(32'h38a16c64),
	.w6(32'h3862b397),
	.w7(32'h38f8f62a),
	.w8(32'h37c1151a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9946313),
	.w1(32'h39e5ec13),
	.w2(32'hbab42fa4),
	.w3(32'hb892adf6),
	.w4(32'hba0d2d05),
	.w5(32'hbb59afde),
	.w6(32'h3aadaafc),
	.w7(32'h3b554c53),
	.w8(32'h3ad0f4b2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881dcd8),
	.w1(32'h3909610e),
	.w2(32'h377e7342),
	.w3(32'hb87a9620),
	.w4(32'h3739ad2d),
	.w5(32'hb7e698b6),
	.w6(32'hb8c9d4fd),
	.w7(32'hb8361881),
	.w8(32'hb88cf906),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02f902),
	.w1(32'h3bb663ba),
	.w2(32'h393bc001),
	.w3(32'hbb853105),
	.w4(32'h3a1a1027),
	.w5(32'hbbb1f9ce),
	.w6(32'h3ba1de2a),
	.w7(32'h3c017e9a),
	.w8(32'h3b2946f6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1351e5),
	.w1(32'h3b41d124),
	.w2(32'hba7e2d09),
	.w3(32'hbab3aaea),
	.w4(32'h3ba8eb24),
	.w5(32'hbbd27739),
	.w6(32'h3c0a142c),
	.w7(32'h3c516c8c),
	.w8(32'h3bdbe4ab),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad87a0a),
	.w1(32'hbaabda00),
	.w2(32'hbac01fd0),
	.w3(32'h3a430dc3),
	.w4(32'hba11b7de),
	.w5(32'h3b224336),
	.w6(32'hbb2e24e5),
	.w7(32'hbb4d401c),
	.w8(32'hbafef8f3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ee58),
	.w1(32'h3a97eb05),
	.w2(32'h3a92069a),
	.w3(32'hba32c8be),
	.w4(32'hbb1b8a78),
	.w5(32'hbb427b46),
	.w6(32'h3a6157bf),
	.w7(32'h3a2dd9c6),
	.w8(32'h393784e7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae99e95),
	.w1(32'h3ba25b01),
	.w2(32'hbb2d1180),
	.w3(32'hbb87168b),
	.w4(32'h3a02b6d7),
	.w5(32'hbb91d165),
	.w6(32'hbb037394),
	.w7(32'h3a494fa6),
	.w8(32'hbbb58937),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae86e0b),
	.w1(32'hbb244cf3),
	.w2(32'hbac1bebb),
	.w3(32'h3aabd303),
	.w4(32'hba2b6a73),
	.w5(32'hba395491),
	.w6(32'hba2d6bd2),
	.w7(32'h3ac901ea),
	.w8(32'h39e0a53c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b4ef8),
	.w1(32'h3ac763d6),
	.w2(32'hb9c351a4),
	.w3(32'hbae9d210),
	.w4(32'hb99ffb53),
	.w5(32'hbb2929a4),
	.w6(32'h3b8680c6),
	.w7(32'h3bb35ccc),
	.w8(32'h3b35ba73),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38291b1f),
	.w1(32'h38126506),
	.w2(32'h376c4f06),
	.w3(32'h380de4ae),
	.w4(32'h380b5a69),
	.w5(32'h36e1e09e),
	.w6(32'h36fe697e),
	.w7(32'h36fde619),
	.w8(32'hb740635e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e704f1),
	.w1(32'hb809bbaa),
	.w2(32'hb7c492f7),
	.w3(32'hb849731d),
	.w4(32'hb85a047d),
	.w5(32'h36da791a),
	.w6(32'hb88bbe54),
	.w7(32'hb8381d5e),
	.w8(32'hb784f2e9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5fc26),
	.w1(32'hb8c079d4),
	.w2(32'hb94a4b0e),
	.w3(32'hb95ffdb5),
	.w4(32'hb9061365),
	.w5(32'hb8e31202),
	.w6(32'hb98bde9e),
	.w7(32'hb91e1adb),
	.w8(32'hb933f43d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba808b29),
	.w1(32'hb97ec913),
	.w2(32'h36bfe986),
	.w3(32'hb9f680b7),
	.w4(32'h3866954a),
	.w5(32'h399c6649),
	.w6(32'hba8e88f4),
	.w7(32'hb9bc9c54),
	.w8(32'hb9824d6b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99c0af),
	.w1(32'h3ac5acc0),
	.w2(32'hb80b8444),
	.w3(32'h3ac80265),
	.w4(32'h39ed4d42),
	.w5(32'h3ad11e0c),
	.w6(32'hbb0d4fdc),
	.w7(32'hba778699),
	.w8(32'hbb09120a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a4d4),
	.w1(32'hb9189e56),
	.w2(32'hb9db28e4),
	.w3(32'hb6e24e2a),
	.w4(32'hb8525938),
	.w5(32'hb9ea45e8),
	.w6(32'hb9ab0bbc),
	.w7(32'hba008b42),
	.w8(32'hba1f53db),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa4309),
	.w1(32'h39b17c12),
	.w2(32'hbb010b4e),
	.w3(32'h3ac5aec3),
	.w4(32'h39db83e2),
	.w5(32'h3b04bed5),
	.w6(32'hb9b66cc1),
	.w7(32'h3a5fe6f8),
	.w8(32'h3b22f10d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb249bb9),
	.w1(32'h3b47dfe3),
	.w2(32'hba8be0d6),
	.w3(32'h3b5960ad),
	.w4(32'h3b0d3bd9),
	.w5(32'hbbddc75f),
	.w6(32'h3c591c21),
	.w7(32'h3c5e5f40),
	.w8(32'h3bec170a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd057e),
	.w1(32'hbbb14ccc),
	.w2(32'hbb3927d1),
	.w3(32'hbb23067d),
	.w4(32'hbb345ea0),
	.w5(32'h3ae61459),
	.w6(32'hbb61d0dd),
	.w7(32'hbb328cda),
	.w8(32'hb7dc58f5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9b49),
	.w1(32'h3b8c9437),
	.w2(32'hbb8452bc),
	.w3(32'hbc28fa7c),
	.w4(32'hbbcefbec),
	.w5(32'hbc0e5e97),
	.w6(32'h3c10802a),
	.w7(32'h3abf04a8),
	.w8(32'hbc2336a0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb224468),
	.w1(32'h39b8297d),
	.w2(32'hbaeba1fb),
	.w3(32'h3af8cf7c),
	.w4(32'h3bb962c6),
	.w5(32'h3bb25c71),
	.w6(32'h3b838ee0),
	.w7(32'h3bca7109),
	.w8(32'h3bc2dadd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c367033),
	.w1(32'h3bb5b6c4),
	.w2(32'h3ba2d154),
	.w3(32'h3b124f95),
	.w4(32'hbb64b8e9),
	.w5(32'hbbefeff7),
	.w6(32'h3bcdb2a8),
	.w7(32'h3aad6401),
	.w8(32'h3aa2d9f6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7d397),
	.w1(32'h37f9bb06),
	.w2(32'hba2b2b9d),
	.w3(32'hba482043),
	.w4(32'hbb9d4f40),
	.w5(32'hbac698c1),
	.w6(32'hbb0ad2f0),
	.w7(32'hbb7d84e7),
	.w8(32'hbbb887d5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa28fe3),
	.w1(32'h3a841458),
	.w2(32'h3b55fdc6),
	.w3(32'h3a61779e),
	.w4(32'h3a939251),
	.w5(32'h3b4c0694),
	.w6(32'hbbbe545c),
	.w7(32'hbbab63a1),
	.w8(32'hbb95fb93),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ced82a),
	.w1(32'hba941e77),
	.w2(32'hb9cbeb01),
	.w3(32'hba3f5022),
	.w4(32'hba73d120),
	.w5(32'h38c7d5a4),
	.w6(32'hbaa4c154),
	.w7(32'hba2636f3),
	.w8(32'hb8e71c7b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e3768),
	.w1(32'hba772917),
	.w2(32'hbacf603d),
	.w3(32'hb84a2322),
	.w4(32'hb9ffbe00),
	.w5(32'hbb95a547),
	.w6(32'h3c011028),
	.w7(32'h3c0b6184),
	.w8(32'h3b97f6b6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e2bfe),
	.w1(32'h3c4bc29c),
	.w2(32'hba31523a),
	.w3(32'hbbcd2aad),
	.w4(32'hb88a33fd),
	.w5(32'hbbce4029),
	.w6(32'h3b8865e2),
	.w7(32'h3bc25b87),
	.w8(32'h38d3420e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7f809),
	.w1(32'h3bcffaac),
	.w2(32'hbc1be7d9),
	.w3(32'hbc1e3f72),
	.w4(32'h3bc2c1bb),
	.w5(32'hbb845a0b),
	.w6(32'h39afe3dc),
	.w7(32'h3c228c1d),
	.w8(32'hba13e88a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54cd5f),
	.w1(32'h3ab5045b),
	.w2(32'h3b7d01c3),
	.w3(32'h3a70604b),
	.w4(32'h3a0b32dc),
	.w5(32'h3b9b6887),
	.w6(32'hbba9a439),
	.w7(32'hbb50e59c),
	.w8(32'h390e1208),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801bf6),
	.w1(32'hbb243ebf),
	.w2(32'hbb0d3d62),
	.w3(32'h3b10fabb),
	.w4(32'h3a6eb530),
	.w5(32'h3b93a978),
	.w6(32'hba84fa90),
	.w7(32'hb8fd5ee6),
	.w8(32'h3aaea07a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc028ef0),
	.w1(32'h3c0f4c41),
	.w2(32'hbbab1527),
	.w3(32'hbc5b59d0),
	.w4(32'hbb596044),
	.w5(32'hbc216a62),
	.w6(32'hbad56f8f),
	.w7(32'h3b1edbb9),
	.w8(32'hbbaa7859),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81220d),
	.w1(32'hbabd2b3e),
	.w2(32'hbab54c6d),
	.w3(32'hba5b5c5a),
	.w4(32'hbac293b8),
	.w5(32'hbb1b17c9),
	.w6(32'hba742cbb),
	.w7(32'hbadb6533),
	.w8(32'hbae7f1f3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3517fc),
	.w1(32'h3c363bb4),
	.w2(32'h3bc3a6bf),
	.w3(32'hbc35a8f9),
	.w4(32'h3c1dac33),
	.w5(32'h3922fa7e),
	.w6(32'h3a55fce5),
	.w7(32'h3c4d91c5),
	.w8(32'h3b668fb0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf9f7f),
	.w1(32'hb9efc3ca),
	.w2(32'h3a474936),
	.w3(32'hbc0996da),
	.w4(32'hbad47349),
	.w5(32'hbafd7269),
	.w6(32'hb9a14122),
	.w7(32'h3aa022bd),
	.w8(32'hbac4cbbf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8acccb2),
	.w1(32'h38064e1f),
	.w2(32'h38dd26c1),
	.w3(32'hb9a70617),
	.w4(32'hb945df08),
	.w5(32'h36ad264a),
	.w6(32'hba43e8f0),
	.w7(32'hb9daffe1),
	.w8(32'hb964b752),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6a11b),
	.w1(32'hba788c4b),
	.w2(32'h38d0a29e),
	.w3(32'h3a9ea8a3),
	.w4(32'hb9208e07),
	.w5(32'h3affd5a2),
	.w6(32'h3aed74e0),
	.w7(32'hba76e9bf),
	.w8(32'h39c262e8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb344dc6),
	.w1(32'hbb2d93f2),
	.w2(32'hbb8792cb),
	.w3(32'hbaf0c48f),
	.w4(32'hba2240b2),
	.w5(32'hbb56a27c),
	.w6(32'h3b8977a6),
	.w7(32'h3b8c4b88),
	.w8(32'h3953cca5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabeb870),
	.w1(32'hbb0421d4),
	.w2(32'hb97cea2e),
	.w3(32'h3aeccbc7),
	.w4(32'h3a21e7e4),
	.w5(32'h3b891e5a),
	.w6(32'hbb28e92a),
	.w7(32'hbb0fb7c5),
	.w8(32'hb9d33d71),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7397b8),
	.w1(32'hbb459cac),
	.w2(32'h3adf4c84),
	.w3(32'h3947428f),
	.w4(32'hbaf2859d),
	.w5(32'h3b0f5957),
	.w6(32'hbb6e37fb),
	.w7(32'hbb0f69bd),
	.w8(32'hba84a11e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd13f3),
	.w1(32'hba368a69),
	.w2(32'h3a051758),
	.w3(32'h39b0b656),
	.w4(32'hba95190b),
	.w5(32'h3ae79abf),
	.w6(32'hbaa29ef6),
	.w7(32'hbaf0bf0c),
	.w8(32'h3a479e98),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadace13),
	.w1(32'hb9f94b8c),
	.w2(32'hbbd0194c),
	.w3(32'h3ba87a08),
	.w4(32'h3af5d731),
	.w5(32'hbbba32b1),
	.w6(32'h3c066d21),
	.w7(32'h3b6db2e9),
	.w8(32'h3b29beef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10a6d8),
	.w1(32'hbad88f72),
	.w2(32'hb97dbcf4),
	.w3(32'hbafc7b48),
	.w4(32'hbba3abff),
	.w5(32'hbbb278a0),
	.w6(32'hb9d4fb34),
	.w7(32'hbbae65c5),
	.w8(32'hbbe4f939),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c3fc0),
	.w1(32'hba338dce),
	.w2(32'hbae99cbb),
	.w3(32'h3a84f501),
	.w4(32'h3a67178b),
	.w5(32'h3a83537e),
	.w6(32'h3a27194a),
	.w7(32'h3a4623f7),
	.w8(32'h39d3cc89),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39648b0d),
	.w1(32'h3910cb0b),
	.w2(32'h389e9640),
	.w3(32'h395623dd),
	.w4(32'h3936e93c),
	.w5(32'h38e70d33),
	.w6(32'h38f71b8f),
	.w7(32'h383c46c1),
	.w8(32'h38bed8e8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0e6f3),
	.w1(32'hba0aac55),
	.w2(32'h372d216c),
	.w3(32'hba160ce5),
	.w4(32'hbac59331),
	.w5(32'hb9cf8f8b),
	.w6(32'hb9893d61),
	.w7(32'hba48e22f),
	.w8(32'hb9cdb689),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7934f08),
	.w1(32'h370988b1),
	.w2(32'hb72c2556),
	.w3(32'h37a4c649),
	.w4(32'h37fc4d4e),
	.w5(32'h370040b0),
	.w6(32'hb74f37bd),
	.w7(32'h355a8fef),
	.w8(32'hb67606ac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22835a),
	.w1(32'hba263b1e),
	.w2(32'hba7f38a3),
	.w3(32'hba04df08),
	.w4(32'hba5800c1),
	.w5(32'hba7d0f64),
	.w6(32'hb9d28f35),
	.w7(32'hb9d037dc),
	.w8(32'hb99c42c4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89ab15),
	.w1(32'hbb3a7fc6),
	.w2(32'hbb76418c),
	.w3(32'hb9c33870),
	.w4(32'hba1c9934),
	.w5(32'h396a9564),
	.w6(32'hb8b3eac5),
	.w7(32'h394f5ac6),
	.w8(32'hba0877eb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9921547),
	.w1(32'h390e30cb),
	.w2(32'h3976cda8),
	.w3(32'hb9e695ef),
	.w4(32'hba27fcd6),
	.w5(32'hba0c3e6d),
	.w6(32'hba332cb4),
	.w7(32'hba5b6be2),
	.w8(32'hba0d95ba),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39959458),
	.w1(32'h3b5c61cc),
	.w2(32'hba4dbee5),
	.w3(32'hbaf943ba),
	.w4(32'h3a2c39d6),
	.w5(32'hbb5ae795),
	.w6(32'h3b7907c4),
	.w7(32'h3bae5526),
	.w8(32'h3b227cba),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a4b92),
	.w1(32'hba33ad17),
	.w2(32'h3adbf64c),
	.w3(32'h3ac3e483),
	.w4(32'hb981947c),
	.w5(32'h3b9fa65f),
	.w6(32'hbbb750c4),
	.w7(32'hbbaca844),
	.w8(32'hbb0cb900),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849918b),
	.w1(32'hb8559b6d),
	.w2(32'h383298c2),
	.w3(32'hb80f30b5),
	.w4(32'hb86951bc),
	.w5(32'h3800e2e6),
	.w6(32'hb8aec5a3),
	.w7(32'hb84034a6),
	.w8(32'hb8b6a258),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37deef75),
	.w1(32'hb90be0c3),
	.w2(32'hb91dc58a),
	.w3(32'hb885693f),
	.w4(32'hb951ca58),
	.w5(32'hb62981ef),
	.w6(32'hb8fdf76a),
	.w7(32'hb924aba4),
	.w8(32'h3921adf8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c9e19),
	.w1(32'h37140585),
	.w2(32'hb87fd8be),
	.w3(32'hb80883cf),
	.w4(32'hb769b353),
	.w5(32'hb888fa1e),
	.w6(32'hb865d075),
	.w7(32'hb810b51d),
	.w8(32'hb8afc84c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e6a92),
	.w1(32'hbb4def0f),
	.w2(32'hba326f07),
	.w3(32'hba01373b),
	.w4(32'hbb04541a),
	.w5(32'hba466669),
	.w6(32'hbaa35bb8),
	.w7(32'hb995cacc),
	.w8(32'hba84b31a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc448200),
	.w1(32'hbad237a6),
	.w2(32'hbc31b2c0),
	.w3(32'hba9dce05),
	.w4(32'h3ba062fe),
	.w5(32'hbc2d82a5),
	.w6(32'h3c77f57f),
	.w7(32'h3c3eef6d),
	.w8(32'h3c291eb9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eee25b),
	.w1(32'h3a0d19f5),
	.w2(32'h3b11cdae),
	.w3(32'h3ac962fa),
	.w4(32'hbb35382b),
	.w5(32'hbbf92a48),
	.w6(32'h3bfa6dd7),
	.w7(32'h3c54f31a),
	.w8(32'h3c15e5e6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066806),
	.w1(32'h3ab0ff3c),
	.w2(32'h3b05c28f),
	.w3(32'h3b387bd3),
	.w4(32'h3a34f884),
	.w5(32'h3a339325),
	.w6(32'h3b05f27b),
	.w7(32'h3b1f497c),
	.w8(32'h399849c2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e2ecd),
	.w1(32'h3a058d90),
	.w2(32'hbb22b629),
	.w3(32'h3b2af009),
	.w4(32'h3ad88ac6),
	.w5(32'hb973254b),
	.w6(32'h3ac3b577),
	.w7(32'h3a764ef6),
	.w8(32'h39ca90ef),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0bd37),
	.w1(32'h3a9e9630),
	.w2(32'hba38d9e2),
	.w3(32'h3ac1337d),
	.w4(32'h3b7a0e9c),
	.w5(32'h3b041311),
	.w6(32'h3b1dac0f),
	.w7(32'hba5f397c),
	.w8(32'hbb2ade87),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a0f6e),
	.w1(32'h3ba48cd6),
	.w2(32'h3b8e8a00),
	.w3(32'hb9f0d175),
	.w4(32'h3b8d5145),
	.w5(32'h3b011c6a),
	.w6(32'h3be5ce47),
	.w7(32'h3b56c3fe),
	.w8(32'h3a6aa09f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1743d8),
	.w1(32'h3b5cae48),
	.w2(32'h3b161c5d),
	.w3(32'h3bbe6812),
	.w4(32'h3a59429c),
	.w5(32'h39bda06b),
	.w6(32'hbaeaefc4),
	.w7(32'hbb853563),
	.w8(32'hbb42cb45),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbcef3),
	.w1(32'h3bfb5e5e),
	.w2(32'h3b00cd3f),
	.w3(32'hbb277159),
	.w4(32'h38aa9aad),
	.w5(32'hbbf13cce),
	.w6(32'h3c427343),
	.w7(32'h3c654761),
	.w8(32'h3b046bea),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684ced),
	.w1(32'h3b0d1e25),
	.w2(32'h39f4b507),
	.w3(32'h3b139bd8),
	.w4(32'h3b2cba09),
	.w5(32'h3b156883),
	.w6(32'hbb005a99),
	.w7(32'hbb111eb5),
	.w8(32'hba5e860e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24b69),
	.w1(32'h39512e5d),
	.w2(32'hbaaeaf63),
	.w3(32'h3ae64fc1),
	.w4(32'hba8425e1),
	.w5(32'hbb349093),
	.w6(32'h3bb76a01),
	.w7(32'hbaba69fa),
	.w8(32'h39a02d53),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42410a),
	.w1(32'h3b7c9f54),
	.w2(32'h3a9f57a9),
	.w3(32'h3a87e31e),
	.w4(32'h397ce3e7),
	.w5(32'hbbcb7339),
	.w6(32'h3c0d1e40),
	.w7(32'h3c07aee7),
	.w8(32'h3b55bf23),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9359a6),
	.w1(32'hbad88d72),
	.w2(32'hbb89a9fa),
	.w3(32'h3b3146e6),
	.w4(32'h3b176f85),
	.w5(32'h3aa1fa87),
	.w6(32'hb8aebda2),
	.w7(32'h38f5f713),
	.w8(32'hbacd8bcf),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba970d98),
	.w1(32'h3b20bcf6),
	.w2(32'hba8dcf5c),
	.w3(32'hbb3e082b),
	.w4(32'hbaccfca2),
	.w5(32'hbb9a0679),
	.w6(32'h3c0066ad),
	.w7(32'h3bc387fe),
	.w8(32'h396bb823),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eea1cf),
	.w1(32'hba7cf4f9),
	.w2(32'hba80f23b),
	.w3(32'h39613141),
	.w4(32'h3a00b9dd),
	.w5(32'h39a9c62f),
	.w6(32'hba05e1df),
	.w7(32'hba2192c3),
	.w8(32'hb9b480a0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9a45),
	.w1(32'h3a0139a5),
	.w2(32'h3b3eb1ae),
	.w3(32'hbb98a523),
	.w4(32'h3b1514c8),
	.w5(32'h3bef35cb),
	.w6(32'hbc12ff1d),
	.w7(32'hbaea5bd5),
	.w8(32'h3bb82fc4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b912673),
	.w1(32'h3baa4c01),
	.w2(32'h3c1203cc),
	.w3(32'h3b812cbb),
	.w4(32'h3b6f0b03),
	.w5(32'h3bc4e7df),
	.w6(32'h3c2aaf7d),
	.w7(32'h3bc21e8d),
	.w8(32'h38951686),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34686a),
	.w1(32'h39d1a4bc),
	.w2(32'hbac49d63),
	.w3(32'h3b085faf),
	.w4(32'h3a95363a),
	.w5(32'hba36d30c),
	.w6(32'h3986361f),
	.w7(32'hba9009e3),
	.w8(32'h38b5e6a9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b80ef),
	.w1(32'hbaa03e23),
	.w2(32'h3adb6f98),
	.w3(32'h3968a87c),
	.w4(32'hbb44aac3),
	.w5(32'hb9be2ab3),
	.w6(32'hbadd313b),
	.w7(32'h3aa39d42),
	.w8(32'hba632463),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f07fb6),
	.w1(32'h3b1e2521),
	.w2(32'h3b5e42dc),
	.w3(32'hbb685d7a),
	.w4(32'h3ace8ce9),
	.w5(32'h3ac29de2),
	.w6(32'hb9b2ae21),
	.w7(32'h39c72182),
	.w8(32'h39e61df6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24be17),
	.w1(32'h3ac08327),
	.w2(32'h3b6bc0cb),
	.w3(32'h3ade01d1),
	.w4(32'h3b174b2c),
	.w5(32'h3aaaa8ae),
	.w6(32'h3a39d5f6),
	.w7(32'hb94b716d),
	.w8(32'h3a8c44a2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3946b4),
	.w1(32'hba83d5ff),
	.w2(32'hbba56035),
	.w3(32'hbaa34cc8),
	.w4(32'hba12c389),
	.w5(32'hbb84c45f),
	.w6(32'h3a22ea63),
	.w7(32'h3a6f8f79),
	.w8(32'h3a797ca5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38841667),
	.w1(32'hba7adcf4),
	.w2(32'hbb4ef039),
	.w3(32'h39a7bb47),
	.w4(32'h38fa56ae),
	.w5(32'hbb08cd0f),
	.w6(32'h39a24204),
	.w7(32'hbaf4b82a),
	.w8(32'hbaf16b46),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90a073),
	.w1(32'h3b6f130d),
	.w2(32'hbb9388a9),
	.w3(32'hbb7ff6aa),
	.w4(32'h3b144252),
	.w5(32'hbb2a60e8),
	.w6(32'h3b037be4),
	.w7(32'h3c13f48c),
	.w8(32'h3b0bed7d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ef19a),
	.w1(32'h3aa5035a),
	.w2(32'h3ae238f7),
	.w3(32'hb6f8d617),
	.w4(32'h3b5ae2f5),
	.w5(32'h3b491140),
	.w6(32'h3b91c3ba),
	.w7(32'h3beac184),
	.w8(32'h3b33ae71),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51e89f),
	.w1(32'h3b73a55c),
	.w2(32'hbb32ec82),
	.w3(32'hbba81c89),
	.w4(32'hbb3fcf32),
	.w5(32'hbbb429ff),
	.w6(32'h3c06d566),
	.w7(32'h3bb3a974),
	.w8(32'h3ab5a2c5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6937),
	.w1(32'h3b1554b5),
	.w2(32'h3b0313b3),
	.w3(32'h3baae0a8),
	.w4(32'h3bab1e03),
	.w5(32'h3c3a451f),
	.w6(32'hbb13731e),
	.w7(32'hba8d87ae),
	.w8(32'h3af0914d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25ad5),
	.w1(32'h38ad07e8),
	.w2(32'h3b540379),
	.w3(32'hba6bdcbe),
	.w4(32'hbb6d6076),
	.w5(32'hb994edcb),
	.w6(32'hbb1c857b),
	.w7(32'hbb7b63e7),
	.w8(32'hbb10c7f2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf75223),
	.w1(32'h39d63d3f),
	.w2(32'hbaf147be),
	.w3(32'hbb504f7d),
	.w4(32'hba4ce8ad),
	.w5(32'hbb143fee),
	.w6(32'hbab10af3),
	.w7(32'hbb1d66a5),
	.w8(32'hbaca71cb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3323f2),
	.w1(32'hba71b388),
	.w2(32'hba775e82),
	.w3(32'h3b06e980),
	.w4(32'h3b192930),
	.w5(32'h3b2edf55),
	.w6(32'h3ad278a7),
	.w7(32'h3a73f670),
	.w8(32'h3b1c66a0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ac08),
	.w1(32'h3a4c51f2),
	.w2(32'hba518f2f),
	.w3(32'h3b0d45b8),
	.w4(32'hb997afe5),
	.w5(32'hbac50b93),
	.w6(32'h3a87e8b6),
	.w7(32'h3a46bf85),
	.w8(32'hb9d732b8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafda1ab),
	.w1(32'hbb327650),
	.w2(32'hbb112cd5),
	.w3(32'hbac5d10b),
	.w4(32'hbb6b840c),
	.w5(32'hbada7ade),
	.w6(32'hbbce40c2),
	.w7(32'hbb8c856b),
	.w8(32'hbb724e7c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf547e6),
	.w1(32'h3a951247),
	.w2(32'hbad08f23),
	.w3(32'hbb69ab4c),
	.w4(32'h3895c798),
	.w5(32'hbb111a53),
	.w6(32'h3b356d97),
	.w7(32'h3a815d57),
	.w8(32'h39748a7c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9ef8a),
	.w1(32'hb9a5e39c),
	.w2(32'hba333bf2),
	.w3(32'hba976e72),
	.w4(32'hb8979b4a),
	.w5(32'h38ec5ebe),
	.w6(32'hb8873bb8),
	.w7(32'hba25f9cd),
	.w8(32'hb9352ca7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bbfb2),
	.w1(32'h3a82da79),
	.w2(32'h39d04cc8),
	.w3(32'hb9a89d24),
	.w4(32'h3a16907f),
	.w5(32'hbb96eac9),
	.w6(32'h3bacc751),
	.w7(32'h3b2726ce),
	.w8(32'hb9a05add),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94027d),
	.w1(32'hbb6d2d24),
	.w2(32'h3c608e94),
	.w3(32'hbb940988),
	.w4(32'hbb768368),
	.w5(32'h3c18cd39),
	.w6(32'hbb079445),
	.w7(32'h3c22b67a),
	.w8(32'hb98b8470),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f0e67),
	.w1(32'hb9b1cb4c),
	.w2(32'h3b01ab62),
	.w3(32'h3b451e6f),
	.w4(32'h3b40de13),
	.w5(32'h3b2e7e3d),
	.w6(32'h3abe500d),
	.w7(32'h3acc57aa),
	.w8(32'h3b8e04a3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395af78f),
	.w1(32'h3a58fbee),
	.w2(32'h37f2626d),
	.w3(32'h3990dcdb),
	.w4(32'h3a89ba48),
	.w5(32'hba19faa2),
	.w6(32'h3a83da7b),
	.w7(32'hb916aa74),
	.w8(32'hb96f790b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc021099),
	.w1(32'h3aeba87b),
	.w2(32'h3b3a025e),
	.w3(32'hbbd68a5d),
	.w4(32'h3a8f4c3e),
	.w5(32'hbadd397a),
	.w6(32'h3ad92546),
	.w7(32'h3bb96b14),
	.w8(32'h3b8b58b1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9197b2),
	.w1(32'hb8a90096),
	.w2(32'h3ac1113c),
	.w3(32'h3a7b96a1),
	.w4(32'h391aec91),
	.w5(32'h3a931ffd),
	.w6(32'h3a0956ac),
	.w7(32'h3a952892),
	.w8(32'hba8534ce),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a6ccb),
	.w1(32'h3a0cda79),
	.w2(32'hba320930),
	.w3(32'h38fb87d2),
	.w4(32'h3a843945),
	.w5(32'h377fbb19),
	.w6(32'h3a2a112b),
	.w7(32'hb8d876bb),
	.w8(32'h3a951f84),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a064de9),
	.w1(32'h3977ec8b),
	.w2(32'h3b4ddfa0),
	.w3(32'h3b10d8ac),
	.w4(32'h3a850f70),
	.w5(32'h3b524c52),
	.w6(32'hb970470f),
	.w7(32'hbaa9d05f),
	.w8(32'hbaffe794),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc246588),
	.w1(32'hbba70b8a),
	.w2(32'hbbf03c59),
	.w3(32'h3b3d80d5),
	.w4(32'h3b3ad15f),
	.w5(32'hbae6eb3f),
	.w6(32'h3c444cae),
	.w7(32'h3c86090b),
	.w8(32'h3c0c06ff),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20440c),
	.w1(32'h3a83f86e),
	.w2(32'h380ae6e7),
	.w3(32'hbb7bf9a8),
	.w4(32'h3a96d039),
	.w5(32'hba1ced2d),
	.w6(32'h3a1aab51),
	.w7(32'hb99a1158),
	.w8(32'hb9abb131),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921c4c7),
	.w1(32'hbafb8bb0),
	.w2(32'h3a968fc6),
	.w3(32'h3a752ab7),
	.w4(32'hba5b2709),
	.w5(32'h3b48ca99),
	.w6(32'hbb64f6a7),
	.w7(32'hbb6cdb23),
	.w8(32'hb98951b8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36acce4e),
	.w1(32'hba2be6cd),
	.w2(32'h3ac1b665),
	.w3(32'hb821ef30),
	.w4(32'hbaaced09),
	.w5(32'h3725025d),
	.w6(32'hbb33b6b5),
	.w7(32'hba40eca2),
	.w8(32'hbb10ba07),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd86b25),
	.w1(32'hbb9d22e3),
	.w2(32'hbba85831),
	.w3(32'h3b089e4c),
	.w4(32'hbb629589),
	.w5(32'hbc10bcf7),
	.w6(32'h3a13c31f),
	.w7(32'h3af8bcdd),
	.w8(32'hbb3386e3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66810f),
	.w1(32'hba4681c4),
	.w2(32'h3ab99ecf),
	.w3(32'hba836914),
	.w4(32'hbb1d7519),
	.w5(32'hba44a816),
	.w6(32'hb9ff7026),
	.w7(32'hb9da0b24),
	.w8(32'h3a9fafef),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31fefd),
	.w1(32'h3b342ccc),
	.w2(32'h3b2fe81f),
	.w3(32'h3b93b94c),
	.w4(32'h3b620964),
	.w5(32'hbae23712),
	.w6(32'h3c7051b4),
	.w7(32'h3c418fec),
	.w8(32'h3b74ad63),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab59839),
	.w1(32'hbab9767a),
	.w2(32'h3acfcffb),
	.w3(32'h3b186ce3),
	.w4(32'hbaae3945),
	.w5(32'h3aab99a3),
	.w6(32'h3a1e8f1d),
	.w7(32'h3b2f020f),
	.w8(32'h3a0f9bef),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87155b),
	.w1(32'h38fcbec8),
	.w2(32'h3a17533d),
	.w3(32'hba37d0c3),
	.w4(32'hbb497b48),
	.w5(32'hbb086054),
	.w6(32'hbb01e99e),
	.w7(32'hbb4e563e),
	.w8(32'hbb4e373c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f78ea7),
	.w1(32'h3a560ba6),
	.w2(32'hba574ea8),
	.w3(32'h388e98a6),
	.w4(32'h3a6f9c12),
	.w5(32'hb953f1e9),
	.w6(32'h3aa663a8),
	.w7(32'h397e63f4),
	.w8(32'h3a9a4173),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab56431),
	.w1(32'hba130568),
	.w2(32'h3ac6a9cc),
	.w3(32'h3ac2c11b),
	.w4(32'hba1d1c73),
	.w5(32'h39385db0),
	.w6(32'h3b0fb1f3),
	.w7(32'h3b5994db),
	.w8(32'h3ada8a44),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad643a2),
	.w1(32'hbab39d6e),
	.w2(32'h39c6b06c),
	.w3(32'h3b396d3c),
	.w4(32'hb9fbb880),
	.w5(32'h3b10461e),
	.w6(32'h39fd3e39),
	.w7(32'h3a877f73),
	.w8(32'h3c3578d9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c608600),
	.w1(32'hb8a78a9c),
	.w2(32'hba0b5ed1),
	.w3(32'h3b1a5788),
	.w4(32'hbb49d9e7),
	.w5(32'hbb4f2cd6),
	.w6(32'h3ab12589),
	.w7(32'hbb3c780f),
	.w8(32'hbb9952b2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae84027),
	.w1(32'h3be60b60),
	.w2(32'h3ba16ada),
	.w3(32'hba448bc8),
	.w4(32'h3bd1d6cf),
	.w5(32'h3b88ec58),
	.w6(32'h3bf39fd5),
	.w7(32'h3a9df779),
	.w8(32'hb9101bb8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b3ad6),
	.w1(32'hba585c61),
	.w2(32'h3a89f584),
	.w3(32'h3b340d55),
	.w4(32'hba8d38cc),
	.w5(32'hb9bafa90),
	.w6(32'hba435703),
	.w7(32'h39450885),
	.w8(32'hbad9e699),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a89f2),
	.w1(32'h3a5325e1),
	.w2(32'hbba07d21),
	.w3(32'h3a9a8f69),
	.w4(32'h3b6188bd),
	.w5(32'hbb4f6ca1),
	.w6(32'h3b3a5b96),
	.w7(32'hba4ffb99),
	.w8(32'h3a68c032),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb045798),
	.w1(32'hbb2ba146),
	.w2(32'hbb99c051),
	.w3(32'hbc499117),
	.w4(32'hbb8e56f6),
	.w5(32'hb9b460d1),
	.w6(32'hbb7ca382),
	.w7(32'h3b9b901f),
	.w8(32'hbaaa75f0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354881),
	.w1(32'h3c287578),
	.w2(32'h3bfe8905),
	.w3(32'hbbc342b0),
	.w4(32'h3bbf9d8b),
	.w5(32'hb89f1728),
	.w6(32'h3bb636ca),
	.w7(32'h3bd210c3),
	.w8(32'h3b1a1c4f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194e45),
	.w1(32'h3af88276),
	.w2(32'h3b17f4ec),
	.w3(32'h3bc538aa),
	.w4(32'h3a8e5d2a),
	.w5(32'h3b200c6b),
	.w6(32'h3ad6e171),
	.w7(32'h3b275172),
	.w8(32'h3abf4e3d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ab729),
	.w1(32'hba921532),
	.w2(32'hbb99f0e7),
	.w3(32'hb89f7d0b),
	.w4(32'h3b32871c),
	.w5(32'hbbb46b74),
	.w6(32'h3c40cbd6),
	.w7(32'h3c33404c),
	.w8(32'h3c2338ba),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87b88e),
	.w1(32'h3ae4c5ef),
	.w2(32'h3b014d71),
	.w3(32'h3be64058),
	.w4(32'hbb6e96de),
	.w5(32'h39ae6673),
	.w6(32'hbbded343),
	.w7(32'hba22aaf1),
	.w8(32'hbb6c34a7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d878b),
	.w1(32'h3b228067),
	.w2(32'hbabee122),
	.w3(32'hbaeb46cc),
	.w4(32'h3a51b9e8),
	.w5(32'hbac25143),
	.w6(32'h3b0725b9),
	.w7(32'h3b55f1bf),
	.w8(32'h3b001fb2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1a339),
	.w1(32'hbae108c8),
	.w2(32'h3acfa1f9),
	.w3(32'h3aa62a82),
	.w4(32'hbb4830f2),
	.w5(32'hba73eec4),
	.w6(32'hbad1819e),
	.w7(32'h3a89994b),
	.w8(32'h3b2b0e26),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b752f),
	.w1(32'hb8e2b93d),
	.w2(32'h3a82d7f6),
	.w3(32'hba013114),
	.w4(32'hb9a9d561),
	.w5(32'h39df5d33),
	.w6(32'h3a745ac2),
	.w7(32'h3a9a3d2f),
	.w8(32'h3a8e1c4f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b917dc),
	.w1(32'h39bd3874),
	.w2(32'h3a85dba7),
	.w3(32'h3a04b305),
	.w4(32'h3a822325),
	.w5(32'h39b851a5),
	.w6(32'h3a826920),
	.w7(32'h3913d00d),
	.w8(32'h385d4383),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb4ea),
	.w1(32'h3a062278),
	.w2(32'h3afbc5f9),
	.w3(32'hbb72bb25),
	.w4(32'hba9ce9d7),
	.w5(32'hbaee2acf),
	.w6(32'h3b8e245e),
	.w7(32'h3bfbdeaf),
	.w8(32'h3b21e0e7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9abca8),
	.w1(32'h3a74f393),
	.w2(32'hba87d5d9),
	.w3(32'h3b5a9d5d),
	.w4(32'hb8f4d405),
	.w5(32'hbb146b58),
	.w6(32'h3b09b34a),
	.w7(32'h3b8bb195),
	.w8(32'h3a543aa0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb592701),
	.w1(32'hbab199e0),
	.w2(32'h3bc8ecd5),
	.w3(32'hbb173869),
	.w4(32'hbac92617),
	.w5(32'h3bd8269f),
	.w6(32'hbbece882),
	.w7(32'h3acd6883),
	.w8(32'hbbdd4cc5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3794a3),
	.w1(32'h3a04f381),
	.w2(32'hbadbdb56),
	.w3(32'hbb130d8f),
	.w4(32'h3adc21dd),
	.w5(32'h3782b3dd),
	.w6(32'h3ae39aec),
	.w7(32'h3984bfa2),
	.w8(32'h3a19dc18),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb383d1a),
	.w1(32'hbb49a1bb),
	.w2(32'h398a5ac4),
	.w3(32'hba93932a),
	.w4(32'hbb190814),
	.w5(32'hbb12b608),
	.w6(32'h3beb8595),
	.w7(32'h3bec8f37),
	.w8(32'h3ba3ef7b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22449b),
	.w1(32'hbaa58cef),
	.w2(32'h38d0112c),
	.w3(32'h3b04cb91),
	.w4(32'h3ac2892f),
	.w5(32'h3b1e6337),
	.w6(32'hbaf0efbe),
	.w7(32'h3a65b8ad),
	.w8(32'h3a8d15ad),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d98842),
	.w1(32'h39400904),
	.w2(32'hb9ab0d60),
	.w3(32'h3a68f9f3),
	.w4(32'h3a8c4690),
	.w5(32'hb94ae5c4),
	.w6(32'h39ea8c72),
	.w7(32'hb983964c),
	.w8(32'h391fa232),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cc486),
	.w1(32'h3b0824bb),
	.w2(32'hba96ab0c),
	.w3(32'hb98cf1ee),
	.w4(32'hbad0b84d),
	.w5(32'hbb12e60b),
	.w6(32'h3a589fa8),
	.w7(32'hba372d2d),
	.w8(32'h3a4c39ed),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2dbca),
	.w1(32'h398bf742),
	.w2(32'hba61ab19),
	.w3(32'h3a7b2849),
	.w4(32'h3a255116),
	.w5(32'hba36d98d),
	.w6(32'h3a0095a9),
	.w7(32'hba14183d),
	.w8(32'hb9881b5c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae59fd5),
	.w1(32'h39974c16),
	.w2(32'h3982fa04),
	.w3(32'h3a4e149b),
	.w4(32'h3ab786da),
	.w5(32'h38cca402),
	.w6(32'h3b831563),
	.w7(32'h3b3c8866),
	.w8(32'h3ac72666),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeb027),
	.w1(32'h3b03598e),
	.w2(32'h38299157),
	.w3(32'h3b28d4f0),
	.w4(32'hbb385476),
	.w5(32'h3a1490e3),
	.w6(32'h3ad12123),
	.w7(32'hbaaaa18d),
	.w8(32'hb942de86),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d7173),
	.w1(32'h38455c61),
	.w2(32'hbb150fe1),
	.w3(32'hbb0871c6),
	.w4(32'h3a906c1b),
	.w5(32'h3a274773),
	.w6(32'h39ac70d7),
	.w7(32'hba27432a),
	.w8(32'h3ac04f4f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49451a),
	.w1(32'hbb05d647),
	.w2(32'hbad4e7c5),
	.w3(32'h3a67ef99),
	.w4(32'hbb1c44ef),
	.w5(32'hbae8649b),
	.w6(32'hbade4752),
	.w7(32'hba8de546),
	.w8(32'h3a3e8914),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2430a3),
	.w1(32'hbaca74d9),
	.w2(32'h3b4ca639),
	.w3(32'hba4764cf),
	.w4(32'hba981532),
	.w5(32'h3b4d9095),
	.w6(32'hbba2a14d),
	.w7(32'hbb4abc9d),
	.w8(32'hbb1966f6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68838ee),
	.w1(32'h3a324b5a),
	.w2(32'hbb4348aa),
	.w3(32'hbabeb6de),
	.w4(32'hb6904a9e),
	.w5(32'hbba47f5e),
	.w6(32'h3b928353),
	.w7(32'h3ad4ce5a),
	.w8(32'hbab0681a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d5b79),
	.w1(32'hbaba3e81),
	.w2(32'h3ad0fde8),
	.w3(32'hbafda9b4),
	.w4(32'h3a8eab18),
	.w5(32'h3af926e6),
	.w6(32'h3b06275c),
	.w7(32'h3c3c470f),
	.w8(32'hbac9e482),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ced65),
	.w1(32'h3ad8d0aa),
	.w2(32'h3b23ec10),
	.w3(32'hbb05afcc),
	.w4(32'h3ae00213),
	.w5(32'h3b2c3e3e),
	.w6(32'h3b2410a6),
	.w7(32'h3b448a78),
	.w8(32'h3a53e2b8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9680b6),
	.w1(32'hb9a033cc),
	.w2(32'hba4fbfdd),
	.w3(32'h3ae34d90),
	.w4(32'hb98373c4),
	.w5(32'hba60f0f3),
	.w6(32'h37f3c242),
	.w7(32'hba274288),
	.w8(32'h38564329),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff30a3),
	.w1(32'hbb5c7746),
	.w2(32'hbc1fc03b),
	.w3(32'h3b02aff0),
	.w4(32'h3bb8a212),
	.w5(32'hb900b73e),
	.w6(32'h3b2da878),
	.w7(32'h3bf2716e),
	.w8(32'h3b4467b2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189493),
	.w1(32'hbbc76511),
	.w2(32'h3b354d6c),
	.w3(32'h3ab9f414),
	.w4(32'h3a189ea8),
	.w5(32'h3c037a2f),
	.w6(32'h3bdc5ec3),
	.w7(32'h3c6690bf),
	.w8(32'h3ba2c8a1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c6497),
	.w1(32'hbb4e1fce),
	.w2(32'hbbb65315),
	.w3(32'h393e0c45),
	.w4(32'hba9a125b),
	.w5(32'hba5c2406),
	.w6(32'hbad713a9),
	.w7(32'hba7485a6),
	.w8(32'hbb398282),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d820),
	.w1(32'h3bf00a3f),
	.w2(32'hbb59484a),
	.w3(32'hbc03f6f6),
	.w4(32'hbb5ed1ed),
	.w5(32'hbbf715a1),
	.w6(32'hbc04c344),
	.w7(32'hbaabcf47),
	.w8(32'hbc005a6a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8e00),
	.w1(32'hb9891754),
	.w2(32'hba8ab690),
	.w3(32'h3ab80a2f),
	.w4(32'hba174b74),
	.w5(32'hba827f1d),
	.w6(32'h3ab75631),
	.w7(32'hbaa5bbeb),
	.w8(32'hbae275a0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37b558),
	.w1(32'hbace54c0),
	.w2(32'hba97167a),
	.w3(32'h3a03f417),
	.w4(32'hba7e1f61),
	.w5(32'hbaafcecb),
	.w6(32'hb9d92a01),
	.w7(32'hba7e7830),
	.w8(32'hbb10aaed),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d967c),
	.w1(32'h3baa4272),
	.w2(32'hbc2f755d),
	.w3(32'hbbe57ced),
	.w4(32'h3c0f4f3a),
	.w5(32'hbb7884cd),
	.w6(32'h3b7fe00c),
	.w7(32'h3ca551fe),
	.w8(32'h3c1c2e46),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52a58d),
	.w1(32'h3a380fe0),
	.w2(32'hbb9cf1f3),
	.w3(32'h3b411001),
	.w4(32'h3b50c95f),
	.w5(32'hbbde50e9),
	.w6(32'h3c4e3423),
	.w7(32'h3c27a7f4),
	.w8(32'h3bd4057c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc264b30),
	.w1(32'h3b406512),
	.w2(32'hb765caaf),
	.w3(32'hbbf14bad),
	.w4(32'h37e37cb9),
	.w5(32'hbbb3b597),
	.w6(32'h3b91792f),
	.w7(32'h3b867731),
	.w8(32'hb9d57d98),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d51eda),
	.w1(32'h3a320882),
	.w2(32'h3ab57fb3),
	.w3(32'h3b284b52),
	.w4(32'h3b29d5ee),
	.w5(32'h3bb44759),
	.w6(32'hba0d91c5),
	.w7(32'hba3308df),
	.w8(32'hb95ad0b1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b314798),
	.w1(32'hba510f8f),
	.w2(32'h3b8a9f4e),
	.w3(32'h3b193900),
	.w4(32'h39bd1803),
	.w5(32'h3bd3c2d2),
	.w6(32'hba190c32),
	.w7(32'h3b210037),
	.w8(32'hbb776135),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb066e39),
	.w1(32'h39d0f304),
	.w2(32'h39a6c496),
	.w3(32'hbaca38c6),
	.w4(32'h3aad56b3),
	.w5(32'h3973dd6e),
	.w6(32'h38f75a76),
	.w7(32'hb99238b5),
	.w8(32'hb8b0db2b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba048d50),
	.w1(32'h3b6322a9),
	.w2(32'hba60e794),
	.w3(32'h388c015b),
	.w4(32'h3b4e4f27),
	.w5(32'h3a03e525),
	.w6(32'h3b47f3e1),
	.w7(32'h3a970c3d),
	.w8(32'hb9c9d131),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb577cfb),
	.w1(32'h3988d5bb),
	.w2(32'h3ba90c7b),
	.w3(32'hbaa62cf7),
	.w4(32'hbb18e5d4),
	.w5(32'hbac0fd46),
	.w6(32'h3b8ae5d4),
	.w7(32'h3c10eb15),
	.w8(32'h3b6697c3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ed6c2),
	.w1(32'hbb3ec5aa),
	.w2(32'h39d387bc),
	.w3(32'hba17bc68),
	.w4(32'hbb32835c),
	.w5(32'hbacc990e),
	.w6(32'hbac6f247),
	.w7(32'hb98f25b1),
	.w8(32'h3b38547b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65bb15),
	.w1(32'hbaa5d70b),
	.w2(32'hb98e2322),
	.w3(32'hbb0e67b1),
	.w4(32'hba635734),
	.w5(32'hbac9ac05),
	.w6(32'h3b4e11ee),
	.w7(32'h3b931407),
	.w8(32'h39ff9dbe),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8108e),
	.w1(32'hbafb4d25),
	.w2(32'hbb78942c),
	.w3(32'h3aa5abce),
	.w4(32'h3ab7e404),
	.w5(32'h3a10d082),
	.w6(32'h3bba41bb),
	.w7(32'h3b1c3f5f),
	.w8(32'h39ccb6ed),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05cb43),
	.w1(32'hbb7759a6),
	.w2(32'h3c46c9a8),
	.w3(32'hba8c2a0a),
	.w4(32'hba5504c6),
	.w5(32'h3b7468f3),
	.w6(32'h3bb5e479),
	.w7(32'h3bf23367),
	.w8(32'h3aae7b07),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc037c),
	.w1(32'h3b50d9ce),
	.w2(32'hb89cb4af),
	.w3(32'h3bdaed9e),
	.w4(32'h3b15a284),
	.w5(32'h3a1168fd),
	.w6(32'h3b8bb05c),
	.w7(32'h3aa905c6),
	.w8(32'hba7abe78),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1922d4),
	.w1(32'h3bd37580),
	.w2(32'hbc33fa0e),
	.w3(32'hbbc8bbd8),
	.w4(32'hb88ae9b6),
	.w5(32'hbc46ad17),
	.w6(32'h3c2f9cb0),
	.w7(32'h3c32fb68),
	.w8(32'h3ba1562e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a421817),
	.w1(32'h3af9c35b),
	.w2(32'hb9adac44),
	.w3(32'h3b3d1f51),
	.w4(32'h3b0ed3bc),
	.w5(32'hbb1a1234),
	.w6(32'h3bc5f781),
	.w7(32'h3b988d69),
	.w8(32'h3a8e80ac),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399872bb),
	.w1(32'h3a1ff112),
	.w2(32'hba95f1f8),
	.w3(32'h3aac5784),
	.w4(32'h3a70ac24),
	.w5(32'hb9e48b33),
	.w6(32'h3aa8d1c4),
	.w7(32'hb925aaa6),
	.w8(32'h3ab1f373),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994208f),
	.w1(32'h3b1e3755),
	.w2(32'hbb551727),
	.w3(32'h3b34bff1),
	.w4(32'h3ad87afa),
	.w5(32'hbba460ba),
	.w6(32'h3be3c877),
	.w7(32'h3bbc090e),
	.w8(32'h3b50f577),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b5102),
	.w1(32'h39f3fdcd),
	.w2(32'h38a830a6),
	.w3(32'hba1204da),
	.w4(32'h3ab2db78),
	.w5(32'h3a6e5f2c),
	.w6(32'h3a3638d7),
	.w7(32'h3989ef94),
	.w8(32'hb926be75),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b8de7),
	.w1(32'hbae68418),
	.w2(32'hbb8f5d67),
	.w3(32'h3abd74e7),
	.w4(32'h398ff74e),
	.w5(32'hbada3229),
	.w6(32'h3a266ddb),
	.w7(32'hba4a4647),
	.w8(32'hba9f39a8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb184c5a),
	.w1(32'h3a273018),
	.w2(32'hba930997),
	.w3(32'hbaba1d99),
	.w4(32'h3a502f5f),
	.w5(32'hb9f76b8e),
	.w6(32'h3a987dd4),
	.w7(32'hb7df64ff),
	.w8(32'h3a9185b4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f287f),
	.w1(32'h3915acbb),
	.w2(32'h3a95acf1),
	.w3(32'h3a933e6f),
	.w4(32'h39a705fa),
	.w5(32'h399cf23c),
	.w6(32'h3a315f9e),
	.w7(32'h3acbf7b8),
	.w8(32'h3b024b3d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97cb3),
	.w1(32'h3a9f53e4),
	.w2(32'hbacd0cfd),
	.w3(32'h3b5050cf),
	.w4(32'h3ae805a1),
	.w5(32'h3aa13ee6),
	.w6(32'h3aa7fcfc),
	.w7(32'h3942b56d),
	.w8(32'h3b28fa24),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeb37f),
	.w1(32'hb9cf7fcb),
	.w2(32'h3b0eb1da),
	.w3(32'hbb4c4358),
	.w4(32'hbbdb352a),
	.w5(32'hbbb9460b),
	.w6(32'h39e4a56e),
	.w7(32'h3b79b0c8),
	.w8(32'h3b8e9255),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7013),
	.w1(32'h3b71c86b),
	.w2(32'hba9f886e),
	.w3(32'h3b64724f),
	.w4(32'h3afd1099),
	.w5(32'hbb8f56f8),
	.w6(32'h3be29250),
	.w7(32'h3b971057),
	.w8(32'h3b0a50aa),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae447e),
	.w1(32'h3b985941),
	.w2(32'h3a1227d3),
	.w3(32'hb9dbe850),
	.w4(32'hb9a2826f),
	.w5(32'hbbfdf619),
	.w6(32'h3bbe7db7),
	.w7(32'h3bef9415),
	.w8(32'h394b8c3e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b9da1),
	.w1(32'h39d4632b),
	.w2(32'hb925d3dc),
	.w3(32'h3ae0bdd8),
	.w4(32'h39e23fb3),
	.w5(32'hb790d873),
	.w6(32'hb9ea27f0),
	.w7(32'hba5c3552),
	.w8(32'h3a79046b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6c9c4),
	.w1(32'h3a599068),
	.w2(32'hbae519e3),
	.w3(32'hba2d00f5),
	.w4(32'h39879dd1),
	.w5(32'hbad95568),
	.w6(32'h3aad2453),
	.w7(32'hba3bf7d3),
	.w8(32'h3abddadc),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa176c1),
	.w1(32'h3a93dff3),
	.w2(32'hba187ebe),
	.w3(32'h3ae6608a),
	.w4(32'h3adf5a92),
	.w5(32'h3804b7d3),
	.w6(32'h3a6140d2),
	.w7(32'hba128905),
	.w8(32'h39fd99a4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05268c),
	.w1(32'h3ac54a32),
	.w2(32'hba690b05),
	.w3(32'h3a917fb8),
	.w4(32'h3b0996a2),
	.w5(32'hb921d216),
	.w6(32'h3ac2784c),
	.w7(32'hba633bfb),
	.w8(32'h3a275b86),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6688f7),
	.w1(32'h3a24504a),
	.w2(32'hba9c2afc),
	.w3(32'h39e49276),
	.w4(32'hb90eb210),
	.w5(32'hbb07d5e1),
	.w6(32'hbac8a233),
	.w7(32'h3a2c9121),
	.w8(32'h3a683af8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eadcf),
	.w1(32'h38ee1397),
	.w2(32'h3b3e6a6e),
	.w3(32'h3acceb91),
	.w4(32'h39dc5d41),
	.w5(32'h3b01e4ee),
	.w6(32'h3a9c115d),
	.w7(32'h3abd3ee7),
	.w8(32'h3a347ec9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad98f33),
	.w1(32'h3a3fcdf0),
	.w2(32'hbab67ff2),
	.w3(32'hba7e20b2),
	.w4(32'h3aad8427),
	.w5(32'hbb07bfed),
	.w6(32'hb98e3f88),
	.w7(32'hbb44a767),
	.w8(32'hbb3954fd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37137e),
	.w1(32'hb8832062),
	.w2(32'hbb08cb6a),
	.w3(32'hba859931),
	.w4(32'hbb02739e),
	.w5(32'hbb24fac5),
	.w6(32'hbb4fd928),
	.w7(32'hbb60e016),
	.w8(32'hb90e178f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba548bcc),
	.w1(32'h3a48405a),
	.w2(32'hba22aa71),
	.w3(32'hba4a300d),
	.w4(32'h3a9c7b5b),
	.w5(32'h39bad389),
	.w6(32'h3a62647a),
	.w7(32'h37518c58),
	.w8(32'h3ab98123),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e8df7),
	.w1(32'h3a0403b9),
	.w2(32'hbba13490),
	.w3(32'h3a17c119),
	.w4(32'h3a6e8b48),
	.w5(32'hba9ae71d),
	.w6(32'h3ac46ba3),
	.w7(32'h3b4be6f4),
	.w8(32'h3a6a0bd5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87e2be),
	.w1(32'h3afe7c9e),
	.w2(32'h3a72bab7),
	.w3(32'h3a869963),
	.w4(32'h3ad8fa72),
	.w5(32'h3abb0a38),
	.w6(32'h3a9f10ac),
	.w7(32'hb98e4657),
	.w8(32'hbaeedac5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f78a4),
	.w1(32'h3ae80629),
	.w2(32'hbb929252),
	.w3(32'h3afccb76),
	.w4(32'hbc0efde9),
	.w5(32'hbc7a2021),
	.w6(32'hbb5a2e0a),
	.w7(32'hbba75812),
	.w8(32'hbbeeff8c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac347e2),
	.w1(32'hb81dbfab),
	.w2(32'hb83b832e),
	.w3(32'hba1f3026),
	.w4(32'hb9163023),
	.w5(32'hb9350bed),
	.w6(32'hb9386427),
	.w7(32'hb8ab536e),
	.w8(32'h38352487),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c8d6f),
	.w1(32'hb8a86b01),
	.w2(32'hbbc35670),
	.w3(32'h3be738f4),
	.w4(32'h3b9c9f9b),
	.w5(32'h3a31062e),
	.w6(32'h3b8b48bf),
	.w7(32'h3b28a616),
	.w8(32'h3ba865b9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule