module layer_8_featuremap_181(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c700c1c),
	.w1(32'hbab1ca82),
	.w2(32'h3baef37d),
	.w3(32'h3c3d7213),
	.w4(32'hba44d46f),
	.w5(32'hb956fb3b),
	.w6(32'h3bed961f),
	.w7(32'h3c548568),
	.w8(32'h3c019c98),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c2b48),
	.w1(32'h3c022c7e),
	.w2(32'h3c2fafc9),
	.w3(32'h3b5c35ae),
	.w4(32'h3bdbd147),
	.w5(32'h3c37a919),
	.w6(32'h3b4d3908),
	.w7(32'h3bc26d6c),
	.w8(32'h3a49dc5b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9e255),
	.w1(32'hbcb57fea),
	.w2(32'hbcf43f61),
	.w3(32'h3bd1a234),
	.w4(32'hbca3ad9d),
	.w5(32'hbcc69cdf),
	.w6(32'hbbd4b67f),
	.w7(32'hbc3543f2),
	.w8(32'hbc5ee88b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb74579),
	.w1(32'hbbf91a9e),
	.w2(32'hbbef8b73),
	.w3(32'hbc882975),
	.w4(32'hbc48dbf3),
	.w5(32'hbc94c589),
	.w6(32'h3b318ae1),
	.w7(32'h3c35950f),
	.w8(32'h3c013e5d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c67c94),
	.w1(32'hbc6706d9),
	.w2(32'hbc22ccaa),
	.w3(32'hbc45f203),
	.w4(32'hbc48e6d9),
	.w5(32'hbbf680ad),
	.w6(32'hbc888379),
	.w7(32'hbc6687bf),
	.w8(32'hbc64fba5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e02bd),
	.w1(32'hbb349d25),
	.w2(32'hbcc65bf0),
	.w3(32'hbc009fea),
	.w4(32'hbc33a20e),
	.w5(32'hbcdf04ad),
	.w6(32'h3b816f1c),
	.w7(32'hbb9335b7),
	.w8(32'hbbb90a72),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb92200),
	.w1(32'hbc03d92b),
	.w2(32'hbc2747a4),
	.w3(32'hbcb9314e),
	.w4(32'hbbd09369),
	.w5(32'hbc3e747a),
	.w6(32'hbb8dbe27),
	.w7(32'hbbd21073),
	.w8(32'hbb6442dc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a27b3),
	.w1(32'hb9c5b537),
	.w2(32'h3b080288),
	.w3(32'hbbf5fb65),
	.w4(32'h3a89fa39),
	.w5(32'h3c0605ab),
	.w6(32'h3b26233f),
	.w7(32'hb9383aaf),
	.w8(32'h3b783794),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c247111),
	.w1(32'h3cbbfd51),
	.w2(32'h3d14b82f),
	.w3(32'h3bda82b5),
	.w4(32'h3cb9fe89),
	.w5(32'h3d08ac0e),
	.w6(32'h3c8a6388),
	.w7(32'h3cd5ef5d),
	.w8(32'h3cb2aba5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb88c2),
	.w1(32'hbc4934ec),
	.w2(32'hbc189dd6),
	.w3(32'h3ce20f39),
	.w4(32'h3bf4a42a),
	.w5(32'h3c13ed78),
	.w6(32'hbc506a41),
	.w7(32'hbbe7df6b),
	.w8(32'hbad39fe9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc355e24),
	.w1(32'hbc05a5da),
	.w2(32'h3c40d1cb),
	.w3(32'h3a088513),
	.w4(32'hbc2a655b),
	.w5(32'h3b23e8cb),
	.w6(32'hbbe1293e),
	.w7(32'h3bf213ba),
	.w8(32'h3c89d20c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dee1d),
	.w1(32'hbb12e6b4),
	.w2(32'hbc74263c),
	.w3(32'h3c437ee2),
	.w4(32'hbb6a6dc1),
	.w5(32'hbc1a986c),
	.w6(32'hbab6aa3a),
	.w7(32'hbc14bb72),
	.w8(32'h3abe6308),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a859520),
	.w1(32'h3a7f774f),
	.w2(32'hbb463871),
	.w3(32'hba7cf70d),
	.w4(32'h3b656dc5),
	.w5(32'h3a49cb14),
	.w6(32'h3b225774),
	.w7(32'h3b727a17),
	.w8(32'h3bf74ab9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb412f18),
	.w1(32'hbcd32632),
	.w2(32'hbd24657e),
	.w3(32'hbb8e9562),
	.w4(32'hbc8a82d2),
	.w5(32'hbd059f61),
	.w6(32'hbc9b000a),
	.w7(32'hbcd7967c),
	.w8(32'hbc65894e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbac223),
	.w1(32'hbb23f295),
	.w2(32'hbbff69bd),
	.w3(32'hbcb6a626),
	.w4(32'h3a8f5bb2),
	.w5(32'hbbc8c0c2),
	.w6(32'h3ba1af1e),
	.w7(32'h3a60e721),
	.w8(32'h3b15b178),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6240f),
	.w1(32'hbba11d5f),
	.w2(32'h3aac5da9),
	.w3(32'hbb33ee17),
	.w4(32'hba1f9491),
	.w5(32'h3a8602f7),
	.w6(32'hbbe0478b),
	.w7(32'h3bcf8f6a),
	.w8(32'h3bdcb028),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49a604),
	.w1(32'h3c681511),
	.w2(32'h3cd61895),
	.w3(32'h3c0ff655),
	.w4(32'h3c4327b9),
	.w5(32'h3cc62b44),
	.w6(32'h3c015421),
	.w7(32'h3c431eb1),
	.w8(32'h3b9c4cee),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb920ef),
	.w1(32'hbbc8658b),
	.w2(32'hbc96dc51),
	.w3(32'h3cbb20ac),
	.w4(32'hbb6abb2c),
	.w5(32'hbc67b318),
	.w6(32'hbbecb963),
	.w7(32'hbc133283),
	.w8(32'hbbb87b8b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187a56),
	.w1(32'h3c2740f8),
	.w2(32'hbbd6aa9d),
	.w3(32'hbc1f79e6),
	.w4(32'h3c0a9378),
	.w5(32'hbc48d504),
	.w6(32'hbb422026),
	.w7(32'hbbc97481),
	.w8(32'hbb436642),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4b4f1),
	.w1(32'h3b8d38fd),
	.w2(32'h3af95ada),
	.w3(32'hbc100ac0),
	.w4(32'h3b749666),
	.w5(32'hb85f5155),
	.w6(32'h3c1bafac),
	.w7(32'h3bc0b8b1),
	.w8(32'h3c2ed83b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2593cc),
	.w1(32'hbb5905b1),
	.w2(32'hbc68449a),
	.w3(32'h3b70d4e1),
	.w4(32'hba20d245),
	.w5(32'hbc870778),
	.w6(32'hbb2ae142),
	.w7(32'hbc4afe52),
	.w8(32'hbc06a208),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc696679),
	.w1(32'hbc0bd5af),
	.w2(32'hbc998f67),
	.w3(32'hbc80c867),
	.w4(32'hbc3d1168),
	.w5(32'hbc6c7a67),
	.w6(32'hba48ce79),
	.w7(32'hbbae77be),
	.w8(32'hbc498901),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89c0b6),
	.w1(32'hbc8d75d8),
	.w2(32'hbcd48d43),
	.w3(32'hbbed38a1),
	.w4(32'hbcc1b8e1),
	.w5(32'hbc81e1f6),
	.w6(32'hbba8ccf3),
	.w7(32'hbcc80608),
	.w8(32'hbc80bab8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba31df7),
	.w1(32'h3a95a092),
	.w2(32'hbb6a35c3),
	.w3(32'h3c376c98),
	.w4(32'hbba86e18),
	.w5(32'h3b1f7693),
	.w6(32'h3aae5863),
	.w7(32'hbaa6b4ed),
	.w8(32'hbbd9b565),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69e61),
	.w1(32'h3b96b0de),
	.w2(32'hbb4c55c7),
	.w3(32'hbb23437e),
	.w4(32'hbba7688b),
	.w5(32'hbbe10ae3),
	.w6(32'h3b6f98f9),
	.w7(32'h3a3756b6),
	.w8(32'hbb16c330),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa2ba6),
	.w1(32'h3b615b26),
	.w2(32'hbc26f54b),
	.w3(32'hbac9a728),
	.w4(32'h3b94b704),
	.w5(32'hbadf6430),
	.w6(32'hbb2c34a3),
	.w7(32'hbc07e4c7),
	.w8(32'h39567239),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6535ae),
	.w1(32'h3c7c89cb),
	.w2(32'h3c4398f0),
	.w3(32'hbc2d6c8e),
	.w4(32'h3b964528),
	.w5(32'hb7f34a51),
	.w6(32'h3c26c947),
	.w7(32'h3c3d1293),
	.w8(32'h3bf35192),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc97dea),
	.w1(32'hbbfa3a93),
	.w2(32'hbbd837de),
	.w3(32'hbb12bf67),
	.w4(32'hbbd8b0f7),
	.w5(32'hbb6de9e3),
	.w6(32'h3a67fc7a),
	.w7(32'h3b306ffd),
	.w8(32'h3bcb5c8b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5b2df),
	.w1(32'h3b841298),
	.w2(32'h3c0aaa60),
	.w3(32'hbb2c04ab),
	.w4(32'h3b1cb9ce),
	.w5(32'h3bff2cb6),
	.w6(32'h3b0e5d69),
	.w7(32'h3bfc5976),
	.w8(32'hbac2c725),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49c113),
	.w1(32'hbb214e30),
	.w2(32'h39e85e46),
	.w3(32'hbb21c550),
	.w4(32'hbbbd1077),
	.w5(32'hbb506fa7),
	.w6(32'hbb9f02a7),
	.w7(32'hbbb25f7b),
	.w8(32'h3c0c7c46),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63ce41),
	.w1(32'h3bc1e026),
	.w2(32'h3bf58145),
	.w3(32'h3c421266),
	.w4(32'h3b59fb41),
	.w5(32'h3c250234),
	.w6(32'hba678a83),
	.w7(32'h3b89e778),
	.w8(32'h3b4e8fe1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b7bea),
	.w1(32'h3c27e01a),
	.w2(32'h3c4d27bf),
	.w3(32'h3c017583),
	.w4(32'h3bcfb5e5),
	.w5(32'h3c217f4a),
	.w6(32'h3b9046ce),
	.w7(32'h3bd758f8),
	.w8(32'h3beab2da),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54f817),
	.w1(32'hbc796839),
	.w2(32'hbc9ff860),
	.w3(32'h3bde0e33),
	.w4(32'hbc588a67),
	.w5(32'hbc729789),
	.w6(32'hbc074021),
	.w7(32'hbc342b1c),
	.w8(32'hbba19958),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8da3ee),
	.w1(32'h3c315b5e),
	.w2(32'h3c49b0d7),
	.w3(32'hbc3bef3f),
	.w4(32'h3b7ad226),
	.w5(32'h3c2735db),
	.w6(32'h3b9a9c95),
	.w7(32'h3c1a8c28),
	.w8(32'h3b829dc6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c48a4),
	.w1(32'h3be434a6),
	.w2(32'h3cb3f91a),
	.w3(32'h3c38f062),
	.w4(32'h3ca9bec3),
	.w5(32'h3d1fd18d),
	.w6(32'h3c48c3db),
	.w7(32'h3cd328f5),
	.w8(32'h3ca1623f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a09e8),
	.w1(32'hbc9418e2),
	.w2(32'hbcf0fd96),
	.w3(32'h3cf24c0d),
	.w4(32'hbbabc8d4),
	.w5(32'hbc0ac582),
	.w6(32'hbbd2b417),
	.w7(32'hbbe7220b),
	.w8(32'hb9d5480d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb18b4e),
	.w1(32'h3c02892e),
	.w2(32'h3c853f98),
	.w3(32'hbbc27e07),
	.w4(32'h3bfb8520),
	.w5(32'h3c4f9bb2),
	.w6(32'h3bfcec07),
	.w7(32'h3c7ccc31),
	.w8(32'h3c750a15),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c870dca),
	.w1(32'h3b0cae0e),
	.w2(32'h3b810408),
	.w3(32'h3c4ade64),
	.w4(32'h3b9511f2),
	.w5(32'h3baf365f),
	.w6(32'h3b6de50c),
	.w7(32'h3b7cc714),
	.w8(32'h3b58820f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38e44a),
	.w1(32'hbc2fd7ff),
	.w2(32'hbd04feb8),
	.w3(32'h3b95c459),
	.w4(32'hbb7eb7e3),
	.w5(32'hbcdbfa3d),
	.w6(32'hbb8568fa),
	.w7(32'hbca4d215),
	.w8(32'hbc2be12d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a7493),
	.w1(32'h3ad4c673),
	.w2(32'h3af01cdf),
	.w3(32'hbc4d75ab),
	.w4(32'hb8f57d13),
	.w5(32'h3b52ce59),
	.w6(32'h3a8932f7),
	.w7(32'h3b862111),
	.w8(32'hba5f42ab),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcaf39),
	.w1(32'h3d02f447),
	.w2(32'h3d514162),
	.w3(32'hbae4672b),
	.w4(32'h3ce406ff),
	.w5(32'h3d3d8429),
	.w6(32'h3c9d295a),
	.w7(32'h3d149b51),
	.w8(32'h3cc6b140),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c8e6f),
	.w1(32'h3b30ca74),
	.w2(32'h37c96bb7),
	.w3(32'h3d067f32),
	.w4(32'h3b1f1f54),
	.w5(32'hb9c15f88),
	.w6(32'h3b52d43f),
	.w7(32'h39fcd1d8),
	.w8(32'h3b8ce0f7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87958c),
	.w1(32'hbc023f85),
	.w2(32'hbadf92d2),
	.w3(32'h3be7faad),
	.w4(32'hbb9dca7a),
	.w5(32'hbb9f4c3d),
	.w6(32'hbb5b0eb3),
	.w7(32'h3a207d51),
	.w8(32'h3ba4f93a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3857b),
	.w1(32'hbc967417),
	.w2(32'hbd38fc34),
	.w3(32'h3beb9408),
	.w4(32'hbc6e3d3a),
	.w5(32'hbd1ee24c),
	.w6(32'hbc877a76),
	.w7(32'hbcf5410f),
	.w8(32'hbca4a859),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd77420),
	.w1(32'hbc8e0449),
	.w2(32'hbc779212),
	.w3(32'hbc9fda1b),
	.w4(32'hbc87df5e),
	.w5(32'hbc5f77a3),
	.w6(32'hbb47b2fd),
	.w7(32'hbb87931d),
	.w8(32'hba65017d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62a875),
	.w1(32'h3bcfb6ca),
	.w2(32'h3c52e751),
	.w3(32'hbc2924dd),
	.w4(32'h3b9b531b),
	.w5(32'h3c243911),
	.w6(32'h3bd93a40),
	.w7(32'h3c4ea9fb),
	.w8(32'h3c2615ec),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf60001),
	.w1(32'hbd75e8af),
	.w2(32'hbd9fc2df),
	.w3(32'h3be3136f),
	.w4(32'hbd3e395c),
	.w5(32'hbd8a3446),
	.w6(32'hbd0c8220),
	.w7(32'hbd5ad5c4),
	.w8(32'hbd33ded4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8745a3),
	.w1(32'h3b81b288),
	.w2(32'hbb59e43e),
	.w3(32'hbd5cacfd),
	.w4(32'hbc10c42e),
	.w5(32'hbc7be137),
	.w6(32'h3c03c57f),
	.w7(32'h3a68a2a1),
	.w8(32'h3a6f5b46),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07b1bd),
	.w1(32'hbcacfe6e),
	.w2(32'hbd154d8e),
	.w3(32'hbc31be9e),
	.w4(32'hbca982c4),
	.w5(32'hbcde2505),
	.w6(32'h399eea11),
	.w7(32'hbc7f3546),
	.w8(32'hbc60f933),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb29ea),
	.w1(32'hbcaf36ac),
	.w2(32'hbd2227cd),
	.w3(32'hbc5bd360),
	.w4(32'hbc065f17),
	.w5(32'hbd0010b0),
	.w6(32'hbc8ea352),
	.w7(32'hbcddbfa4),
	.w8(32'hbc27e977),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca5629),
	.w1(32'h3bb482dc),
	.w2(32'h3c3e7808),
	.w3(32'hbd01aff5),
	.w4(32'hbb125f14),
	.w5(32'h3b3722f4),
	.w6(32'hbaa213ee),
	.w7(32'h3b78e6e8),
	.w8(32'hbb42082a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1bd51),
	.w1(32'h3c3b6c3a),
	.w2(32'hbb33d743),
	.w3(32'hbb37d1ea),
	.w4(32'h3b7513fe),
	.w5(32'hbb3f8421),
	.w6(32'h3c533b12),
	.w7(32'h3bc71c93),
	.w8(32'h3bb7b528),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90275),
	.w1(32'hbb4fcd05),
	.w2(32'h3bc489a1),
	.w3(32'h3a755899),
	.w4(32'hbbb03f08),
	.w5(32'h3b2b1399),
	.w6(32'hbace80af),
	.w7(32'h3b398c3d),
	.w8(32'hbb9e6b21),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5c36b),
	.w1(32'h3c4dd3ee),
	.w2(32'h3c0910cf),
	.w3(32'hbbaed412),
	.w4(32'h3c1f0ec7),
	.w5(32'h3c1be16a),
	.w6(32'h3c047ab9),
	.w7(32'h3bb3cd3d),
	.w8(32'hbb6931a4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c08c),
	.w1(32'h3b081f74),
	.w2(32'hbc0daa6a),
	.w3(32'hbbaf8bc1),
	.w4(32'h3b96d21d),
	.w5(32'hbbd4bcd2),
	.w6(32'hbbd354ff),
	.w7(32'hbc0f748b),
	.w8(32'hbc40c9f8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0136b3),
	.w1(32'hbc4ae399),
	.w2(32'hbc9852f9),
	.w3(32'hbc1317d9),
	.w4(32'hbc120508),
	.w5(32'hbca9997f),
	.w6(32'hbc073c3b),
	.w7(32'hbc6fa037),
	.w8(32'hbbaf3b84),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc695ec1),
	.w1(32'hbc2f8482),
	.w2(32'hbc5f8c38),
	.w3(32'hbc847ec2),
	.w4(32'hbc8fd22b),
	.w5(32'hbc09446e),
	.w6(32'hbb215538),
	.w7(32'hbc065e06),
	.w8(32'hbb37dac0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc9f9d),
	.w1(32'h3bd30f27),
	.w2(32'h3c2d11e6),
	.w3(32'h3c3d615c),
	.w4(32'h3c1a5e46),
	.w5(32'h3c2eeb07),
	.w6(32'h3bb93fe6),
	.w7(32'h3c259d16),
	.w8(32'h3bc272e2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c279558),
	.w1(32'hba8d5aa4),
	.w2(32'hbaba9242),
	.w3(32'h3c26d03d),
	.w4(32'hbb31fa8e),
	.w5(32'hbb8cf048),
	.w6(32'hba483ba3),
	.w7(32'hbaa81bb0),
	.w8(32'hba97fd0e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36c6ab),
	.w1(32'h3b3c5a66),
	.w2(32'hbc4ceee7),
	.w3(32'hbaf8e5d3),
	.w4(32'hbc47b217),
	.w5(32'hbc06cd01),
	.w6(32'h3c13abf8),
	.w7(32'hbb4770c3),
	.w8(32'hbc3fd41d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82d450),
	.w1(32'hba099843),
	.w2(32'hbc7bbb54),
	.w3(32'hbbfb6566),
	.w4(32'hbc19b46d),
	.w5(32'hbc856113),
	.w6(32'h3c1e653e),
	.w7(32'h3ae6f7b1),
	.w8(32'hbb9b4e31),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc499f32),
	.w1(32'h3bde0ede),
	.w2(32'h3c3d2e8b),
	.w3(32'hbba01066),
	.w4(32'h3b3b37df),
	.w5(32'h3c01027d),
	.w6(32'h3c20d71c),
	.w7(32'h3c8c5fd3),
	.w8(32'h3c142037),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcff6f6),
	.w1(32'h3cc822ef),
	.w2(32'h3d515620),
	.w3(32'h3b33a690),
	.w4(32'h3cb5f45d),
	.w5(32'h3d35a711),
	.w6(32'h3c15cf74),
	.w7(32'h3ce1a7bf),
	.w8(32'h3cde26d4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d360629),
	.w1(32'hbb953ac7),
	.w2(32'hbba5e209),
	.w3(32'h3d160c30),
	.w4(32'hbbedff39),
	.w5(32'hbbddef7f),
	.w6(32'hbbad284e),
	.w7(32'hbbcc0c82),
	.w8(32'hbc0263d4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf62e9a),
	.w1(32'h3c5e7c27),
	.w2(32'h3c83dc24),
	.w3(32'hbc0280c7),
	.w4(32'h3c2a82e1),
	.w5(32'h3c3d294c),
	.w6(32'h3c33e022),
	.w7(32'h3c509a21),
	.w8(32'h3c57ce58),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c800e5c),
	.w1(32'h3b7ad2a4),
	.w2(32'h3b22bb43),
	.w3(32'h3c2c02e9),
	.w4(32'h3b3c24cd),
	.w5(32'h3acebfc7),
	.w6(32'h3adadc25),
	.w7(32'h3b64bd46),
	.w8(32'h3add7093),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b298694),
	.w1(32'h3be10533),
	.w2(32'hbbcad06f),
	.w3(32'hba30a208),
	.w4(32'h3b8e693e),
	.w5(32'h3acdbf87),
	.w6(32'h3bddb74c),
	.w7(32'h3b17f9bf),
	.w8(32'h3b5cda27),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca587),
	.w1(32'hbcfbddcc),
	.w2(32'hbd4e5606),
	.w3(32'hb9480a88),
	.w4(32'hbca516a5),
	.w5(32'hbce7be6d),
	.w6(32'hbbffec9e),
	.w7(32'hbca198e6),
	.w8(32'hbcac5ca7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd24b859),
	.w1(32'hbc242dd9),
	.w2(32'hbc54d3f0),
	.w3(32'hbcc93aee),
	.w4(32'h3b20cf10),
	.w5(32'hbc0d104f),
	.w6(32'hba9f8e52),
	.w7(32'hbbcc18a6),
	.w8(32'hbbe02a22),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6497dc),
	.w1(32'hbc8c9e0f),
	.w2(32'hbcb0a574),
	.w3(32'hbc488ead),
	.w4(32'hbc8d6d8d),
	.w5(32'hbcd3cc7f),
	.w6(32'hbaa43929),
	.w7(32'hbc1cd3cc),
	.w8(32'hbc662ad6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1ead9),
	.w1(32'h3b6bcae2),
	.w2(32'h3b47b99c),
	.w3(32'hbc55ba74),
	.w4(32'h3ad65020),
	.w5(32'h3b8caf18),
	.w6(32'hbb0a3089),
	.w7(32'hba833f06),
	.w8(32'h3b000b27),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ddb0b),
	.w1(32'hbd1c8fb6),
	.w2(32'hbd2d24af),
	.w3(32'h3b905a4e),
	.w4(32'hbc5d7b58),
	.w5(32'hbcc120b6),
	.w6(32'hbc09e656),
	.w7(32'hbc885404),
	.w8(32'hbc0b3094),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf90b9b),
	.w1(32'hbcb79668),
	.w2(32'hbd11e35e),
	.w3(32'hbca5b9a5),
	.w4(32'hbc95cc3f),
	.w5(32'hbd05f9e7),
	.w6(32'hbb4cfb15),
	.w7(32'hbc6ab3b4),
	.w8(32'hbbad240e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd08c55),
	.w1(32'h3b5ea917),
	.w2(32'h3b571277),
	.w3(32'hbc96e0d1),
	.w4(32'h3a9724e8),
	.w5(32'hba5cc2ea),
	.w6(32'h3af418a6),
	.w7(32'h3a54874f),
	.w8(32'h3b2dd9df),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884dc8),
	.w1(32'h3babae8a),
	.w2(32'hba4c2ceb),
	.w3(32'h3a3c1796),
	.w4(32'h3b7ce8ea),
	.w5(32'hbb12a61b),
	.w6(32'h3c0f2477),
	.w7(32'h3b97945b),
	.w8(32'h3bd336c4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cefb6),
	.w1(32'hbc3277d2),
	.w2(32'hbc93468d),
	.w3(32'h3bda053b),
	.w4(32'hbc6a0433),
	.w5(32'hbccd3098),
	.w6(32'hbc2583da),
	.w7(32'hbc854dc5),
	.w8(32'hbc02baba),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3d67f),
	.w1(32'hbb37e11f),
	.w2(32'hbb542c91),
	.w3(32'hba1bc249),
	.w4(32'hbb998e78),
	.w5(32'hbb9c9efc),
	.w6(32'h3a587846),
	.w7(32'h399de355),
	.w8(32'hbaf075eb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf36e3c),
	.w1(32'hbc22bf04),
	.w2(32'hbc196fd9),
	.w3(32'h3a017a49),
	.w4(32'hbc0d1b37),
	.w5(32'hbc33385b),
	.w6(32'hbb8585a0),
	.w7(32'hbb02c6d0),
	.w8(32'hbb8acf9a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbb663),
	.w1(32'hbb1867f3),
	.w2(32'hbbe2bc43),
	.w3(32'hbbbca5db),
	.w4(32'hbb10c315),
	.w5(32'h38a0f98a),
	.w6(32'hbbac6bc3),
	.w7(32'h3add9699),
	.w8(32'h3b52508a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb588b6a),
	.w1(32'hbc35ae84),
	.w2(32'hbc62492d),
	.w3(32'h3b1be489),
	.w4(32'hbc02ce64),
	.w5(32'hbc3b3ef0),
	.w6(32'hbbd432dc),
	.w7(32'hbad85c22),
	.w8(32'hb9afe339),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba909961),
	.w1(32'hbcd5b9f1),
	.w2(32'hbd0115f8),
	.w3(32'hbbba5ace),
	.w4(32'hbbdd695f),
	.w5(32'hbcb20377),
	.w6(32'hbc2364a2),
	.w7(32'hbc908359),
	.w8(32'hbc478d3d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1cb10),
	.w1(32'hb9fd015f),
	.w2(32'hbbc2a309),
	.w3(32'hbc6b9def),
	.w4(32'hbb6afa9d),
	.w5(32'hbbcf1ccb),
	.w6(32'h3a6d22c9),
	.w7(32'hbb7f2d08),
	.w8(32'h3ba86509),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac10776),
	.w1(32'hbbda4123),
	.w2(32'hbc03f92f),
	.w3(32'hbb0f481f),
	.w4(32'hbc6cee9c),
	.w5(32'hbc71d9e1),
	.w6(32'hbbfaa227),
	.w7(32'hbbff86d4),
	.w8(32'hbbb4cfd8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07c0d),
	.w1(32'h3c113053),
	.w2(32'h3ba99f1b),
	.w3(32'hbb8aecdd),
	.w4(32'h3c059fb1),
	.w5(32'hbb5623f3),
	.w6(32'h3beb5e4a),
	.w7(32'h3c4565c2),
	.w8(32'h3bf99c30),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b916b31),
	.w1(32'hbcd72f2a),
	.w2(32'hbcf9973c),
	.w3(32'hbb120122),
	.w4(32'hbc8ee729),
	.w5(32'hbce1269c),
	.w6(32'hbc90e58c),
	.w7(32'hbc86baa4),
	.w8(32'hbc61e029),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d0aca),
	.w1(32'h3c8483cb),
	.w2(32'h3c5b0fb2),
	.w3(32'hbcae2e94),
	.w4(32'h3c22d31c),
	.w5(32'h3bec7448),
	.w6(32'h3c350195),
	.w7(32'h3c134ae8),
	.w8(32'h3c01f05f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39058b),
	.w1(32'h3bee3c2f),
	.w2(32'h3c3f48ea),
	.w3(32'h3b8e233c),
	.w4(32'h3c64603c),
	.w5(32'h3c957767),
	.w6(32'h39b4d018),
	.w7(32'h3b7a11da),
	.w8(32'h3b8b46f8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c576e04),
	.w1(32'h3b456780),
	.w2(32'h3b83b44f),
	.w3(32'h3c4a3428),
	.w4(32'hb9ce200c),
	.w5(32'h3b7fb62a),
	.w6(32'h3c03d130),
	.w7(32'h3c2c9896),
	.w8(32'h3c4eacdb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c036be5),
	.w1(32'h3b671880),
	.w2(32'h39caa46e),
	.w3(32'h3bff7586),
	.w4(32'h3b8622a6),
	.w5(32'h3a977b80),
	.w6(32'h3ac93ec2),
	.w7(32'hb9211e5d),
	.w8(32'h3ab40628),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96229b),
	.w1(32'hbc94cf25),
	.w2(32'hbcea2282),
	.w3(32'h3aeb3532),
	.w4(32'hbc5b942d),
	.w5(32'hbcb91ebd),
	.w6(32'hbc3d4c7a),
	.w7(32'hbc7b29f6),
	.w8(32'hbbbacd69),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9680d3),
	.w1(32'hbca02e1b),
	.w2(32'hbd08c7a1),
	.w3(32'hbc499727),
	.w4(32'hbc97b3ff),
	.w5(32'hbcec91aa),
	.w6(32'hbc10b5ee),
	.w7(32'hbc67a189),
	.w8(32'hbc077047),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca60ee9),
	.w1(32'hba354d8e),
	.w2(32'h3bd5e365),
	.w3(32'hbc94e5ac),
	.w4(32'hbab98986),
	.w5(32'h3bbfae4c),
	.w6(32'h3a9e37c5),
	.w7(32'h3ba019a7),
	.w8(32'hbaab3349),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4aebe6),
	.w1(32'h3b9cc081),
	.w2(32'h3b9c105d),
	.w3(32'h3b315f65),
	.w4(32'h3bba0622),
	.w5(32'h3bf88a35),
	.w6(32'h3a4d1208),
	.w7(32'h3b2c51be),
	.w8(32'h3b5e6035),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddd2fc),
	.w1(32'hbbcb31d7),
	.w2(32'hbc425ea8),
	.w3(32'h3bf024b0),
	.w4(32'hbbcee2e8),
	.w5(32'hbc18157d),
	.w6(32'hbba5c77c),
	.w7(32'hbc07fa13),
	.w8(32'hbc0be98c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f9079),
	.w1(32'h3c44e51d),
	.w2(32'hbadb00ab),
	.w3(32'hbc1a8eeb),
	.w4(32'h3be9faed),
	.w5(32'hb9676946),
	.w6(32'h3c687271),
	.w7(32'hbb21871e),
	.w8(32'hbba1679b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc249406),
	.w1(32'h3c288f39),
	.w2(32'h3c50b65a),
	.w3(32'hbc3c28c6),
	.w4(32'h3c336a0b),
	.w5(32'h3c65359a),
	.w6(32'h3b850ba6),
	.w7(32'h3bce13f8),
	.w8(32'h3bfb8783),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81895c),
	.w1(32'hbc485dd6),
	.w2(32'hbc8e4c97),
	.w3(32'h3c821912),
	.w4(32'hbc590e70),
	.w5(32'hbc8e22d2),
	.w6(32'hbb8a667d),
	.w7(32'hbbeba46c),
	.w8(32'hbc2bee25),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ed747),
	.w1(32'hbc1b3e4e),
	.w2(32'hbce5a7b4),
	.w3(32'hbbfb1959),
	.w4(32'hbbd21f35),
	.w5(32'hbcdbb941),
	.w6(32'hbb9b6839),
	.w7(32'hbca48129),
	.w8(32'hbc93674d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91f16c),
	.w1(32'hbc83c6f7),
	.w2(32'hbd1d680b),
	.w3(32'hbc80f7d5),
	.w4(32'hbc675b13),
	.w5(32'hbcf3cb83),
	.w6(32'hbbdde90f),
	.w7(32'hbcae628e),
	.w8(32'hbc56c453),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9623f1),
	.w1(32'hbbca8b3a),
	.w2(32'h3bdc7e35),
	.w3(32'hbc9c260f),
	.w4(32'hbc34fd78),
	.w5(32'h3bceb53d),
	.w6(32'hbbd3ce0a),
	.w7(32'h3bcfa0dd),
	.w8(32'h3c2277a0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76d028),
	.w1(32'h3b82a139),
	.w2(32'h3b87b6dc),
	.w3(32'h3c24f7f4),
	.w4(32'h3c1400fe),
	.w5(32'h3c0c42be),
	.w6(32'h39fa5747),
	.w7(32'h3bd4c922),
	.w8(32'hbb8792c2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ee17),
	.w1(32'h3c153c9b),
	.w2(32'h3c18ebd2),
	.w3(32'h3912ae99),
	.w4(32'h3c2d87db),
	.w5(32'h3c56e442),
	.w6(32'h3b819b4f),
	.w7(32'h3beff855),
	.w8(32'h3c40d162),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0b12),
	.w1(32'hbc2d2704),
	.w2(32'hbc3bb39a),
	.w3(32'h3bf882c0),
	.w4(32'hbafa627f),
	.w5(32'hbc04b139),
	.w6(32'hb9a0a714),
	.w7(32'h3aed6739),
	.w8(32'h3b81fa1e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bd935),
	.w1(32'hbc90be8f),
	.w2(32'hbcac774f),
	.w3(32'hbc210e80),
	.w4(32'hbc5bddf2),
	.w5(32'hbb407f41),
	.w6(32'hbbd471da),
	.w7(32'hbc637574),
	.w8(32'hbc21c092),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2df7),
	.w1(32'h3bd4b407),
	.w2(32'h3c81be0c),
	.w3(32'h3bc8b817),
	.w4(32'h39b7c2cc),
	.w5(32'h3c2fd415),
	.w6(32'h3c1bc7eb),
	.w7(32'h3bc2b33e),
	.w8(32'h3c17a76c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c863cd3),
	.w1(32'hbba0c566),
	.w2(32'hbada6016),
	.w3(32'h3c7e542b),
	.w4(32'hbb554a1d),
	.w5(32'hbb2080ca),
	.w6(32'h3b3a07a8),
	.w7(32'h3b276566),
	.w8(32'h3ae82fc0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc204ae),
	.w1(32'hbb91b75a),
	.w2(32'hbc21bea8),
	.w3(32'hbb9a7ccd),
	.w4(32'hbc08ce28),
	.w5(32'hbbc76a7d),
	.w6(32'hbb0faa4b),
	.w7(32'hbbaf6d83),
	.w8(32'hbb59e1a6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5328e),
	.w1(32'h396b5c48),
	.w2(32'h3a716fba),
	.w3(32'hbba0cb7b),
	.w4(32'h3b486b6a),
	.w5(32'hbaeb95ff),
	.w6(32'h3a586f9c),
	.w7(32'hb865ccd0),
	.w8(32'h3bba1f39),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4f861),
	.w1(32'h3c099558),
	.w2(32'h3cb2c679),
	.w3(32'h3b879d1b),
	.w4(32'h3c211984),
	.w5(32'h3ca50a15),
	.w6(32'hbb7ea9a7),
	.w7(32'h3bd1c7f2),
	.w8(32'h3bb4fdc1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8502b2),
	.w1(32'hbaef3949),
	.w2(32'h3b7cb2af),
	.w3(32'h3c51b3d6),
	.w4(32'hbb4af30d),
	.w5(32'h3b3580ac),
	.w6(32'hbb94b45a),
	.w7(32'hba9f9249),
	.w8(32'hbb3a9d64),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dd7a5),
	.w1(32'hbc3257c9),
	.w2(32'hbc7a1a60),
	.w3(32'h3aa9b8f4),
	.w4(32'hbbe68b09),
	.w5(32'hbc46d7f5),
	.w6(32'hbb453450),
	.w7(32'hbbb9d001),
	.w8(32'hbbc9b0fd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2a1ed),
	.w1(32'hba0b8ab7),
	.w2(32'h3b42f746),
	.w3(32'hbc013bde),
	.w4(32'hbb15cbeb),
	.w5(32'h3ae45833),
	.w6(32'hbaa983de),
	.w7(32'h3ad1c057),
	.w8(32'h3abcd604),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c47e),
	.w1(32'h3b4dc5fd),
	.w2(32'h3c3bb5b3),
	.w3(32'hba3bdd5e),
	.w4(32'h3bf292d0),
	.w5(32'h3be054be),
	.w6(32'h3b679103),
	.w7(32'h3c54ddd8),
	.w8(32'h3c32a41a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c008c1a),
	.w1(32'h3ab392b7),
	.w2(32'hbae0ac6f),
	.w3(32'h3bed5059),
	.w4(32'hba853cb4),
	.w5(32'h3b783e86),
	.w6(32'hbb00d5b5),
	.w7(32'hbb14fc4d),
	.w8(32'h3a0efdf2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be79c82),
	.w1(32'h3bfd50ff),
	.w2(32'h3bc4fe43),
	.w3(32'hb9fde43e),
	.w4(32'h3c485931),
	.w5(32'h3bd763bc),
	.w6(32'h3b351657),
	.w7(32'h3b97db70),
	.w8(32'h3c42bf31),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c354dc7),
	.w1(32'h3a36c5da),
	.w2(32'h3bd8bccd),
	.w3(32'h3bba2bec),
	.w4(32'hba1abff1),
	.w5(32'h3b7004cf),
	.w6(32'hb9a402f2),
	.w7(32'h3b218af9),
	.w8(32'h3ade4d84),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf1e20),
	.w1(32'h3ceff648),
	.w2(32'h3d10cb77),
	.w3(32'h3b523654),
	.w4(32'h3c66b139),
	.w5(32'h3cbb9cb2),
	.w6(32'h3c7ebf8a),
	.w7(32'h3cdab03e),
	.w8(32'h3c786060),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3ee75),
	.w1(32'h3beda24e),
	.w2(32'h3b9b56c0),
	.w3(32'h3c403ba1),
	.w4(32'h3b8e2bb3),
	.w5(32'h3b2de82a),
	.w6(32'h3b710436),
	.w7(32'hbb02ce28),
	.w8(32'h3b1eb276),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08f796),
	.w1(32'hbcc8f7db),
	.w2(32'hbcb6b755),
	.w3(32'h3c1cd849),
	.w4(32'hbb163ae1),
	.w5(32'hbc723302),
	.w6(32'hbbf384ae),
	.w7(32'hbb7fbe0c),
	.w8(32'hba1ce23e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7018fc),
	.w1(32'hbb0c74af),
	.w2(32'hbbae3a45),
	.w3(32'hbc79f7ad),
	.w4(32'hbb46b049),
	.w5(32'hbb45e2f5),
	.w6(32'hbb96a5e6),
	.w7(32'h37df2b2e),
	.w8(32'hba3a1e79),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a084f),
	.w1(32'hbbd1ae50),
	.w2(32'hbb891d54),
	.w3(32'hbace899f),
	.w4(32'hbad40ef2),
	.w5(32'hbbb2c24c),
	.w6(32'hbbeea066),
	.w7(32'h3bc17ed5),
	.w8(32'hbb79c18d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad74553),
	.w1(32'hbc6d5163),
	.w2(32'hbc94203d),
	.w3(32'hbb8dc2ab),
	.w4(32'hbc9e5559),
	.w5(32'hbc8ca208),
	.w6(32'hbbc57bd6),
	.w7(32'hbbfbcb2d),
	.w8(32'hbc38bcc8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e09c8),
	.w1(32'h3bedebbc),
	.w2(32'h3c35c569),
	.w3(32'hbc35b83c),
	.w4(32'h3b711359),
	.w5(32'h3c360c3b),
	.w6(32'hb979c7d2),
	.w7(32'h3b62781d),
	.w8(32'h3a5d7526),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a66ad),
	.w1(32'h3b9e7bf5),
	.w2(32'h3c537c72),
	.w3(32'h3bb12814),
	.w4(32'h3c1139bb),
	.w5(32'h3c4d555d),
	.w6(32'h3bc02889),
	.w7(32'h3bab060d),
	.w8(32'h3bd23aa7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8d195),
	.w1(32'h3af9a8af),
	.w2(32'hbc02a7f3),
	.w3(32'h3c7065a5),
	.w4(32'h3c5fd106),
	.w5(32'h3c0695fe),
	.w6(32'h39e3eded),
	.w7(32'hb9d5f51c),
	.w8(32'hbb3eacd4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08eae8),
	.w1(32'h39d93412),
	.w2(32'hbc3cf1e5),
	.w3(32'hb9a76135),
	.w4(32'hbc5290be),
	.w5(32'hbc5c2d58),
	.w6(32'h3bfe1a5f),
	.w7(32'h3ba1bbb0),
	.w8(32'hbb1f14f7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3612c8),
	.w1(32'hba27a261),
	.w2(32'h3b0dc0fe),
	.w3(32'hbbb726c1),
	.w4(32'h3a0507ca),
	.w5(32'hb806ed34),
	.w6(32'h3a871e23),
	.w7(32'h39d80aeb),
	.w8(32'h3a4701df),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85763eb),
	.w1(32'hbc037443),
	.w2(32'hbbd40b63),
	.w3(32'hb9e2e2f5),
	.w4(32'hbae6fd30),
	.w5(32'hba19e5a2),
	.w6(32'hbb8c6ab7),
	.w7(32'hbb178483),
	.w8(32'h3b4ac49a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule