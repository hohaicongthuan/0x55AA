module layer_10_featuremap_502(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b788ff8),
	.w1(32'h3a0e974a),
	.w2(32'hbae9ecb4),
	.w3(32'h3a89a63a),
	.w4(32'hba7587dc),
	.w5(32'hbbae31cb),
	.w6(32'hbbf7b513),
	.w7(32'hbb42ce7f),
	.w8(32'hbb635dfb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37770a),
	.w1(32'hbb7f6860),
	.w2(32'hbb3a264d),
	.w3(32'hbae95fda),
	.w4(32'hba9f5c5d),
	.w5(32'h3a42cbec),
	.w6(32'hbb959181),
	.w7(32'hb9c1cf9c),
	.w8(32'hbb8d3d1d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d1a4d),
	.w1(32'hba41f0dd),
	.w2(32'h3ad89ad3),
	.w3(32'h3ab647e9),
	.w4(32'h3b08fef6),
	.w5(32'h3c3e52f7),
	.w6(32'hb973d809),
	.w7(32'hbb4f382e),
	.w8(32'h3bb5156a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ab863),
	.w1(32'h3af6b811),
	.w2(32'h3b38bc0b),
	.w3(32'hbbf09dfd),
	.w4(32'hbb604d1e),
	.w5(32'hbb127aa0),
	.w6(32'h3bc5d27b),
	.w7(32'hba47e23a),
	.w8(32'hbb5a1ccc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02c49),
	.w1(32'h36e92130),
	.w2(32'h39e8cf08),
	.w3(32'hb9a22c9e),
	.w4(32'hb992cbbb),
	.w5(32'h3a8b9651),
	.w6(32'h3b58c914),
	.w7(32'h3b4790c6),
	.w8(32'h39789ae6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf1e09),
	.w1(32'h39f10cf2),
	.w2(32'hbbab3bf3),
	.w3(32'hbb683922),
	.w4(32'hbb43486f),
	.w5(32'hbbbec2d7),
	.w6(32'hbb02b116),
	.w7(32'h3b4b2581),
	.w8(32'hbbc76276),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb44019),
	.w1(32'hbabe359e),
	.w2(32'hbb33ccd5),
	.w3(32'hbb990a8c),
	.w4(32'hb7d5ab10),
	.w5(32'hbb113d26),
	.w6(32'hbbea90c4),
	.w7(32'hbc01b5e6),
	.w8(32'hbc02ff40),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74b2e),
	.w1(32'hbb45a290),
	.w2(32'hbaa462d8),
	.w3(32'hbac7f0a0),
	.w4(32'hbb46bb97),
	.w5(32'hbc0ec0a3),
	.w6(32'hbbf680a4),
	.w7(32'h3ad89a8f),
	.w8(32'hbaf2722a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37008d96),
	.w1(32'h3a94207d),
	.w2(32'hbb06e9d3),
	.w3(32'hbb168186),
	.w4(32'hbb6a53de),
	.w5(32'hbb8ed6df),
	.w6(32'hbb369a84),
	.w7(32'hbb3ae014),
	.w8(32'hbbbeec13),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc098ea8),
	.w1(32'hba140548),
	.w2(32'h3c0f7acc),
	.w3(32'hbbb8a03e),
	.w4(32'hbc0b7963),
	.w5(32'hb9cd04a3),
	.w6(32'hbb6396d4),
	.w7(32'hbb863fd8),
	.w8(32'h3b468c7e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2219cb),
	.w1(32'hbac785d2),
	.w2(32'hb8a45158),
	.w3(32'h378a0bed),
	.w4(32'h3ab40c77),
	.w5(32'h3c0b5180),
	.w6(32'h3bfc24e1),
	.w7(32'hb9d99ce5),
	.w8(32'h3b174dda),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b83f9b),
	.w1(32'hbb007f8a),
	.w2(32'hbbdcdad0),
	.w3(32'h3c1d5ecf),
	.w4(32'h3bbbb080),
	.w5(32'hbbfea2a5),
	.w6(32'h3bc7ff0f),
	.w7(32'h3b9fde14),
	.w8(32'hbbffc245),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a69d73),
	.w1(32'h3b2231a7),
	.w2(32'h3b7dad73),
	.w3(32'h3a8efd8d),
	.w4(32'hb92d794a),
	.w5(32'h3a99754e),
	.w6(32'hbb1230e3),
	.w7(32'hbbca9298),
	.w8(32'hbacb59db),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd6827),
	.w1(32'hbbd0257d),
	.w2(32'h39b85c65),
	.w3(32'h3ba4a9c3),
	.w4(32'h3b3b0beb),
	.w5(32'h3c4f1918),
	.w6(32'h398a3b90),
	.w7(32'hbbddfe9b),
	.w8(32'h3bf096d4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb769352),
	.w1(32'h3b23fec6),
	.w2(32'h3b85ed05),
	.w3(32'hbaa4e8f5),
	.w4(32'h3aa921ca),
	.w5(32'h3c512865),
	.w6(32'h3b3ebf03),
	.w7(32'hbbb0242d),
	.w8(32'hb9cb4d2e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2e8f1),
	.w1(32'h3b20c6ee),
	.w2(32'hba78dfbc),
	.w3(32'h3b3d1c97),
	.w4(32'hb9af9f43),
	.w5(32'h3a8b11b9),
	.w6(32'h3a890d82),
	.w7(32'hbbc9be62),
	.w8(32'hbb02ccdb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a719930),
	.w1(32'hbb2d0d51),
	.w2(32'hbb77cb7b),
	.w3(32'h3b58f7a7),
	.w4(32'h3ae55305),
	.w5(32'h3ac4d0e1),
	.w6(32'h3a4a5528),
	.w7(32'hba65860c),
	.w8(32'hb9d690fe),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ddcca),
	.w1(32'hbb8b99b2),
	.w2(32'hbb86bf65),
	.w3(32'hbb7f7c29),
	.w4(32'hbb80a787),
	.w5(32'hbb27787b),
	.w6(32'hbc3fff1e),
	.w7(32'hbb9a88d3),
	.w8(32'h3b3130f7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc386306),
	.w1(32'h3a04c3b9),
	.w2(32'h3bd42d07),
	.w3(32'hbb22442c),
	.w4(32'hbb449c5c),
	.w5(32'h3ae67a8c),
	.w6(32'hbb9e4730),
	.w7(32'hbbc535d2),
	.w8(32'hbc17f629),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ae70),
	.w1(32'h3a6ed976),
	.w2(32'h3bfe0410),
	.w3(32'h3bb1d0c9),
	.w4(32'hbb5292c5),
	.w5(32'h3c2671c4),
	.w6(32'hba3de175),
	.w7(32'hbafcc480),
	.w8(32'hbb5bb5d4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae89fec),
	.w1(32'h3b77d6ae),
	.w2(32'hbb98362b),
	.w3(32'h3c1dc45f),
	.w4(32'h3bb5e5b1),
	.w5(32'hbb86fd21),
	.w6(32'h3c132954),
	.w7(32'h3c3db3a5),
	.w8(32'h3a859439),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4109fb),
	.w1(32'h3a5e2e8c),
	.w2(32'h3bbb1fef),
	.w3(32'hbb927cdf),
	.w4(32'hbbac1dcc),
	.w5(32'hbc02dd25),
	.w6(32'hb9ae4424),
	.w7(32'hbb2221e5),
	.w8(32'hbb0d8630),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1329ff),
	.w1(32'h3b25b050),
	.w2(32'h3bb64975),
	.w3(32'hbc55fab5),
	.w4(32'hbc0c8c87),
	.w5(32'hbbc378a7),
	.w6(32'hbc472d8b),
	.w7(32'hbc896ca1),
	.w8(32'hbbd1a3b8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde9de3),
	.w1(32'h3bbc6808),
	.w2(32'h3c04a420),
	.w3(32'hbb5e02d7),
	.w4(32'hbb812bd8),
	.w5(32'h3a9594c4),
	.w6(32'hbb8aa41a),
	.w7(32'hbb9cfead),
	.w8(32'hbb804038),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c052dc6),
	.w1(32'hbac50786),
	.w2(32'hb9066ea3),
	.w3(32'h3ae98fd0),
	.w4(32'h39cfcbe9),
	.w5(32'hb70fec4a),
	.w6(32'hbb13991d),
	.w7(32'hbb325339),
	.w8(32'h3abdbacc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82b9c2),
	.w1(32'h3bd648d2),
	.w2(32'h3bb1e266),
	.w3(32'hbb6ab224),
	.w4(32'hbbb10049),
	.w5(32'hbbd552c0),
	.w6(32'h37579b61),
	.w7(32'h3b9ff76c),
	.w8(32'hbb0c9485),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba77a49),
	.w1(32'h3c1b9b87),
	.w2(32'h39bed1ae),
	.w3(32'h3b3fd0bf),
	.w4(32'h3c58f9a8),
	.w5(32'h39804d99),
	.w6(32'h3afd034d),
	.w7(32'hbb88cd05),
	.w8(32'hbbe12b8f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be5f6),
	.w1(32'hba3ef2bc),
	.w2(32'hbb836f46),
	.w3(32'h3cef9243),
	.w4(32'hbb86f2f4),
	.w5(32'hbc05e9b1),
	.w6(32'h3be84b3f),
	.w7(32'hbba6ea30),
	.w8(32'hba9be134),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1544eb),
	.w1(32'hbb6b030b),
	.w2(32'h39374b1a),
	.w3(32'hbb65a037),
	.w4(32'hba9a776a),
	.w5(32'hbb3d41f7),
	.w6(32'h3ad92fe7),
	.w7(32'hbb102147),
	.w8(32'hbb874040),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba270270),
	.w1(32'h38e6710f),
	.w2(32'hbb80b9e3),
	.w3(32'h3ba7fefb),
	.w4(32'h3bf0acfe),
	.w5(32'h3a9649f7),
	.w6(32'h3a5055fb),
	.w7(32'h3c1054df),
	.w8(32'h3b9b54df),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68dfd),
	.w1(32'h3a93cf14),
	.w2(32'hbba9b021),
	.w3(32'hbb9058f9),
	.w4(32'h3baa5933),
	.w5(32'hb95ab2af),
	.w6(32'hbbb14367),
	.w7(32'hb99c2781),
	.w8(32'hbaac9c99),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba1ebd),
	.w1(32'h3a03dc5f),
	.w2(32'h3b344a43),
	.w3(32'hb6948f96),
	.w4(32'h3b5fe3ee),
	.w5(32'h3c1ac154),
	.w6(32'h39b9925b),
	.w7(32'hba781201),
	.w8(32'h3b262ffc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59c63f),
	.w1(32'hbb640f2a),
	.w2(32'h3ba419f8),
	.w3(32'h3b76f48a),
	.w4(32'hbb977cab),
	.w5(32'h3a4d743b),
	.w6(32'h3b446bd6),
	.w7(32'h3b1fd099),
	.w8(32'hbb5c2912),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c494235),
	.w1(32'h3b36fa68),
	.w2(32'h3b89643c),
	.w3(32'h3a6456b8),
	.w4(32'hbbb10ebe),
	.w5(32'hbb1f1556),
	.w6(32'h3c06680f),
	.w7(32'h3a6f9a6a),
	.w8(32'h3b8075be),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb021d),
	.w1(32'hb810423b),
	.w2(32'h3a1ef59a),
	.w3(32'hba59e993),
	.w4(32'h3b0a4858),
	.w5(32'h3913ae36),
	.w6(32'h3bd359cc),
	.w7(32'h3b2b509d),
	.w8(32'h3b823923),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0fe5),
	.w1(32'hbb1a167b),
	.w2(32'h391696fd),
	.w3(32'hb940c934),
	.w4(32'h39de2ae0),
	.w5(32'hbb938098),
	.w6(32'hbae13e59),
	.w7(32'h3b542476),
	.w8(32'h3a71f658),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2bedf),
	.w1(32'h3b94ed0d),
	.w2(32'h3b249540),
	.w3(32'hbc1379ae),
	.w4(32'h3c3c4d68),
	.w5(32'h3c71c3ec),
	.w6(32'hbc1a4cd3),
	.w7(32'hba714fb7),
	.w8(32'hbb478841),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba979e5),
	.w1(32'hbb1b7fb4),
	.w2(32'hbbab5b52),
	.w3(32'h3b2b27b8),
	.w4(32'hba97bc55),
	.w5(32'h3ba5707b),
	.w6(32'h3b67ff2f),
	.w7(32'hbc0800e2),
	.w8(32'hbc0ce28a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb408e6f),
	.w1(32'hbb412daa),
	.w2(32'hb7e05a04),
	.w3(32'h3a72247e),
	.w4(32'hbbb0cf38),
	.w5(32'hbc04f44e),
	.w6(32'hbabed894),
	.w7(32'hbb627736),
	.w8(32'hbc0ed182),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a66eb),
	.w1(32'h3bdf5089),
	.w2(32'h3baeb899),
	.w3(32'hbb17d5da),
	.w4(32'hba4b3600),
	.w5(32'h3b17aeb2),
	.w6(32'hba9e116a),
	.w7(32'hbb39b8c8),
	.w8(32'h3b1bfd34),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1661de),
	.w1(32'hbb1ad7f1),
	.w2(32'hb9a87751),
	.w3(32'h3b091947),
	.w4(32'hbc1114f5),
	.w5(32'hbbd785d2),
	.w6(32'h3b29b128),
	.w7(32'hbc0d07b6),
	.w8(32'hbae319b2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf549d2),
	.w1(32'h3b88a4db),
	.w2(32'hba8fecae),
	.w3(32'h39c26c88),
	.w4(32'h3b27f998),
	.w5(32'hbb6ba04b),
	.w6(32'h3a0412a2),
	.w7(32'h3bec40a4),
	.w8(32'h3aee7c8a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdfe78),
	.w1(32'h3aa74d67),
	.w2(32'h3beb3af5),
	.w3(32'hbb8d8810),
	.w4(32'hbbdb6ba8),
	.w5(32'h3b3e2cc5),
	.w6(32'hbacf7232),
	.w7(32'hbbb990af),
	.w8(32'hbb6f67e4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc2626),
	.w1(32'h3badc610),
	.w2(32'h3aae3c4d),
	.w3(32'h3c05108a),
	.w4(32'h3ae3a32a),
	.w5(32'hbb417220),
	.w6(32'h3a9c6a23),
	.w7(32'hba391293),
	.w8(32'hbb374bd8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a8858),
	.w1(32'h3a4bb984),
	.w2(32'h3cae76f4),
	.w3(32'h3c354de6),
	.w4(32'hbb9b09ca),
	.w5(32'h3c3070f0),
	.w6(32'h3be6fd1c),
	.w7(32'hbbc4aa43),
	.w8(32'h3c12e9d1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39b38e),
	.w1(32'h39aefc80),
	.w2(32'h3b25032d),
	.w3(32'h3bdc9fd0),
	.w4(32'hb8cb909e),
	.w5(32'h3ba7a83d),
	.w6(32'h3c14428d),
	.w7(32'hbb797683),
	.w8(32'h3b2662c7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70ab00),
	.w1(32'h3b0a71f4),
	.w2(32'h3bd7bc74),
	.w3(32'hba12e8e0),
	.w4(32'hb9be0b8f),
	.w5(32'hbb05ae05),
	.w6(32'hbb47be03),
	.w7(32'hbb83fa32),
	.w8(32'hbaaa90e7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27f349),
	.w1(32'hbbb89ae7),
	.w2(32'h3b10b605),
	.w3(32'h3b02f428),
	.w4(32'hb9152f6f),
	.w5(32'hba929caf),
	.w6(32'hbbd1ef56),
	.w7(32'hb99a83ea),
	.w8(32'hbab61e3f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5f134),
	.w1(32'h3b9c5a74),
	.w2(32'hbb52d175),
	.w3(32'hbacacb82),
	.w4(32'h3bdcc3e7),
	.w5(32'hbb98af25),
	.w6(32'hbb19d9f1),
	.w7(32'h3c27c782),
	.w8(32'h3bd7789e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d82c),
	.w1(32'hba924fad),
	.w2(32'hbaf14943),
	.w3(32'hbb59619f),
	.w4(32'h3baae946),
	.w5(32'hbc3fd16d),
	.w6(32'h3bc101a5),
	.w7(32'h3c193e47),
	.w8(32'hbb63e13c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dd645),
	.w1(32'h39ff995c),
	.w2(32'h3b81a6d2),
	.w3(32'hbb2eb787),
	.w4(32'hbbc4bff8),
	.w5(32'hbabe641b),
	.w6(32'hbab42eec),
	.w7(32'hbc09240c),
	.w8(32'hbb8eeea5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb74ab6),
	.w1(32'hbb994555),
	.w2(32'h39e86b97),
	.w3(32'h3bcaf560),
	.w4(32'hbba14b03),
	.w5(32'hbb95e5d8),
	.w6(32'hb8087591),
	.w7(32'h3b8ab630),
	.w8(32'hbc071aa1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a3f15),
	.w1(32'h3b25e107),
	.w2(32'hbb2b4ee0),
	.w3(32'hba6534f2),
	.w4(32'h3bd736e9),
	.w5(32'hbb3a3f7c),
	.w6(32'hbb742a9c),
	.w7(32'h3c773463),
	.w8(32'h3c1515f4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c413),
	.w1(32'hba9c0cbd),
	.w2(32'h3ae7e5b7),
	.w3(32'hbbe61622),
	.w4(32'hbade2811),
	.w5(32'hb7594536),
	.w6(32'hbb1e3187),
	.w7(32'h3bb59b4d),
	.w8(32'h3b9baabe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857e94),
	.w1(32'h3bcc30cc),
	.w2(32'h3bf9196b),
	.w3(32'hbb94f9eb),
	.w4(32'h3b3ff814),
	.w5(32'h3cbdfe1f),
	.w6(32'hbb35fe59),
	.w7(32'hbc20b88e),
	.w8(32'h3c01c8ef),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1b12),
	.w1(32'h3b6ab2fd),
	.w2(32'h3b9697a6),
	.w3(32'h3c3e9d6f),
	.w4(32'hbb3a8eab),
	.w5(32'h3c5863f8),
	.w6(32'h3bb01c0a),
	.w7(32'hbbfa2898),
	.w8(32'hba087a04),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b02b9),
	.w1(32'h3a04b53b),
	.w2(32'h38cb77aa),
	.w3(32'h3aaf3308),
	.w4(32'h3a8bee23),
	.w5(32'hba827d92),
	.w6(32'h39b2ac4d),
	.w7(32'hbbb7e0b6),
	.w8(32'hbba958ca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba60dd0),
	.w1(32'hbb80f46d),
	.w2(32'hbb3cba22),
	.w3(32'h3bd2cbe8),
	.w4(32'hbba50030),
	.w5(32'h3a8ab4bb),
	.w6(32'hbb07d828),
	.w7(32'h3a824222),
	.w8(32'hbb366697),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6569d),
	.w1(32'hba912577),
	.w2(32'hb9377c01),
	.w3(32'h39570683),
	.w4(32'hbb1cb66e),
	.w5(32'hbb870c29),
	.w6(32'h3b5288a1),
	.w7(32'hbbb02b8f),
	.w8(32'hbbeae8f2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fad32),
	.w1(32'h3a2b10fd),
	.w2(32'h3c26a110),
	.w3(32'hbb1871c9),
	.w4(32'h3b617552),
	.w5(32'h3c4a7f1c),
	.w6(32'hbc03e2d7),
	.w7(32'hbb2d3cd8),
	.w8(32'h3affabeb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed4db0),
	.w1(32'h375771ff),
	.w2(32'h3b808fbe),
	.w3(32'h3c3d52a2),
	.w4(32'hbc16723a),
	.w5(32'h3b6916f4),
	.w6(32'h3b9a8a0f),
	.w7(32'hbc13ca90),
	.w8(32'hbbea9889),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f6d4),
	.w1(32'h3a9989bc),
	.w2(32'h3bd123b3),
	.w3(32'h3cab7c61),
	.w4(32'hbc05b3c8),
	.w5(32'h3c021cde),
	.w6(32'h3a6e4c34),
	.w7(32'hbc2b636b),
	.w8(32'h3b2fdb5a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dc3a1),
	.w1(32'hba8ca58b),
	.w2(32'h3bbfaa19),
	.w3(32'h3b36229b),
	.w4(32'hbb8dd966),
	.w5(32'h3b42f9cf),
	.w6(32'hb89eef1e),
	.w7(32'hbbc67a99),
	.w8(32'hbb0cd6cd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5670c5),
	.w1(32'h3b1f1f9f),
	.w2(32'h3ba0fc4c),
	.w3(32'hba3509a5),
	.w4(32'hba96a785),
	.w5(32'h3b1bd7d8),
	.w6(32'hbbafdd20),
	.w7(32'hbb998aff),
	.w8(32'hbb3df024),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c163bb2),
	.w1(32'h3b27fcfe),
	.w2(32'h39db3406),
	.w3(32'h3c062da8),
	.w4(32'h39d5222e),
	.w5(32'hbb7afb98),
	.w6(32'h3ac086e6),
	.w7(32'h3a879014),
	.w8(32'h39791e8f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c924e),
	.w1(32'h3b29bd32),
	.w2(32'hbb1bd21a),
	.w3(32'h3b4daf05),
	.w4(32'h3b1e769e),
	.w5(32'hbbabcebe),
	.w6(32'h3b3f3f06),
	.w7(32'h3bfa9b0a),
	.w8(32'h39f1754a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd39a2),
	.w1(32'h3ba8d9d7),
	.w2(32'h3b8211ed),
	.w3(32'hb9e81d9f),
	.w4(32'h3c027f40),
	.w5(32'h3bf1a6f7),
	.w6(32'hbb7f6214),
	.w7(32'h3b173e5f),
	.w8(32'h3bdb345f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba22550),
	.w1(32'h3aaa97a6),
	.w2(32'hbb6a105a),
	.w3(32'h3b15690b),
	.w4(32'hbbdc649a),
	.w5(32'h3acd9897),
	.w6(32'h3afbac08),
	.w7(32'hbb9d47cd),
	.w8(32'hbb45ff5f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cb049),
	.w1(32'hbc1d00e9),
	.w2(32'h3b5de0cd),
	.w3(32'hbc5c3d74),
	.w4(32'hbbde8dd4),
	.w5(32'hbb0a7cab),
	.w6(32'hbc29482e),
	.w7(32'hbb814bbf),
	.w8(32'hbb8854bc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e32ae),
	.w1(32'h3abfd07d),
	.w2(32'h3c898801),
	.w3(32'hbbb48dce),
	.w4(32'h3c08df1e),
	.w5(32'hbb234027),
	.w6(32'hbbf2991d),
	.w7(32'hba080492),
	.w8(32'h3a7ae46a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf44f73),
	.w1(32'h3c036c7e),
	.w2(32'h3b2b7837),
	.w3(32'hbb31667d),
	.w4(32'h3c217e77),
	.w5(32'hbad58b14),
	.w6(32'h3b745f17),
	.w7(32'h3b3975ba),
	.w8(32'h3b8241db),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2239fa),
	.w1(32'h3c387a72),
	.w2(32'h3a6760ce),
	.w3(32'h3bcaae89),
	.w4(32'h3bd2fa1b),
	.w5(32'hbb638c56),
	.w6(32'hbab9baa8),
	.w7(32'h3b7c0a15),
	.w8(32'h3b173b1a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98a7e2),
	.w1(32'h3c0f9b7c),
	.w2(32'hbb28219c),
	.w3(32'h3a67cf55),
	.w4(32'h3c1e4592),
	.w5(32'hbc8049ac),
	.w6(32'h3b68d04d),
	.w7(32'h3c3060e9),
	.w8(32'hbb4d35f2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ec0d4),
	.w1(32'h3a1637f5),
	.w2(32'hbafb53a2),
	.w3(32'hbab3385a),
	.w4(32'hbb294b80),
	.w5(32'hbb49f64e),
	.w6(32'hbb2e5583),
	.w7(32'hbbb54ea0),
	.w8(32'hb9b488b1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed196a),
	.w1(32'h3bad5dc2),
	.w2(32'h3b2d49b0),
	.w3(32'h3af0ba16),
	.w4(32'h3942f2b4),
	.w5(32'h3b9cba8d),
	.w6(32'h3a22f975),
	.w7(32'h3b004998),
	.w8(32'hbaaff9d9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4a534),
	.w1(32'hbbd98a93),
	.w2(32'hbbaa0a8a),
	.w3(32'h3b8fc8f7),
	.w4(32'h398f625e),
	.w5(32'hbbc1942c),
	.w6(32'hba19af8a),
	.w7(32'h3ba30181),
	.w8(32'h3c02ea6e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6720f),
	.w1(32'h3a9106f8),
	.w2(32'h3b2416c9),
	.w3(32'h3b12c57c),
	.w4(32'h3b1fd209),
	.w5(32'h3c609c5f),
	.w6(32'hbab8f144),
	.w7(32'h3b19df96),
	.w8(32'hb97074d1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d6f10),
	.w1(32'h3b6dd263),
	.w2(32'h3bdc698c),
	.w3(32'h388834d1),
	.w4(32'h3b3263e0),
	.w5(32'hbc22f22c),
	.w6(32'h3b729270),
	.w7(32'h3bceaaea),
	.w8(32'h3bc4ee76),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb456e73),
	.w1(32'hbb9df7d0),
	.w2(32'h3b29c0be),
	.w3(32'h3b91c912),
	.w4(32'hbc018138),
	.w5(32'h3bd084ed),
	.w6(32'h3bdb431d),
	.w7(32'hbbc6358d),
	.w8(32'h3aa6acef),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7188ac),
	.w1(32'hba5ae56b),
	.w2(32'h3bdfb0cc),
	.w3(32'hbb0f6f15),
	.w4(32'h3bc25102),
	.w5(32'h3bf85f9c),
	.w6(32'hbba6c239),
	.w7(32'h3bf80e51),
	.w8(32'h3bda022c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a663fe8),
	.w1(32'hbc26b7fb),
	.w2(32'h3a7b2e78),
	.w3(32'h3b4a5abb),
	.w4(32'h3b8e52a4),
	.w5(32'h3c8d2496),
	.w6(32'h3b7de028),
	.w7(32'hbbdec745),
	.w8(32'hbb81f267),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1115c8),
	.w1(32'h3b551195),
	.w2(32'hbbd68621),
	.w3(32'hba979f06),
	.w4(32'h3bf8dd78),
	.w5(32'hbc1f9874),
	.w6(32'hbadc79d2),
	.w7(32'h3b68cf46),
	.w8(32'hbbb42de4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3ec9),
	.w1(32'h3aed6c7c),
	.w2(32'hba75be87),
	.w3(32'hbb9200b4),
	.w4(32'hbb873f56),
	.w5(32'hbbff6855),
	.w6(32'hba582628),
	.w7(32'h3ad97a4b),
	.w8(32'hbb85688f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc580b7),
	.w1(32'h3b417607),
	.w2(32'h3c0b8270),
	.w3(32'h3b785288),
	.w4(32'h3bee74d4),
	.w5(32'hbc3d10a7),
	.w6(32'hb9933b6f),
	.w7(32'h3c1822bb),
	.w8(32'h3bba694c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81849b),
	.w1(32'h3bfcb20b),
	.w2(32'hbb9b262c),
	.w3(32'hbab50791),
	.w4(32'h3c1479f3),
	.w5(32'hbc865cc2),
	.w6(32'hbc0db5df),
	.w7(32'h3c4046af),
	.w8(32'h39d45a6b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20e53),
	.w1(32'h3b0cd77c),
	.w2(32'h3b7b3544),
	.w3(32'hbc15a475),
	.w4(32'hbbf7653d),
	.w5(32'h3c94a98f),
	.w6(32'hbb7dd47e),
	.w7(32'h3c11fc22),
	.w8(32'h3c518ce1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb8add),
	.w1(32'h3b85fc37),
	.w2(32'hbb3cd98f),
	.w3(32'h3b2fe947),
	.w4(32'h3b6b93db),
	.w5(32'hbb57ab58),
	.w6(32'h3b24bd43),
	.w7(32'hb8ee57c0),
	.w8(32'h3b5be1b1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af65194),
	.w1(32'hbaf1bd82),
	.w2(32'hbaee8444),
	.w3(32'h3b0de73a),
	.w4(32'hbac882e8),
	.w5(32'hbb9559f4),
	.w6(32'h3ae2342c),
	.w7(32'hba5146ab),
	.w8(32'hba6fa6f8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f5cac),
	.w1(32'hba6e7a57),
	.w2(32'h3bf027b1),
	.w3(32'hbb3382ce),
	.w4(32'h3b488ef7),
	.w5(32'h39b95343),
	.w6(32'h3a3663a5),
	.w7(32'h3c4f2088),
	.w8(32'h3b2b910b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e446f),
	.w1(32'hba12e73f),
	.w2(32'hb988be38),
	.w3(32'h3b514316),
	.w4(32'hbbc409a4),
	.w5(32'hba565b21),
	.w6(32'h3af37118),
	.w7(32'hbbbab1ef),
	.w8(32'hbb9e711c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918903d),
	.w1(32'h3be112b8),
	.w2(32'h3b12e585),
	.w3(32'hbb52a2ee),
	.w4(32'h3c40afcd),
	.w5(32'hbc9f4aca),
	.w6(32'hbaccbc0a),
	.w7(32'h3bcfb113),
	.w8(32'hbba9fbff),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1edd05),
	.w1(32'h3a829035),
	.w2(32'hba5341e4),
	.w3(32'h3bdb1fed),
	.w4(32'hbb3a5acb),
	.w5(32'hbb4244bd),
	.w6(32'h3b84e752),
	.w7(32'hbb159c5e),
	.w8(32'h3ae5fbe1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa7c6e),
	.w1(32'hba3e5b64),
	.w2(32'hbb7f9189),
	.w3(32'h3aaed68c),
	.w4(32'hbb84ac76),
	.w5(32'hbc1938f9),
	.w6(32'h3b8f9acb),
	.w7(32'hbbc2f735),
	.w8(32'hbc3bb3ad),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ceb15),
	.w1(32'h3b6ba3a4),
	.w2(32'h3b50721d),
	.w3(32'hbc2449cc),
	.w4(32'hbb091661),
	.w5(32'hbb2e9457),
	.w6(32'hbc7b2091),
	.w7(32'hbb83a831),
	.w8(32'hba8949e1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea4d7c),
	.w1(32'h3c095881),
	.w2(32'h3c08c751),
	.w3(32'hbb3da3ea),
	.w4(32'h3b71a9b4),
	.w5(32'hba8ba331),
	.w6(32'h3a534f65),
	.w7(32'h3bee87bc),
	.w8(32'h3c0c1987),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc638ee),
	.w1(32'h3bc7c12d),
	.w2(32'h3c3f14be),
	.w3(32'h3b82c465),
	.w4(32'h3b819123),
	.w5(32'hbbe4fc85),
	.w6(32'h3c6eb038),
	.w7(32'h3a6a004f),
	.w8(32'h3ac3a3e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be190d9),
	.w1(32'h3be46fc5),
	.w2(32'hb9a6de09),
	.w3(32'h3a7d340e),
	.w4(32'hbab3e9e7),
	.w5(32'hbc35f811),
	.w6(32'h3bdf5023),
	.w7(32'hb9e5a382),
	.w8(32'hbbc6660a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6650ce),
	.w1(32'h3b9b83ef),
	.w2(32'hbaf9667f),
	.w3(32'hbb9b5832),
	.w4(32'h3b6782fd),
	.w5(32'hbb6edd56),
	.w6(32'hbbfe6f27),
	.w7(32'h3b9925e1),
	.w8(32'hbc1ccac7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf9eb7),
	.w1(32'h3b972759),
	.w2(32'hbbaa3570),
	.w3(32'hbb0c8f72),
	.w4(32'h3ba9a81e),
	.w5(32'hbcb2bcb3),
	.w6(32'hbbf26de0),
	.w7(32'h3b8187a5),
	.w8(32'hbc3e584b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86bf70),
	.w1(32'h3b21fb0b),
	.w2(32'hbaf43ec4),
	.w3(32'hbcc18b21),
	.w4(32'hbb45c3c8),
	.w5(32'hbacacc3b),
	.w6(32'hbca5a50d),
	.w7(32'hbb039cba),
	.w8(32'h3ba4463b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa1507),
	.w1(32'h3c2fcef2),
	.w2(32'h3b9465a3),
	.w3(32'h3b35ffd4),
	.w4(32'h3b56a74f),
	.w5(32'hbbc428e0),
	.w6(32'h39e3555b),
	.w7(32'hbbaec757),
	.w8(32'hbb20ce72),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7853e),
	.w1(32'h3babfbef),
	.w2(32'hbb96658d),
	.w3(32'h3a596fe9),
	.w4(32'hb8bd1f08),
	.w5(32'hbbb8e054),
	.w6(32'hb8b2cb09),
	.w7(32'h3b77bf27),
	.w8(32'hbc1a687c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd9ca),
	.w1(32'hbb69a789),
	.w2(32'h3917ef38),
	.w3(32'hbc3c6277),
	.w4(32'h384a5618),
	.w5(32'hbc9bd755),
	.w6(32'hbc436903),
	.w7(32'hbac17acf),
	.w8(32'hbc36e12d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24479),
	.w1(32'h3b63c1a1),
	.w2(32'hbbe90548),
	.w3(32'hbc489554),
	.w4(32'hb90280d9),
	.w5(32'hbc8ec567),
	.w6(32'hbc0095e1),
	.w7(32'h3bedfd13),
	.w8(32'hbb67ee8e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dfd66),
	.w1(32'hbbb45a64),
	.w2(32'h378cab93),
	.w3(32'hbccc43b9),
	.w4(32'hbb14b557),
	.w5(32'hbbbaf7b5),
	.w6(32'hbc78f4db),
	.w7(32'hbb809abd),
	.w8(32'hbabac17b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51663c),
	.w1(32'hba761287),
	.w2(32'hbc117ce8),
	.w3(32'h3bd83c57),
	.w4(32'h3b109ca4),
	.w5(32'hbba6209e),
	.w6(32'h3bd751e1),
	.w7(32'h3bc2a665),
	.w8(32'hbba29691),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e529b),
	.w1(32'hb9270f05),
	.w2(32'h3b2da3ca),
	.w3(32'hbb846145),
	.w4(32'hbaf0f34d),
	.w5(32'h3b102160),
	.w6(32'hbafa7479),
	.w7(32'h39edac8e),
	.w8(32'h3a15eca7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbe87b),
	.w1(32'h3be22432),
	.w2(32'h3afc478b),
	.w3(32'h3bd5a913),
	.w4(32'h3c95dc73),
	.w5(32'hbca427c3),
	.w6(32'h3b1a8878),
	.w7(32'h3c3af363),
	.w8(32'hba996537),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aa6a8),
	.w1(32'h3c1e9566),
	.w2(32'h3bc704cb),
	.w3(32'h3b1f744f),
	.w4(32'h3bd8ab9a),
	.w5(32'hbc419238),
	.w6(32'h3b31d8de),
	.w7(32'h3b40fb01),
	.w8(32'hb9f8a345),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af893),
	.w1(32'h3a4ffda1),
	.w2(32'hb840a9ad),
	.w3(32'h3a8b8e62),
	.w4(32'h3bb6f37d),
	.w5(32'hbc249958),
	.w6(32'h3b84eee6),
	.w7(32'h3b9ecaf0),
	.w8(32'h3b125e3d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5a732),
	.w1(32'hbbfabb55),
	.w2(32'hbc121781),
	.w3(32'hbb2af9b8),
	.w4(32'hbb50410d),
	.w5(32'hbb86c294),
	.w6(32'hbb7f19ed),
	.w7(32'h3a5d6d90),
	.w8(32'h3a5a24ec),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3ca62),
	.w1(32'h3bd9f8db),
	.w2(32'h3be89d33),
	.w3(32'hbb748889),
	.w4(32'hbc122b69),
	.w5(32'h3b379853),
	.w6(32'h3a17a094),
	.w7(32'h3a290054),
	.w8(32'h3b64fcea),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7a0fc),
	.w1(32'h3c4fa6ad),
	.w2(32'h3b920e8c),
	.w3(32'hbb34a834),
	.w4(32'h3be94cd2),
	.w5(32'hbc06d4b7),
	.w6(32'hbbdb758b),
	.w7(32'h3bdeda87),
	.w8(32'hbbdbd4ef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc227fe0),
	.w1(32'hbb91509d),
	.w2(32'hba96f347),
	.w3(32'hbc218b8a),
	.w4(32'h3bb3dd54),
	.w5(32'h3c115e4c),
	.w6(32'hbb9d5b59),
	.w7(32'hbbac9268),
	.w8(32'hbb6ec263),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb696c),
	.w1(32'h3c4769d0),
	.w2(32'hbacfb292),
	.w3(32'hbc04bc98),
	.w4(32'hba6b37ac),
	.w5(32'hbb1993fb),
	.w6(32'hbaabb72e),
	.w7(32'h3c0e61d9),
	.w8(32'hbb4c1673),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b4a3),
	.w1(32'h3bc5ca1a),
	.w2(32'h3af4c05c),
	.w3(32'hbb0921dd),
	.w4(32'h3b36dc19),
	.w5(32'h3bd57b21),
	.w6(32'hbbe171de),
	.w7(32'h3b8b706c),
	.w8(32'h3b6b0be8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd35b5),
	.w1(32'h3c607789),
	.w2(32'h3b1dfa8f),
	.w3(32'h3b5736e5),
	.w4(32'h3a271b31),
	.w5(32'hbc805020),
	.w6(32'hbbc6922e),
	.w7(32'h3c3ee669),
	.w8(32'h3addf245),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab90f0d),
	.w1(32'h3b3a7919),
	.w2(32'hbaaeaec0),
	.w3(32'h3ad5aea9),
	.w4(32'hbbda2173),
	.w5(32'hbbbb10c1),
	.w6(32'hbaed371c),
	.w7(32'hbb03f5f6),
	.w8(32'h3b0d119f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7dcf2),
	.w1(32'hbb9c4cc3),
	.w2(32'hbad07d6d),
	.w3(32'hbad04c1f),
	.w4(32'hbbb82eb4),
	.w5(32'hbb091574),
	.w6(32'h3a88228b),
	.w7(32'hbb9b97bf),
	.w8(32'hbaf9977c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11b6c7),
	.w1(32'h3be398c2),
	.w2(32'hbad0a712),
	.w3(32'h3b3e6ce7),
	.w4(32'h3c1fe61f),
	.w5(32'hbc5dc1b6),
	.w6(32'h3ba08e0f),
	.w7(32'h3bcd33cd),
	.w8(32'hbb843b45),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b737a0),
	.w1(32'h3b9b27b4),
	.w2(32'h3bb3b798),
	.w3(32'hbbd5d5d0),
	.w4(32'h3aff22fd),
	.w5(32'h3bd75304),
	.w6(32'hbb9e3249),
	.w7(32'h3b3427ed),
	.w8(32'h3b81f6ae),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8459ed),
	.w1(32'hbaebc77f),
	.w2(32'h3c64bfe4),
	.w3(32'h3cb0ee34),
	.w4(32'h3c48cc50),
	.w5(32'hbbc905a2),
	.w6(32'h3c35f723),
	.w7(32'hbad36fae),
	.w8(32'hbbd65a84),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4e79d),
	.w1(32'h3b975d89),
	.w2(32'h3b9afabf),
	.w3(32'hba29b9d5),
	.w4(32'h3a86a24c),
	.w5(32'h3b478fa4),
	.w6(32'h3b7ba9d5),
	.w7(32'h3bedab6c),
	.w8(32'h3935db80),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b283a8e),
	.w1(32'hbb74bbae),
	.w2(32'hbb50403c),
	.w3(32'h3c3361cc),
	.w4(32'hbbbb9a1b),
	.w5(32'hbb67eb4b),
	.w6(32'h3b664514),
	.w7(32'hbbc0761f),
	.w8(32'hbc0da297),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f30b7),
	.w1(32'h3b062499),
	.w2(32'h39799ec9),
	.w3(32'h3b3fdcf9),
	.w4(32'h3ade89f4),
	.w5(32'hbb261242),
	.w6(32'h3b1106e4),
	.w7(32'hbb43eeea),
	.w8(32'h3bba7c0e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65b756),
	.w1(32'h3bba774d),
	.w2(32'hbadc5893),
	.w3(32'h3be33fb4),
	.w4(32'h3bb6f5e3),
	.w5(32'hbc1683ac),
	.w6(32'h3a3e27ed),
	.w7(32'h3bac6150),
	.w8(32'hbbbd50b8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe3bcd),
	.w1(32'hba5a9ec3),
	.w2(32'hbaa770de),
	.w3(32'hbbe9a96d),
	.w4(32'hbc5d52ba),
	.w5(32'hbc2e8fe2),
	.w6(32'hbc04ea1d),
	.w7(32'hbb166fb6),
	.w8(32'h3a85544c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab02bbc),
	.w1(32'h3c4d499d),
	.w2(32'h3c157c87),
	.w3(32'h3ad91ebb),
	.w4(32'h3c1de001),
	.w5(32'hbb287aca),
	.w6(32'hbba1bcf0),
	.w7(32'h3b43f2fa),
	.w8(32'h3b347e58),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dcad2),
	.w1(32'hb8a93c55),
	.w2(32'h3bdc810b),
	.w3(32'h3a973ad0),
	.w4(32'h3be19b50),
	.w5(32'h3c4c8189),
	.w6(32'hbb029200),
	.w7(32'h3ae927bb),
	.w8(32'hbaeeaede),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2a874),
	.w1(32'h3bfbbe68),
	.w2(32'h399f914f),
	.w3(32'h3a9b6d45),
	.w4(32'h3b84e20d),
	.w5(32'hbbd46d37),
	.w6(32'h3a0538d3),
	.w7(32'h3bdb559d),
	.w8(32'hbb809850),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dc28a),
	.w1(32'hba2bfc8e),
	.w2(32'hbbfd8421),
	.w3(32'hba2a05e2),
	.w4(32'hbbc36177),
	.w5(32'hbc99c275),
	.w6(32'hbbea06a1),
	.w7(32'hb9d54679),
	.w8(32'hbc34511a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3688e),
	.w1(32'hbbcec17c),
	.w2(32'h3bc6698b),
	.w3(32'hbbf0b438),
	.w4(32'h3b971fbe),
	.w5(32'hbbb7c3c7),
	.w6(32'hbad9c54c),
	.w7(32'h3b2ff196),
	.w8(32'hba039009),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3570a3),
	.w1(32'h3b4f3038),
	.w2(32'hbaf4666d),
	.w3(32'h3c161b37),
	.w4(32'h3a8673bc),
	.w5(32'h3952f533),
	.w6(32'hb9a1d731),
	.w7(32'hb9c7cdf1),
	.w8(32'hbbbe6b00),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56835d),
	.w1(32'h3b949b5b),
	.w2(32'hb91b45e4),
	.w3(32'hba1d8a44),
	.w4(32'hbbdd5838),
	.w5(32'h3b34855c),
	.w6(32'hbafb4995),
	.w7(32'hbaae4b59),
	.w8(32'hbb77e400),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265dd1),
	.w1(32'hbb272f67),
	.w2(32'h3b070cce),
	.w3(32'hbb941a38),
	.w4(32'h3b8a7a67),
	.w5(32'h3aa2a5ac),
	.w6(32'hbba680e7),
	.w7(32'h3b2d3bbc),
	.w8(32'h3b146204),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03786e),
	.w1(32'h3ab08d07),
	.w2(32'h3aa484d2),
	.w3(32'h398110cd),
	.w4(32'hb9d2370b),
	.w5(32'hba00bb0b),
	.w6(32'h3af4320f),
	.w7(32'h3a1fbd3c),
	.w8(32'hbba03c9d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea801b),
	.w1(32'h3a42601b),
	.w2(32'hba1f1eda),
	.w3(32'hbbc4138f),
	.w4(32'h395f23d1),
	.w5(32'hbc374176),
	.w6(32'hba92134f),
	.w7(32'hb985b445),
	.w8(32'hbad640bb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a209),
	.w1(32'h3c3d9ee6),
	.w2(32'h3bb5d8b9),
	.w3(32'hbbb65c2a),
	.w4(32'h3c310607),
	.w5(32'hbbac0b05),
	.w6(32'hbb1b1145),
	.w7(32'h3bd57d46),
	.w8(32'hbb91457a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a824fe5),
	.w1(32'h3c06ba86),
	.w2(32'h3c0d8b2b),
	.w3(32'hbba1819d),
	.w4(32'hbab94de7),
	.w5(32'hbb71f5c5),
	.w6(32'hbc2e0cf8),
	.w7(32'hbba65542),
	.w8(32'h3af6c57c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04bd21),
	.w1(32'hba940cbc),
	.w2(32'h39383143),
	.w3(32'h3ab8a025),
	.w4(32'hbb7ae05f),
	.w5(32'h3c68ac0f),
	.w6(32'hbb66b60d),
	.w7(32'hbaeb5aed),
	.w8(32'hba66e4f1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a1b64),
	.w1(32'h3b53ed3b),
	.w2(32'hbaa38960),
	.w3(32'h3c0d09e6),
	.w4(32'h3998a626),
	.w5(32'hbc512831),
	.w6(32'h3b1454a2),
	.w7(32'h3b3f873a),
	.w8(32'hbb215c02),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ea2ac),
	.w1(32'h3b43ce5c),
	.w2(32'h3b397358),
	.w3(32'h3b483004),
	.w4(32'hbbc3e742),
	.w5(32'hbc1b152a),
	.w6(32'h3c077898),
	.w7(32'h3ba7f103),
	.w8(32'hbaaf3677),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd52c2),
	.w1(32'h3bc2c225),
	.w2(32'hbaadbc42),
	.w3(32'hbbcd9606),
	.w4(32'h3bfd8f55),
	.w5(32'hbba1d7f0),
	.w6(32'hbbbacefb),
	.w7(32'h3c1bd631),
	.w8(32'h3b498b1a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9833159),
	.w1(32'h3b1001e8),
	.w2(32'h3b91f8ac),
	.w3(32'h3bedd2fc),
	.w4(32'h3b8cb561),
	.w5(32'h3c1dc6f4),
	.w6(32'h3b826ddf),
	.w7(32'hbb20831e),
	.w8(32'h3bbbd6ab),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beabf8d),
	.w1(32'h3bc23156),
	.w2(32'h3ba3c9b9),
	.w3(32'h3c3afe0c),
	.w4(32'hbb0f4f09),
	.w5(32'hbb0ef592),
	.w6(32'h3b95d2b6),
	.w7(32'h3a16341b),
	.w8(32'hba8c98f0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41612d),
	.w1(32'h3b0e445c),
	.w2(32'h3a782630),
	.w3(32'h3b66a18f),
	.w4(32'hbb9b66b9),
	.w5(32'h3b98ecfb),
	.w6(32'hbac7cbd6),
	.w7(32'h3b3ac03b),
	.w8(32'hbb1a3274),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba858f49),
	.w1(32'h3b7f00b7),
	.w2(32'h3ab40a97),
	.w3(32'hbba9687a),
	.w4(32'h392c96f8),
	.w5(32'hbc0ad8bb),
	.w6(32'hbad780f7),
	.w7(32'h39ddb0c0),
	.w8(32'hb9d73283),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95e9e4),
	.w1(32'h3c0c98af),
	.w2(32'h395a6f2f),
	.w3(32'h3af07734),
	.w4(32'h3c2b164f),
	.w5(32'hbc4907b9),
	.w6(32'hbbb7e867),
	.w7(32'h3c079117),
	.w8(32'h3ba31f91),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2f5e),
	.w1(32'h3a3adfde),
	.w2(32'hb9c41331),
	.w3(32'h3bfa5e8c),
	.w4(32'hbba01416),
	.w5(32'h3a783894),
	.w6(32'hbb1b2198),
	.w7(32'hbb3bb30d),
	.w8(32'hba220d7f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dc3ca),
	.w1(32'h3bbc416f),
	.w2(32'h3bea8992),
	.w3(32'h3c07bc56),
	.w4(32'h3b1200e6),
	.w5(32'h3b8e10f0),
	.w6(32'h3bb6d35e),
	.w7(32'h3b526de5),
	.w8(32'h3b626962),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8585cd),
	.w1(32'h3c3dce70),
	.w2(32'h3c6b4a53),
	.w3(32'h3a99e7f2),
	.w4(32'h3c1c6152),
	.w5(32'hbbb63d6b),
	.w6(32'h3acd84c7),
	.w7(32'hbb8d34c8),
	.w8(32'hbb889935),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3c9ac),
	.w1(32'h393c514b),
	.w2(32'hbc19de87),
	.w3(32'hba5821f7),
	.w4(32'h3b6f5f76),
	.w5(32'hbb9ee84f),
	.w6(32'hbbad48a7),
	.w7(32'hbb0daef3),
	.w8(32'hbc45a493),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc845b0),
	.w1(32'h3c807ddd),
	.w2(32'h3bebbcac),
	.w3(32'hbae3f93b),
	.w4(32'hb933e3bf),
	.w5(32'hbc834a9b),
	.w6(32'hbb80b7d8),
	.w7(32'h3c316a86),
	.w8(32'h3c022baa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df473),
	.w1(32'hbb9466f8),
	.w2(32'hba062c52),
	.w3(32'hb8efecfe),
	.w4(32'hbc3a25b7),
	.w5(32'hbc6577df),
	.w6(32'hbb9ada48),
	.w7(32'hbc10d717),
	.w8(32'hbc01bf86),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a9285),
	.w1(32'hb9864c17),
	.w2(32'h3b52b506),
	.w3(32'hbbd99b9b),
	.w4(32'h3b533991),
	.w5(32'hbbd95195),
	.w6(32'hbc13459d),
	.w7(32'hba9dfdc4),
	.w8(32'hbb96270a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf02064),
	.w1(32'h3c0bcec1),
	.w2(32'h3bc1c8a3),
	.w3(32'hbc8a76fb),
	.w4(32'h3c572f57),
	.w5(32'hbc7b27fd),
	.w6(32'hbad6fffb),
	.w7(32'h3c2f21e0),
	.w8(32'hb9c02260),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba53ca8),
	.w1(32'h3be9e9b8),
	.w2(32'h3c2cdb43),
	.w3(32'hbbd478a4),
	.w4(32'hbb40eb61),
	.w5(32'h3b09e95a),
	.w6(32'hbb0c6238),
	.w7(32'hbb139b2a),
	.w8(32'hbb5fbca7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f94f4),
	.w1(32'hb8af52aa),
	.w2(32'hbaf71ab2),
	.w3(32'hbb5a4fdf),
	.w4(32'hbb661b47),
	.w5(32'h3b465d41),
	.w6(32'hbb05c776),
	.w7(32'hbb9d19b9),
	.w8(32'hbc07e8fd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b8bc),
	.w1(32'h3a5b9036),
	.w2(32'h3b1542ce),
	.w3(32'hbbcee059),
	.w4(32'hbb93d836),
	.w5(32'h3c14f1bf),
	.w6(32'hba766027),
	.w7(32'hba80c807),
	.w8(32'h3bdd4c35),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d1e22),
	.w1(32'hba59da44),
	.w2(32'hbb2a8f40),
	.w3(32'h3b1487b8),
	.w4(32'h3b362757),
	.w5(32'hbbc82b9f),
	.w6(32'h3bda8767),
	.w7(32'h3b887d9c),
	.w8(32'hbad83505),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ff932),
	.w1(32'h3bedca16),
	.w2(32'h3bf951bc),
	.w3(32'hbb8255dd),
	.w4(32'h3c44b102),
	.w5(32'hbbe96d3d),
	.w6(32'hb9888bfc),
	.w7(32'h3a2ca859),
	.w8(32'hba5cca3d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6dc69),
	.w1(32'h3ad087ac),
	.w2(32'h3b3381ee),
	.w3(32'hbc1269a0),
	.w4(32'h3bf8bd6e),
	.w5(32'hbc983b1a),
	.w6(32'hbb4d65d6),
	.w7(32'h3a94d347),
	.w8(32'hbc070818),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba855b),
	.w1(32'hb89b3b07),
	.w2(32'hbb68d83d),
	.w3(32'hbc14f683),
	.w4(32'hbb4768ca),
	.w5(32'hbb58afec),
	.w6(32'hbb7af68f),
	.w7(32'h3a523d0a),
	.w8(32'hbb8522b6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2103d5),
	.w1(32'hba87d5dc),
	.w2(32'h3c1bf634),
	.w3(32'hbbf7eea6),
	.w4(32'h3b3f2023),
	.w5(32'h3c3194ad),
	.w6(32'hbc214da8),
	.w7(32'h38b7d034),
	.w8(32'h3b438022),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396bca22),
	.w1(32'hbb7cd3b2),
	.w2(32'hbbae9e24),
	.w3(32'h3b188675),
	.w4(32'hbbf15e25),
	.w5(32'hbc8e435e),
	.w6(32'hb9b1160a),
	.w7(32'hbc0be4da),
	.w8(32'hbbd7c424),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18acb7),
	.w1(32'h3b7500e5),
	.w2(32'h399e7379),
	.w3(32'hbb927755),
	.w4(32'h3b6af146),
	.w5(32'hbbeb3289),
	.w6(32'h3a53f16a),
	.w7(32'h3bce1652),
	.w8(32'h3b60345b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7faa8),
	.w1(32'hbb0218cb),
	.w2(32'h3b08582d),
	.w3(32'h3ba02022),
	.w4(32'h3b9161fe),
	.w5(32'hbba028b6),
	.w6(32'h3b3810bd),
	.w7(32'h3aa91d35),
	.w8(32'h3b28a27a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07acfd),
	.w1(32'h3c11c183),
	.w2(32'h3bd71f05),
	.w3(32'hbb16ab78),
	.w4(32'h3c59cdbc),
	.w5(32'hbbda00b8),
	.w6(32'hbb393998),
	.w7(32'h3c01e640),
	.w8(32'h3ac5918a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87a0e2),
	.w1(32'hbb623c29),
	.w2(32'hbb86326c),
	.w3(32'hbc089bcb),
	.w4(32'h3bbebf42),
	.w5(32'h3c13a95e),
	.w6(32'hbc3e9a53),
	.w7(32'hba862346),
	.w8(32'hbc445b78),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd885d7),
	.w1(32'hba91cce7),
	.w2(32'hbb2ff1cf),
	.w3(32'hbbacdcd5),
	.w4(32'hbb4e8bff),
	.w5(32'hbbe234bb),
	.w6(32'hbbba1083),
	.w7(32'hba9dd0e3),
	.w8(32'hbbd5653d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22da0a),
	.w1(32'hbb4f20cb),
	.w2(32'hbb72b22d),
	.w3(32'hbb554720),
	.w4(32'hba90acc8),
	.w5(32'hbc1767d1),
	.w6(32'hbb8296bc),
	.w7(32'hbb9fd23b),
	.w8(32'hbc2ab000),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cf589),
	.w1(32'h3a9b6f0a),
	.w2(32'h3bfc89c3),
	.w3(32'hbbe42d6b),
	.w4(32'h3b9056b6),
	.w5(32'h3c7c0e98),
	.w6(32'hbbe89779),
	.w7(32'h3b1794b6),
	.w8(32'h3b38c13e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aaa68),
	.w1(32'h3c718135),
	.w2(32'hb9886742),
	.w3(32'h3bf4b8a2),
	.w4(32'h3c968250),
	.w5(32'hbbc06cc0),
	.w6(32'hbae233b1),
	.w7(32'h3bfccf43),
	.w8(32'hbbb0675d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ee18d),
	.w1(32'h3b828b46),
	.w2(32'h3bd28a91),
	.w3(32'h3a16fdfa),
	.w4(32'h3ba0067f),
	.w5(32'h3ca89d1f),
	.w6(32'hbbc69a3e),
	.w7(32'hba74d2ff),
	.w8(32'h3bba682e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc48c8),
	.w1(32'h3aaa7419),
	.w2(32'h39ee721a),
	.w3(32'h3ba5039c),
	.w4(32'hbad68658),
	.w5(32'hbbf0e2a7),
	.w6(32'hbb2e0ec1),
	.w7(32'h3a956ac2),
	.w8(32'h3b575d51),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0652a),
	.w1(32'hbac0a6b9),
	.w2(32'h3ac91b59),
	.w3(32'h3a0f5ba8),
	.w4(32'h3ba2a8c9),
	.w5(32'hbbb94b89),
	.w6(32'h39eb034f),
	.w7(32'h3aa2a3e1),
	.w8(32'h3a8c44ab),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0b0f8),
	.w1(32'hbb823fbf),
	.w2(32'h3b73ec68),
	.w3(32'h39eb319e),
	.w4(32'hba358f8a),
	.w5(32'h3b05041c),
	.w6(32'h3b1afc71),
	.w7(32'h3b005a3a),
	.w8(32'h3b4d2cb9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9308df),
	.w1(32'hbc08fedc),
	.w2(32'h3b02d87d),
	.w3(32'hbb8b8515),
	.w4(32'hbbf908bd),
	.w5(32'h3aa5e8e7),
	.w6(32'h3bb211e5),
	.w7(32'hbb579252),
	.w8(32'hbae1bfad),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99175fb),
	.w1(32'h3b4a1f88),
	.w2(32'hbb8ec267),
	.w3(32'hbbd72848),
	.w4(32'hbb9db4fe),
	.w5(32'h3c07d984),
	.w6(32'hb9d61aa0),
	.w7(32'hba724ef9),
	.w8(32'hb952659d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9504d),
	.w1(32'hbb0a5c02),
	.w2(32'hbb82e7ab),
	.w3(32'hbbea6dd1),
	.w4(32'h3c135a01),
	.w5(32'h3989778a),
	.w6(32'hbb924406),
	.w7(32'hb99bcbfd),
	.w8(32'h3b5e30f2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f1f578),
	.w1(32'hbac1b642),
	.w2(32'hbb9c1086),
	.w3(32'hbb90186d),
	.w4(32'hbbd6623a),
	.w5(32'hbb559cd8),
	.w6(32'hbaf92b29),
	.w7(32'h38e7f67b),
	.w8(32'h389c90e3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6584),
	.w1(32'h3a70ed0b),
	.w2(32'h39d2e575),
	.w3(32'hbb9309d9),
	.w4(32'hb7f1cac7),
	.w5(32'hbbb43fb9),
	.w6(32'h3b7207c1),
	.w7(32'h3b019322),
	.w8(32'hba83e19b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffc302),
	.w1(32'h3c9b103c),
	.w2(32'hbb82548a),
	.w3(32'hbc1ee855),
	.w4(32'h3ccfb8cd),
	.w5(32'hbc4d0975),
	.w6(32'hbbc860d4),
	.w7(32'h3cb17dcc),
	.w8(32'hbae0ba0a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe07415),
	.w1(32'h3bc601d4),
	.w2(32'hbbbee027),
	.w3(32'hbb98b86d),
	.w4(32'h3b807141),
	.w5(32'hbc86c610),
	.w6(32'hbb6d2fec),
	.w7(32'h3c0ed4d5),
	.w8(32'hbb841b0b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac60243),
	.w1(32'h391e9fa0),
	.w2(32'h3b02bab6),
	.w3(32'hbc238cbb),
	.w4(32'h3a77e94a),
	.w5(32'h3c2b2d5b),
	.w6(32'hbb677bcb),
	.w7(32'hbacb205e),
	.w8(32'hba683cf7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3124f4),
	.w1(32'h3ac00f8b),
	.w2(32'h3b4f0b8d),
	.w3(32'hbb4b5f32),
	.w4(32'hbc19ad0b),
	.w5(32'h3bc232b5),
	.w6(32'hbbb4fd57),
	.w7(32'hbac1cff9),
	.w8(32'hbb203687),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e3dc),
	.w1(32'hbb7c97ce),
	.w2(32'hbb02e6f4),
	.w3(32'h3a9fd75a),
	.w4(32'hbb6213b4),
	.w5(32'hbac92249),
	.w6(32'hbbefd600),
	.w7(32'hbb5b34e5),
	.w8(32'hbbf63c13),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099387),
	.w1(32'h3c7f5f8b),
	.w2(32'h3a4b7eec),
	.w3(32'hbb659aaa),
	.w4(32'h3c8c40c0),
	.w5(32'hbc308fd2),
	.w6(32'hbb1bbfc9),
	.w7(32'h3c7158b0),
	.w8(32'h3c30b2d2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a380),
	.w1(32'h3be6f0cc),
	.w2(32'h3b1151ab),
	.w3(32'h3be92ef7),
	.w4(32'h3babef21),
	.w5(32'hbc0f7321),
	.w6(32'h3bd80ec8),
	.w7(32'h3c087bfa),
	.w8(32'hbb81219c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4221a7),
	.w1(32'h3c860e8e),
	.w2(32'hbb0f74ed),
	.w3(32'hbc636cde),
	.w4(32'h3cba5b59),
	.w5(32'hbcaadcd5),
	.w6(32'hbc008ae7),
	.w7(32'h3c944da0),
	.w8(32'hbba64663),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf194ce),
	.w1(32'h3b6fbdfe),
	.w2(32'h3a93781f),
	.w3(32'hbc30b333),
	.w4(32'h3b95e00e),
	.w5(32'hbc25be23),
	.w6(32'hbb9d440e),
	.w7(32'h3a9f3826),
	.w8(32'hbbc8d8df),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855e8a),
	.w1(32'hba938652),
	.w2(32'h3a24f459),
	.w3(32'h3acf9bd6),
	.w4(32'hb8b43a31),
	.w5(32'h3c38fb35),
	.w6(32'hb9eb4e88),
	.w7(32'h3adc19fc),
	.w8(32'hb99d106e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaec31e),
	.w1(32'hbc0ab166),
	.w2(32'h3b28a03e),
	.w3(32'h3be5787b),
	.w4(32'hbb44d915),
	.w5(32'h3bc83e6d),
	.w6(32'hbaafe9dd),
	.w7(32'hbbbdb055),
	.w8(32'hba721d94),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cfbd1),
	.w1(32'hbba4a45a),
	.w2(32'h3afb2077),
	.w3(32'h3bf1490e),
	.w4(32'hbb870c5e),
	.w5(32'hbbd19bf6),
	.w6(32'h3bcedde0),
	.w7(32'hbbb878ef),
	.w8(32'hbb172f21),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38050c),
	.w1(32'h3b89bcdf),
	.w2(32'hbb60c735),
	.w3(32'hbbb3da46),
	.w4(32'hbaa2791e),
	.w5(32'hbb80433e),
	.w6(32'h3a4dc16d),
	.w7(32'hbafabd95),
	.w8(32'hbaffb5e5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba406463),
	.w1(32'h3c4e9e7d),
	.w2(32'h3a8d8daf),
	.w3(32'h3938fe6d),
	.w4(32'h3c265e8d),
	.w5(32'hbc98680a),
	.w6(32'h3a035284),
	.w7(32'h3c735f6d),
	.w8(32'h3b276257),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390d0a),
	.w1(32'hbab821e9),
	.w2(32'h3a96eeee),
	.w3(32'h3b11cb61),
	.w4(32'hbc122be3),
	.w5(32'hbb8574f4),
	.w6(32'h3c2de701),
	.w7(32'h3a9b5b06),
	.w8(32'h3b3ad2d9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb52572),
	.w1(32'h3b088097),
	.w2(32'h3a1e6fa0),
	.w3(32'h3bf0153e),
	.w4(32'h3b3d9b4c),
	.w5(32'h39b23a15),
	.w6(32'h3bf40e76),
	.w7(32'h3a1967bc),
	.w8(32'hba671d42),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1acd1),
	.w1(32'hb9c8eb5c),
	.w2(32'hb974c7d1),
	.w3(32'h3a21eb7d),
	.w4(32'h3a5c37d4),
	.w5(32'h3931ca56),
	.w6(32'h3a03a8a0),
	.w7(32'h3a1867e2),
	.w8(32'hba1d8c9e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63c1e1c),
	.w1(32'h35488d57),
	.w2(32'h37be9678),
	.w3(32'h375074e0),
	.w4(32'h3725015f),
	.w5(32'h37df37a5),
	.w6(32'h382542bd),
	.w7(32'h38176623),
	.w8(32'h385ae7d0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3e44c),
	.w1(32'hba6ce1ce),
	.w2(32'hb90d23c4),
	.w3(32'hba878237),
	.w4(32'h3a511419),
	.w5(32'h3aa974b7),
	.w6(32'hbae5bca5),
	.w7(32'hb9d4e077),
	.w8(32'h3ac1edbe),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75cafd5),
	.w1(32'hb7b659ed),
	.w2(32'h38669975),
	.w3(32'h3635fd8f),
	.w4(32'hb78fa3ad),
	.w5(32'h38786ec6),
	.w6(32'h38727248),
	.w7(32'h3810cf35),
	.w8(32'h38b3c2b4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5810f4),
	.w1(32'hba34a44d),
	.w2(32'hbabe0580),
	.w3(32'hba6862a5),
	.w4(32'h3997fb0a),
	.w5(32'hb9e54d73),
	.w6(32'hba1b79f6),
	.w7(32'hba72aa98),
	.w8(32'h3a2cd038),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d959d),
	.w1(32'h39c746e5),
	.w2(32'h3af25263),
	.w3(32'h3a0ed5cf),
	.w4(32'hba0515ea),
	.w5(32'h3a84fc96),
	.w6(32'hbab80ca1),
	.w7(32'hbb2e2703),
	.w8(32'hbb22c9c7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba1fe0),
	.w1(32'h3ab88f70),
	.w2(32'h3a91f581),
	.w3(32'h3a8cf944),
	.w4(32'h3a25a287),
	.w5(32'h39f6519c),
	.w6(32'h3895418d),
	.w7(32'hba061a18),
	.w8(32'hba7d649c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8f643),
	.w1(32'h39aadb57),
	.w2(32'hb9ee7810),
	.w3(32'h39733770),
	.w4(32'h392b5fd0),
	.w5(32'hb9f8dea5),
	.w6(32'hb93e5f61),
	.w7(32'hb975c8de),
	.w8(32'hba6827f6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1056bf),
	.w1(32'h3ac62a82),
	.w2(32'h3acc0ad2),
	.w3(32'h3ac8cf79),
	.w4(32'h3943d504),
	.w5(32'h3a7d2ac8),
	.w6(32'h3a3f51b2),
	.w7(32'hba80cdae),
	.w8(32'hb8e0fc9e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f716e5),
	.w1(32'h3a894045),
	.w2(32'h3ac2c679),
	.w3(32'h3904c918),
	.w4(32'h3aa98d45),
	.w5(32'h3af269e9),
	.w6(32'h39235b98),
	.w7(32'h3a386a2e),
	.w8(32'h3ab3a006),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0c317),
	.w1(32'h3ad4ccba),
	.w2(32'h3ad68631),
	.w3(32'h3b6f1c4f),
	.w4(32'h3b6537de),
	.w5(32'h3af30ed1),
	.w6(32'h3b811f90),
	.w7(32'h3b3494c1),
	.w8(32'hba3a3c95),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62125b5),
	.w1(32'hb71a4efc),
	.w2(32'h3762e206),
	.w3(32'h366a090c),
	.w4(32'h364352ed),
	.w5(32'h3761f7fe),
	.w6(32'h378d984c),
	.w7(32'h3730045d),
	.w8(32'h376e9986),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8659c85),
	.w1(32'hb8ca14ae),
	.w2(32'h368d9480),
	.w3(32'hb8924102),
	.w4(32'hb89ff91c),
	.w5(32'hb85a6794),
	.w6(32'hb7ba95c4),
	.w7(32'hb8bee4e7),
	.w8(32'hb80c190f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c67b6),
	.w1(32'h3b2f8b1e),
	.w2(32'h39f7a8e2),
	.w3(32'hb85b71c6),
	.w4(32'h3af15b4e),
	.w5(32'hb80a1bbc),
	.w6(32'hbae4d4aa),
	.w7(32'h3987b395),
	.w8(32'hbb2592dd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacfbfe),
	.w1(32'h39509adc),
	.w2(32'h3a2d4861),
	.w3(32'hbb501248),
	.w4(32'hba7a4e55),
	.w5(32'h39d3a65d),
	.w6(32'hbb4e6329),
	.w7(32'hbb0a38f3),
	.w8(32'hbae2cd04),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add55c6),
	.w1(32'h3b358185),
	.w2(32'h3b233141),
	.w3(32'h3a9b6cae),
	.w4(32'h3ad94580),
	.w5(32'h3b2f0a6d),
	.w6(32'h3ac13d6d),
	.w7(32'h3aa903b8),
	.w8(32'h3a30ba7e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc41b2),
	.w1(32'h3a8c5771),
	.w2(32'h3ac2f17d),
	.w3(32'h3b29dc81),
	.w4(32'h3b2b0b50),
	.w5(32'h3949742f),
	.w6(32'hb81b9474),
	.w7(32'hb98b0d4e),
	.w8(32'hb9faad6e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935b887),
	.w1(32'h38bfb3a6),
	.w2(32'h382cbdcc),
	.w3(32'h374f921b),
	.w4(32'hb96d5994),
	.w5(32'h393b5226),
	.w6(32'hb93cfced),
	.w7(32'hb99f2153),
	.w8(32'h38e7beb7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d7c5a),
	.w1(32'h3921e388),
	.w2(32'h39aa58dd),
	.w3(32'hba30afce),
	.w4(32'hb85acc51),
	.w5(32'h3a2eaa66),
	.w6(32'hba23fe5c),
	.w7(32'hb9b3e3ea),
	.w8(32'h39baec95),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad0479),
	.w1(32'h3ad3b631),
	.w2(32'hba12b2b5),
	.w3(32'hba2bc593),
	.w4(32'h3b15884d),
	.w5(32'hbaaa6c3a),
	.w6(32'hbb8e4109),
	.w7(32'hbb53f7e9),
	.w8(32'hbb0be310),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05fce4),
	.w1(32'hbaad7ed7),
	.w2(32'hb9101653),
	.w3(32'h3b023dc6),
	.w4(32'h3ac30fb2),
	.w5(32'h3aaf416b),
	.w6(32'h38b3ccd8),
	.w7(32'h38fedca3),
	.w8(32'hb9397f56),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148ad7),
	.w1(32'h37eda6e7),
	.w2(32'hb92e11fe),
	.w3(32'hbb5dddd9),
	.w4(32'h3a0536a2),
	.w5(32'h3925f3c4),
	.w6(32'hbbdddb5e),
	.w7(32'hbb21db15),
	.w8(32'hbabcecad),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c52b50),
	.w1(32'h39d86bf2),
	.w2(32'h3a7adca5),
	.w3(32'h3937bbe9),
	.w4(32'hba5d11e1),
	.w5(32'hb92166dd),
	.w6(32'hb975cb2b),
	.w7(32'hbab7accc),
	.w8(32'hbae10ba5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d7fae),
	.w1(32'hb8d3b66c),
	.w2(32'h3aa15799),
	.w3(32'h380eed6e),
	.w4(32'hba6258ef),
	.w5(32'h3a11ba69),
	.w6(32'h3accaeeb),
	.w7(32'hba0d7d97),
	.w8(32'hb8bd2247),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370bc81e),
	.w1(32'h36bc12f9),
	.w2(32'h37541b04),
	.w3(32'h3793b8b6),
	.w4(32'h370f3e35),
	.w5(32'h379585d5),
	.w6(32'h37c00b24),
	.w7(32'h37469dd4),
	.w8(32'h379dd5f2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b8403b),
	.w1(32'h374079f3),
	.w2(32'h37343123),
	.w3(32'h37b63929),
	.w4(32'h3756393c),
	.w5(32'h37579d4f),
	.w6(32'h37d52edb),
	.w7(32'h37a7bc9f),
	.w8(32'h37a37c09),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867387),
	.w1(32'h3a6132c3),
	.w2(32'h3a08700e),
	.w3(32'h39b20518),
	.w4(32'hba2cb555),
	.w5(32'hbaee0947),
	.w6(32'hba19365e),
	.w7(32'hba2b080b),
	.w8(32'hbaa5341e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365ea166),
	.w1(32'h37148053),
	.w2(32'h37cf6d24),
	.w3(32'h37c165e2),
	.w4(32'h36ec0428),
	.w5(32'h379f9f11),
	.w6(32'h37d08842),
	.w7(32'h379b1329),
	.w8(32'h380a476a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a607f90),
	.w1(32'hba643785),
	.w2(32'hbac50474),
	.w3(32'h3a80b578),
	.w4(32'hb97edac4),
	.w5(32'hbaf32bb1),
	.w6(32'h38a26c6a),
	.w7(32'hb90cf46d),
	.w8(32'hbabb9b31),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ed3ad),
	.w1(32'h3ae9a797),
	.w2(32'h3b0397f4),
	.w3(32'hbb48d5e3),
	.w4(32'hb9ffe13f),
	.w5(32'h3ac99920),
	.w6(32'hbad6f430),
	.w7(32'hbaf0084c),
	.w8(32'h3a848967),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3583c),
	.w1(32'h3ac17151),
	.w2(32'h3a705bd3),
	.w3(32'h3a828b13),
	.w4(32'h3a3f7da6),
	.w5(32'h3a30d684),
	.w6(32'hb927bdc7),
	.w7(32'hb90f9bb2),
	.w8(32'hba44fc64),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381dd4de),
	.w1(32'h37928130),
	.w2(32'h375261f6),
	.w3(32'h3849ed3f),
	.w4(32'h383be97e),
	.w5(32'h38086e44),
	.w6(32'h388aa154),
	.w7(32'h38632c08),
	.w8(32'h38069e28),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53f9be),
	.w1(32'hb911df49),
	.w2(32'hba465b67),
	.w3(32'hbb392350),
	.w4(32'h3ad7ce4e),
	.w5(32'hbab33ebb),
	.w6(32'hbbe66be8),
	.w7(32'hbad33637),
	.w8(32'hbb079fa5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5a69),
	.w1(32'hba0c6fdc),
	.w2(32'hb8ed0aec),
	.w3(32'hb9a27eba),
	.w4(32'h38a9c6fd),
	.w5(32'h373bb4e9),
	.w6(32'hbaa8660c),
	.w7(32'hba6e0950),
	.w8(32'hba7e6ba9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9290f0a),
	.w1(32'hb91ea96d),
	.w2(32'hb91947cd),
	.w3(32'hb8ea4a5b),
	.w4(32'hb93b7545),
	.w5(32'hb902e8d5),
	.w6(32'hb8bc5358),
	.w7(32'hb8f61dbd),
	.w8(32'hb888e650),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f857a),
	.w1(32'hba1919b7),
	.w2(32'hba45b096),
	.w3(32'h37b17880),
	.w4(32'h39ec8223),
	.w5(32'hba143d52),
	.w6(32'hbabd7932),
	.w7(32'hba1b498c),
	.w8(32'hba7846b3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793cdd8),
	.w1(32'hb474c1c5),
	.w2(32'h38d31478),
	.w3(32'hb8bd1a37),
	.w4(32'h36313a02),
	.w5(32'h38dc66a3),
	.w6(32'hb7a9f887),
	.w7(32'h3865886a),
	.w8(32'h39130ab0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a185eb7),
	.w1(32'h39b03361),
	.w2(32'h36ed24f9),
	.w3(32'h39e31c24),
	.w4(32'h38019eb0),
	.w5(32'hb9231796),
	.w6(32'h3984eddb),
	.w7(32'hb8c23c2a),
	.w8(32'hb968048b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36eb3194),
	.w1(32'hb66cf8b8),
	.w2(32'h379bf70f),
	.w3(32'h37a8c34c),
	.w4(32'h36dca810),
	.w5(32'h378c3373),
	.w6(32'h382a4bc5),
	.w7(32'h37eecef3),
	.w8(32'hb5657f08),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380fa655),
	.w1(32'hb44f5190),
	.w2(32'h35f10205),
	.w3(32'h37d7aafa),
	.w4(32'h36d97c31),
	.w5(32'h375c9617),
	.w6(32'h37cdb2d6),
	.w7(32'h3788f60a),
	.w8(32'h3801cc93),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e33f78),
	.w1(32'h39359d00),
	.w2(32'hb9b185f0),
	.w3(32'h3a346936),
	.w4(32'h39bcacfd),
	.w5(32'hb9bfd204),
	.w6(32'h39e2a774),
	.w7(32'h397e72c9),
	.w8(32'hba252b49),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0853ae),
	.w1(32'h3a4f91c9),
	.w2(32'hb9ddde4a),
	.w3(32'h3aceab80),
	.w4(32'h3a63ff2b),
	.w5(32'hb9d65b07),
	.w6(32'h39dfd7f9),
	.w7(32'hba444796),
	.w8(32'hb9b61a47),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf78f9),
	.w1(32'hba89a63f),
	.w2(32'h3a5b9e3c),
	.w3(32'hba1924fa),
	.w4(32'hb93b7722),
	.w5(32'h3a14a22b),
	.w6(32'hbabc70b7),
	.w7(32'hba1992cf),
	.w8(32'hb8773090),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27fbc0),
	.w1(32'h3a3727f7),
	.w2(32'hb84b41ac),
	.w3(32'h3afb114e),
	.w4(32'h3abf48ab),
	.w5(32'h39ac7534),
	.w6(32'h3a58d7f7),
	.w7(32'hb96d1f17),
	.w8(32'hb9270eed),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05be13),
	.w1(32'h3a01729b),
	.w2(32'h38cbd7dd),
	.w3(32'h3a097206),
	.w4(32'h39f0d706),
	.w5(32'h3903cb74),
	.w6(32'h399b0a2b),
	.w7(32'h39929500),
	.w8(32'h39121008),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea1cf6),
	.w1(32'h38e3c57e),
	.w2(32'hb6d3e346),
	.w3(32'hb9852fe8),
	.w4(32'hb91955bc),
	.w5(32'hb682c12c),
	.w6(32'hb811c07b),
	.w7(32'h385d7f80),
	.w8(32'h39621661),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb745f069),
	.w1(32'hb790b440),
	.w2(32'hb7083d0b),
	.w3(32'hb662430a),
	.w4(32'hb74e9792),
	.w5(32'hb6a79156),
	.w6(32'h36f8d4d9),
	.w7(32'h3421a73f),
	.w8(32'h368f64ba),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b03bda),
	.w1(32'h37a946b1),
	.w2(32'h37913246),
	.w3(32'h372dc436),
	.w4(32'hb74898aa),
	.w5(32'hb8162d6d),
	.w6(32'h38196b9d),
	.w7(32'h3753d570),
	.w8(32'hb839bd9e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70d95d),
	.w1(32'h3890e390),
	.w2(32'h38fe20c9),
	.w3(32'hba407a90),
	.w4(32'hba7b517a),
	.w5(32'h3a4a1213),
	.w6(32'hbabb1e79),
	.w7(32'hbaca4ba9),
	.w8(32'h3905fbd8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c3550f),
	.w1(32'h383caf30),
	.w2(32'h37cde8d8),
	.w3(32'hb888d935),
	.w4(32'hb755b50a),
	.w5(32'h3713b6aa),
	.w6(32'hb9094a6e),
	.w7(32'hb7a705fc),
	.w8(32'hb7b9908f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e50ee1),
	.w1(32'h3a03c239),
	.w2(32'hb9debae4),
	.w3(32'h3a297ef8),
	.w4(32'h3a04605c),
	.w5(32'hba17fa2d),
	.w6(32'hb902e81a),
	.w7(32'h399b3512),
	.w8(32'hba56ebd6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e328b7),
	.w1(32'hba10d919),
	.w2(32'hba04c94b),
	.w3(32'hb9f8baf0),
	.w4(32'h3907f616),
	.w5(32'h39e74582),
	.w6(32'hba317ed6),
	.w7(32'h39b3c5ae),
	.w8(32'h39f8f982),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bd1ee9),
	.w1(32'hb70a556a),
	.w2(32'hb50da7ac),
	.w3(32'hb6d24641),
	.w4(32'h35cbd549),
	.w5(32'hb5ac2568),
	.w6(32'hb5d86091),
	.w7(32'h34b87a8a),
	.w8(32'h37411881),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ffa00),
	.w1(32'h3a44e938),
	.w2(32'h39c4856c),
	.w3(32'h3ab22029),
	.w4(32'h3aaa1fa7),
	.w5(32'h3a404508),
	.w6(32'h3a81c88a),
	.w7(32'h3a2eff37),
	.w8(32'h396a0151),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d27d28),
	.w1(32'h38c8927c),
	.w2(32'h38414990),
	.w3(32'hb912c3d2),
	.w4(32'hb7bf8071),
	.w5(32'h3790fd0f),
	.w6(32'h38e0357f),
	.w7(32'h38dc953a),
	.w8(32'h39544c7c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c859),
	.w1(32'h39af3c26),
	.w2(32'hba1ae22c),
	.w3(32'h3a382cf9),
	.w4(32'hb986a5b0),
	.w5(32'h3a0da3f7),
	.w6(32'hbb19b78e),
	.w7(32'hbb6b0808),
	.w8(32'h3aff8679),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c6ff5),
	.w1(32'hb8d8e5fa),
	.w2(32'hb919f031),
	.w3(32'hb8a473f0),
	.w4(32'hb95b6787),
	.w5(32'hb957c691),
	.w6(32'hb882d160),
	.w7(32'hb90c6998),
	.w8(32'hb90ac37b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ccf4b),
	.w1(32'h3ae30d5d),
	.w2(32'h3b132a1c),
	.w3(32'hba97295c),
	.w4(32'h3a037f8c),
	.w5(32'h3a920147),
	.w6(32'hbb3d3c1b),
	.w7(32'hbafd053c),
	.w8(32'hbadc0082),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule