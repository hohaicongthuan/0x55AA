module layer_10_featuremap_278(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa795f9),
	.w1(32'h3b974380),
	.w2(32'h3bfad5c5),
	.w3(32'hbbcde019),
	.w4(32'hbbae3de2),
	.w5(32'hbbd61fc4),
	.w6(32'hbc836668),
	.w7(32'hbbea84c1),
	.w8(32'hb9858b24),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56e752),
	.w1(32'h3bc10346),
	.w2(32'h3b6b90a3),
	.w3(32'hbab726b4),
	.w4(32'h3b8c4e44),
	.w5(32'hb9d3f1fe),
	.w6(32'hbb976c38),
	.w7(32'h3a92ee48),
	.w8(32'h3a1a20ba),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5bc6),
	.w1(32'hbc02249b),
	.w2(32'hbc02136e),
	.w3(32'h3b1dc970),
	.w4(32'hbb907d2b),
	.w5(32'hba33e3f4),
	.w6(32'hbb83367c),
	.w7(32'hbbcc8413),
	.w8(32'hbb25fe1b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19a4b2),
	.w1(32'h3ba5a5f1),
	.w2(32'h3b2d24be),
	.w3(32'hbaaddad5),
	.w4(32'hba1f09e1),
	.w5(32'hbaa91f0f),
	.w6(32'h3af9500c),
	.w7(32'hb6f55c62),
	.w8(32'h3bfe9102),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c258),
	.w1(32'h3b9f238c),
	.w2(32'hbbe4c841),
	.w3(32'h3ac5d3de),
	.w4(32'hbb6fb7a0),
	.w5(32'h3b4a6647),
	.w6(32'h3b4aad8d),
	.w7(32'h3a9e6c32),
	.w8(32'h3b8568a8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd037a),
	.w1(32'h3c08ee7f),
	.w2(32'h3c196167),
	.w3(32'h3a7c0220),
	.w4(32'h3b5e64b8),
	.w5(32'h3b96fdde),
	.w6(32'h3c2f6d17),
	.w7(32'h3c1d5ab8),
	.w8(32'h39eafd5f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5052d),
	.w1(32'h3be64a59),
	.w2(32'h3c0be466),
	.w3(32'h3bea4bc2),
	.w4(32'h3c2c674c),
	.w5(32'h3c960f70),
	.w6(32'hbb318b4b),
	.w7(32'h3b3d4016),
	.w8(32'h3bfb28a3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b870e91),
	.w1(32'h3c53e983),
	.w2(32'h3c212642),
	.w3(32'h3c947124),
	.w4(32'h3c10c694),
	.w5(32'h3c153482),
	.w6(32'h3b856e3b),
	.w7(32'h3ba0d594),
	.w8(32'h3b83fdae),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8d882),
	.w1(32'h3b338a93),
	.w2(32'h3a73617a),
	.w3(32'h3b5e7bfc),
	.w4(32'h399a65ce),
	.w5(32'h3922306b),
	.w6(32'h3bb6c7b3),
	.w7(32'h3a97780f),
	.w8(32'h3ade8677),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f10d4),
	.w1(32'h3c1deb07),
	.w2(32'h3c4ce438),
	.w3(32'h3c11d776),
	.w4(32'h3b88b98d),
	.w5(32'h3abfa3d8),
	.w6(32'h3c5f7c0e),
	.w7(32'h3c043b4c),
	.w8(32'h3b0c8428),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b834957),
	.w1(32'h3bb1082f),
	.w2(32'h3bae4e21),
	.w3(32'hbb61c465),
	.w4(32'hbb2f9efc),
	.w5(32'hbb8da207),
	.w6(32'hbb4fe54e),
	.w7(32'hbb17a611),
	.w8(32'h3bbfae18),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb734c7),
	.w1(32'hbb7dba39),
	.w2(32'hbaeb12ec),
	.w3(32'h3b315dc8),
	.w4(32'hbab80fbc),
	.w5(32'h3ad6c572),
	.w6(32'h3c0208a6),
	.w7(32'h3ba53c7d),
	.w8(32'h3bc8c80b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33b0b5),
	.w1(32'h3a0a2655),
	.w2(32'h3bba9442),
	.w3(32'h3b740c61),
	.w4(32'hbbee2da1),
	.w5(32'h3aa1b765),
	.w6(32'h3b779552),
	.w7(32'hb9b27d89),
	.w8(32'h3b801b6a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a64c),
	.w1(32'h3b13c89a),
	.w2(32'h3b436c0f),
	.w3(32'h3b63e1b3),
	.w4(32'h3b687822),
	.w5(32'hb9cb0dfc),
	.w6(32'hbb2bb323),
	.w7(32'h3b7c4398),
	.w8(32'hbbb51094),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296566),
	.w1(32'hbb4a4d22),
	.w2(32'hbb4dd799),
	.w3(32'hbb845cb0),
	.w4(32'hbc1bd5a6),
	.w5(32'hbb450f0c),
	.w6(32'hbba08645),
	.w7(32'hbbccce46),
	.w8(32'h3b3049cb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c070a27),
	.w1(32'h3bac2e66),
	.w2(32'h3bb2d065),
	.w3(32'h3c01a6f6),
	.w4(32'h3accec60),
	.w5(32'hbb89a29c),
	.w6(32'h3bdd300e),
	.w7(32'h3bacaf0c),
	.w8(32'h3994fad9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3c26d),
	.w1(32'h3ab9eceb),
	.w2(32'hba80beb7),
	.w3(32'hbb588d43),
	.w4(32'hbb650ed7),
	.w5(32'hba05d19e),
	.w6(32'h3b9814fb),
	.w7(32'h3976df51),
	.w8(32'h39638949),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c9655),
	.w1(32'h3ad97d06),
	.w2(32'h3ac22a9e),
	.w3(32'h3c118376),
	.w4(32'h3a59b655),
	.w5(32'h3aaa01e9),
	.w6(32'h3b893810),
	.w7(32'hbb87ae01),
	.w8(32'h3b369e0a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ddf01),
	.w1(32'h39cadf26),
	.w2(32'h3a91aad7),
	.w3(32'h3b21eb85),
	.w4(32'hba84beff),
	.w5(32'h3c083961),
	.w6(32'h3b8368c9),
	.w7(32'h3b2fbc97),
	.w8(32'h3bc2bc7e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba089b17),
	.w1(32'h3b0da8fe),
	.w2(32'h3aa3cfbb),
	.w3(32'h3b9390c5),
	.w4(32'h3a542911),
	.w5(32'h3a8d1f04),
	.w6(32'h3bab1652),
	.w7(32'h3b448dc9),
	.w8(32'h3ba2ac2d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6235d8),
	.w1(32'h3c1355b1),
	.w2(32'h3b93568c),
	.w3(32'h3b5568c9),
	.w4(32'h3b635965),
	.w5(32'h3a208179),
	.w6(32'h3b3edd2f),
	.w7(32'h3b80d1ae),
	.w8(32'h3a5365bd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967706),
	.w1(32'h3afbbbab),
	.w2(32'h3b77ad50),
	.w3(32'h3aae06ea),
	.w4(32'h3ab19b61),
	.w5(32'hba8532a9),
	.w6(32'h3b9e90a6),
	.w7(32'h3a841f4b),
	.w8(32'h3b120876),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab5f0d),
	.w1(32'hb899efe7),
	.w2(32'hba88628c),
	.w3(32'h3c63360a),
	.w4(32'h3b4620ea),
	.w5(32'h3bf0334e),
	.w6(32'h3c7e4736),
	.w7(32'hb9cdbbf0),
	.w8(32'h3c0fcbf7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d895d),
	.w1(32'h3beb0be4),
	.w2(32'h3c08d80f),
	.w3(32'h3c42712f),
	.w4(32'h38c8f3cf),
	.w5(32'hbb669bf3),
	.w6(32'h3abaa04a),
	.w7(32'h3acf4b75),
	.w8(32'h3be96ef7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c804f4d),
	.w1(32'h3bcb1f39),
	.w2(32'h3be1bdd2),
	.w3(32'h3b91843d),
	.w4(32'hbbdf8bd7),
	.w5(32'hbb2f16f2),
	.w6(32'h3c9e1647),
	.w7(32'h3b76857f),
	.w8(32'hbc5f6781),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086174),
	.w1(32'h3b01b122),
	.w2(32'h3b12b29d),
	.w3(32'hba31d179),
	.w4(32'h3b545dcc),
	.w5(32'h3ae2240b),
	.w6(32'hbc29beb0),
	.w7(32'hbbd98624),
	.w8(32'h3b2f04f9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c0856),
	.w1(32'hbbae15d2),
	.w2(32'hbb45247a),
	.w3(32'hbad5f3ea),
	.w4(32'hba87c5a1),
	.w5(32'h3ab65f3c),
	.w6(32'h3a3a1e1e),
	.w7(32'hb99c5f5f),
	.w8(32'h3b832c1f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebc9f6),
	.w1(32'h3c10c86c),
	.w2(32'h3c28cbeb),
	.w3(32'h3b09d458),
	.w4(32'h3a671af4),
	.w5(32'hbbce79ef),
	.w6(32'h3c16841e),
	.w7(32'h3b5e0d85),
	.w8(32'h37bc41bb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bb843),
	.w1(32'h3ad866c1),
	.w2(32'h3b130bb6),
	.w3(32'hbb3dd016),
	.w4(32'hbb9dcb10),
	.w5(32'hb9555908),
	.w6(32'h38a156c8),
	.w7(32'hbbbcf4e8),
	.w8(32'hb9c86aab),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc92dba),
	.w1(32'h3b08c9cf),
	.w2(32'h3af75331),
	.w3(32'h3c20012d),
	.w4(32'h3a791626),
	.w5(32'h3bc2260d),
	.w6(32'h3bacb683),
	.w7(32'h3ba8e101),
	.w8(32'h3ad76324),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9620e4),
	.w1(32'h3beff328),
	.w2(32'h3b9491dd),
	.w3(32'h3bf4b1a4),
	.w4(32'h3c18c235),
	.w5(32'hbba0a60a),
	.w6(32'hbb26845f),
	.w7(32'h3be46bcb),
	.w8(32'h38caa7ec),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69973f),
	.w1(32'hbab2a43e),
	.w2(32'hbb1498b7),
	.w3(32'hba650605),
	.w4(32'hbb022231),
	.w5(32'h39a013e7),
	.w6(32'h3b8b14f2),
	.w7(32'h3bb622be),
	.w8(32'hb9a94867),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32b75d),
	.w1(32'h3bd297e2),
	.w2(32'h3bad81c5),
	.w3(32'h3bebc2e2),
	.w4(32'h3a112202),
	.w5(32'h3ad5cac4),
	.w6(32'h3b6a9d8c),
	.w7(32'h3b1ac01a),
	.w8(32'h3b9ae42d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6e900),
	.w1(32'h39288764),
	.w2(32'hbb1e2ea9),
	.w3(32'h3a82f796),
	.w4(32'hba2c4f6c),
	.w5(32'hbacc6370),
	.w6(32'hba9e1905),
	.w7(32'hbabcc8d2),
	.w8(32'h3b5126ae),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e7716),
	.w1(32'h3b333339),
	.w2(32'h3b13babe),
	.w3(32'hbb2b14dd),
	.w4(32'hbba60128),
	.w5(32'h3bc75102),
	.w6(32'h3ae4bad7),
	.w7(32'hb9e86ba7),
	.w8(32'h3c10cbd6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b260682),
	.w1(32'h3aa5b77f),
	.w2(32'h3a84bc2c),
	.w3(32'h3ba73b8d),
	.w4(32'h3a4fcf83),
	.w5(32'h3b96f71d),
	.w6(32'h3ba3c85e),
	.w7(32'hbb234357),
	.w8(32'hb9f231f9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42f00a),
	.w1(32'h3aea8f1e),
	.w2(32'hbb555fce),
	.w3(32'h3c5a5049),
	.w4(32'h3b4ef58a),
	.w5(32'hbc012f5f),
	.w6(32'h3bbf29dd),
	.w7(32'h3a6708ed),
	.w8(32'hbc10dfd7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb87f5e),
	.w1(32'h3adabb48),
	.w2(32'h3beb1133),
	.w3(32'h3be5642d),
	.w4(32'hbb2a1e69),
	.w5(32'hbc61a552),
	.w6(32'h3c493da2),
	.w7(32'h3bc8ed41),
	.w8(32'hbc76aecb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64cb7f),
	.w1(32'hbbf9fe79),
	.w2(32'hbb872e28),
	.w3(32'h3aea391c),
	.w4(32'hbc521db9),
	.w5(32'hbc80e51d),
	.w6(32'hb9ca1e55),
	.w7(32'hbc210435),
	.w8(32'hbbf6234e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f71b8),
	.w1(32'h3aa4fc1e),
	.w2(32'h3acfc687),
	.w3(32'hbc0c72d0),
	.w4(32'hbc08dff7),
	.w5(32'h3b10a748),
	.w6(32'h3a206684),
	.w7(32'hbaf56172),
	.w8(32'h3b8709ed),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e1c42),
	.w1(32'hb98b5013),
	.w2(32'hb994d913),
	.w3(32'h3b944712),
	.w4(32'h3b5f44c8),
	.w5(32'hbaab7969),
	.w6(32'h3bf02202),
	.w7(32'h3a6997e4),
	.w8(32'hbc4b92d6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a724569),
	.w1(32'h3b1eb094),
	.w2(32'h3aad5aa1),
	.w3(32'hbb61456d),
	.w4(32'hb8e5e55d),
	.w5(32'hbb8f8f10),
	.w6(32'hbc50058b),
	.w7(32'hbc2f2d25),
	.w8(32'hbb51a9fc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc34a8f),
	.w1(32'h3b33a1a7),
	.w2(32'hbb9e26a9),
	.w3(32'h3bea854a),
	.w4(32'h3ac434cf),
	.w5(32'hbbbd326b),
	.w6(32'h3a988fcc),
	.w7(32'hbb86491e),
	.w8(32'h3b8ea1f2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49b80a),
	.w1(32'h3a8a12b0),
	.w2(32'h3ae105da),
	.w3(32'h3c9266c7),
	.w4(32'h3b3fe6e1),
	.w5(32'hbada404a),
	.w6(32'h3cf59488),
	.w7(32'h3c2c266d),
	.w8(32'hbbce37e4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b506fb7),
	.w1(32'hbbb9f868),
	.w2(32'hbbc5a507),
	.w3(32'h3b3351dd),
	.w4(32'hbbb4cda3),
	.w5(32'h3c474ce5),
	.w6(32'hbbafae12),
	.w7(32'hbc61195a),
	.w8(32'hbbb848c2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2cac1),
	.w1(32'h3c1d0ee1),
	.w2(32'h3c224e77),
	.w3(32'h3cae527b),
	.w4(32'h3bafe2d0),
	.w5(32'h3ab87812),
	.w6(32'hbaadeab1),
	.w7(32'hbc8538aa),
	.w8(32'h3ac2acf4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c115d),
	.w1(32'h3b323cc5),
	.w2(32'h3b00750d),
	.w3(32'h3c1222e7),
	.w4(32'hba65206d),
	.w5(32'hbbc6a7b7),
	.w6(32'h3c14abac),
	.w7(32'hba9e9a7c),
	.w8(32'h3b20fc15),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21dcda),
	.w1(32'h3ba357da),
	.w2(32'h3bbe6987),
	.w3(32'hbaed89d2),
	.w4(32'h39eb9873),
	.w5(32'h3b8c2ffc),
	.w6(32'h3bd3eb10),
	.w7(32'h38f71cc5),
	.w8(32'hbbe42c1b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398efa2d),
	.w1(32'h3b312ac4),
	.w2(32'h3b9ed78e),
	.w3(32'hbc12002e),
	.w4(32'hbc060a54),
	.w5(32'hba0a0dac),
	.w6(32'hbc848069),
	.w7(32'hbb7c997e),
	.w8(32'hbb06ec7a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b549b3e),
	.w1(32'h3b6ce83a),
	.w2(32'h3b7011da),
	.w3(32'hb94203cc),
	.w4(32'h3b1941c6),
	.w5(32'hb92ea980),
	.w6(32'hbb54a08b),
	.w7(32'h3ae68bf9),
	.w8(32'h3bcc7b80),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821350),
	.w1(32'h3a980b37),
	.w2(32'hbb1b4552),
	.w3(32'h395f8ef1),
	.w4(32'h3a8f397f),
	.w5(32'hba35ea63),
	.w6(32'h3b90a6a8),
	.w7(32'h3b16f539),
	.w8(32'h3b37754b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dda27),
	.w1(32'h39f67f9f),
	.w2(32'h39878dc3),
	.w3(32'h3bd723cc),
	.w4(32'h3a7efccc),
	.w5(32'h3a4dc1c6),
	.w6(32'h3c047173),
	.w7(32'h3a1f51d8),
	.w8(32'hbb2e248c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc46b),
	.w1(32'h3b3bf77a),
	.w2(32'h3b9062bb),
	.w3(32'h3b22e71a),
	.w4(32'hbb303e9e),
	.w5(32'h3a81dfaa),
	.w6(32'hbb50ed67),
	.w7(32'hbba7fdda),
	.w8(32'hba6c142c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7961d8),
	.w1(32'h3bee5189),
	.w2(32'h3c3b915c),
	.w3(32'h3c365525),
	.w4(32'h3ba9e371),
	.w5(32'h3bb12379),
	.w6(32'h3bae6ec8),
	.w7(32'hb9a473a1),
	.w8(32'h3af41d6e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a78c),
	.w1(32'h3a406d01),
	.w2(32'hbafeba77),
	.w3(32'h3b8fb14f),
	.w4(32'hbaebd9b7),
	.w5(32'hbbcb39a3),
	.w6(32'h3bb60686),
	.w7(32'hb84043fb),
	.w8(32'hbb1a28b4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc177),
	.w1(32'hbb08e6a3),
	.w2(32'hbac2b401),
	.w3(32'hbb927ed4),
	.w4(32'h3a61975f),
	.w5(32'h3b9a6fb9),
	.w6(32'hbbd7623f),
	.w7(32'hbaeab017),
	.w8(32'h3b874269),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b501569),
	.w1(32'h3a5feadc),
	.w2(32'h3a51426f),
	.w3(32'h3bac52fe),
	.w4(32'h3bca9890),
	.w5(32'hbb21c5ff),
	.w6(32'h3c3380c2),
	.w7(32'h3bb53564),
	.w8(32'hbb5d6215),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c7d83),
	.w1(32'h3a9810d3),
	.w2(32'h3b643861),
	.w3(32'hbb2718c4),
	.w4(32'hbb35b736),
	.w5(32'hba8adad0),
	.w6(32'hbb753fe0),
	.w7(32'hbb7cfa6f),
	.w8(32'hba97e3ba),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc48a5),
	.w1(32'h394f1d68),
	.w2(32'hba17c1f2),
	.w3(32'hb8859fd2),
	.w4(32'h3ac4dad3),
	.w5(32'hbb1ab215),
	.w6(32'hbb73b68a),
	.w7(32'hbb059631),
	.w8(32'h3938d8e1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3b8c0),
	.w1(32'hbb5bd700),
	.w2(32'h3ae24c2b),
	.w3(32'hba42ada8),
	.w4(32'hbb2eb3ec),
	.w5(32'hb9d44a38),
	.w6(32'h3b73b236),
	.w7(32'h3ab1c384),
	.w8(32'hbb9b2ba0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbab994),
	.w1(32'hb732874e),
	.w2(32'h3b27ff6f),
	.w3(32'h3ba23340),
	.w4(32'h39c8dc81),
	.w5(32'h3bfb2765),
	.w6(32'hbb36b4ad),
	.w7(32'hbb4a62e6),
	.w8(32'hbb80f1e9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80af34),
	.w1(32'h3c465622),
	.w2(32'h3c30d56b),
	.w3(32'h3c498cd9),
	.w4(32'h3bea1cf2),
	.w5(32'hbbbce059),
	.w6(32'hbb74ea9b),
	.w7(32'hbaf8b08a),
	.w8(32'h3bb595ff),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bfaa4),
	.w1(32'h3b6a1536),
	.w2(32'hbb521ee6),
	.w3(32'hbbac035a),
	.w4(32'hbbc8dde0),
	.w5(32'h3a75c8af),
	.w6(32'hb91d2e8c),
	.w7(32'h3970dee2),
	.w8(32'h3ae7b076),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2577b2),
	.w1(32'hbb5ea3f3),
	.w2(32'hbab87eb1),
	.w3(32'hbafc57d9),
	.w4(32'hba9a37d2),
	.w5(32'h37354fb7),
	.w6(32'hbab143a4),
	.w7(32'h3787b391),
	.w8(32'hbb22003d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9462e16),
	.w1(32'hba72c3b6),
	.w2(32'h3ac60a49),
	.w3(32'hb9ce4e36),
	.w4(32'hb9ff0e9e),
	.w5(32'hbbb03e57),
	.w6(32'hbbb77d0f),
	.w7(32'hb9594507),
	.w8(32'hba4fdf1e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990ff4),
	.w1(32'h3acc7ad1),
	.w2(32'hb8d5ad07),
	.w3(32'hbbc36097),
	.w4(32'hbbe10c4a),
	.w5(32'h3c031b83),
	.w6(32'hbb15a906),
	.w7(32'hba03e7d7),
	.w8(32'hbb685de0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba51de9),
	.w1(32'h3ba11cd4),
	.w2(32'h3bb09d4a),
	.w3(32'h3c2ce6c7),
	.w4(32'hbb64e8d2),
	.w5(32'hbba4263d),
	.w6(32'hbb85c0bd),
	.w7(32'hbb3c0c05),
	.w8(32'h3b82ed58),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b2a42),
	.w1(32'h3b226516),
	.w2(32'h3915bf94),
	.w3(32'h3bc1fa2a),
	.w4(32'hbbc8a4b3),
	.w5(32'hbaab5c30),
	.w6(32'h3c7d659d),
	.w7(32'hbb98d8cf),
	.w8(32'hbbd4f986),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5f56),
	.w1(32'h3b090ffb),
	.w2(32'h3b401273),
	.w3(32'h3bf4ace1),
	.w4(32'hbba7156f),
	.w5(32'hba996382),
	.w6(32'h3c05af87),
	.w7(32'hbb1c56da),
	.w8(32'h3b96c882),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74916a),
	.w1(32'h3ae13907),
	.w2(32'h3b2ed0ab),
	.w3(32'h3c8d6cd4),
	.w4(32'hbb3d33c9),
	.w5(32'hbbb3d893),
	.w6(32'h3cd4d157),
	.w7(32'h394810e5),
	.w8(32'hbb480258),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d89b1f),
	.w1(32'hba6e1ff9),
	.w2(32'hbad58bd0),
	.w3(32'h399cd284),
	.w4(32'hba9200cf),
	.w5(32'h3ad69940),
	.w6(32'h3936f6e9),
	.w7(32'hb9c7b1fd),
	.w8(32'h3b5ab6e4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b1c87),
	.w1(32'h3afba932),
	.w2(32'h3be91367),
	.w3(32'hbaf6a58d),
	.w4(32'h39dbd3d1),
	.w5(32'hbb702516),
	.w6(32'hbb2f81e1),
	.w7(32'h3b3f87d4),
	.w8(32'hbc343625),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25667c),
	.w1(32'hbba9b096),
	.w2(32'h3b2a58e7),
	.w3(32'hbc3f07ed),
	.w4(32'hbc012ae9),
	.w5(32'hbb3ea092),
	.w6(32'hbc9766c1),
	.w7(32'hbc570e45),
	.w8(32'h3b216785),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf834),
	.w1(32'h3b80dd6d),
	.w2(32'hbade5f59),
	.w3(32'hbaec7d2f),
	.w4(32'h3a23b312),
	.w5(32'hbb26678f),
	.w6(32'hb98a1c3c),
	.w7(32'hbb726969),
	.w8(32'hbb483985),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a0ee9),
	.w1(32'h38b3b36d),
	.w2(32'h3b73c416),
	.w3(32'hbbb5b524),
	.w4(32'hbb94564b),
	.w5(32'hbb95a7c9),
	.w6(32'hbb8479f9),
	.w7(32'hb89ef4e5),
	.w8(32'h3ae5299d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18352),
	.w1(32'h3870e9e9),
	.w2(32'hba6badd5),
	.w3(32'hbb945fb3),
	.w4(32'hbb34e095),
	.w5(32'h3aab4f27),
	.w6(32'hba5bb627),
	.w7(32'hbab99f5e),
	.w8(32'hbab62e09),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf15262),
	.w1(32'h3ac166e1),
	.w2(32'h3aa45334),
	.w3(32'h3bfbb0bd),
	.w4(32'h3a7a2117),
	.w5(32'hba8e4979),
	.w6(32'h3c0dfec2),
	.w7(32'h3b890085),
	.w8(32'hbaa62df6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61af42),
	.w1(32'hba917edf),
	.w2(32'hbb76149b),
	.w3(32'h3ab5ec23),
	.w4(32'hbbc4258e),
	.w5(32'hb95d3961),
	.w6(32'h3a62dbf8),
	.w7(32'hbbc26615),
	.w8(32'hba189d86),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd1e4),
	.w1(32'h39cfc69f),
	.w2(32'h3b72c82d),
	.w3(32'h3a8a8c4e),
	.w4(32'hbba7bec2),
	.w5(32'h3bb3756b),
	.w6(32'h3abbbd74),
	.w7(32'h3a74959e),
	.w8(32'h3b31be67),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2b140),
	.w1(32'h3bd3674e),
	.w2(32'h3bba4b10),
	.w3(32'h3ab63ee2),
	.w4(32'hba3ae9e0),
	.w5(32'hba3f58aa),
	.w6(32'h3b70646d),
	.w7(32'hb5f0700e),
	.w8(32'h3c0b4275),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5a62f),
	.w1(32'h3a6a37db),
	.w2(32'hb9883799),
	.w3(32'h3bb47b80),
	.w4(32'hbb08a9f0),
	.w5(32'hba9f712f),
	.w6(32'h3c88e8c0),
	.w7(32'h3c25353c),
	.w8(32'h39b79cd2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34b4e),
	.w1(32'h3b3216ef),
	.w2(32'h3b2f11ae),
	.w3(32'hb9da5859),
	.w4(32'h3a88fa6f),
	.w5(32'h3b83f1cc),
	.w6(32'hbba9c1af),
	.w7(32'hbb1e0b50),
	.w8(32'h3a4c0288),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bd306),
	.w1(32'h3bb74ab2),
	.w2(32'h3c0a3752),
	.w3(32'hba8d0b55),
	.w4(32'h3af1fa6e),
	.w5(32'hbbdf9904),
	.w6(32'hba2dd0b1),
	.w7(32'h3bc8cb3a),
	.w8(32'hbb91e9ff),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb282),
	.w1(32'hbb22ec62),
	.w2(32'hbb2508ec),
	.w3(32'hbbfdf6f8),
	.w4(32'hbc09a475),
	.w5(32'hba620e94),
	.w6(32'hbac61b65),
	.w7(32'hbb86571b),
	.w8(32'h3a2376cb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e94cf2),
	.w1(32'hbb15c640),
	.w2(32'h3a2c0bc2),
	.w3(32'hba866c15),
	.w4(32'hba975bb6),
	.w5(32'hbaec2da3),
	.w6(32'hbad49a1f),
	.w7(32'hba4f640a),
	.w8(32'hbc29cfa6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c194eb6),
	.w1(32'h3c00e7e6),
	.w2(32'h3c3f94df),
	.w3(32'hbc049571),
	.w4(32'hbbae35ff),
	.w5(32'hbabac49b),
	.w6(32'hbc9bf026),
	.w7(32'hbc4327b6),
	.w8(32'hbad27467),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16e17c),
	.w1(32'h3bd12d47),
	.w2(32'hbaf8902f),
	.w3(32'h3c467d5b),
	.w4(32'hb8c89fac),
	.w5(32'hbbd6dae5),
	.w6(32'h3be8536d),
	.w7(32'hbaebdb1d),
	.w8(32'hbb0bb8e2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fdfaa),
	.w1(32'h3b6b3a40),
	.w2(32'h3ad7e33a),
	.w3(32'hbb81f6b2),
	.w4(32'hbafbe383),
	.w5(32'h3b0fc0da),
	.w6(32'hb9cd384b),
	.w7(32'h3a86356c),
	.w8(32'h3b12dc14),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cd01b),
	.w1(32'h3bcc5260),
	.w2(32'h3bd17a39),
	.w3(32'h3c31b338),
	.w4(32'h3b8624f6),
	.w5(32'hbabdae11),
	.w6(32'h3c31f5df),
	.w7(32'h3b6dbbfd),
	.w8(32'hbb8921d7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d9dd),
	.w1(32'h3bd1c475),
	.w2(32'h3bce78f9),
	.w3(32'h3bd17972),
	.w4(32'h3bf36f6e),
	.w5(32'h3c0a27e9),
	.w6(32'h3b52e1f6),
	.w7(32'h3c1c249c),
	.w8(32'h3c2718e8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a0f5d),
	.w1(32'h3985c1f6),
	.w2(32'h38180613),
	.w3(32'h3bd71bc3),
	.w4(32'h379b47fc),
	.w5(32'hba6edcb3),
	.w6(32'h3bab6fe2),
	.w7(32'hbaf91997),
	.w8(32'hb96c0b24),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03b929),
	.w1(32'h3bddb557),
	.w2(32'h3b005941),
	.w3(32'h3ba49467),
	.w4(32'h3bb744a3),
	.w5(32'hbb3bd249),
	.w6(32'h3bcf031a),
	.w7(32'h3b9b1dbe),
	.w8(32'h3b3f0fb0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d15fc),
	.w1(32'hb9cf096a),
	.w2(32'hbbcec22d),
	.w3(32'h3b64ff8e),
	.w4(32'hbb39babe),
	.w5(32'hbbc10d5b),
	.w6(32'h3b84b593),
	.w7(32'h3ad21472),
	.w8(32'hb9802976),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f43d3),
	.w1(32'h394f09e2),
	.w2(32'hbbaaeaad),
	.w3(32'h3be98abd),
	.w4(32'hbb57534e),
	.w5(32'h3a555fab),
	.w6(32'h3c3e1b3d),
	.w7(32'h3a90f320),
	.w8(32'hbaf9e8d0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2731c1),
	.w1(32'h3c0a6003),
	.w2(32'h3c6b1b70),
	.w3(32'h3aac5977),
	.w4(32'h3b3fcbf8),
	.w5(32'h3a1e2df5),
	.w6(32'hbad0cc24),
	.w7(32'h3b0d58de),
	.w8(32'hbad76ef8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b73e8),
	.w1(32'hbb8b6030),
	.w2(32'hbaad5e9b),
	.w3(32'h3c237a45),
	.w4(32'h3adcc492),
	.w5(32'hbc2f19da),
	.w6(32'h3bcc70a6),
	.w7(32'hb8dbe396),
	.w8(32'hbbbab4ef),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa40d21),
	.w1(32'hbb23121f),
	.w2(32'hbb468f26),
	.w3(32'hbc18c5c2),
	.w4(32'hbbafbacb),
	.w5(32'hbb82a080),
	.w6(32'hbaa582e6),
	.w7(32'hbb2126b3),
	.w8(32'hbbdd9931),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43b52f),
	.w1(32'h3b7bef3c),
	.w2(32'h3ba6a7d2),
	.w3(32'h3bf24f6e),
	.w4(32'h3ad86423),
	.w5(32'hb9dcc729),
	.w6(32'h3be894f9),
	.w7(32'h3a9a5a6e),
	.w8(32'h3ab9ae56),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6602),
	.w1(32'hbb0a5b7d),
	.w2(32'hb9651477),
	.w3(32'h3a8c918b),
	.w4(32'hbb2ad2b4),
	.w5(32'hbb8b3306),
	.w6(32'h3b01f114),
	.w7(32'hba84eb4e),
	.w8(32'h381f6e11),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b18ea),
	.w1(32'h3b67da48),
	.w2(32'h3b5908cf),
	.w3(32'h3b8a7542),
	.w4(32'hb97839b0),
	.w5(32'hbbb26c55),
	.w6(32'h3b91f4ce),
	.w7(32'hbb08ecfc),
	.w8(32'hbc01378a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b026f),
	.w1(32'h3aa396ab),
	.w2(32'hbc02af10),
	.w3(32'h3c2453ac),
	.w4(32'hbb7b2d67),
	.w5(32'hbc45cbcb),
	.w6(32'h3c04570a),
	.w7(32'h3ab21ad4),
	.w8(32'hbbde895e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d27e),
	.w1(32'h3a9d12fc),
	.w2(32'h3b7f41ac),
	.w3(32'h3c0088ef),
	.w4(32'hba64bc5e),
	.w5(32'h3a9a6bc9),
	.w6(32'h3bbf4e47),
	.w7(32'hba2355ea),
	.w8(32'h3a5cf44f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b2069),
	.w1(32'h3ac20351),
	.w2(32'hbb26252c),
	.w3(32'h3b6960e2),
	.w4(32'h3b31e0c2),
	.w5(32'hbb5ca6c3),
	.w6(32'h3b20dd4b),
	.w7(32'h3a443594),
	.w8(32'hba80ac52),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a381ef9),
	.w1(32'h3a284cd5),
	.w2(32'h3a5904bc),
	.w3(32'h385db413),
	.w4(32'h3a25fa95),
	.w5(32'hb9857371),
	.w6(32'h39cc32cc),
	.w7(32'h3ac6acf9),
	.w8(32'h3a556350),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bfa3a),
	.w1(32'h3c0f4acb),
	.w2(32'h3ab5be9d),
	.w3(32'h3b0aa1f3),
	.w4(32'h3b406682),
	.w5(32'hbbaa3b5e),
	.w6(32'h3a5864a1),
	.w7(32'h3affa3dc),
	.w8(32'hbbeb8a0f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5da5),
	.w1(32'h3a4715e8),
	.w2(32'hbb367f7d),
	.w3(32'h3ae81f91),
	.w4(32'h3b056b20),
	.w5(32'hbafa81b2),
	.w6(32'h3b1c5a53),
	.w7(32'h3b8e9b3b),
	.w8(32'hbb023dce),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370a841d),
	.w1(32'hb7c38dd6),
	.w2(32'h395c0374),
	.w3(32'hb90c0706),
	.w4(32'hb95d2947),
	.w5(32'hb8aaae6a),
	.w6(32'hb88e033e),
	.w7(32'hb90c3c52),
	.w8(32'h379f6ea5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7c36c),
	.w1(32'h3a7a68ee),
	.w2(32'h3aa46251),
	.w3(32'h3a2f871e),
	.w4(32'hb8da285e),
	.w5(32'hba32ef0b),
	.w6(32'h3aee10e2),
	.w7(32'h3a3829a9),
	.w8(32'hba09fe78),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9981f),
	.w1(32'h3ad75baf),
	.w2(32'h3b3e7be8),
	.w3(32'h3b90161d),
	.w4(32'h3b1de1a9),
	.w5(32'h3b87797f),
	.w6(32'h3ba739e1),
	.w7(32'h3b7f771a),
	.w8(32'h3b8f47ea),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7fc5e),
	.w1(32'h39281f36),
	.w2(32'h3aec85c6),
	.w3(32'h3bd721c4),
	.w4(32'hb7e31565),
	.w5(32'h39b4a400),
	.w6(32'h3baf082f),
	.w7(32'h38fee6af),
	.w8(32'h3aa1a499),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2949b),
	.w1(32'hb8bcd94d),
	.w2(32'hba823bb9),
	.w3(32'h392462d9),
	.w4(32'hbae26d09),
	.w5(32'hbaeb34b5),
	.w6(32'h3b0aaa7f),
	.w7(32'hbaa27bd5),
	.w8(32'hba9483f3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac4c21),
	.w1(32'h3a03f71b),
	.w2(32'h39ea717d),
	.w3(32'h3b2651f8),
	.w4(32'hbab40fbb),
	.w5(32'hba86763f),
	.w6(32'h3ae24895),
	.w7(32'hba3598e8),
	.w8(32'h39b61255),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac66e8),
	.w1(32'hba95ce80),
	.w2(32'hbb0813e0),
	.w3(32'h3b6ba5b3),
	.w4(32'hbb89ef82),
	.w5(32'hbb9c254f),
	.w6(32'h3bb88272),
	.w7(32'hbb5081e0),
	.w8(32'hbbaa54b6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebd532),
	.w1(32'h3ac61f86),
	.w2(32'h3b73ff20),
	.w3(32'h3b982aae),
	.w4(32'h3a3c530d),
	.w5(32'hba39ec16),
	.w6(32'h3b8cd550),
	.w7(32'h3ab92191),
	.w8(32'h3a49f186),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb844b5),
	.w1(32'h39b3097a),
	.w2(32'h390c49ec),
	.w3(32'h3ba3be7f),
	.w4(32'hb984e806),
	.w5(32'hb92fab73),
	.w6(32'h3b86e94f),
	.w7(32'hb9822795),
	.w8(32'h39c3d0e3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374e8be6),
	.w1(32'h38723587),
	.w2(32'h3876a785),
	.w3(32'h382aa849),
	.w4(32'h3874c464),
	.w5(32'h369a7496),
	.w6(32'h3831d7a3),
	.w7(32'h38e70bb8),
	.w8(32'h381f999d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25bc4c),
	.w1(32'h39bb79df),
	.w2(32'h388e9381),
	.w3(32'h39a1e674),
	.w4(32'hb72baba8),
	.w5(32'hb99b6ca0),
	.w6(32'h394c58a3),
	.w7(32'hb91bd2d8),
	.w8(32'hb968234c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1f0b1),
	.w1(32'hb914cff2),
	.w2(32'hb7c8bb37),
	.w3(32'h390503cc),
	.w4(32'hb9115eec),
	.w5(32'hb8b4d7ec),
	.w6(32'h391fce9d),
	.w7(32'hb8d4adc4),
	.w8(32'hb8822a64),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f34b8),
	.w1(32'hb978833d),
	.w2(32'h38a7264e),
	.w3(32'hb8989baa),
	.w4(32'h373d671d),
	.w5(32'h39897e43),
	.w6(32'hb918850a),
	.w7(32'h35bbbc29),
	.w8(32'hb88357e9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becacd9),
	.w1(32'hb9a6692b),
	.w2(32'h39925ad6),
	.w3(32'h3bc40fac),
	.w4(32'hbad053c5),
	.w5(32'hb9d7804c),
	.w6(32'h3ba4965c),
	.w7(32'hba8d2acb),
	.w8(32'h39a8cd87),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a534987),
	.w1(32'h39c362e5),
	.w2(32'h399807ae),
	.w3(32'h39ce5239),
	.w4(32'h390fdd0e),
	.w5(32'h39bba047),
	.w6(32'hb8490a6b),
	.w7(32'hb76a7d3c),
	.w8(32'h3a1cbfbb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c5e1f),
	.w1(32'h39e138fd),
	.w2(32'h3a047ece),
	.w3(32'h3a82b1c4),
	.w4(32'h3a4159c8),
	.w5(32'hba099e4f),
	.w6(32'hba317e52),
	.w7(32'hba157f41),
	.w8(32'hba884425),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06db87),
	.w1(32'h3b2ec9b2),
	.w2(32'h3b641c4a),
	.w3(32'h3ba3e754),
	.w4(32'hbb1288ff),
	.w5(32'hbb05e4ab),
	.w6(32'h3bbfaea9),
	.w7(32'hba2944a2),
	.w8(32'hb99e71ed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93875b8),
	.w1(32'hb86837fb),
	.w2(32'h37d41acb),
	.w3(32'hb916f921),
	.w4(32'hb888b1f4),
	.w5(32'hb8051f7e),
	.w6(32'hb95094f8),
	.w7(32'hb90195c3),
	.w8(32'hb8a2023d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985a825),
	.w1(32'h38585737),
	.w2(32'h39699285),
	.w3(32'hb9518eb3),
	.w4(32'hb8a191b4),
	.w5(32'hb8dbe48b),
	.w6(32'hb959ad36),
	.w7(32'hb6f61acc),
	.w8(32'h38a5f7be),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b23374),
	.w1(32'hb7e1a174),
	.w2(32'hb7a67c73),
	.w3(32'hb88c13d4),
	.w4(32'hb7cf4461),
	.w5(32'hb79e6bba),
	.w6(32'hb84eda5d),
	.w7(32'hb863b56f),
	.w8(32'hb8067684),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c78dab),
	.w1(32'h38f912f3),
	.w2(32'h3a01ede8),
	.w3(32'h389b7e4b),
	.w4(32'hba069ad4),
	.w5(32'hb9860b5c),
	.w6(32'h391008c7),
	.w7(32'hb90ed326),
	.w8(32'h3893f855),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4210a7),
	.w1(32'h3b5fa4a5),
	.w2(32'h3b0c194d),
	.w3(32'h3a826085),
	.w4(32'hba321a64),
	.w5(32'h3ac5e54f),
	.w6(32'h3b0085fc),
	.w7(32'hbae84d6b),
	.w8(32'hba7ae735),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf33b7b),
	.w1(32'h39fec297),
	.w2(32'h3b63bb2a),
	.w3(32'h3bbf828b),
	.w4(32'h3a36bf3d),
	.w5(32'h3ae983bc),
	.w6(32'h3ba6d7c9),
	.w7(32'hb898decf),
	.w8(32'h3b18c6bd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6129),
	.w1(32'h3a207986),
	.w2(32'hb7c24f6d),
	.w3(32'h3971acc2),
	.w4(32'h3a3aab92),
	.w5(32'hba0540d5),
	.w6(32'h3927ffa7),
	.w7(32'h39a99fc9),
	.w8(32'hb93c9ce8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0a7ce),
	.w1(32'h39ba0925),
	.w2(32'h383f5fe6),
	.w3(32'h3b196b43),
	.w4(32'h38f2f466),
	.w5(32'h39847b54),
	.w6(32'h3b28d827),
	.w7(32'h37d26384),
	.w8(32'h36c4d473),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018993),
	.w1(32'h399de27d),
	.w2(32'h3a248112),
	.w3(32'h3ab7a618),
	.w4(32'hba1c87be),
	.w5(32'hb9f6191e),
	.w6(32'h3ab84dd7),
	.w7(32'hb9a928f0),
	.w8(32'hb9ee1cc8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881235),
	.w1(32'h39c5d4a0),
	.w2(32'h39693a45),
	.w3(32'h3b748c73),
	.w4(32'h3a200890),
	.w5(32'hb9bee6e3),
	.w6(32'h3b823b4b),
	.w7(32'h3a591bdf),
	.w8(32'hb9a4efda),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d0a6),
	.w1(32'h3a2d585d),
	.w2(32'h3b0cf0d8),
	.w3(32'h3b1725fb),
	.w4(32'hbb3e4673),
	.w5(32'hbb21f5ad),
	.w6(32'h3b0e90e7),
	.w7(32'hbb135a4c),
	.w8(32'hbb14c977),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce5f33),
	.w1(32'h3981bea8),
	.w2(32'h3b1b0b3e),
	.w3(32'h3b7063f7),
	.w4(32'h3a8b241b),
	.w5(32'hb8fd4986),
	.w6(32'h3b36cb78),
	.w7(32'hbaba51e0),
	.w8(32'h3b313d58),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a313),
	.w1(32'h3a8eb961),
	.w2(32'h3a2575a0),
	.w3(32'h3bad5ed7),
	.w4(32'hb99b8393),
	.w5(32'hba29d719),
	.w6(32'h3ba3cd19),
	.w7(32'h39baa6a3),
	.w8(32'h39df0e7c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc45b4),
	.w1(32'h3ae41f1c),
	.w2(32'h3a6cee40),
	.w3(32'h3b18b110),
	.w4(32'hb9bd0402),
	.w5(32'hbb0b8b6e),
	.w6(32'h3b23b9c0),
	.w7(32'h39d2f12f),
	.w8(32'h38c0bc3a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15b63d),
	.w1(32'hba8226e9),
	.w2(32'h3b112454),
	.w3(32'h3bcaae1d),
	.w4(32'h388dbd79),
	.w5(32'h3b0c4964),
	.w6(32'h3b88c193),
	.w7(32'hbb75f8e4),
	.w8(32'h3b1da853),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcadab0),
	.w1(32'h3b2c4a7d),
	.w2(32'hb9002484),
	.w3(32'h3b80eb6a),
	.w4(32'h38817f87),
	.w5(32'hbb020ff0),
	.w6(32'h3b9359b0),
	.w7(32'hb8837a5e),
	.w8(32'hbad6de7a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc04b4f),
	.w1(32'h3aa771c2),
	.w2(32'h3ad3d085),
	.w3(32'h3b75c183),
	.w4(32'h3b05bc43),
	.w5(32'h3af2eaaf),
	.w6(32'h3b4bd65e),
	.w7(32'h3b174806),
	.w8(32'h3b60e71d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10d8fa),
	.w1(32'h39395e56),
	.w2(32'h399a38d2),
	.w3(32'h3ade4cb1),
	.w4(32'hb9d01283),
	.w5(32'hb9b7f167),
	.w6(32'h3ae2a001),
	.w7(32'h36a86000),
	.w8(32'h37ba58dc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f0a8),
	.w1(32'hbacce0c5),
	.w2(32'h3abe574a),
	.w3(32'h3ba6d93c),
	.w4(32'hbb87bf72),
	.w5(32'h39bc843d),
	.w6(32'h3bbf4d38),
	.w7(32'hbb104aad),
	.w8(32'h3ab7a6e1),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72f2a8),
	.w1(32'h39d2547f),
	.w2(32'hba86de39),
	.w3(32'h3b22a0a4),
	.w4(32'hba1cf215),
	.w5(32'hbab2eea6),
	.w6(32'h3b2372b6),
	.w7(32'h384632c4),
	.w8(32'hbaba04ec),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369d41d1),
	.w1(32'h375fb2ad),
	.w2(32'h370da40c),
	.w3(32'h389e5309),
	.w4(32'h38efb07e),
	.w5(32'h39203faf),
	.w6(32'h3870eb0f),
	.w7(32'h3895bdc8),
	.w8(32'h389ddd72),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2466a),
	.w1(32'h34bc9e6f),
	.w2(32'h3874ccc1),
	.w3(32'h37af5e20),
	.w4(32'h382d79e8),
	.w5(32'h389c8bb2),
	.w6(32'hb7a745e5),
	.w7(32'hb7878a5a),
	.w8(32'hb66b8f10),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fcede),
	.w1(32'h3a196970),
	.w2(32'hba46025f),
	.w3(32'h3b0a1337),
	.w4(32'h3a23f807),
	.w5(32'hbad58773),
	.w6(32'h3abc7dad),
	.w7(32'h3a5f9259),
	.w8(32'hbad90d04),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff546f),
	.w1(32'h3b41faa9),
	.w2(32'h3ae78f01),
	.w3(32'h3b267845),
	.w4(32'hba77b07b),
	.w5(32'h3a881e1f),
	.w6(32'h3b20323e),
	.w7(32'h3aa09e19),
	.w8(32'h39ce796f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be47c),
	.w1(32'h39c2f06f),
	.w2(32'h3b3d6c08),
	.w3(32'h3c0ad419),
	.w4(32'hba7083ec),
	.w5(32'h3a9ae02d),
	.w6(32'h3be88460),
	.w7(32'hbaa653bd),
	.w8(32'h3aed5006),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f3513),
	.w1(32'hb8499503),
	.w2(32'h36c34127),
	.w3(32'hb82c7ea9),
	.w4(32'h37827823),
	.w5(32'h371f886a),
	.w6(32'hb68cd2ef),
	.w7(32'h380b99d4),
	.w8(32'h372a46ca),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f862b),
	.w1(32'h3aabba0e),
	.w2(32'h3b21037d),
	.w3(32'h3be7f271),
	.w4(32'h399a08b6),
	.w5(32'h3af5a396),
	.w6(32'h3bd52f4c),
	.w7(32'h3ac32056),
	.w8(32'h3b32c8c2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba652c8),
	.w1(32'h3a9ad666),
	.w2(32'h3b08112f),
	.w3(32'h3b655f82),
	.w4(32'hb93d37c9),
	.w5(32'hb8f98d80),
	.w6(32'h3b664b0a),
	.w7(32'h38d233b0),
	.w8(32'h37e6ff59),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6ce12),
	.w1(32'h3afefb15),
	.w2(32'h3b853f36),
	.w3(32'h3b0b6b5a),
	.w4(32'h3a78460e),
	.w5(32'hb90f7454),
	.w6(32'h3a9529aa),
	.w7(32'h3a4cc2bf),
	.w8(32'h3b251fae),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829287),
	.w1(32'hbab97337),
	.w2(32'h3b0eafa3),
	.w3(32'h3b163d9d),
	.w4(32'hbba10d49),
	.w5(32'hba73cb0e),
	.w6(32'h3b484d94),
	.w7(32'hbbb6ff47),
	.w8(32'hbab47b54),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b305ff5),
	.w1(32'h3acea080),
	.w2(32'h399134fc),
	.w3(32'h3aab6e67),
	.w4(32'h39bc1bc4),
	.w5(32'hba1e9abe),
	.w6(32'h3abd2731),
	.w7(32'hb81feb91),
	.w8(32'h39392edd),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa00ee3),
	.w1(32'h3a974308),
	.w2(32'h3a90357d),
	.w3(32'h3a20b191),
	.w4(32'h3987b20c),
	.w5(32'h3a5d2817),
	.w6(32'h3a0ba621),
	.w7(32'h3a428eda),
	.w8(32'h39818e80),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7a09e),
	.w1(32'hba532c1a),
	.w2(32'hbabed7c6),
	.w3(32'h3ba4029e),
	.w4(32'hbad645a7),
	.w5(32'hba96543e),
	.w6(32'h3b953105),
	.w7(32'hbab6fb3f),
	.w8(32'h3a06445c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5da24),
	.w1(32'hbabbe3e4),
	.w2(32'hbb1d36f7),
	.w3(32'h3b460a23),
	.w4(32'hbba0a9b0),
	.w5(32'hbb916bb9),
	.w6(32'h3b42dc0d),
	.w7(32'hbb155706),
	.w8(32'hbaac32d3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376a6a),
	.w1(32'hbb0ccdff),
	.w2(32'hbaaf5382),
	.w3(32'h3b0f8df1),
	.w4(32'hbb79eff4),
	.w5(32'hbb5f9a3e),
	.w6(32'h3b70ccc7),
	.w7(32'hbb23a47c),
	.w8(32'hbb0cc82a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7ca13),
	.w1(32'hb7fbe4db),
	.w2(32'hb8420c54),
	.w3(32'h3a3a3608),
	.w4(32'h3a276104),
	.w5(32'h39b9bb72),
	.w6(32'h3a464f39),
	.w7(32'h38e28c0e),
	.w8(32'h39abf1c3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960f113),
	.w1(32'hb81212bf),
	.w2(32'h39067647),
	.w3(32'h380e0e37),
	.w4(32'hb911a5e7),
	.w5(32'hb93298f8),
	.w6(32'h39beb65d),
	.w7(32'h39232785),
	.w8(32'h35ed5e54),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda7399),
	.w1(32'h3abed6bf),
	.w2(32'h3b2e8e98),
	.w3(32'h3b815882),
	.w4(32'hb9850299),
	.w5(32'hb9ea6938),
	.w6(32'h3b8649a2),
	.w7(32'h3834aa39),
	.w8(32'h395a81cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383122ea),
	.w1(32'h397d8f3b),
	.w2(32'h3a1578f3),
	.w3(32'hb951fab5),
	.w4(32'hb79b5a98),
	.w5(32'h39e42b5b),
	.w6(32'hb9b1dbcb),
	.w7(32'hb844703a),
	.w8(32'hb8e1b236),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d99d),
	.w1(32'h39eaa18f),
	.w2(32'hb921864e),
	.w3(32'h3b5bc78b),
	.w4(32'h39a756ef),
	.w5(32'hb9fbdeb7),
	.w6(32'h3b549d7a),
	.w7(32'hb96add32),
	.w8(32'hb962aacd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921569f),
	.w1(32'hb90a3193),
	.w2(32'h361475b1),
	.w3(32'hb9d98ce9),
	.w4(32'hb9bc76f9),
	.w5(32'hb9392079),
	.w6(32'hb860f2ca),
	.w7(32'hb9a1adf8),
	.w8(32'hb92e2a3c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5edb),
	.w1(32'hbaf6b2e2),
	.w2(32'h37baf0c2),
	.w3(32'h3b336b1e),
	.w4(32'hbb30395d),
	.w5(32'hbac3ac23),
	.w6(32'h3baf6a6a),
	.w7(32'hbabe80ef),
	.w8(32'hba560ff4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef1510),
	.w1(32'h396970c9),
	.w2(32'h3980c262),
	.w3(32'hb960dc67),
	.w4(32'h39149972),
	.w5(32'h398edab0),
	.w6(32'hb9453718),
	.w7(32'h38a0ebbb),
	.w8(32'h397ec3ec),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ebf02),
	.w1(32'h38d63b07),
	.w2(32'hb887f5d1),
	.w3(32'h38f687bb),
	.w4(32'hb94e43a1),
	.w5(32'hb8c2e701),
	.w6(32'hb82de0a6),
	.w7(32'hb9e98cb3),
	.w8(32'h388b0500),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a72ee),
	.w1(32'h3b0700a3),
	.w2(32'h3aafee35),
	.w3(32'h3b493ffe),
	.w4(32'h3a464e1d),
	.w5(32'h3aa5e2b6),
	.w6(32'h3b2ebbf7),
	.w7(32'h3a4adda8),
	.w8(32'h3ab9e326),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46fd2a),
	.w1(32'h3b0cdea5),
	.w2(32'h3ada3b46),
	.w3(32'h3c2c0103),
	.w4(32'h3a95aac3),
	.w5(32'h3b6a607a),
	.w6(32'h3c276e18),
	.w7(32'hb7f28c80),
	.w8(32'h3a27730c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b433e27),
	.w1(32'hbaf9318c),
	.w2(32'hbaf7983b),
	.w3(32'h3b2a050a),
	.w4(32'hbb4e8c6f),
	.w5(32'hbb5a185a),
	.w6(32'h3b915dc3),
	.w7(32'hba9e2a03),
	.w8(32'hbaea3071),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be51138),
	.w1(32'h3aba6dc4),
	.w2(32'h3b047cf7),
	.w3(32'h3ba9e078),
	.w4(32'h39063f49),
	.w5(32'h3a30a6bd),
	.w6(32'h3b9a14df),
	.w7(32'h3a1807dd),
	.w8(32'h3a9a9255),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39915eab),
	.w1(32'hb9597c28),
	.w2(32'h386b433e),
	.w3(32'hb8690e2d),
	.w4(32'hba796dd5),
	.w5(32'hba9d04a0),
	.w6(32'hb75d64dc),
	.w7(32'hba8990ae),
	.w8(32'hbacd8646),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55d6a2),
	.w1(32'h3a31563e),
	.w2(32'h3bbda7e5),
	.w3(32'h3c260279),
	.w4(32'hb93e4894),
	.w5(32'h39bb45d9),
	.w6(32'h3c46dbf8),
	.w7(32'h3b2edaef),
	.w8(32'h3ba68e89),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024867),
	.w1(32'h3aa3fd0e),
	.w2(32'h3b08fc37),
	.w3(32'h3bb6e6ad),
	.w4(32'hba9b2928),
	.w5(32'hbad4e841),
	.w6(32'h3badc66f),
	.w7(32'hbaa8085d),
	.w8(32'hbaa14584),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff2304),
	.w1(32'hb976c5fe),
	.w2(32'h3b52f492),
	.w3(32'h3be08484),
	.w4(32'h39ef61b8),
	.w5(32'h3b2779bd),
	.w6(32'h3bbbcf4c),
	.w7(32'hb8c22a94),
	.w8(32'h3b3814d6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908c477),
	.w1(32'h39892be9),
	.w2(32'hb88feab3),
	.w3(32'h39a58308),
	.w4(32'h392a17f9),
	.w5(32'h37b18e58),
	.w6(32'h39b2a7a0),
	.w7(32'h391a16b4),
	.w8(32'h384787d9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8588de),
	.w1(32'hba381096),
	.w2(32'h3adf77f4),
	.w3(32'h3b4ce3d8),
	.w4(32'hba4106b1),
	.w5(32'h3a4fd5a4),
	.w6(32'h3b2e433d),
	.w7(32'hba9c22f5),
	.w8(32'h3a2c5072),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932fd36),
	.w1(32'hb85fbddd),
	.w2(32'hb7737e06),
	.w3(32'hb90e7eef),
	.w4(32'hb7a49f1a),
	.w5(32'h3734b7ec),
	.w6(32'hb918d32f),
	.w7(32'hb8312755),
	.w8(32'hb7375a61),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7a78b),
	.w1(32'h39b8e196),
	.w2(32'h3a60557e),
	.w3(32'h3a6f083f),
	.w4(32'hb7966518),
	.w5(32'h39767009),
	.w6(32'h3a7977e8),
	.w7(32'hb9d6c4b1),
	.w8(32'h3941ca64),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3d766),
	.w1(32'h39fe12ae),
	.w2(32'h39ed6421),
	.w3(32'h3acd8fc8),
	.w4(32'hb992310c),
	.w5(32'h391173e6),
	.w6(32'h3aa8988d),
	.w7(32'h385c8db8),
	.w8(32'h39e1c70d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdab99),
	.w1(32'h39f20e6a),
	.w2(32'h3b46ee9d),
	.w3(32'h3b7531f7),
	.w4(32'hba03e582),
	.w5(32'h3873b3db),
	.w6(32'h3b8de99a),
	.w7(32'hb900ca64),
	.w8(32'h3accdc35),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8778a0c),
	.w1(32'hb78e5e5f),
	.w2(32'hb65426cf),
	.w3(32'hb8621969),
	.w4(32'h36e916a8),
	.w5(32'h37a6517a),
	.w6(32'hb88829ba),
	.w7(32'hb74a474f),
	.w8(32'hb70037ef),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381314d2),
	.w1(32'hb72cd61c),
	.w2(32'hb8087a59),
	.w3(32'hb825afd7),
	.w4(32'hb68daa27),
	.w5(32'h37d847a4),
	.w6(32'hb9058651),
	.w7(32'hb8087825),
	.w8(32'h38006c7f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d39a8),
	.w1(32'h3999bafb),
	.w2(32'h39bf70a8),
	.w3(32'h3aa5604a),
	.w4(32'hbad5fa5c),
	.w5(32'hbaf82381),
	.w6(32'h3a5a5355),
	.w7(32'hbafe1d16),
	.w8(32'hba9b1e43),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1edfd),
	.w1(32'hba511ac7),
	.w2(32'hbae7f46a),
	.w3(32'h3b9aa382),
	.w4(32'hba5ef0b8),
	.w5(32'hbbc03082),
	.w6(32'h3b8e1529),
	.w7(32'hbaec329b),
	.w8(32'hbb5270a1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836ccd),
	.w1(32'h3a1661db),
	.w2(32'hbb49514f),
	.w3(32'h3aef49a9),
	.w4(32'hb9a6226c),
	.w5(32'hbb065de5),
	.w6(32'h3a3b9466),
	.w7(32'hba4ae1c4),
	.w8(32'hbb66569e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3856dfe0),
	.w1(32'hba409715),
	.w2(32'hb9daa8bd),
	.w3(32'h3a4cc807),
	.w4(32'hb9393a17),
	.w5(32'hb8e44a31),
	.w6(32'h3a98e5e1),
	.w7(32'hb901b9a3),
	.w8(32'h3a399066),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ed8c2),
	.w1(32'h3b66276c),
	.w2(32'h3c25007f),
	.w3(32'h3c836400),
	.w4(32'h3ba2575b),
	.w5(32'h3c025dab),
	.w6(32'h3c47d541),
	.w7(32'hb9bc2e76),
	.w8(32'h3be6fc79),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ff619),
	.w1(32'hb9eda9ec),
	.w2(32'h3a40d1c9),
	.w3(32'h3c1eb9ed),
	.w4(32'hbbaa3bc5),
	.w5(32'hbbb18ba2),
	.w6(32'h3c26652c),
	.w7(32'hbb9e7a6f),
	.w8(32'hbb809b6c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949bb4e),
	.w1(32'h3a1ab341),
	.w2(32'hb92c6e45),
	.w3(32'hb976a986),
	.w4(32'h39b12786),
	.w5(32'h3a2e06a8),
	.w6(32'h38a35386),
	.w7(32'h3a97b150),
	.w8(32'h3a844e9b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88232f4),
	.w1(32'h37fde570),
	.w2(32'h381310cc),
	.w3(32'hb8589dcc),
	.w4(32'h382dac38),
	.w5(32'h389222d4),
	.w6(32'hb8e7f0ed),
	.w7(32'h3891787c),
	.w8(32'h388d0a84),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39490064),
	.w1(32'hb86ea0bd),
	.w2(32'hb8e29dac),
	.w3(32'hb883b82f),
	.w4(32'hb8ca11b2),
	.w5(32'hb91fe820),
	.w6(32'hb8babdb4),
	.w7(32'hb9037411),
	.w8(32'hb832c9e1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb6939),
	.w1(32'hb7b00d50),
	.w2(32'hb735b354),
	.w3(32'hb8cded0a),
	.w4(32'h36195999),
	.w5(32'h3730d7f7),
	.w6(32'hb8d6a8d9),
	.w7(32'hb79a6fde),
	.w8(32'hb79e5393),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a829d43),
	.w1(32'h3a3928d6),
	.w2(32'h39b7fed9),
	.w3(32'h3a3fc2fa),
	.w4(32'h3aa6ff0c),
	.w5(32'h3a01d5e7),
	.w6(32'h3a860445),
	.w7(32'h3ae6c8eb),
	.w8(32'h399968cb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfa418),
	.w1(32'h3adf1a11),
	.w2(32'h3658c1fb),
	.w3(32'h3b4412df),
	.w4(32'hbac01ecf),
	.w5(32'hbb655f52),
	.w6(32'h3b7d9a8d),
	.w7(32'h3a2edd6e),
	.w8(32'h3a3a93aa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cdcda),
	.w1(32'h3b49a7b0),
	.w2(32'h3bb3e084),
	.w3(32'h3be6737b),
	.w4(32'hbaac678a),
	.w5(32'h3a07a854),
	.w6(32'h3bd8e48f),
	.w7(32'hba6cebdd),
	.w8(32'hba6088de),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95c051),
	.w1(32'hba484bb0),
	.w2(32'hb9987796),
	.w3(32'h3a6359a8),
	.w4(32'hba8f00d1),
	.w5(32'hba969ae2),
	.w6(32'h3a9844bf),
	.w7(32'hba711500),
	.w8(32'hba331db5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cecc1),
	.w1(32'h3b28fd18),
	.w2(32'h3b6b1290),
	.w3(32'h3b9b347f),
	.w4(32'h3b2c7d49),
	.w5(32'h3a9c4072),
	.w6(32'h3b90e557),
	.w7(32'h3ad03a4b),
	.w8(32'h3b0925c4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99e510),
	.w1(32'hba018b5a),
	.w2(32'hbadd421f),
	.w3(32'h3a02e80d),
	.w4(32'hb9af0e91),
	.w5(32'hbab6fb76),
	.w6(32'h3aa6c51a),
	.w7(32'h396075db),
	.w8(32'hbae7534d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926dae7),
	.w1(32'hb83d68ec),
	.w2(32'hb8546f58),
	.w3(32'hb90fefd6),
	.w4(32'hb7a7ba9d),
	.w5(32'hb7765bfb),
	.w6(32'hb9280599),
	.w7(32'hb82708c0),
	.w8(32'hb8464f85),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95d97),
	.w1(32'h39b7e706),
	.w2(32'hb91e69f6),
	.w3(32'h3a663add),
	.w4(32'h3ac36bf3),
	.w5(32'hbab93296),
	.w6(32'h39c2d70b),
	.w7(32'hba3643bd),
	.w8(32'hbb1bd435),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd0a08),
	.w1(32'hb8d6266b),
	.w2(32'hb8a7591f),
	.w3(32'hb9a14605),
	.w4(32'hb7c12e68),
	.w5(32'h3822f409),
	.w6(32'hb9b369f9),
	.w7(32'hb8b9c6ba),
	.w8(32'hb8460e3b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be07506),
	.w1(32'h3a8ac6f9),
	.w2(32'h3a94de48),
	.w3(32'h3ba80184),
	.w4(32'hb7a2e30b),
	.w5(32'hbac968ac),
	.w6(32'h3ba57b5a),
	.w7(32'hba20a9a3),
	.w8(32'hbaaff035),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be08ef2),
	.w1(32'hb9c3ff96),
	.w2(32'hbaf13964),
	.w3(32'h3b9021ff),
	.w4(32'hbb98f6c3),
	.w5(32'hbb9eef6e),
	.w6(32'h3be131b0),
	.w7(32'hbaf03947),
	.w8(32'hbb3c639c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befd36b),
	.w1(32'h3af9251b),
	.w2(32'h3b02398c),
	.w3(32'h3bab0833),
	.w4(32'hb940f285),
	.w5(32'hb8f6e0e1),
	.w6(32'h3ba89e9d),
	.w7(32'h397b7f38),
	.w8(32'h3a0fc4e9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a492502),
	.w1(32'hba79cbd7),
	.w2(32'hbaf62dad),
	.w3(32'h3a48b875),
	.w4(32'hba5fcaa6),
	.w5(32'hbaf2c8f1),
	.w6(32'h3aac95c0),
	.w7(32'hb89804e3),
	.w8(32'hba3f8fa3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa0db9),
	.w1(32'h3aa1464d),
	.w2(32'h3b5c49fa),
	.w3(32'h3bae8b15),
	.w4(32'hbaffceac),
	.w5(32'hbabc817e),
	.w6(32'h3bbee985),
	.w7(32'hba5de901),
	.w8(32'hba348e12),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa75a0),
	.w1(32'h3a419f28),
	.w2(32'h3a8486d5),
	.w3(32'h3b8e509b),
	.w4(32'h3a7d8166),
	.w5(32'hb88c0da2),
	.w6(32'h3b868b4d),
	.w7(32'h3ad50c2c),
	.w8(32'h3a8a2a96),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c252023),
	.w1(32'hb8e6e1a7),
	.w2(32'h3b2bb9e4),
	.w3(32'h3bfbd4ed),
	.w4(32'hbb79a1f9),
	.w5(32'hbaa56a56),
	.w6(32'h3bec3cb5),
	.w7(32'hbb237fce),
	.w8(32'h3a59c9fa),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f243c2),
	.w1(32'h36ad810e),
	.w2(32'hb71e67d3),
	.w3(32'hb84f1330),
	.w4(32'hb79c543f),
	.w5(32'h37de11d3),
	.w6(32'hb912b121),
	.w7(32'hb83a8a5d),
	.w8(32'hb89f60f5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934859c),
	.w1(32'hb98f0aee),
	.w2(32'hb90b5233),
	.w3(32'hb900ca83),
	.w4(32'hb9030f51),
	.w5(32'hb7753b58),
	.w6(32'h37b26696),
	.w7(32'hb945ea76),
	.w8(32'h36ceb277),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2a3dc),
	.w1(32'h3aa7fb77),
	.w2(32'hb96b36e7),
	.w3(32'h3b944e7d),
	.w4(32'hbb21f764),
	.w5(32'hbb5e35b9),
	.w6(32'h3bbb03b5),
	.w7(32'hbae6924e),
	.w8(32'hbb810fde),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e4f2f),
	.w1(32'h3a2c0cd6),
	.w2(32'h3a9fcff3),
	.w3(32'h3c1c4df2),
	.w4(32'h3a7ca104),
	.w5(32'h3a8faacc),
	.w6(32'h3c1084a0),
	.w7(32'hbae4ba71),
	.w8(32'hbaa3e594),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d1321),
	.w1(32'h3ada9829),
	.w2(32'h3b209796),
	.w3(32'h3bd5b5fa),
	.w4(32'hbb1367cd),
	.w5(32'hbaa0b2ac),
	.w6(32'h3bb53d62),
	.w7(32'hbb05b39f),
	.w8(32'hb997ab61),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc94a5),
	.w1(32'hb9004a8c),
	.w2(32'h390b10dc),
	.w3(32'h391706e7),
	.w4(32'h3a8ff182),
	.w5(32'hb921ec1c),
	.w6(32'hba818436),
	.w7(32'hbaa95c01),
	.w8(32'h3b365fd2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e267ef),
	.w1(32'h39341283),
	.w2(32'h39fcb5e4),
	.w3(32'h38b7cc89),
	.w4(32'h39c3d2d7),
	.w5(32'h39ee6ae1),
	.w6(32'h3863169c),
	.w7(32'h399f0978),
	.w8(32'h39ca9ef2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5425af),
	.w1(32'h3a5e0427),
	.w2(32'h39b7004d),
	.w3(32'h3a4c47e2),
	.w4(32'h3a32269f),
	.w5(32'h39a7f62a),
	.w6(32'h3a0c84e8),
	.w7(32'h399ea875),
	.w8(32'hb92b366c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e8dd),
	.w1(32'h3a0c4eb8),
	.w2(32'hbaae5981),
	.w3(32'h3aa402fe),
	.w4(32'h3afb1206),
	.w5(32'h399c6b01),
	.w6(32'h3b190279),
	.w7(32'h3b323607),
	.w8(32'hbb5e246c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c297bef),
	.w1(32'h3af2ffff),
	.w2(32'h3b83068e),
	.w3(32'h3c1a7227),
	.w4(32'h3b8a4e72),
	.w5(32'h384c7e17),
	.w6(32'h3bfce498),
	.w7(32'hb891a383),
	.w8(32'h3b498aa5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba40c50),
	.w1(32'h3b425ed9),
	.w2(32'hb932495d),
	.w3(32'hba2e3d9b),
	.w4(32'h3b194224),
	.w5(32'h397f4f90),
	.w6(32'h3a84e62e),
	.w7(32'h3a17e68b),
	.w8(32'hbb1e4f97),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d16f),
	.w1(32'hbb210968),
	.w2(32'hbaa15ee2),
	.w3(32'h3b4a8b8c),
	.w4(32'hbb8cb38e),
	.w5(32'hbb854a46),
	.w6(32'h3b95eb6a),
	.w7(32'hbb01562d),
	.w8(32'hbb2d62eb),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf104cd),
	.w1(32'h3aaec618),
	.w2(32'h3b0e3148),
	.w3(32'h3bc9be5f),
	.w4(32'hbb094b08),
	.w5(32'hbb271275),
	.w6(32'h3bdf71e3),
	.w7(32'hbacf31e7),
	.w8(32'hbaa1f1d9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89ede87),
	.w1(32'hb7cb339c),
	.w2(32'hb7b3ed8a),
	.w3(32'hb880a636),
	.w4(32'hb7987ae1),
	.w5(32'hb714d9cf),
	.w6(32'hb88a8c79),
	.w7(32'hb7fe973a),
	.w8(32'hb7dbe76b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d39813),
	.w1(32'hb8119b74),
	.w2(32'hb7f02ecf),
	.w3(32'hb8b349ce),
	.w4(32'hb799229c),
	.w5(32'hb7813a0d),
	.w6(32'hb8c92dc4),
	.w7(32'hb80ecfef),
	.w8(32'hb7c4da95),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9162f97),
	.w1(32'hb8187d77),
	.w2(32'hb93bd064),
	.w3(32'hba85fd6c),
	.w4(32'hb9ecaa45),
	.w5(32'hb8b40595),
	.w6(32'hb9d780f4),
	.w7(32'hb7ba1633),
	.w8(32'hb916d86d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d2c16),
	.w1(32'hb6e39aaf),
	.w2(32'h37242537),
	.w3(32'hb8f60811),
	.w4(32'h37af0ce6),
	.w5(32'hba022bc3),
	.w6(32'hb91c2c8c),
	.w7(32'hb5ecf959),
	.w8(32'hb9e60038),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40dc5f),
	.w1(32'h3a8b2b0b),
	.w2(32'h3a5ae5f6),
	.w3(32'hba2bcfb9),
	.w4(32'h398ae909),
	.w5(32'hb86a5b99),
	.w6(32'h39016df5),
	.w7(32'h3a486318),
	.w8(32'hb8ce1d3f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095d26),
	.w1(32'h3ad02089),
	.w2(32'h3aa79616),
	.w3(32'h3bd4c0d9),
	.w4(32'h3af27d7c),
	.w5(32'h3a1be75d),
	.w6(32'h3bc7c361),
	.w7(32'h398b92a4),
	.w8(32'h3a8478f2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd083d9),
	.w1(32'h3abe7cec),
	.w2(32'h3acbd2e9),
	.w3(32'h3ba2983a),
	.w4(32'h3a3e9395),
	.w5(32'h3a715053),
	.w6(32'h3b631fd4),
	.w7(32'h3a91b102),
	.w8(32'h39dc9baa),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00ede8),
	.w1(32'hba329f1a),
	.w2(32'hb94fb78e),
	.w3(32'h39274965),
	.w4(32'h3a0bd187),
	.w5(32'hb897910a),
	.w6(32'h39feffaa),
	.w7(32'h399a0dd1),
	.w8(32'h3807be8b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a7422),
	.w1(32'h3b6f23a8),
	.w2(32'hb9f69d0c),
	.w3(32'h3b661938),
	.w4(32'h3b119588),
	.w5(32'h383f0a65),
	.w6(32'h3b047b27),
	.w7(32'hbb2ce6f7),
	.w8(32'hbb338e57),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad09461),
	.w1(32'hba90cb4e),
	.w2(32'h37d2e56b),
	.w3(32'h3ad93917),
	.w4(32'hb9b27998),
	.w5(32'h3a1ad246),
	.w6(32'h3ae4fcb4),
	.w7(32'hba657ec9),
	.w8(32'h38d7ea6b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9818859),
	.w1(32'hba55b1e4),
	.w2(32'hba0d9de8),
	.w3(32'hba3ef20b),
	.w4(32'hba2646b4),
	.w5(32'hbaa48373),
	.w6(32'hba5cb932),
	.w7(32'hba8c8d2e),
	.w8(32'hba818f32),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b064d7f),
	.w1(32'hb923efe1),
	.w2(32'h3a316c5c),
	.w3(32'h3a94479b),
	.w4(32'h3a5dfa4d),
	.w5(32'hb95ad6fa),
	.w6(32'h3a714a55),
	.w7(32'h3a6ff047),
	.w8(32'h3a04a97c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afa7a8),
	.w1(32'hba26ab2f),
	.w2(32'hba6e7268),
	.w3(32'hba96f5b4),
	.w4(32'hb9630409),
	.w5(32'h38d9c7e9),
	.w6(32'hbaa25705),
	.w7(32'hb9fac6b0),
	.w8(32'hb8117cb7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e91532),
	.w1(32'h398e0527),
	.w2(32'h3999391c),
	.w3(32'h3a271019),
	.w4(32'h3953926a),
	.w5(32'hbaa59a9e),
	.w6(32'h3a81a92f),
	.w7(32'h396b5f61),
	.w8(32'hba7a6e91),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c7a99),
	.w1(32'hba568531),
	.w2(32'hba485914),
	.w3(32'hbac507fe),
	.w4(32'hba8b04b7),
	.w5(32'hba3e698f),
	.w6(32'hba80d0e6),
	.w7(32'hba6a235f),
	.w8(32'hba3f7a25),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c0176),
	.w1(32'hb9eca9e3),
	.w2(32'hb9a90a2d),
	.w3(32'hba16d50e),
	.w4(32'hb9c3981c),
	.w5(32'h3a2f0538),
	.w6(32'hba0bea95),
	.w7(32'hb9858923),
	.w8(32'h3a43d56f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed0bca),
	.w1(32'hb9df0dba),
	.w2(32'hba43a24c),
	.w3(32'h3b0922b9),
	.w4(32'h3a00c255),
	.w5(32'hba6f6967),
	.w6(32'h3b3dbbc1),
	.w7(32'h3a87ec4d),
	.w8(32'hba3c020c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12517e),
	.w1(32'hba0712eb),
	.w2(32'h3b645e5a),
	.w3(32'h3c013f4e),
	.w4(32'h3a5c0939),
	.w5(32'h3b18f99c),
	.w6(32'h3bf53d84),
	.w7(32'h3af9ef68),
	.w8(32'h3bae5142),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06b930),
	.w1(32'h3acc6e18),
	.w2(32'h3af4a805),
	.w3(32'h3be8540e),
	.w4(32'h3b2ff542),
	.w5(32'h3ae2378e),
	.w6(32'h3bae9aa3),
	.w7(32'h3aadecad),
	.w8(32'h3aa9ee95),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca4fb0),
	.w1(32'h3a6a5ae9),
	.w2(32'h3b941b51),
	.w3(32'h3ba77ebd),
	.w4(32'h3aef8fb9),
	.w5(32'h3b2fc51b),
	.w6(32'h3b905abf),
	.w7(32'h3aaf23d5),
	.w8(32'h3b7ee216),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c0937),
	.w1(32'hba21b441),
	.w2(32'hb8ce6915),
	.w3(32'h3994df32),
	.w4(32'hb9ebd22d),
	.w5(32'hb9a4cebb),
	.w6(32'h3948cf21),
	.w7(32'hb9a08a8b),
	.w8(32'hb9f47812),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90941d8),
	.w1(32'hb933b0fc),
	.w2(32'hb8a4b359),
	.w3(32'h394b6967),
	.w4(32'h393bfaa7),
	.w5(32'hba1f4047),
	.w6(32'hb910d901),
	.w7(32'h38795458),
	.w8(32'hba2f9ed0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04ebfe),
	.w1(32'hb8db5703),
	.w2(32'hb903aff8),
	.w3(32'hb98ac58f),
	.w4(32'hb9752c14),
	.w5(32'h38ae3da9),
	.w6(32'hb803e1e7),
	.w7(32'hb8451444),
	.w8(32'hb9881cdf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56ec0a),
	.w1(32'hba9bbf4f),
	.w2(32'h3791af67),
	.w3(32'hba42692a),
	.w4(32'hba057d33),
	.w5(32'hb9c4e971),
	.w6(32'hba38d0da),
	.w7(32'hb961a4aa),
	.w8(32'hb9e23424),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c223af9),
	.w1(32'h3b3cdf1a),
	.w2(32'h3bbc4f9f),
	.w3(32'h3be24299),
	.w4(32'h3b069c08),
	.w5(32'h3ad67811),
	.w6(32'h3baace7a),
	.w7(32'h3722e64b),
	.w8(32'hba234cde),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09efe1),
	.w1(32'hbb33510f),
	.w2(32'hbb1c1e52),
	.w3(32'hbb1a8ef3),
	.w4(32'hbb08bcc8),
	.w5(32'h3a3a5059),
	.w6(32'hbb2686c6),
	.w7(32'hbafa8fa9),
	.w8(32'h3a4e5a2c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d731),
	.w1(32'hba9fab1e),
	.w2(32'hba52bbb4),
	.w3(32'h3ac2778c),
	.w4(32'hbaab2d93),
	.w5(32'hb9a7d092),
	.w6(32'h3b120f8d),
	.w7(32'hb996e62a),
	.w8(32'h3a423628),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349f8a),
	.w1(32'h3a0a9f24),
	.w2(32'h38b6e0cc),
	.w3(32'h3b367e96),
	.w4(32'h3957d63e),
	.w5(32'hbaa11dfc),
	.w6(32'h3b245650),
	.w7(32'h3941a72f),
	.w8(32'hb98f1752),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ec680),
	.w1(32'h3a1a04ac),
	.w2(32'h3a11951c),
	.w3(32'h3893a3f2),
	.w4(32'h3906eeda),
	.w5(32'h3a69d31d),
	.w6(32'h39d02022),
	.w7(32'h39f46e0b),
	.w8(32'h3a7198a3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1971dc),
	.w1(32'h3a99a2da),
	.w2(32'h3aeab5ad),
	.w3(32'h3af8c491),
	.w4(32'h3a874c0b),
	.w5(32'h3a566c46),
	.w6(32'h3aaa8853),
	.w7(32'h3a3a08d1),
	.w8(32'h3aaed5b4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a951976),
	.w1(32'h3a9b5ed5),
	.w2(32'h3a94cc92),
	.w3(32'h3a11a803),
	.w4(32'h3a23ba5a),
	.w5(32'h39aefe6a),
	.w6(32'h3a2586c4),
	.w7(32'h3a4cfd67),
	.w8(32'h37854284),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c151e07),
	.w1(32'h3b691b69),
	.w2(32'h3ba3d3e8),
	.w3(32'h3bc6f602),
	.w4(32'h3b6c5a6b),
	.w5(32'h38b18f9c),
	.w6(32'h3c003351),
	.w7(32'h3b1467a8),
	.w8(32'h3ac2f839),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f95a35),
	.w1(32'h397de378),
	.w2(32'h390ca080),
	.w3(32'h3916b526),
	.w4(32'h38280280),
	.w5(32'hb997c926),
	.w6(32'h3a735c7f),
	.w7(32'h39e305cc),
	.w8(32'hba0ea991),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46bd6b),
	.w1(32'hbb32ff83),
	.w2(32'hbbb89cbf),
	.w3(32'h3b462e8e),
	.w4(32'hbb9b9839),
	.w5(32'hbba6d84b),
	.w6(32'h3b1b1f40),
	.w7(32'hbbc11777),
	.w8(32'hbbfdef5a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule