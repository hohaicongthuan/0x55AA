module layer_10_featuremap_341(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82d3df),
	.w1(32'hbb3ba6d5),
	.w2(32'hbb8f0d31),
	.w3(32'hbb3d9510),
	.w4(32'hbb644647),
	.w5(32'h3b081a7b),
	.w6(32'hba53c613),
	.w7(32'hbb18163b),
	.w8(32'hba1d77e1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcc79f),
	.w1(32'h3afac016),
	.w2(32'h3be3dd04),
	.w3(32'h3bea5063),
	.w4(32'hbb1bd751),
	.w5(32'hbb3fe722),
	.w6(32'h3bc74de3),
	.w7(32'hba21826a),
	.w8(32'h3b3ada71),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998279c),
	.w1(32'h3a8f68c3),
	.w2(32'hb99da374),
	.w3(32'hba8074b9),
	.w4(32'h39abb643),
	.w5(32'h3b0364c5),
	.w6(32'hb9dc2309),
	.w7(32'hba092604),
	.w8(32'h3b1352f6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395022d1),
	.w1(32'h3aa5172e),
	.w2(32'h3a049351),
	.w3(32'h3b08247a),
	.w4(32'h3b3f215c),
	.w5(32'h3a61a671),
	.w6(32'h3b2b6463),
	.w7(32'h3b18bdfd),
	.w8(32'hbab5ad83),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02b758),
	.w1(32'h39ada564),
	.w2(32'h3bd1403d),
	.w3(32'hb920ef9a),
	.w4(32'h3be11bc5),
	.w5(32'hb98fefac),
	.w6(32'hbb57bee9),
	.w7(32'h3b161caf),
	.w8(32'h3a7f4388),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d607d3),
	.w1(32'h3ae51d2b),
	.w2(32'h3b0c398a),
	.w3(32'h39ca3b59),
	.w4(32'h3a57b3e2),
	.w5(32'h3bd54499),
	.w6(32'h3aa28722),
	.w7(32'h3ae60936),
	.w8(32'h3bd30aef),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb906e),
	.w1(32'h3c530e75),
	.w2(32'h3ca14869),
	.w3(32'h3bd72124),
	.w4(32'h3c6d0a4f),
	.w5(32'h3c67c937),
	.w6(32'h3bacf5f9),
	.w7(32'h3c56300c),
	.w8(32'h3c70979c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97838a),
	.w1(32'h3c4e95a3),
	.w2(32'h3bdb0057),
	.w3(32'h3c857899),
	.w4(32'h3c5db5d6),
	.w5(32'h3c20327a),
	.w6(32'h3c934c65),
	.w7(32'h3bdf39c3),
	.w8(32'h3c27eb13),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae52444),
	.w1(32'hba67aeca),
	.w2(32'h3b1213f9),
	.w3(32'h3afe44c4),
	.w4(32'h3a82abcc),
	.w5(32'h385197bd),
	.w6(32'h3b0f8583),
	.w7(32'h3b1b07bf),
	.w8(32'h3b427ef0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65b8c2),
	.w1(32'h3bc4e436),
	.w2(32'h3cb7b529),
	.w3(32'h3c2ebdf0),
	.w4(32'h3ac2567f),
	.w5(32'h3c7fbb7b),
	.w6(32'h3c6d49d4),
	.w7(32'h3bc4c8be),
	.w8(32'h3ca2c274),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28bbc1),
	.w1(32'h3b298602),
	.w2(32'h3b374fd8),
	.w3(32'h3aa10cdb),
	.w4(32'h3ac164a5),
	.w5(32'hba2c54e2),
	.w6(32'h3b3286c2),
	.w7(32'h3b443500),
	.w8(32'h3a0a1434),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38b962),
	.w1(32'hbb6eb9b8),
	.w2(32'h3b9d9ea5),
	.w3(32'h3b612d51),
	.w4(32'h3a901bd2),
	.w5(32'h3b951c32),
	.w6(32'h3b96c84b),
	.w7(32'hba9f2962),
	.w8(32'h3c041108),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14f5cf),
	.w1(32'h3b957ee9),
	.w2(32'h3cb177b1),
	.w3(32'h3bc61f45),
	.w4(32'h3b4b115b),
	.w5(32'h3ca1edad),
	.w6(32'h3b8ff465),
	.w7(32'h3b8f09ef),
	.w8(32'h3c9d583b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8d996),
	.w1(32'h3c229e15),
	.w2(32'h3c86a0b1),
	.w3(32'h3b006c0c),
	.w4(32'h3bfc8e8d),
	.w5(32'h3c203260),
	.w6(32'h3b63e141),
	.w7(32'h3bfab6cd),
	.w8(32'h3c1e500c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c316bd7),
	.w1(32'h3a3a3491),
	.w2(32'h3ba44691),
	.w3(32'h3b875309),
	.w4(32'hbbe630c5),
	.w5(32'hbbb9d0f6),
	.w6(32'h3c1bbfae),
	.w7(32'hbab8f955),
	.w8(32'hba055e94),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c327e22),
	.w1(32'h3b78f8aa),
	.w2(32'h3c9644c4),
	.w3(32'h3bb23fef),
	.w4(32'hbaeae08c),
	.w5(32'h3c0affd1),
	.w6(32'h3be99602),
	.w7(32'h3bf5d554),
	.w8(32'h3c610c78),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03bb6),
	.w1(32'hb9c14c73),
	.w2(32'h389dc8eb),
	.w3(32'h38ca0f09),
	.w4(32'h390b0a31),
	.w5(32'hba988df5),
	.w6(32'h398223bf),
	.w7(32'hb91d2329),
	.w8(32'hbacc1dc9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fe212),
	.w1(32'h3ba4040a),
	.w2(32'h3c513e78),
	.w3(32'h3c0818a4),
	.w4(32'h3b0c1af9),
	.w5(32'h3c88076c),
	.w6(32'h3c2fc587),
	.w7(32'h3b95465e),
	.w8(32'h3c9d86d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef7967),
	.w1(32'h3bb20a8d),
	.w2(32'h3c3ffb75),
	.w3(32'h3b140986),
	.w4(32'h3b829c1b),
	.w5(32'h3c3bc630),
	.w6(32'h3bb69f2f),
	.w7(32'h3bd30754),
	.w8(32'h3c28dd03),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d4170),
	.w1(32'hbb281582),
	.w2(32'hba20050a),
	.w3(32'hb8ac2039),
	.w4(32'h39c4718b),
	.w5(32'hbb7056f0),
	.w6(32'hba2b6d0d),
	.w7(32'h39f925d9),
	.w8(32'hbb6a935d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37b1e8),
	.w1(32'hbb537696),
	.w2(32'hb83a4f47),
	.w3(32'hbb2ceddf),
	.w4(32'hb9d79745),
	.w5(32'h3b3ef117),
	.w6(32'hbb6fe119),
	.w7(32'hba777489),
	.w8(32'h3b2524e9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2503c0),
	.w1(32'hba841465),
	.w2(32'h3ba0d62e),
	.w3(32'h3aa80f54),
	.w4(32'hbb85fbba),
	.w5(32'hbab5c04d),
	.w6(32'h3b8c23cd),
	.w7(32'hbae94532),
	.w8(32'h3a59bd1b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cececb0),
	.w1(32'h3a8db106),
	.w2(32'h3c1ff42e),
	.w3(32'h3c9ae4c8),
	.w4(32'hbb9dd65d),
	.w5(32'h3c2d630f),
	.w6(32'h3cc878fa),
	.w7(32'h3c201480),
	.w8(32'h3cf2c1d8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c292d7f),
	.w1(32'hbad2b5e6),
	.w2(32'h3c88c916),
	.w3(32'h3b6d7b48),
	.w4(32'hbb9b2aea),
	.w5(32'h3c083cf2),
	.w6(32'h3c1e2b3f),
	.w7(32'hb9db037a),
	.w8(32'h3c582cfe),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb93c9c),
	.w1(32'h3a584130),
	.w2(32'h3c66bcfd),
	.w3(32'h3c7c2bc5),
	.w4(32'hbc0e3b1e),
	.w5(32'h3b73c03e),
	.w6(32'h3cc5ae50),
	.w7(32'hbb113f86),
	.w8(32'h3c546416),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0687d0),
	.w1(32'h3b8a96c6),
	.w2(32'h3b9ea9cd),
	.w3(32'h3af1216a),
	.w4(32'h3b43c739),
	.w5(32'h3ba16382),
	.w6(32'h3b86f499),
	.w7(32'h3bb68116),
	.w8(32'h3bc41ff0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842af8),
	.w1(32'h3bb44ba8),
	.w2(32'h3bef571f),
	.w3(32'h3b815f30),
	.w4(32'h3bcab2d7),
	.w5(32'hbad2bfb2),
	.w6(32'h3b9d29a1),
	.w7(32'h3bf33e6a),
	.w8(32'hbb32509e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fafc9),
	.w1(32'hbc303676),
	.w2(32'h3acd9e30),
	.w3(32'hbb54485e),
	.w4(32'hbc15fee1),
	.w5(32'hbb1b5531),
	.w6(32'hbb09b883),
	.w7(32'hbb573a70),
	.w8(32'h3acaa537),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc68041),
	.w1(32'hb9d98c41),
	.w2(32'h3b0df57a),
	.w3(32'h3b55c04d),
	.w4(32'hbb7ded03),
	.w5(32'hbad4c5bd),
	.w6(32'h3bc1ef35),
	.w7(32'hbae3237b),
	.w8(32'hba825956),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad84145),
	.w1(32'hbc24947b),
	.w2(32'h3b4a7d7e),
	.w3(32'h3b4121de),
	.w4(32'hbbf8bc26),
	.w5(32'h3aa1ca2a),
	.w6(32'h3bbcd377),
	.w7(32'hbb64313d),
	.w8(32'h3ba09cd8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28cf0f),
	.w1(32'hbb2e3c5c),
	.w2(32'hbac0cbc6),
	.w3(32'hbb03e0f0),
	.w4(32'hbaf5da75),
	.w5(32'hba37e99d),
	.w6(32'hbba4adb7),
	.w7(32'hbb45615c),
	.w8(32'hba39f93c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443cf7),
	.w1(32'hbab5291b),
	.w2(32'h3abab492),
	.w3(32'hb905011b),
	.w4(32'h3b36e3b2),
	.w5(32'h3a5610db),
	.w6(32'hba4db1ed),
	.w7(32'h3a4e463b),
	.w8(32'h3a33d922),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815147),
	.w1(32'hbacd1e5b),
	.w2(32'h3c2136e5),
	.w3(32'h3abcfc0d),
	.w4(32'hbb193c2f),
	.w5(32'h3ae2fc2d),
	.w6(32'h3b849677),
	.w7(32'h3aae9b4f),
	.w8(32'h3b40a170),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85bbd3),
	.w1(32'hbb0a44a4),
	.w2(32'hba8346c1),
	.w3(32'h3b7d3158),
	.w4(32'hbba9bdb2),
	.w5(32'h3a3ceaa9),
	.w6(32'h3bae1e0c),
	.w7(32'hbb33d3d7),
	.w8(32'h3b34126b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1561e6),
	.w1(32'h3b010212),
	.w2(32'h3b18ba87),
	.w3(32'h3b257fd2),
	.w4(32'h3b3b4a8e),
	.w5(32'hbb92bf72),
	.w6(32'h3b3508c6),
	.w7(32'h3b6631d4),
	.w8(32'hbb7e5f1c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2862ca),
	.w1(32'hbacc15b0),
	.w2(32'h3b09e421),
	.w3(32'hbbb13401),
	.w4(32'h3a239ac2),
	.w5(32'h3b553cb1),
	.w6(32'hbbb1df2b),
	.w7(32'hb9ee1dff),
	.w8(32'h3b42f2b5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7fd6ba),
	.w1(32'h3b7911f9),
	.w2(32'h3c9043c4),
	.w3(32'h3bad65de),
	.w4(32'hbbc47f9e),
	.w5(32'h3c1d177e),
	.w6(32'h3a63d613),
	.w7(32'hbc1b37b4),
	.w8(32'h3c8bb105),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d056609),
	.w1(32'hbbd86f60),
	.w2(32'h3bc109cf),
	.w3(32'h3cba349d),
	.w4(32'hbc794231),
	.w5(32'hbc259306),
	.w6(32'h3d1d6e08),
	.w7(32'hb89d99e2),
	.w8(32'h3b9a27b2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0605a9),
	.w1(32'hbc859a75),
	.w2(32'hbba7a998),
	.w3(32'h3c9134ec),
	.w4(32'hbc3da1ef),
	.w5(32'hbb4aa33b),
	.w6(32'h3ce10b7f),
	.w7(32'hbb056654),
	.w8(32'h3c067cf1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad214a0),
	.w1(32'hbbf14850),
	.w2(32'hbb9ad30d),
	.w3(32'hba000c3b),
	.w4(32'hbc001ba7),
	.w5(32'h3a068e0c),
	.w6(32'h39bd7f5f),
	.w7(32'hbb8e9cca),
	.w8(32'h3b6f583a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46d347),
	.w1(32'h3b14a351),
	.w2(32'h3b0926e4),
	.w3(32'h3ad2c5cc),
	.w4(32'h3a98fe26),
	.w5(32'h3b268e6b),
	.w6(32'h3acf5c92),
	.w7(32'h3aa3dd15),
	.w8(32'h3b98b942),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b087a85),
	.w1(32'h3b804a3b),
	.w2(32'h3b986b6f),
	.w3(32'h3b2c73da),
	.w4(32'h3b81c218),
	.w5(32'hbb671843),
	.w6(32'h3b8df3d9),
	.w7(32'h3bad557a),
	.w8(32'hbb24f55d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f2884),
	.w1(32'hbbdea53f),
	.w2(32'hbb8975cc),
	.w3(32'hba2456a9),
	.w4(32'hbbdfc276),
	.w5(32'hb9adaeba),
	.w6(32'h39965c97),
	.w7(32'hbb33e9ee),
	.w8(32'h3ab6b7ec),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c97cd),
	.w1(32'h3be8d608),
	.w2(32'h3ca5c9d9),
	.w3(32'h3c3cd1f3),
	.w4(32'h3ba8c2a1),
	.w5(32'h3c70de72),
	.w6(32'h3c83d949),
	.w7(32'h3c8f4ba9),
	.w8(32'h3cd7327d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c637e7d),
	.w1(32'hba5f15a5),
	.w2(32'h3c849b00),
	.w3(32'h3bb42be7),
	.w4(32'hbc231910),
	.w5(32'h3b80be9e),
	.w6(32'h3c7b2c37),
	.w7(32'hba27ed54),
	.w8(32'h3c434a06),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90300b),
	.w1(32'h3a5aceb4),
	.w2(32'h3c750be6),
	.w3(32'h3bf04a84),
	.w4(32'hbc152660),
	.w5(32'h3bd25860),
	.w6(32'h3ca2c620),
	.w7(32'h397224b2),
	.w8(32'h3c53f95c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42a1c0),
	.w1(32'hbb65eea3),
	.w2(32'h3b8cb385),
	.w3(32'h3c19e25e),
	.w4(32'hbbd2fff5),
	.w5(32'h3b965142),
	.w6(32'h3c4bcf12),
	.w7(32'hbad48f89),
	.w8(32'h3c1fce07),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4385b1),
	.w1(32'h3c00b761),
	.w2(32'h3c7c2911),
	.w3(32'h3c02b85f),
	.w4(32'h3c3704f6),
	.w5(32'h3c8b1ff8),
	.w6(32'h3bf1dbe1),
	.w7(32'h3c216215),
	.w8(32'h3c838a0a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbfba4),
	.w1(32'hbaf87914),
	.w2(32'hbb48110c),
	.w3(32'hba61dd59),
	.w4(32'hbab6a011),
	.w5(32'h3b98672f),
	.w6(32'hbab2d274),
	.w7(32'hbaee88bd),
	.w8(32'h3bb61f40),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad65c8),
	.w1(32'h3b83705f),
	.w2(32'h3b7590a3),
	.w3(32'h3b68f41f),
	.w4(32'h3b8129c4),
	.w5(32'h3b4c68a7),
	.w6(32'h3ba1cf74),
	.w7(32'h3bae223a),
	.w8(32'h3b50dc0c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4babe9),
	.w1(32'hbaeb97af),
	.w2(32'h39ebcdb2),
	.w3(32'hb9a8ab31),
	.w4(32'h3a77d60d),
	.w5(32'hb9148c36),
	.w6(32'hbb582e9b),
	.w7(32'hb9ab5a40),
	.w8(32'hba6a1278),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c114ef9),
	.w1(32'h3b2fa835),
	.w2(32'h3c50275a),
	.w3(32'h3b85437b),
	.w4(32'hba9af2bf),
	.w5(32'h3be82f18),
	.w6(32'h3bb01e07),
	.w7(32'h3a9fe063),
	.w8(32'h3bb951ab),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb2acd),
	.w1(32'hb99533b0),
	.w2(32'h3b653a69),
	.w3(32'h39f03799),
	.w4(32'hb9c1d57b),
	.w5(32'h3b2d857d),
	.w6(32'h3a49d5f0),
	.w7(32'h37a9c42d),
	.w8(32'h3b41a8ad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f51f6),
	.w1(32'h3bd80590),
	.w2(32'h3c9598bf),
	.w3(32'h3bf6eb9a),
	.w4(32'h3b472742),
	.w5(32'h3c4b5c3a),
	.w6(32'h3bf251cf),
	.w7(32'h3b6aa94c),
	.w8(32'h3c1dd5da),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58b988),
	.w1(32'hbb8fe98e),
	.w2(32'h39937293),
	.w3(32'h3aa51934),
	.w4(32'h3b4603bf),
	.w5(32'h3b31c8db),
	.w6(32'h3a4e3c53),
	.w7(32'h3b056351),
	.w8(32'h3b1eab86),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a622797),
	.w1(32'hb9329259),
	.w2(32'h3af2efcb),
	.w3(32'hbaa160f2),
	.w4(32'hba9ff881),
	.w5(32'h3ac7160d),
	.w6(32'hb8e73b61),
	.w7(32'hb69d2e02),
	.w8(32'h3a4adce0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2950ce),
	.w1(32'h3b046376),
	.w2(32'h3ab7bbd4),
	.w3(32'h3a4b5c78),
	.w4(32'h386b8d23),
	.w5(32'h3a14bd67),
	.w6(32'h3aa0e6ae),
	.w7(32'h3995c802),
	.w8(32'h3a9ccc80),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b7e0f),
	.w1(32'hbb23a7dc),
	.w2(32'h3850297a),
	.w3(32'hba9b2fdf),
	.w4(32'hbabe11b8),
	.w5(32'h3ba938a3),
	.w6(32'hbae85a67),
	.w7(32'hb9bb89a1),
	.w8(32'h3bd03e3f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9038a6),
	.w1(32'h3aa509ca),
	.w2(32'h3baa3cc3),
	.w3(32'h3b1a7dc1),
	.w4(32'h3ad10899),
	.w5(32'h39a7792f),
	.w6(32'h3bc7df2f),
	.w7(32'h3b9d7a3d),
	.w8(32'h3b7b994d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82622d),
	.w1(32'h3b94143a),
	.w2(32'h3b18a444),
	.w3(32'h3a634f1e),
	.w4(32'hbaf27ed0),
	.w5(32'hbab83623),
	.w6(32'h3b5c8b85),
	.w7(32'h3a83f0b5),
	.w8(32'hb89018d2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c061ff6),
	.w1(32'h3a79174f),
	.w2(32'h3b39af6e),
	.w3(32'h3b9a8415),
	.w4(32'h3acf5c0b),
	.w5(32'h3bfe3548),
	.w6(32'h3b1b9f7f),
	.w7(32'h3ab33bbf),
	.w8(32'h3c1de39b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d6203),
	.w1(32'h3b99127d),
	.w2(32'h3bf90f1f),
	.w3(32'h3c04f1d9),
	.w4(32'h3b95de75),
	.w5(32'h3be611d3),
	.w6(32'h3c094861),
	.w7(32'h3c0b3860),
	.w8(32'h3c11f5d7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa84d1e),
	.w1(32'h3ad74bbf),
	.w2(32'h3b1348b6),
	.w3(32'h3b4c3492),
	.w4(32'h3b969fb6),
	.w5(32'h3a8417d2),
	.w6(32'h3ad0b58c),
	.w7(32'h3b2ef265),
	.w8(32'h3a069b93),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf020e),
	.w1(32'hb92a0b66),
	.w2(32'h3a3da188),
	.w3(32'h389d8784),
	.w4(32'h39a4f568),
	.w5(32'hb9abfdca),
	.w6(32'hb884c7f0),
	.w7(32'h3a3c4168),
	.w8(32'hba595214),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a4319),
	.w1(32'hbb14612a),
	.w2(32'h3a8e8abb),
	.w3(32'hbab159dd),
	.w4(32'h3b4b75b8),
	.w5(32'h39f6171d),
	.w6(32'hbb19d7f1),
	.w7(32'h3b0c4bb4),
	.w8(32'hba9821c4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb651172),
	.w1(32'hbb01fcb9),
	.w2(32'hba4b29aa),
	.w3(32'h3af9c05d),
	.w4(32'h3b5508e7),
	.w5(32'hbaffd8da),
	.w6(32'hba5c61d7),
	.w7(32'h39892a80),
	.w8(32'h3a2e1e0f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8d197),
	.w1(32'h3c094ab1),
	.w2(32'h3c3de53a),
	.w3(32'h3c0ea897),
	.w4(32'h3bffcdfc),
	.w5(32'h3bc50838),
	.w6(32'h3bcfef9b),
	.w7(32'h3c0759fd),
	.w8(32'h3c18a194),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c655e06),
	.w1(32'hbab0be75),
	.w2(32'h3c6f91a3),
	.w3(32'h3bead6ec),
	.w4(32'h39cdbd3a),
	.w5(32'h3c739f5a),
	.w6(32'h3c7158be),
	.w7(32'h3b28310f),
	.w8(32'h3c8a3ded),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a1370),
	.w1(32'hbbca60ed),
	.w2(32'h3c629d5a),
	.w3(32'h3c144be9),
	.w4(32'hbafeb24d),
	.w5(32'h3b800c0b),
	.w6(32'h3c8443f9),
	.w7(32'h3c0d82c0),
	.w8(32'h3c5ae0b7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac00d9),
	.w1(32'hbc3bb532),
	.w2(32'h3c87a353),
	.w3(32'h3c32a157),
	.w4(32'hbcc1b404),
	.w5(32'h3a2374fa),
	.w6(32'h3ce4ce4a),
	.w7(32'hbc223777),
	.w8(32'h3c8d715e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ad854),
	.w1(32'h3aa17951),
	.w2(32'h3abc4f75),
	.w3(32'h385f6bca),
	.w4(32'h3a950476),
	.w5(32'hbb804c98),
	.w6(32'h3ad49b6e),
	.w7(32'h3b1c05a2),
	.w8(32'hbb52368c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d556),
	.w1(32'hbb80f450),
	.w2(32'hbb61dba8),
	.w3(32'hbb58cde5),
	.w4(32'hbad99016),
	.w5(32'hbb0f22fb),
	.w6(32'hbb80f788),
	.w7(32'hbb2307ec),
	.w8(32'hbabb370d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76cc68),
	.w1(32'hbb2982fb),
	.w2(32'hbb3634b5),
	.w3(32'hb9d66668),
	.w4(32'h39eec30c),
	.w5(32'hba86a291),
	.w6(32'hba006fb1),
	.w7(32'hb91c15fd),
	.w8(32'hbae598b8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ba307),
	.w1(32'hbadbeed7),
	.w2(32'h3936671f),
	.w3(32'h3a012a59),
	.w4(32'hbb25d304),
	.w5(32'h395648ea),
	.w6(32'hb8b053d5),
	.w7(32'hbaab5178),
	.w8(32'h3a9d63d9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14b326),
	.w1(32'hbaa3f2cb),
	.w2(32'hba93c677),
	.w3(32'hba6dae34),
	.w4(32'h397f8b72),
	.w5(32'hbb45826d),
	.w6(32'hbaa324af),
	.w7(32'h3a335ef4),
	.w8(32'hbb6b5431),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b80624),
	.w1(32'hbb1138ba),
	.w2(32'hb9bcda37),
	.w3(32'h3a73d73e),
	.w4(32'h3a07caaf),
	.w5(32'h3b857ed5),
	.w6(32'hb9fe06bc),
	.w7(32'hbaa2574d),
	.w8(32'h3b6b549c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c590800),
	.w1(32'h3ba31c3f),
	.w2(32'h3c3a6e4b),
	.w3(32'h3c0bd7e2),
	.w4(32'h3a8bc128),
	.w5(32'h3b8a8ebd),
	.w6(32'h3c3660d2),
	.w7(32'h3bda2ee1),
	.w8(32'h3c42c77d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ce6d5),
	.w1(32'h3b487b75),
	.w2(32'h3c53ca1e),
	.w3(32'h3bd322e2),
	.w4(32'hbb77cc29),
	.w5(32'h3b736cfe),
	.w6(32'h3c16e62e),
	.w7(32'hba13ea9b),
	.w8(32'h3bc8af40),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8a209),
	.w1(32'hba006399),
	.w2(32'h3b8d8862),
	.w3(32'h3b480792),
	.w4(32'hbb60ee24),
	.w5(32'h3b971d8f),
	.w6(32'h3bca1505),
	.w7(32'hbaac29db),
	.w8(32'h3bca5984),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43153),
	.w1(32'hb8852f7f),
	.w2(32'h3babf72f),
	.w3(32'h3abe3f9e),
	.w4(32'h3aefe779),
	.w5(32'h3b17d698),
	.w6(32'hbb2a13d4),
	.w7(32'hbb3f581a),
	.w8(32'h3b31229c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0348c),
	.w1(32'hbab1e8b5),
	.w2(32'h3b43df8d),
	.w3(32'h3aaebeca),
	.w4(32'hbaf44e32),
	.w5(32'h3ad33aa3),
	.w6(32'h3b817d8c),
	.w7(32'hba87aded),
	.w8(32'h3b6db02d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a636460),
	.w1(32'h3a470053),
	.w2(32'h3bbeec90),
	.w3(32'h39e3aa8c),
	.w4(32'h3ac3a713),
	.w5(32'h3c0cb17e),
	.w6(32'h3ada7a38),
	.w7(32'h3a53d6e5),
	.w8(32'h3bed3a08),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6ec28),
	.w1(32'hbb431676),
	.w2(32'hb874bf8e),
	.w3(32'hbaf10ef1),
	.w4(32'hb79b9a8d),
	.w5(32'hb9bcb998),
	.w6(32'hbb61682e),
	.w7(32'hba331b9e),
	.w8(32'hbb5a4918),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85c962),
	.w1(32'hba40589a),
	.w2(32'h3a1d5785),
	.w3(32'h3b596a43),
	.w4(32'h3b92fe3d),
	.w5(32'hba570d8a),
	.w6(32'hb9f01f66),
	.w7(32'h3b05316a),
	.w8(32'hbaaac207),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66fe6),
	.w1(32'hbab1d9be),
	.w2(32'hba9b98ee),
	.w3(32'hba6d2990),
	.w4(32'hba8c215f),
	.w5(32'hbb4f17ef),
	.w6(32'hbaa58b6e),
	.w7(32'hbabb2149),
	.w8(32'hb9ac1755),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d4c5e),
	.w1(32'hbac8cfb5),
	.w2(32'hbae81084),
	.w3(32'hba9ec9ac),
	.w4(32'hbab67f9d),
	.w5(32'h39b02e5b),
	.w6(32'h3a82cbaf),
	.w7(32'h39092e7e),
	.w8(32'h3b1df88b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e89c4),
	.w1(32'hbb94b80c),
	.w2(32'hba9fd4a2),
	.w3(32'h3c1ecc22),
	.w4(32'hbba971bc),
	.w5(32'hbbffad15),
	.w6(32'h3c3b555b),
	.w7(32'hbb8b0c01),
	.w8(32'hbb770050),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb027d02),
	.w1(32'hbb29790a),
	.w2(32'hba604a7b),
	.w3(32'h3a3cb7f4),
	.w4(32'hb9f9ba8b),
	.w5(32'h3b910537),
	.w6(32'h3b00f26b),
	.w7(32'hba4ce01e),
	.w8(32'h3bb6d839),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61ca1c),
	.w1(32'h3c06deea),
	.w2(32'h3c7f96f9),
	.w3(32'h3c083310),
	.w4(32'h3b75ea84),
	.w5(32'h3b83725c),
	.w6(32'h3c4d37cb),
	.w7(32'h3ba76f8b),
	.w8(32'h3b77d684),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f36dd),
	.w1(32'hb99bdb50),
	.w2(32'h3bd3b7d5),
	.w3(32'h3c3b098a),
	.w4(32'h3b031e59),
	.w5(32'h3bd7d132),
	.w6(32'h3c84d38b),
	.w7(32'h3c009c7c),
	.w8(32'h3c133bae),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e6110f),
	.w1(32'hbc109157),
	.w2(32'hbb60fe5d),
	.w3(32'h3b84af36),
	.w4(32'hbbd98060),
	.w5(32'h394b3b2e),
	.w6(32'h3bd90277),
	.w7(32'hbbd0d320),
	.w8(32'h3b23d6ad),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cc235),
	.w1(32'h3bcac8bc),
	.w2(32'h3c2da4cc),
	.w3(32'h3bdd385c),
	.w4(32'hbb353e17),
	.w5(32'h3bcf82fb),
	.w6(32'h3b1e3bbc),
	.w7(32'h3b25ba12),
	.w8(32'h3c7a7bba),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addeb46),
	.w1(32'hbbb02881),
	.w2(32'h3c00c32e),
	.w3(32'h3ae0a7f9),
	.w4(32'hbb15782e),
	.w5(32'h3a332ef8),
	.w6(32'h3b8a6cf8),
	.w7(32'hbb038e7c),
	.w8(32'h3a214daa),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8df1ec),
	.w1(32'h3b94fe9e),
	.w2(32'h3c32b424),
	.w3(32'h3c3f9c13),
	.w4(32'hbad28157),
	.w5(32'h3a7aead7),
	.w6(32'h3c7c2a44),
	.w7(32'h3b161cc1),
	.w8(32'h3c17cbb5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb7bc7),
	.w1(32'hba91f1f4),
	.w2(32'h3b79c36c),
	.w3(32'h3b69105b),
	.w4(32'hbba9937b),
	.w5(32'hbbb861e8),
	.w6(32'h3b5315ee),
	.w7(32'hbb11bc89),
	.w8(32'h3ab1853f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd668d7),
	.w1(32'hbbfba751),
	.w2(32'h3b86e5af),
	.w3(32'h3ba49c22),
	.w4(32'hbc08e1bb),
	.w5(32'h3b209ad8),
	.w6(32'h3c38b26f),
	.w7(32'hbb9b1de3),
	.w8(32'h3b30287a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba447b20),
	.w1(32'hbaf486cc),
	.w2(32'hbb425218),
	.w3(32'hba3c30c9),
	.w4(32'hbac0850d),
	.w5(32'h3aade66a),
	.w6(32'hbae1f66f),
	.w7(32'hbb07d082),
	.w8(32'h3a4410c8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c447a60),
	.w1(32'h3ae0c385),
	.w2(32'h3c76f8e6),
	.w3(32'h3bc94560),
	.w4(32'hbb579b57),
	.w5(32'h3bf4f169),
	.w6(32'h3c403e5f),
	.w7(32'h3b912576),
	.w8(32'h3c7eea29),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb21bc5),
	.w1(32'h3b1b5552),
	.w2(32'h3c11bd36),
	.w3(32'h3be13641),
	.w4(32'hbb23744c),
	.w5(32'h3b0a6bd1),
	.w6(32'h3b338467),
	.w7(32'h3a212a31),
	.w8(32'h3c24302b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8064bf),
	.w1(32'h3a8360ee),
	.w2(32'h3c89dca8),
	.w3(32'hba9f4fed),
	.w4(32'hbbcc4ea8),
	.w5(32'h3bc95c20),
	.w6(32'h3b804768),
	.w7(32'hbbb0ec9d),
	.w8(32'h3c2592f8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb82d4),
	.w1(32'hbc7713b4),
	.w2(32'hbc521e4f),
	.w3(32'h3c8afbe0),
	.w4(32'hbcf16391),
	.w5(32'hbcb77818),
	.w6(32'h3ca9da72),
	.w7(32'hbc8b37e0),
	.w8(32'hbb68ada6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c377fde),
	.w1(32'h3b5e3f38),
	.w2(32'h3c95a245),
	.w3(32'h3b7a0b3f),
	.w4(32'hbc0a4f69),
	.w5(32'h3c2fafc3),
	.w6(32'h3c57fa30),
	.w7(32'h3a96862f),
	.w8(32'h3c45c3b6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22fb34),
	.w1(32'h3bb5ad78),
	.w2(32'h3c321c53),
	.w3(32'h3ba301d9),
	.w4(32'h3ac5c6dc),
	.w5(32'h3c03611d),
	.w6(32'hbb8b607c),
	.w7(32'hbb2fbe90),
	.w8(32'h3c4bcb3b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac4351),
	.w1(32'h3a420657),
	.w2(32'h399bbc23),
	.w3(32'hb9cd96bd),
	.w4(32'h39b7ccfd),
	.w5(32'hbb3d8f74),
	.w6(32'h3990b9e8),
	.w7(32'h3b0e7b57),
	.w8(32'hbb274258),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabead5),
	.w1(32'h3c2fc0aa),
	.w2(32'h3c7db5be),
	.w3(32'h3c088c23),
	.w4(32'hba9c125a),
	.w5(32'h3b91928e),
	.w6(32'h3ac9bb7a),
	.w7(32'hbc02cedc),
	.w8(32'h39d79de2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33b4b2),
	.w1(32'h3aa66305),
	.w2(32'h3b920129),
	.w3(32'h3ac21214),
	.w4(32'h3b2dbefa),
	.w5(32'h3b62daa4),
	.w6(32'h3a8f95f0),
	.w7(32'h3b582a0c),
	.w8(32'h3ba4fcf8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a004),
	.w1(32'hbb0d7eb5),
	.w2(32'hbafccf04),
	.w3(32'hbbc11f4a),
	.w4(32'hbbbdbf46),
	.w5(32'hbabc8980),
	.w6(32'hbb566792),
	.w7(32'hbb7c541f),
	.w8(32'hbb03e31c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa215e8),
	.w1(32'h3a0af883),
	.w2(32'h3b006128),
	.w3(32'hb9d936cd),
	.w4(32'hb94bec05),
	.w5(32'hba393ccb),
	.w6(32'h3b16738b),
	.w7(32'h3aea0896),
	.w8(32'hb9d055f0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb121b6),
	.w1(32'h3b5c0395),
	.w2(32'h3c1fe969),
	.w3(32'h3b71a119),
	.w4(32'h3b04a325),
	.w5(32'h3c369494),
	.w6(32'h3b928d3d),
	.w7(32'h3bfab3c8),
	.w8(32'h3c81cc1f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43a68),
	.w1(32'h3aa46fd0),
	.w2(32'h3c3edd5b),
	.w3(32'h3bb2ed0e),
	.w4(32'hb9189339),
	.w5(32'h3abce62d),
	.w6(32'h3c19bbc2),
	.w7(32'h3b8dac2d),
	.w8(32'h3ba16f2c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54132),
	.w1(32'hb99099e3),
	.w2(32'h3ad0e4d4),
	.w3(32'h3b9a6fa5),
	.w4(32'hbb9c0788),
	.w5(32'h3a6e3f12),
	.w6(32'h3c22740f),
	.w7(32'h3aa511b3),
	.w8(32'h3bc66409),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7e04d),
	.w1(32'h39b765b9),
	.w2(32'h3bb83555),
	.w3(32'h3ba823b8),
	.w4(32'hbaf0f216),
	.w5(32'h3b8aa282),
	.w6(32'h3b972392),
	.w7(32'h39f9ee54),
	.w8(32'h3c133329),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc40243),
	.w1(32'hbb054470),
	.w2(32'h3b4cfb87),
	.w3(32'h3b41d490),
	.w4(32'hbb67d4ad),
	.w5(32'h3aa53e0d),
	.w6(32'h3c33fe90),
	.w7(32'h3ac3f415),
	.w8(32'h3bd3dae1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0519d1),
	.w1(32'h3b35acc1),
	.w2(32'h3be1be11),
	.w3(32'h3b80de72),
	.w4(32'hbb23e8c9),
	.w5(32'hbaf96b95),
	.w6(32'h3b6ccd4e),
	.w7(32'h3a07b545),
	.w8(32'h3bd9f813),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce7e3),
	.w1(32'hb8aa25b0),
	.w2(32'h3b4859aa),
	.w3(32'h3b20790f),
	.w4(32'hbb189672),
	.w5(32'h3b030d75),
	.w6(32'h3bdd35a2),
	.w7(32'h3a875d42),
	.w8(32'h3b931e72),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba954516),
	.w1(32'h3ab87413),
	.w2(32'h3a855f11),
	.w3(32'h3911fed0),
	.w4(32'hba38f106),
	.w5(32'h3a5b2252),
	.w6(32'hba74926e),
	.w7(32'h3a4cc432),
	.w8(32'hb9e41c2f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a9edc),
	.w1(32'h3a53d5d2),
	.w2(32'h3a8265ae),
	.w3(32'h3a4c3763),
	.w4(32'h3a54429c),
	.w5(32'hb91c0411),
	.w6(32'h398b6909),
	.w7(32'h3a1e0a05),
	.w8(32'h3aaeabcc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beb81a),
	.w1(32'hba532f5f),
	.w2(32'hba6a6a3d),
	.w3(32'hb906a290),
	.w4(32'hba347b89),
	.w5(32'h3b1cb19d),
	.w6(32'h3b1f891b),
	.w7(32'hbad7f999),
	.w8(32'h3acc06db),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32849e),
	.w1(32'h3aa8196a),
	.w2(32'h3afe89d8),
	.w3(32'h3aacab00),
	.w4(32'h3a8824b5),
	.w5(32'hbb9f5764),
	.w6(32'h3ab49a87),
	.w7(32'h3a1943a8),
	.w8(32'hbb9dba28),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b437754),
	.w1(32'hbbe155a0),
	.w2(32'h3b1934c8),
	.w3(32'hbb0c7262),
	.w4(32'hbc285654),
	.w5(32'h3b242739),
	.w6(32'h3b429a29),
	.w7(32'hbb976215),
	.w8(32'h3be09909),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb57b0),
	.w1(32'h3af2be85),
	.w2(32'h3b7b3e99),
	.w3(32'h3b27dcb3),
	.w4(32'h3b2cdaf7),
	.w5(32'hb8e97fc3),
	.w6(32'hb9c49473),
	.w7(32'h3b29be0d),
	.w8(32'h390f7274),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adf765),
	.w1(32'h37c82523),
	.w2(32'h3b9a02ce),
	.w3(32'h39768ac3),
	.w4(32'hb9c29443),
	.w5(32'h3bde4d77),
	.w6(32'hbb216798),
	.w7(32'h385ed457),
	.w8(32'h3bcbe70b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c851a),
	.w1(32'h3b4de055),
	.w2(32'h3c1783b4),
	.w3(32'h3c655777),
	.w4(32'hbb2f16f3),
	.w5(32'hb99abd57),
	.w6(32'h3c8f4ef1),
	.w7(32'h3b4ec9b1),
	.w8(32'h3bc8d3dc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba807cdb),
	.w1(32'hbaabcc14),
	.w2(32'hbb164427),
	.w3(32'hba1c543c),
	.w4(32'h38a5e65d),
	.w5(32'h3af8f248),
	.w6(32'hba238e0e),
	.w7(32'hba8d20ff),
	.w8(32'h39b71711),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b843),
	.w1(32'h3b6ff95d),
	.w2(32'h3b8a7429),
	.w3(32'h3b14513f),
	.w4(32'hb93f3203),
	.w5(32'hba197cc0),
	.w6(32'h3a6aa9bc),
	.w7(32'h3a12291d),
	.w8(32'h39002d34),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be16b4),
	.w1(32'hba1172fc),
	.w2(32'h3a4172ed),
	.w3(32'h3aa36fd0),
	.w4(32'h3b114ae2),
	.w5(32'hb9c83a21),
	.w6(32'h3aa782a4),
	.w7(32'h3af85786),
	.w8(32'h39f5ff58),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6e15e),
	.w1(32'h3a9497ab),
	.w2(32'h3a9d966c),
	.w3(32'h3a98afb0),
	.w4(32'h3a8c9a97),
	.w5(32'hba666acc),
	.w6(32'h3b78f55c),
	.w7(32'h3b49fd3a),
	.w8(32'h3ad4f439),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be70cd5),
	.w1(32'h3c178c4d),
	.w2(32'h3be13582),
	.w3(32'hbb1e12d5),
	.w4(32'h3be76e57),
	.w5(32'h3c80a352),
	.w6(32'h3b83f819),
	.w7(32'h3be29013),
	.w8(32'h3c3e86e6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c144a9f),
	.w1(32'h3b514d29),
	.w2(32'h3c6f726e),
	.w3(32'h3b5fb9b1),
	.w4(32'h3ac48da7),
	.w5(32'h3c47c000),
	.w6(32'h3b92ebe8),
	.w7(32'h3bd68448),
	.w8(32'h3c46a6ce),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1bbd4),
	.w1(32'h3a9ef566),
	.w2(32'h3a87d102),
	.w3(32'h3aca2c5d),
	.w4(32'h3ac797ef),
	.w5(32'hbaf4e2dc),
	.w6(32'h3ab2347f),
	.w7(32'hb9c8e8cd),
	.w8(32'hbaa529e1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4db77f),
	.w1(32'h3b0bbfa4),
	.w2(32'h3b926b45),
	.w3(32'h3b3154b8),
	.w4(32'hba02d3e5),
	.w5(32'h3afd2b05),
	.w6(32'h3b898b3b),
	.w7(32'h3aa6861f),
	.w8(32'h3ba22dce),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6676ac),
	.w1(32'hba9ce7d1),
	.w2(32'h3ae48163),
	.w3(32'h3b51ce89),
	.w4(32'hba8b3484),
	.w5(32'h387088c2),
	.w6(32'h3b13806d),
	.w7(32'hbb1e0cc5),
	.w8(32'h3b310abe),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad77b4),
	.w1(32'h39132250),
	.w2(32'h3b0b2d59),
	.w3(32'h3a9e1175),
	.w4(32'hbb4228d0),
	.w5(32'h3b2373dd),
	.w6(32'h3baa8b5d),
	.w7(32'h3a96dd04),
	.w8(32'h3b9ca3a7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c186fbc),
	.w1(32'h3b9b9a41),
	.w2(32'h3c3d4a07),
	.w3(32'h3b8712e6),
	.w4(32'hbb087111),
	.w5(32'h3a222d37),
	.w6(32'h3bc00fa5),
	.w7(32'h3aad966b),
	.w8(32'h3b05c24b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0077f),
	.w1(32'h3b702e4b),
	.w2(32'h3c4565cb),
	.w3(32'h3ba313f6),
	.w4(32'h3b5bbe79),
	.w5(32'h3c2720af),
	.w6(32'h3baa8392),
	.w7(32'h3b6b3c04),
	.w8(32'h3c482f99),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2985e),
	.w1(32'hba36479e),
	.w2(32'h3bc0613e),
	.w3(32'h3b5a392c),
	.w4(32'hbbdd6c3a),
	.w5(32'h3adcf233),
	.w6(32'h3bb67b31),
	.w7(32'hbb38bb72),
	.w8(32'h3bd80a76),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35a87b),
	.w1(32'h3bc07d60),
	.w2(32'h3bf3fcf6),
	.w3(32'h3ba42fe1),
	.w4(32'hba54bb0c),
	.w5(32'h3b5a6f39),
	.w6(32'h3b8bfffb),
	.w7(32'h3b237735),
	.w8(32'h3c04b933),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cde97),
	.w1(32'h3bc3ecc9),
	.w2(32'h3c5fb24d),
	.w3(32'h3c01c4f1),
	.w4(32'h3b934f61),
	.w5(32'h3c2f5be8),
	.w6(32'h3c00e768),
	.w7(32'h3b9125de),
	.w8(32'h3c1f2d52),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24d26f),
	.w1(32'h3b01ba02),
	.w2(32'h3b85b7d4),
	.w3(32'h3bb09a83),
	.w4(32'hbafc7263),
	.w5(32'hbac3378a),
	.w6(32'h3c26fda3),
	.w7(32'h3af0c44f),
	.w8(32'h3ae6e738),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74e39f),
	.w1(32'h3abddece),
	.w2(32'h3bbf761d),
	.w3(32'h3a8af359),
	.w4(32'hbb764b9f),
	.w5(32'h3a15b2b8),
	.w6(32'h3a632512),
	.w7(32'hba40c0fc),
	.w8(32'h3bad368f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8fc7),
	.w1(32'hbaf03570),
	.w2(32'h3a61d157),
	.w3(32'hbb0c8996),
	.w4(32'hbb648297),
	.w5(32'h39ddd412),
	.w6(32'h3a74acd1),
	.w7(32'hba9e0c13),
	.w8(32'h3a4ffd65),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c198c15),
	.w1(32'hbc474a43),
	.w2(32'h3acb402a),
	.w3(32'h3c4edba9),
	.w4(32'hbbd57d7f),
	.w5(32'h3b61e7f6),
	.w6(32'h3c71c578),
	.w7(32'hbb885aaa),
	.w8(32'h3c0f2b27),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c052243),
	.w1(32'hbb3459e6),
	.w2(32'hbba534fe),
	.w3(32'h3ba1ccae),
	.w4(32'hbba4de0b),
	.w5(32'hbbc867d7),
	.w6(32'h3be75103),
	.w7(32'hbb843e16),
	.w8(32'hba9f91c8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ed174),
	.w1(32'h3a1a0070),
	.w2(32'h38f52a2c),
	.w3(32'h38831663),
	.w4(32'h3a29ba67),
	.w5(32'hba0b5311),
	.w6(32'h3abad5be),
	.w7(32'h3a87af12),
	.w8(32'hba89bdac),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77aea70),
	.w1(32'h39069680),
	.w2(32'h3aad4f54),
	.w3(32'hba43cc63),
	.w4(32'h3acd882d),
	.w5(32'h3922f826),
	.w6(32'hb8fa86cf),
	.w7(32'h3a986a5c),
	.w8(32'h3ad55108),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b779a80),
	.w1(32'h3abf9d24),
	.w2(32'h3ad73f1f),
	.w3(32'h3b4fa481),
	.w4(32'hba21cccc),
	.w5(32'h379b5101),
	.w6(32'h3b6c74a6),
	.w7(32'hb99d85bb),
	.w8(32'h3ba5be60),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48a012),
	.w1(32'hbaca8ff0),
	.w2(32'h3ae116ed),
	.w3(32'h3b58c636),
	.w4(32'hbc2506a7),
	.w5(32'hbba48eab),
	.w6(32'h3c00bb3a),
	.w7(32'hbbcedef7),
	.w8(32'h3a083308),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2159f7),
	.w1(32'h3af50a33),
	.w2(32'h3c635e1e),
	.w3(32'h3c41c8c7),
	.w4(32'h3ac9b838),
	.w5(32'h3c1dc487),
	.w6(32'h3c40211d),
	.w7(32'h3b92ac79),
	.w8(32'h3c262280),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8999f3),
	.w1(32'hbac5007c),
	.w2(32'hba65eca1),
	.w3(32'hbab622a9),
	.w4(32'hb7e1ac64),
	.w5(32'h3aca40fb),
	.w6(32'hba0b7d8e),
	.w7(32'hb96f876d),
	.w8(32'h395daf0a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf12ce6),
	.w1(32'h3b09d9df),
	.w2(32'h3c5917c6),
	.w3(32'h3bd4531d),
	.w4(32'h3ae69865),
	.w5(32'h3c24766a),
	.w6(32'h3c11afb3),
	.w7(32'h3b897f0a),
	.w8(32'h3c2f0ea4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba806de),
	.w1(32'h3abff2eb),
	.w2(32'h3bf3cf41),
	.w3(32'h3aec24b3),
	.w4(32'hbb2bcdbe),
	.w5(32'h3b138ef0),
	.w6(32'h3b69fd3b),
	.w7(32'hb9909e2e),
	.w8(32'h3ba2078e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236701),
	.w1(32'h3bc90e0c),
	.w2(32'h3c2eaa6f),
	.w3(32'h3b7da1d5),
	.w4(32'h38bafce5),
	.w5(32'h3c1eac78),
	.w6(32'hbad12adb),
	.w7(32'hba49038a),
	.w8(32'h3c2ba719),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc554c),
	.w1(32'hbc10d910),
	.w2(32'h3c104426),
	.w3(32'h3b164f9f),
	.w4(32'hbc61febb),
	.w5(32'h3a97212f),
	.w6(32'h3c05ad3c),
	.w7(32'hbbd6b8d5),
	.w8(32'h3b811eaf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb13cf6),
	.w1(32'hba06b597),
	.w2(32'hba3bbec5),
	.w3(32'h3b57bef8),
	.w4(32'hbab78308),
	.w5(32'hbb75645d),
	.w6(32'h3bf5333d),
	.w7(32'hba4db2bf),
	.w8(32'hbb081ff2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c379d),
	.w1(32'h3a89bf0f),
	.w2(32'hba3766c7),
	.w3(32'hbb31387b),
	.w4(32'hbb2655b1),
	.w5(32'h3a96b30a),
	.w6(32'hbb003435),
	.w7(32'hbb06be66),
	.w8(32'hb7fcdc3c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb7f8e),
	.w1(32'hbb4b791f),
	.w2(32'h3aff67e4),
	.w3(32'h3b263875),
	.w4(32'hbba243f8),
	.w5(32'hbb59380d),
	.w6(32'h3c19bed9),
	.w7(32'h3abc69b7),
	.w8(32'h3ab7df28),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bd70e),
	.w1(32'hbba3e53f),
	.w2(32'hbb23cae2),
	.w3(32'h3c0133a4),
	.w4(32'hbc04b1c2),
	.w5(32'hbb964254),
	.w6(32'h3c24669c),
	.w7(32'hbb928823),
	.w8(32'h3af054e5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace87b8),
	.w1(32'hbc10e93e),
	.w2(32'hbacd2165),
	.w3(32'h3a892702),
	.w4(32'hbc02330d),
	.w5(32'hbaa51e83),
	.w6(32'h3b9d0878),
	.w7(32'hbbaeea10),
	.w8(32'h3ac1992b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0107),
	.w1(32'h3b1d69e7),
	.w2(32'h3a6233a7),
	.w3(32'h3b019e69),
	.w4(32'h3ac9812e),
	.w5(32'h3aba3962),
	.w6(32'h3b53e201),
	.w7(32'h3afc687f),
	.w8(32'h3b71f0b7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b845525),
	.w1(32'h3b8cb4b6),
	.w2(32'h3b375732),
	.w3(32'h3ad350d4),
	.w4(32'h393cf0e7),
	.w5(32'h39bfd894),
	.w6(32'h3afa4460),
	.w7(32'h3a8c6cf2),
	.w8(32'h3acaf51a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c218fd0),
	.w1(32'h3b34b653),
	.w2(32'h3bc18764),
	.w3(32'h3b99a995),
	.w4(32'hbafc2969),
	.w5(32'h3bb5c0e3),
	.w6(32'h3b970f71),
	.w7(32'h39bf1db0),
	.w8(32'h3bd27af6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a14ec),
	.w1(32'hbac04a5c),
	.w2(32'h38f8571c),
	.w3(32'hbac8bf24),
	.w4(32'hba803f22),
	.w5(32'h3afc58f6),
	.w6(32'hbafb07c1),
	.w7(32'hbad9adaf),
	.w8(32'h3a27cd04),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b922121),
	.w1(32'hbb49dec0),
	.w2(32'h3b8922d7),
	.w3(32'h3ae8539e),
	.w4(32'hbb429a70),
	.w5(32'h3a436b58),
	.w6(32'h3b9086fd),
	.w7(32'hbac9e686),
	.w8(32'hba519318),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c184),
	.w1(32'hbb206419),
	.w2(32'hba5373e6),
	.w3(32'hbb6ccab2),
	.w4(32'hbb680ef9),
	.w5(32'h3a3f7d38),
	.w6(32'hbb4ec8e6),
	.w7(32'hbb341bb1),
	.w8(32'hb9c694a1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b161050),
	.w1(32'h39ca510f),
	.w2(32'h3bd468c5),
	.w3(32'h3b3a7465),
	.w4(32'h3b12565b),
	.w5(32'h3c2ab8cd),
	.w6(32'h3ba7f2b5),
	.w7(32'h3b8030e2),
	.w8(32'h3c5ad82d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c052f),
	.w1(32'h3b63ae98),
	.w2(32'h3b821137),
	.w3(32'h38339bf4),
	.w4(32'h3aa66d29),
	.w5(32'h3aea5872),
	.w6(32'h3b0af775),
	.w7(32'h3b518a79),
	.w8(32'h3a197a7c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996c8f),
	.w1(32'h3af38947),
	.w2(32'h3a8993de),
	.w3(32'h3b72b87a),
	.w4(32'h3b22596b),
	.w5(32'h3a2d43a8),
	.w6(32'h3ac069a1),
	.w7(32'h393764c6),
	.w8(32'hb9c174bb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdadca2),
	.w1(32'hbb76225f),
	.w2(32'h3a694f58),
	.w3(32'h3bcb9d4b),
	.w4(32'hbaf765ee),
	.w5(32'hbac21cc5),
	.w6(32'h3c01e89e),
	.w7(32'h3aa4d130),
	.w8(32'h3b210444),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d347b),
	.w1(32'hbac527f9),
	.w2(32'h3c0b6840),
	.w3(32'h3bd4f71a),
	.w4(32'h3a0b616c),
	.w5(32'h3c8742a2),
	.w6(32'h3c231c9b),
	.w7(32'hb9302519),
	.w8(32'h3c914062),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55b17),
	.w1(32'hbb4fce64),
	.w2(32'h3a96f8e0),
	.w3(32'h3ad3309c),
	.w4(32'hbaec6447),
	.w5(32'h3b80cd64),
	.w6(32'h3ba99a84),
	.w7(32'hba13b121),
	.w8(32'h3bf7eb9d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c20d0),
	.w1(32'h3bc050b9),
	.w2(32'h3c66026c),
	.w3(32'h3bbef188),
	.w4(32'hb79b228b),
	.w5(32'h3b4ff33f),
	.w6(32'h3c49177c),
	.w7(32'h3b6eda6a),
	.w8(32'h3ba911db),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bb2c7),
	.w1(32'hbb622f0b),
	.w2(32'hb8f9ef01),
	.w3(32'hbb585cdd),
	.w4(32'hbb82e43d),
	.w5(32'h3af43096),
	.w6(32'hbb849b15),
	.w7(32'hbb8d84b3),
	.w8(32'h3aa740d4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c958d4a),
	.w1(32'h3a87e10d),
	.w2(32'h3c8ec79e),
	.w3(32'h3c3cc385),
	.w4(32'hbbb13bb5),
	.w5(32'h3c22e951),
	.w6(32'h3c49f837),
	.w7(32'h3b915a47),
	.w8(32'h3c677d5e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9880e),
	.w1(32'h3921094f),
	.w2(32'h3c1a31dc),
	.w3(32'h3bbd04a8),
	.w4(32'hbb31d50c),
	.w5(32'hba6cd812),
	.w6(32'h3c29b448),
	.w7(32'h3a6939bd),
	.w8(32'h3b4e9ea1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43c25c),
	.w1(32'hba06f688),
	.w2(32'h3c2483b7),
	.w3(32'hbb658892),
	.w4(32'hbba6e181),
	.w5(32'h3c489604),
	.w6(32'h3a8eb042),
	.w7(32'hbaf00471),
	.w8(32'h3c512c95),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cef7b),
	.w1(32'h3b136181),
	.w2(32'h3acc0647),
	.w3(32'h3b6d02bc),
	.w4(32'h3b2b9915),
	.w5(32'hbb6b8508),
	.w6(32'h3b05a8ff),
	.w7(32'h3b01c7bb),
	.w8(32'hbb5b7149),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2379c2),
	.w1(32'h3917dc71),
	.w2(32'h3b445262),
	.w3(32'hb9a42c13),
	.w4(32'hbb2a1636),
	.w5(32'h3b8cc47f),
	.w6(32'hb853f234),
	.w7(32'hbb2a7d76),
	.w8(32'h3b896b5f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f3f3a),
	.w1(32'h3b124702),
	.w2(32'h3b0da0e7),
	.w3(32'h3af56f62),
	.w4(32'h3b0bfa43),
	.w5(32'hba45f286),
	.w6(32'h3aa8730c),
	.w7(32'h3ad20e08),
	.w8(32'h3adcaba6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215e56),
	.w1(32'h3b283a30),
	.w2(32'h3b778a52),
	.w3(32'hb959564d),
	.w4(32'hbb0c900b),
	.w5(32'h3b0585c9),
	.w6(32'h3a4ea01c),
	.w7(32'h3a55d4d6),
	.w8(32'h3bc1d99d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bcf5e),
	.w1(32'hba311720),
	.w2(32'h3ac4a888),
	.w3(32'h3b1120e1),
	.w4(32'h39c286b1),
	.w5(32'h3af410ba),
	.w6(32'h3b71edf6),
	.w7(32'hba08dc42),
	.w8(32'h3a8c8547),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7a9be),
	.w1(32'h3a97c36b),
	.w2(32'h3c07da76),
	.w3(32'h3c153657),
	.w4(32'hb9841dad),
	.w5(32'h39963d0a),
	.w6(32'h3c0365b4),
	.w7(32'h3b439bac),
	.w8(32'h3bba6853),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cc164),
	.w1(32'hbbbb9811),
	.w2(32'hbb751d39),
	.w3(32'hbb87ab41),
	.w4(32'hbb837333),
	.w5(32'hbab7c458),
	.w6(32'hbb7a1dad),
	.w7(32'hbb2f3252),
	.w8(32'hb86d7742),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95453c0),
	.w1(32'hba965f62),
	.w2(32'hbaa462f6),
	.w3(32'h38b9fd4e),
	.w4(32'h3aa5537e),
	.w5(32'hba8df8cd),
	.w6(32'h3a58564c),
	.w7(32'h3a02a993),
	.w8(32'h3a15ce0d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f17b5),
	.w1(32'hbb27c4bc),
	.w2(32'hba007a5e),
	.w3(32'h3a75a6ce),
	.w4(32'hbb8f298e),
	.w5(32'hbacc34a8),
	.w6(32'h3b9cd00b),
	.w7(32'h386879bd),
	.w8(32'hb981bc65),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce1bbd),
	.w1(32'hba05ce4b),
	.w2(32'h3b42cc81),
	.w3(32'h3bd0bc14),
	.w4(32'hbb2b7067),
	.w5(32'hb8ab150e),
	.w6(32'h3bf88a4a),
	.w7(32'h3b1252cf),
	.w8(32'h3bbbd3a4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e016b),
	.w1(32'hbb486d61),
	.w2(32'h3a1bd835),
	.w3(32'h3a7c70b4),
	.w4(32'hba2bae4c),
	.w5(32'h3b9559df),
	.w6(32'hbb8325cd),
	.w7(32'hbb8bba42),
	.w8(32'h3ba78e97),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89e1c4),
	.w1(32'h3b515acb),
	.w2(32'h3b69a90a),
	.w3(32'h3b86135e),
	.w4(32'h3b410d4a),
	.w5(32'h3b34b2b3),
	.w6(32'h3b91c156),
	.w7(32'h3b44c27a),
	.w8(32'h3b0d48e6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9e5c1),
	.w1(32'h3c4bdf61),
	.w2(32'h3d0b31e7),
	.w3(32'h3c2a395d),
	.w4(32'h3bf5a53d),
	.w5(32'h3cd359d8),
	.w6(32'h3a1a4412),
	.w7(32'h3c3c1243),
	.w8(32'h3cbc6a5f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba0579),
	.w1(32'h3b399d5a),
	.w2(32'h3c4b55a6),
	.w3(32'h3c9acc8b),
	.w4(32'hbbaf705a),
	.w5(32'h38bf4806),
	.w6(32'h3c80e16e),
	.w7(32'hbb8ffe10),
	.w8(32'h3b924d78),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c08a8),
	.w1(32'h3a95d52b),
	.w2(32'h3aa929c9),
	.w3(32'hba8a9951),
	.w4(32'h3acbbc96),
	.w5(32'h3b69403d),
	.w6(32'hb9ce7063),
	.w7(32'h3a8a0661),
	.w8(32'h3baa6bd8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b33aa9),
	.w1(32'h39db6ee4),
	.w2(32'h3a95a854),
	.w3(32'h3a136cb7),
	.w4(32'h39d50139),
	.w5(32'hba5cee25),
	.w6(32'h3b50ec11),
	.w7(32'h3afe5cba),
	.w8(32'hbac83205),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc8f77),
	.w1(32'hbb161803),
	.w2(32'hba81adc0),
	.w3(32'hbb22be3f),
	.w4(32'hba769b5e),
	.w5(32'hbb14c5a9),
	.w6(32'hbafaa688),
	.w7(32'hba21f80b),
	.w8(32'hbace8cda),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae99cfa),
	.w1(32'hbb4aa26c),
	.w2(32'hbaf57a7e),
	.w3(32'hbad92074),
	.w4(32'h3960be6c),
	.w5(32'h3ae4b420),
	.w6(32'hbaaae014),
	.w7(32'hba1f20ad),
	.w8(32'h3b0a2dfe),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adbe32),
	.w1(32'h3b4252fe),
	.w2(32'h3ba6317c),
	.w3(32'h39da861a),
	.w4(32'h3b4186ea),
	.w5(32'h3b7662cc),
	.w6(32'h3a7eaaab),
	.w7(32'h3b3bf2df),
	.w8(32'h3b89fa29),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30758a),
	.w1(32'h3b36fc46),
	.w2(32'h3baa9a97),
	.w3(32'h3bbb513c),
	.w4(32'hbb64c5de),
	.w5(32'h3b5d64c7),
	.w6(32'h3bd9c91b),
	.w7(32'hba798787),
	.w8(32'h3bf22067),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86b5fe),
	.w1(32'h3b9f69b3),
	.w2(32'h3c37b2a0),
	.w3(32'h3c331701),
	.w4(32'hbba0520d),
	.w5(32'h3b43b548),
	.w6(32'h3c58aaec),
	.w7(32'hbb4ef2db),
	.w8(32'h3ba10d5b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf00f8),
	.w1(32'hb964659e),
	.w2(32'h3a09ca56),
	.w3(32'h3abb4582),
	.w4(32'hbb085329),
	.w5(32'hbb79a161),
	.w6(32'h3b7c0806),
	.w7(32'h3ab94c1f),
	.w8(32'hbaa6e18a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc87870),
	.w1(32'h3b9606cf),
	.w2(32'h3c5d5082),
	.w3(32'hba546b10),
	.w4(32'hbb95b676),
	.w5(32'h3c4e1e71),
	.w6(32'h3be12c2e),
	.w7(32'h3b4cf7b1),
	.w8(32'h3c846d47),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157bf8),
	.w1(32'h3b09dce2),
	.w2(32'h3b039328),
	.w3(32'h3aa6e3e2),
	.w4(32'h3a92367a),
	.w5(32'h3b554e4f),
	.w6(32'h3b41a699),
	.w7(32'h3b206e37),
	.w8(32'h3b191c1c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39283384),
	.w1(32'h3a810b47),
	.w2(32'h3ab2c0f9),
	.w3(32'h3b00de31),
	.w4(32'h3aa196e1),
	.w5(32'h39972f65),
	.w6(32'h3b03a957),
	.w7(32'h3aac0d18),
	.w8(32'h3a2803a1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84d758),
	.w1(32'h3abe542a),
	.w2(32'hb9178c36),
	.w3(32'h3b3f6a38),
	.w4(32'h3b241567),
	.w5(32'hbb46417a),
	.w6(32'h3b7019e1),
	.w7(32'h3b702179),
	.w8(32'hbb031dc0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cd6ae),
	.w1(32'hbafceddc),
	.w2(32'hb9a8ef6b),
	.w3(32'hbabe4dd7),
	.w4(32'hba975d68),
	.w5(32'h3a392404),
	.w6(32'h3a673232),
	.w7(32'h3a0d9546),
	.w8(32'h3aae3694),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c256057),
	.w1(32'h3aae0f34),
	.w2(32'h3b981410),
	.w3(32'h3bcadde8),
	.w4(32'hbaf599e3),
	.w5(32'hbaf7d6b9),
	.w6(32'h3c144d92),
	.w7(32'h3badeee9),
	.w8(32'h3b748eba),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28784e),
	.w1(32'hbbcea22f),
	.w2(32'h3a2c45d5),
	.w3(32'h3bb56636),
	.w4(32'hbc22ea64),
	.w5(32'hba967794),
	.w6(32'h3c7edb28),
	.w7(32'hbb14a58e),
	.w8(32'h3bdd7d17),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c036b1f),
	.w1(32'hb9efd966),
	.w2(32'h3be18638),
	.w3(32'h3bbf1b7a),
	.w4(32'hbb9bea93),
	.w5(32'h3b31085f),
	.w6(32'h3c2429a0),
	.w7(32'h3a438f37),
	.w8(32'h3c1a4195),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b203985),
	.w1(32'hbae5efd8),
	.w2(32'hbad469c2),
	.w3(32'hb91439e2),
	.w4(32'hbaad9981),
	.w5(32'hba6d04ab),
	.w6(32'h3ad025f5),
	.w7(32'h38e26b66),
	.w8(32'h3a9cad16),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b4e2f),
	.w1(32'h3b02b29f),
	.w2(32'h3c243a03),
	.w3(32'h3bce2ac1),
	.w4(32'hbbb6ceec),
	.w5(32'hba52822a),
	.w6(32'h3c44b384),
	.w7(32'h3a7a7c07),
	.w8(32'h3bc59fe3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc965b2),
	.w1(32'h3b2de9f4),
	.w2(32'h3be3a3d4),
	.w3(32'h3b704ecc),
	.w4(32'h3a58f9d3),
	.w5(32'h3ba7f04f),
	.w6(32'h3ba28eec),
	.w7(32'h3b65032e),
	.w8(32'h3bb878b1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c810a53),
	.w1(32'h3b7d6764),
	.w2(32'h3c7e351f),
	.w3(32'h3c747b76),
	.w4(32'hbb3ce340),
	.w5(32'h3c1a17fb),
	.w6(32'h3c5997b0),
	.w7(32'h3ad67858),
	.w8(32'h3c808cdf),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f91c7),
	.w1(32'h3a36bc89),
	.w2(32'h39e69d94),
	.w3(32'h38e01fe8),
	.w4(32'hb98e3cc6),
	.w5(32'hba627448),
	.w6(32'h3af3d1ab),
	.w7(32'h3a78b2fe),
	.w8(32'hbae853a5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a11d7c),
	.w1(32'h3a577721),
	.w2(32'h3b6a158f),
	.w3(32'hba357b15),
	.w4(32'hba44c562),
	.w5(32'h3b17534a),
	.w6(32'hbb428d56),
	.w7(32'h3aa74ee5),
	.w8(32'h3ad2084f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69e6eb),
	.w1(32'h3b28814c),
	.w2(32'h3c38fe1c),
	.w3(32'h3c0a92e8),
	.w4(32'h3ab4499c),
	.w5(32'h3bedeffb),
	.w6(32'h3c6015e3),
	.w7(32'h3ba6d5db),
	.w8(32'h3c348dc3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fac99),
	.w1(32'hbb948376),
	.w2(32'h3c3c08bf),
	.w3(32'h3b87b565),
	.w4(32'hbb93b8d6),
	.w5(32'h3c434eb4),
	.w6(32'h3bfedd95),
	.w7(32'hba9f73e8),
	.w8(32'h3c047aed),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f0427),
	.w1(32'h39787164),
	.w2(32'h3c150ab0),
	.w3(32'h3b5825a2),
	.w4(32'hbbfa0e90),
	.w5(32'hb908e61e),
	.w6(32'h3c222e50),
	.w7(32'hbab6528f),
	.w8(32'h3badc54a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22ea54),
	.w1(32'h39e9a71b),
	.w2(32'h392db974),
	.w3(32'h3a648f2d),
	.w4(32'h3b36f01b),
	.w5(32'h3b5a1738),
	.w6(32'hbc11d08e),
	.w7(32'hbb018fb4),
	.w8(32'h3bb95a81),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925a4ce),
	.w1(32'h3945ec8e),
	.w2(32'h3aef747b),
	.w3(32'h3aa61df5),
	.w4(32'h3add178d),
	.w5(32'h39f319ed),
	.w6(32'h3ac06976),
	.w7(32'h3ae1ccd7),
	.w8(32'h39a722b1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b607f8b),
	.w1(32'h3b250e3c),
	.w2(32'h3aa085c9),
	.w3(32'h3a713ec5),
	.w4(32'h3b0e72cb),
	.w5(32'hbb28956f),
	.w6(32'h3a9a0897),
	.w7(32'h3a9ed699),
	.w8(32'hbac9ebc9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb366955),
	.w1(32'h3af2d4e3),
	.w2(32'h3c2c7770),
	.w3(32'hb9c61822),
	.w4(32'h3c352c04),
	.w5(32'h3c710905),
	.w6(32'hbaa7744b),
	.w7(32'h3b7353d5),
	.w8(32'h3c0ddcb0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f45b6),
	.w1(32'h3ba736be),
	.w2(32'h3c8bfb0e),
	.w3(32'h3c2c76d9),
	.w4(32'h3b062d71),
	.w5(32'h3c66d859),
	.w6(32'h3c0207e0),
	.w7(32'h3bfac520),
	.w8(32'h3c975818),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0110c5),
	.w1(32'h3b1357ea),
	.w2(32'h3b565435),
	.w3(32'h3b15757f),
	.w4(32'h3b9a98ee),
	.w5(32'h3ac0df44),
	.w6(32'h3ac427f1),
	.w7(32'h3ac5e497),
	.w8(32'h3b9fecd5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba88093),
	.w1(32'hbbd12b16),
	.w2(32'hbb597597),
	.w3(32'h3b7bad04),
	.w4(32'hbc2da1a0),
	.w5(32'hba7faabe),
	.w6(32'h3c3f09e5),
	.w7(32'hbb9f525c),
	.w8(32'h3b73a863),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c682126),
	.w1(32'h3b5dca87),
	.w2(32'h3c33c34d),
	.w3(32'h3c3aad43),
	.w4(32'hbb59e94f),
	.w5(32'h3b2b121f),
	.w6(32'h3c80831d),
	.w7(32'h3a51d0da),
	.w8(32'h3bff556d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0325ee),
	.w1(32'h3b372454),
	.w2(32'h3b785e56),
	.w3(32'h3a27006b),
	.w4(32'h3af4900e),
	.w5(32'h3a64d9c1),
	.w6(32'h3acad000),
	.w7(32'h3b190aab),
	.w8(32'h3b63db77),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b736f07),
	.w1(32'h3b736300),
	.w2(32'h3b345c27),
	.w3(32'h3884dfa8),
	.w4(32'h3a01f348),
	.w5(32'h3af6f24c),
	.w6(32'h3b1c31f1),
	.w7(32'h3b025534),
	.w8(32'h39f332b1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba195161),
	.w1(32'hb94c490a),
	.w2(32'h3a5248a9),
	.w3(32'h3abc7cd0),
	.w4(32'h3b6b0264),
	.w5(32'h3b0b0475),
	.w6(32'h3a901e9f),
	.w7(32'h3b602732),
	.w8(32'h3a92da57),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b0347),
	.w1(32'hbaea8bf0),
	.w2(32'hbaccfc77),
	.w3(32'hba9dab06),
	.w4(32'hbb379e58),
	.w5(32'hbb2ab6b6),
	.w6(32'hbb327aae),
	.w7(32'hbad6ea13),
	.w8(32'hbb29a503),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab65ae),
	.w1(32'h3a7497f2),
	.w2(32'hb984282f),
	.w3(32'hbb20eeea),
	.w4(32'h3b0da070),
	.w5(32'h3bef86c9),
	.w6(32'hba922ab9),
	.w7(32'h3b912ef1),
	.w8(32'hbae8544c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c174ee1),
	.w1(32'h3c2a4eed),
	.w2(32'h3c035162),
	.w3(32'h3b72de10),
	.w4(32'hbb3a83b7),
	.w5(32'h3ca023cb),
	.w6(32'h3cb4d0fc),
	.w7(32'h3b72c665),
	.w8(32'h3cc4ae6b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4331cb),
	.w1(32'h3bf147d9),
	.w2(32'h3c9a49c3),
	.w3(32'h3cc85f4e),
	.w4(32'h3c7f1bc6),
	.w5(32'hbb6ff628),
	.w6(32'h3c99b2a8),
	.w7(32'h3c92915e),
	.w8(32'h3beb5f79),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13af5c),
	.w1(32'h3b254aed),
	.w2(32'h3c49fb68),
	.w3(32'h3b932778),
	.w4(32'hba33887c),
	.w5(32'h3b008754),
	.w6(32'h3c0153ef),
	.w7(32'h3b1a6838),
	.w8(32'h3b3d6abb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6989c),
	.w1(32'h3c10ea18),
	.w2(32'h3c6bdebb),
	.w3(32'h3ba75100),
	.w4(32'h3bd813ae),
	.w5(32'h3c80ac44),
	.w6(32'h3c608d54),
	.w7(32'h3b646bf9),
	.w8(32'h3c8750ea),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba6afc),
	.w1(32'h3a8954cd),
	.w2(32'h3b7f2a22),
	.w3(32'h3bc94c3e),
	.w4(32'h3c32afd4),
	.w5(32'h3c56aeff),
	.w6(32'hbb3b5759),
	.w7(32'hba5f0e8f),
	.w8(32'h3b7e20ef),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d00ed),
	.w1(32'h3b5317b4),
	.w2(32'h3c213ef4),
	.w3(32'h3c2753b4),
	.w4(32'h3c044564),
	.w5(32'hbb522434),
	.w6(32'h3c61e77c),
	.w7(32'hbbaedf24),
	.w8(32'h3bf8b6b0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44f947),
	.w1(32'h3bf15807),
	.w2(32'h3c26d58f),
	.w3(32'h3a9ef282),
	.w4(32'hbbf5cef9),
	.w5(32'h3bebd1e3),
	.w6(32'hbb8e2005),
	.w7(32'h3ab56d6d),
	.w8(32'hbb9923ae),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d8bd9),
	.w1(32'hbba6c4c9),
	.w2(32'hbc2fab00),
	.w3(32'hba60705d),
	.w4(32'hb8a239d6),
	.w5(32'h3b872cb7),
	.w6(32'hb6e35644),
	.w7(32'hbae40125),
	.w8(32'hbb5ef2ef),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08f2e6),
	.w1(32'h3c5c7309),
	.w2(32'hbacb4be3),
	.w3(32'h3c57d5d1),
	.w4(32'h3a65e195),
	.w5(32'hbc4dc2be),
	.w6(32'h3cc1c4b1),
	.w7(32'h3b17d65b),
	.w8(32'hbc794644),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc095cb0),
	.w1(32'hbc4028dc),
	.w2(32'hbc5ab16a),
	.w3(32'hbc1863a6),
	.w4(32'hbc145215),
	.w5(32'hbb907122),
	.w6(32'hbc887adc),
	.w7(32'hbc2aa496),
	.w8(32'hbbdeb7b2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfae583),
	.w1(32'hbc069de9),
	.w2(32'hbbbe3587),
	.w3(32'hbb66c499),
	.w4(32'hbaae8275),
	.w5(32'hba1a4b33),
	.w6(32'hbba8ee37),
	.w7(32'h3a1e0d5b),
	.w8(32'h3b80a1d0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6859a2),
	.w1(32'hbbd0f5a0),
	.w2(32'hbb531351),
	.w3(32'h3bd31766),
	.w4(32'hbb047ef3),
	.w5(32'h3b64351e),
	.w6(32'h3cd0766c),
	.w7(32'h3c1b903c),
	.w8(32'hba4b3d18),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1787d),
	.w1(32'h3c0929fc),
	.w2(32'h3c3e2607),
	.w3(32'h3c3a5840),
	.w4(32'h3bbad998),
	.w5(32'h3be483cb),
	.w6(32'h3c3ee5b7),
	.w7(32'h3c05f0a1),
	.w8(32'h3b28aa55),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7ef94),
	.w1(32'h39b9d4ed),
	.w2(32'h3be50f7d),
	.w3(32'hbab8d117),
	.w4(32'hbb626a1a),
	.w5(32'h3b239a3f),
	.w6(32'h3ae26314),
	.w7(32'hba8915c8),
	.w8(32'h3bebed42),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36e567),
	.w1(32'h3b9c59dd),
	.w2(32'h3c5600cd),
	.w3(32'h3b9b0a39),
	.w4(32'h3b859f93),
	.w5(32'h3c92d04e),
	.w6(32'hbad7b5a3),
	.w7(32'h3b9f9456),
	.w8(32'h3c1b15d4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb762473),
	.w1(32'h3c982ba0),
	.w2(32'h3c0a985b),
	.w3(32'hbb4fb87b),
	.w4(32'h3b0ac87a),
	.w5(32'h3b87264f),
	.w6(32'h3c5829d5),
	.w7(32'hba5b95af),
	.w8(32'h3a49c3d8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52f7db),
	.w1(32'h3b7fb936),
	.w2(32'h3872572c),
	.w3(32'h3934195c),
	.w4(32'hba7ef351),
	.w5(32'hbb196ce6),
	.w6(32'hba1cbc1a),
	.w7(32'h3b634ebd),
	.w8(32'hbb90e04d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae86666),
	.w1(32'hbb637f15),
	.w2(32'h3b24885d),
	.w3(32'hbbb5f329),
	.w4(32'hbbcb4aa8),
	.w5(32'h3bdf997d),
	.w6(32'hbb8a9bb3),
	.w7(32'hba721db4),
	.w8(32'h3b62603d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aabd8),
	.w1(32'h3bae4b6a),
	.w2(32'h3c12e098),
	.w3(32'h3c06a07e),
	.w4(32'hbb54ae5d),
	.w5(32'h3aa9dd10),
	.w6(32'h3c4c4089),
	.w7(32'h3c471018),
	.w8(32'h3aa2a1e5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d7d55),
	.w1(32'h3c141f67),
	.w2(32'h3a97d7e4),
	.w3(32'h3b220242),
	.w4(32'hbc141b34),
	.w5(32'hb9de06fe),
	.w6(32'h3c2a9007),
	.w7(32'h3bac5bb2),
	.w8(32'h3a813186),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fe3a9),
	.w1(32'hbbad52c7),
	.w2(32'hbb0d4ae9),
	.w3(32'h3bb68307),
	.w4(32'h3a9fa8e8),
	.w5(32'hbab5e5f6),
	.w6(32'hbc804de9),
	.w7(32'hba49f070),
	.w8(32'hbb8f9d10),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25a9f5),
	.w1(32'hba8b6b3c),
	.w2(32'h39d858d6),
	.w3(32'h387ef145),
	.w4(32'hbab06bad),
	.w5(32'h3ae186e9),
	.w6(32'hbb911d0c),
	.w7(32'hba2e48dd),
	.w8(32'h3974aaa6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6f0f7),
	.w1(32'hbb2b0f1e),
	.w2(32'hbbbf0ee4),
	.w3(32'h3bc05aff),
	.w4(32'hba4bb743),
	.w5(32'hbbb16ffe),
	.w6(32'hb98351a1),
	.w7(32'hbb47523d),
	.w8(32'h3b8424ce),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4198e3),
	.w1(32'hb94e2580),
	.w2(32'hbac1c3ad),
	.w3(32'hbc398a06),
	.w4(32'hbc4c73d4),
	.w5(32'h384fb150),
	.w6(32'h3c0bc349),
	.w7(32'h37fb8a21),
	.w8(32'hbb6b6e64),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad87c61),
	.w1(32'h3b4ca5d0),
	.w2(32'hba4d0962),
	.w3(32'hbb1236d7),
	.w4(32'hbc0e4ef7),
	.w5(32'hbacb64f3),
	.w6(32'h3bad285e),
	.w7(32'hbc44cc6c),
	.w8(32'h3be7efbd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6def8),
	.w1(32'hbb132eb4),
	.w2(32'hbbb2a344),
	.w3(32'hbb812191),
	.w4(32'hb9c20b2e),
	.w5(32'hb99c2074),
	.w6(32'h3bc814c2),
	.w7(32'hb9f00b5e),
	.w8(32'hbb1f36b3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25ff0e),
	.w1(32'h3c081f6d),
	.w2(32'h3c7a6ff9),
	.w3(32'h3c3fbb22),
	.w4(32'hb9706826),
	.w5(32'h3b8b052f),
	.w6(32'h3c5c962e),
	.w7(32'h3bab8520),
	.w8(32'h3b9c8d33),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8344e),
	.w1(32'hbbaef340),
	.w2(32'hbb954b41),
	.w3(32'hbaac09f7),
	.w4(32'hbc040b86),
	.w5(32'h3bbdae98),
	.w6(32'h3c56113a),
	.w7(32'hbb83b5bc),
	.w8(32'h3c8d884b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d74b9),
	.w1(32'h3a97ff1d),
	.w2(32'hbb884055),
	.w3(32'h3bc05485),
	.w4(32'hbb277a49),
	.w5(32'hbb57f6f8),
	.w6(32'hbb81ed29),
	.w7(32'h3a472230),
	.w8(32'hbb967b39),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule