module layer_10_featuremap_423(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c711e),
	.w1(32'h3a917e5d),
	.w2(32'h3ac7a68c),
	.w3(32'hbb5d5fc9),
	.w4(32'hba0a3765),
	.w5(32'hbb0f43de),
	.w6(32'h3b3c1eb9),
	.w7(32'hbb076743),
	.w8(32'hbb72ca2c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56b100),
	.w1(32'h38eb14a8),
	.w2(32'hb919a6df),
	.w3(32'hbc2a28ef),
	.w4(32'hba3c61ed),
	.w5(32'hbb093a52),
	.w6(32'hbc08e2de),
	.w7(32'hba840250),
	.w8(32'hba8209e6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969b39),
	.w1(32'hbb527429),
	.w2(32'hba6cf264),
	.w3(32'h3b80993d),
	.w4(32'hbc38e504),
	.w5(32'hbc2b21ca),
	.w6(32'h3b8f652f),
	.w7(32'hbc6ba65a),
	.w8(32'hbc3e6696),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63825c),
	.w1(32'h3c124f6b),
	.w2(32'h3b639291),
	.w3(32'hbcc6fb79),
	.w4(32'h3c0588d5),
	.w5(32'h3a50e54e),
	.w6(32'hbcd5c567),
	.w7(32'h3bcf34af),
	.w8(32'hbaa95941),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadccc09),
	.w1(32'h3bb83f96),
	.w2(32'h3b0d2c10),
	.w3(32'hbb37de7a),
	.w4(32'h3b6945dc),
	.w5(32'hb99e0be1),
	.w6(32'hbb9d737f),
	.w7(32'h3a05b316),
	.w8(32'hbb587e6c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91456d),
	.w1(32'hb83d56e7),
	.w2(32'h3aaa0230),
	.w3(32'h3b581730),
	.w4(32'h3985a8d4),
	.w5(32'h3b3e9cab),
	.w6(32'h3b22fd6a),
	.w7(32'h3afd7cd8),
	.w8(32'h3a548cb8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec6bdc),
	.w1(32'hbbf0831f),
	.w2(32'hb9643bb1),
	.w3(32'h3be0a6a3),
	.w4(32'hbbdd9a0c),
	.w5(32'hbb78b19e),
	.w6(32'h3be42983),
	.w7(32'hba92ad07),
	.w8(32'h3b6ef0ff),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacb772),
	.w1(32'hba3fc69b),
	.w2(32'hba06f1d3),
	.w3(32'h3bc08d11),
	.w4(32'hbba3e03b),
	.w5(32'h3a806018),
	.w6(32'h3c7729a7),
	.w7(32'hbbf54a92),
	.w8(32'h3bb762ef),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ff0302),
	.w1(32'h3b106cfe),
	.w2(32'hbc37f52d),
	.w3(32'h3af51ccc),
	.w4(32'h3c48ad1f),
	.w5(32'hbb000afe),
	.w6(32'h3c44e4c3),
	.w7(32'h3bb7d026),
	.w8(32'hbbe8938b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bdc72),
	.w1(32'hba901863),
	.w2(32'hbad1bd50),
	.w3(32'h3afecef9),
	.w4(32'hbbcdd41d),
	.w5(32'hbb9f33ff),
	.w6(32'hbaecab03),
	.w7(32'hbab5e6c9),
	.w8(32'hbb0cd1bb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b2663),
	.w1(32'h3b9a7c75),
	.w2(32'h3bd08c97),
	.w3(32'h3af122ac),
	.w4(32'hba950928),
	.w5(32'h3acfbf61),
	.w6(32'h3bc7a4b4),
	.w7(32'h3b830722),
	.w8(32'h3bcbefe4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3c81),
	.w1(32'h3be7916a),
	.w2(32'h3bd42e9e),
	.w3(32'h3c4f0d9f),
	.w4(32'h3be50523),
	.w5(32'h3bfbafdb),
	.w6(32'h3c838e75),
	.w7(32'h3b1d03d5),
	.w8(32'h3b9c90aa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66fe8f),
	.w1(32'hbc4b3fe0),
	.w2(32'hbc23b666),
	.w3(32'h3b5c96f4),
	.w4(32'hbbd311bd),
	.w5(32'hbbadff90),
	.w6(32'h3b98de66),
	.w7(32'hbbe3d792),
	.w8(32'hbbc07ed7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4717c8),
	.w1(32'hbb878ab8),
	.w2(32'hbc32e617),
	.w3(32'hbc7c1e13),
	.w4(32'h380b9a41),
	.w5(32'hbb691743),
	.w6(32'hbc406562),
	.w7(32'hbab3b312),
	.w8(32'hbbeabf3e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4eb80),
	.w1(32'h3ab3187b),
	.w2(32'hbaa5d31c),
	.w3(32'h3b1deccd),
	.w4(32'h3b22c9c9),
	.w5(32'hb98b6808),
	.w6(32'h390335ad),
	.w7(32'h3aa6853f),
	.w8(32'h3ae33de6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a1ff),
	.w1(32'hb9bdd385),
	.w2(32'h3b1b4ae4),
	.w3(32'h398fc550),
	.w4(32'hba838ea6),
	.w5(32'h3b906389),
	.w6(32'hb8e40d1d),
	.w7(32'hbb913d4a),
	.w8(32'h3b354b2f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d4cfd),
	.w1(32'hbb3c9ef3),
	.w2(32'h3b116372),
	.w3(32'h3b9bd8fa),
	.w4(32'hbac28165),
	.w5(32'h3b0f8cfc),
	.w6(32'h3b15ad7c),
	.w7(32'h3b34b9cd),
	.w8(32'h3b930ff3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d5011),
	.w1(32'hbb9e71c1),
	.w2(32'hbb4c8de3),
	.w3(32'hba9bb214),
	.w4(32'hbb91311c),
	.w5(32'hbb5bd1f1),
	.w6(32'h38fd576f),
	.w7(32'hba6f39d3),
	.w8(32'hbb7a7c99),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39926a5d),
	.w1(32'h3a25d158),
	.w2(32'hbba113b8),
	.w3(32'hbb390102),
	.w4(32'h3b682c2c),
	.w5(32'hba5abd3d),
	.w6(32'h3a3892b1),
	.w7(32'h3b585f12),
	.w8(32'h3a0ca3b0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be065ef),
	.w1(32'h39bccc5c),
	.w2(32'h3a1e1b8d),
	.w3(32'h3c3601c4),
	.w4(32'h3c17b54f),
	.w5(32'h39a77642),
	.w6(32'h3c1f7223),
	.w7(32'h3c141ce4),
	.w8(32'h3b7a5e81),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be820b6),
	.w1(32'h3b0bebc4),
	.w2(32'hbabf5870),
	.w3(32'h3bab0be8),
	.w4(32'h3a7c1935),
	.w5(32'hb91a4b53),
	.w6(32'h3ae2ccc3),
	.w7(32'hba585a2c),
	.w8(32'hb9b48898),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf12d33),
	.w1(32'h3bca8e58),
	.w2(32'h3bd25484),
	.w3(32'h3c236e75),
	.w4(32'h3bfd708f),
	.w5(32'h3bdf0efd),
	.w6(32'h3c204148),
	.w7(32'h3b9941b7),
	.w8(32'h3b6ecb8b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf4c4b),
	.w1(32'hbaa6b59b),
	.w2(32'hbc153a82),
	.w3(32'hbad5880d),
	.w4(32'h3ab53588),
	.w5(32'hbbce8db5),
	.w6(32'hbb839ac7),
	.w7(32'h3a616e3f),
	.w8(32'hbb5be969),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8453c1),
	.w1(32'hbab34391),
	.w2(32'hbb37d7ab),
	.w3(32'hbb987027),
	.w4(32'h3b18ef08),
	.w5(32'hbb09b269),
	.w6(32'hba4bd333),
	.w7(32'h3b5d6d9b),
	.w8(32'h3ad7d2f8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c627916),
	.w1(32'h3a7534ad),
	.w2(32'hbc016c30),
	.w3(32'h3c51b22f),
	.w4(32'h3911b65c),
	.w5(32'hbb82a5f5),
	.w6(32'h3c47c313),
	.w7(32'hbb4f15d6),
	.w8(32'hbbc4a9ec),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80083b),
	.w1(32'h3b0babcf),
	.w2(32'hb9f5d4e1),
	.w3(32'h3beede75),
	.w4(32'h3ac92613),
	.w5(32'hbb83e173),
	.w6(32'h3baff3cc),
	.w7(32'h3b74490e),
	.w8(32'hba5c69a3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d7448),
	.w1(32'h3be3f064),
	.w2(32'hb99d6f06),
	.w3(32'hb80bb9a9),
	.w4(32'h3a79ac98),
	.w5(32'hbbce9c9c),
	.w6(32'h3b17db4d),
	.w7(32'h3a6ff5e6),
	.w8(32'hbb96582d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ab27),
	.w1(32'h3b75bdf9),
	.w2(32'hb9b3b621),
	.w3(32'h3998ad74),
	.w4(32'h3b2513b0),
	.w5(32'h3aee736f),
	.w6(32'h3a90aa49),
	.w7(32'hba30fb0d),
	.w8(32'hb9336722),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e500f),
	.w1(32'h3b6e1deb),
	.w2(32'h3b74da2c),
	.w3(32'h3bb125a2),
	.w4(32'h3a9ad15e),
	.w5(32'hba8a4ee6),
	.w6(32'h3b902818),
	.w7(32'h3a5636da),
	.w8(32'h3a06e548),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919d40),
	.w1(32'hbbd00970),
	.w2(32'hbba9fb16),
	.w3(32'hbba18d94),
	.w4(32'hbbd72a5e),
	.w5(32'hbaff30a3),
	.w6(32'hbb4d754d),
	.w7(32'hbb4e6bff),
	.w8(32'hba48287c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81141a),
	.w1(32'hba947a90),
	.w2(32'h3acddc86),
	.w3(32'hbb9ea372),
	.w4(32'h3b96c427),
	.w5(32'h3b5f5033),
	.w6(32'hbb94fd3e),
	.w7(32'h3c1202cf),
	.w8(32'h3bbb8a70),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66ca57),
	.w1(32'hbc8abe6b),
	.w2(32'hb9986e31),
	.w3(32'hb930f394),
	.w4(32'hbca5e714),
	.w5(32'hbc10eff9),
	.w6(32'hb832dde9),
	.w7(32'hbcb0d8a5),
	.w8(32'hbc0529d7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc753149),
	.w1(32'hb99d716c),
	.w2(32'hbad6ce04),
	.w3(32'hbcb16a81),
	.w4(32'hbb295fa2),
	.w5(32'hbb8ecae3),
	.w6(32'hbcc70b70),
	.w7(32'h3a29d733),
	.w8(32'hbb2510e0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc3659),
	.w1(32'h3aa846c8),
	.w2(32'hbaa5bca6),
	.w3(32'hbbf15eed),
	.w4(32'h3bad5502),
	.w5(32'h3a232f86),
	.w6(32'hbb1c467f),
	.w7(32'h3ba9b7c2),
	.w8(32'h3b616aef),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e101e3),
	.w1(32'hbc77f936),
	.w2(32'hbc1d6a7f),
	.w3(32'h3a4b67d5),
	.w4(32'hbb515c5c),
	.w5(32'hb726c9e4),
	.w6(32'h3b060c9a),
	.w7(32'hbbb3537b),
	.w8(32'hbc1930a2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e0e43),
	.w1(32'h3bb0020a),
	.w2(32'h3b96ca4b),
	.w3(32'h3c18a0a8),
	.w4(32'h3b628240),
	.w5(32'h39a56236),
	.w6(32'hba1fa935),
	.w7(32'h3baba9e5),
	.w8(32'hb8e4e60e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd297d),
	.w1(32'hbc648d0d),
	.w2(32'hbbc8ad6e),
	.w3(32'hbb4f9a6d),
	.w4(32'hbc265988),
	.w5(32'hbb414b0f),
	.w6(32'hba635432),
	.w7(32'h3991f133),
	.w8(32'h3aebf464),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8666ee),
	.w1(32'hbc03ded1),
	.w2(32'h3ba51855),
	.w3(32'h3bd555eb),
	.w4(32'hbbfb1d8e),
	.w5(32'h3ae089c2),
	.w6(32'h3a627850),
	.w7(32'hbc3069fe),
	.w8(32'h3acfcd6e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee2085),
	.w1(32'h3bce8876),
	.w2(32'h3bb5c77f),
	.w3(32'h3b0cd551),
	.w4(32'h3bb96cbd),
	.w5(32'h3b6b54f0),
	.w6(32'hbb8cc555),
	.w7(32'hbb8a7e55),
	.w8(32'hbb779bfa),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90f9a8),
	.w1(32'h388d9216),
	.w2(32'hba577287),
	.w3(32'hba9ff352),
	.w4(32'hbb06a548),
	.w5(32'hbb752a1f),
	.w6(32'hbb54fc7c),
	.w7(32'hbab51f8e),
	.w8(32'hbacbeb5a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0892fc),
	.w1(32'h3a2d7b48),
	.w2(32'hbbdd064c),
	.w3(32'hbad8a85d),
	.w4(32'h3ba2830a),
	.w5(32'hbbc1d2e8),
	.w6(32'hbac12345),
	.w7(32'h3acb686f),
	.w8(32'hbc00762b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc568729),
	.w1(32'hbbd03af2),
	.w2(32'hbbe300da),
	.w3(32'hbca3c829),
	.w4(32'hbbd07a78),
	.w5(32'hbbb7b646),
	.w6(32'hbcbba233),
	.w7(32'hbc0a726c),
	.w8(32'hbbd5f56f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023144),
	.w1(32'hbbd1d678),
	.w2(32'hbace952c),
	.w3(32'hbc0addbc),
	.w4(32'hbbc591d0),
	.w5(32'hbb2054ed),
	.w6(32'hbc4141fd),
	.w7(32'hbbabd7eb),
	.w8(32'hbb66e52e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2913aa),
	.w1(32'hbb53e678),
	.w2(32'hbc1afb8c),
	.w3(32'hbc2b19f9),
	.w4(32'hbab43ba3),
	.w5(32'hbbf173d6),
	.w6(32'hbc124173),
	.w7(32'hba9f7f7b),
	.w8(32'hbc0d37e1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebf883),
	.w1(32'h3b331178),
	.w2(32'hbb07e9a8),
	.w3(32'hbbc10fe6),
	.w4(32'h3c12bf94),
	.w5(32'h39b03bee),
	.w6(32'hbbc9d897),
	.w7(32'h3bd188a1),
	.w8(32'hb98d461c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca938d),
	.w1(32'hbb36a007),
	.w2(32'hbb5a399d),
	.w3(32'h3b00e62a),
	.w4(32'hba8911de),
	.w5(32'hbb8ca97e),
	.w6(32'h3ae9e931),
	.w7(32'hbb780e1c),
	.w8(32'hbbc14b81),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fab44),
	.w1(32'hbbc81810),
	.w2(32'hbb3cf5ca),
	.w3(32'hbafe481b),
	.w4(32'hba01c64a),
	.w5(32'hbabb8524),
	.w6(32'hbbac198f),
	.w7(32'h3ab1cf36),
	.w8(32'h3aa693b1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c3d01),
	.w1(32'hbb4f2f6f),
	.w2(32'hbbd85723),
	.w3(32'hba9204ed),
	.w4(32'h393e9f42),
	.w5(32'hbbef92ba),
	.w6(32'h3b22571b),
	.w7(32'h3b52821c),
	.w8(32'hbba647c7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8ea8),
	.w1(32'h3c03a12b),
	.w2(32'h3b2f3d11),
	.w3(32'hbbd205fb),
	.w4(32'h3c6dabe8),
	.w5(32'h3c438fc5),
	.w6(32'hbc042b1b),
	.w7(32'h3c7d163e),
	.w8(32'h3c80f5c8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c867661),
	.w1(32'hbc6f11b2),
	.w2(32'h398456e4),
	.w3(32'h3ce09a5a),
	.w4(32'hbca42055),
	.w5(32'hbbee7ca8),
	.w6(32'h3cefaf8c),
	.w7(32'hbca30289),
	.w8(32'hbbdd9d79),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c3a49),
	.w1(32'h3bbaa323),
	.w2(32'h3a487dbd),
	.w3(32'hbcbb148e),
	.w4(32'h3c13dd2d),
	.w5(32'h3baaf7a8),
	.w6(32'hbcabce85),
	.w7(32'h3b9d7958),
	.w8(32'h3ba608f7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dfefc),
	.w1(32'hbc08df0a),
	.w2(32'hbc389081),
	.w3(32'h3b2c6696),
	.w4(32'hbbb15abb),
	.w5(32'hbc0ec0eb),
	.w6(32'h3ab4a362),
	.w7(32'hbb15ec10),
	.w8(32'hbbf7b6c0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0285c7),
	.w1(32'h3a59c4c8),
	.w2(32'h398542aa),
	.w3(32'h3bba4767),
	.w4(32'h3aff56cd),
	.w5(32'h3b851c36),
	.w6(32'h3b27f1b6),
	.w7(32'h3b972740),
	.w8(32'h3bcb5bf5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e0e10),
	.w1(32'hbb795f3e),
	.w2(32'hbbc3b89b),
	.w3(32'hbbaa5534),
	.w4(32'hbaee9c65),
	.w5(32'h398ee707),
	.w6(32'h3b025141),
	.w7(32'h3be6c6f5),
	.w8(32'h3b38350b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe43023),
	.w1(32'hbb988ac1),
	.w2(32'h3a8f506e),
	.w3(32'h3ac8d46e),
	.w4(32'hbbb74125),
	.w5(32'hbb155203),
	.w6(32'h3ab871b7),
	.w7(32'hbb8e1a5e),
	.w8(32'hbb044d8d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b30cb),
	.w1(32'h3b2f588b),
	.w2(32'hbb8322cc),
	.w3(32'hbb83fa72),
	.w4(32'hbac16a08),
	.w5(32'hbbdc4d45),
	.w6(32'hbbd5bb2b),
	.w7(32'h3b0c9e79),
	.w8(32'hbbc36970),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b692a76),
	.w1(32'hba96554e),
	.w2(32'hbb0b9803),
	.w3(32'h3bae191b),
	.w4(32'hbb13908e),
	.w5(32'hbb5dca2a),
	.w6(32'h3c16b238),
	.w7(32'hbb57e3b6),
	.w8(32'hbbb082d6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f69770),
	.w1(32'h3ba80637),
	.w2(32'h3a7a2786),
	.w3(32'hbb2bf509),
	.w4(32'h3b323f74),
	.w5(32'hbb65357e),
	.w6(32'hbaaf78a2),
	.w7(32'h3b431334),
	.w8(32'hbbba5f91),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9553bd),
	.w1(32'hbb34bfa5),
	.w2(32'hbc406e71),
	.w3(32'h3b55a31e),
	.w4(32'hbb8edb5d),
	.w5(32'hbc5a7f69),
	.w6(32'h3a5ea1da),
	.w7(32'hbbc4bf2b),
	.w8(32'hbc667757),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc307b56),
	.w1(32'h3a8da8ff),
	.w2(32'h38f6f52e),
	.w3(32'hbc3fea1b),
	.w4(32'h3aa19aa3),
	.w5(32'h3b80bf7b),
	.w6(32'hbc28dc96),
	.w7(32'h3b92867e),
	.w8(32'h3b4588cb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77961b),
	.w1(32'h3bc50d6e),
	.w2(32'h3bdfbf96),
	.w3(32'h3b0bb287),
	.w4(32'h3b6e47d7),
	.w5(32'hbbc4f80b),
	.w6(32'h3b7be53c),
	.w7(32'h3b850d09),
	.w8(32'hb98bc0c8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83363a),
	.w1(32'h3b2b2145),
	.w2(32'h3b6cf757),
	.w3(32'hbabc3d4a),
	.w4(32'h3b3d8282),
	.w5(32'h3b4ce20a),
	.w6(32'hbaa45a29),
	.w7(32'h3b4327dd),
	.w8(32'h3bca11cd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf77516),
	.w1(32'hbc679242),
	.w2(32'hbbb24d75),
	.w3(32'h3bcf4e89),
	.w4(32'hbc940ad3),
	.w5(32'hbc2982ea),
	.w6(32'h3bd6fde4),
	.w7(32'hbc8fc560),
	.w8(32'hbc40bdf9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1345b1),
	.w1(32'h39a70e72),
	.w2(32'hbaca7d11),
	.w3(32'hbc780848),
	.w4(32'h3ad24415),
	.w5(32'h3a97d7c9),
	.w6(32'hbc8b7ef2),
	.w7(32'hba6a8f20),
	.w8(32'hb9175e9b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2d055),
	.w1(32'h3bbe84fb),
	.w2(32'h3ae18f3b),
	.w3(32'hbbc4d817),
	.w4(32'h3baac986),
	.w5(32'h3b13f28b),
	.w6(32'hbb2b2884),
	.w7(32'h3b6704dc),
	.w8(32'h394ec91e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13b759),
	.w1(32'h3bbbff88),
	.w2(32'h3b125b15),
	.w3(32'h3adf9652),
	.w4(32'h3c07b164),
	.w5(32'h3b946719),
	.w6(32'h3a410e8a),
	.w7(32'h3bad9b93),
	.w8(32'h3bab2243),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baccf74),
	.w1(32'h3b628d74),
	.w2(32'hba5096cf),
	.w3(32'h3c27d7a9),
	.w4(32'h3bd5157b),
	.w5(32'h3b5a0258),
	.w6(32'h3c102d59),
	.w7(32'hbab13e81),
	.w8(32'hba875a5d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75e944),
	.w1(32'hbb68ce91),
	.w2(32'h3a968f4e),
	.w3(32'hb9a83859),
	.w4(32'hb872be08),
	.w5(32'hba93b9e7),
	.w6(32'hbadd124c),
	.w7(32'h3accb35a),
	.w8(32'h3a9b84f8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b0b67),
	.w1(32'hbb860ce1),
	.w2(32'hbc1442f0),
	.w3(32'h3b38f202),
	.w4(32'hbb712ad6),
	.w5(32'hbbd4a092),
	.w6(32'h3b292d4a),
	.w7(32'hbbd73458),
	.w8(32'hbc0f15ff),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bd4b9),
	.w1(32'h3af93615),
	.w2(32'hbb78aed8),
	.w3(32'h3a91bb02),
	.w4(32'h3b033143),
	.w5(32'hbab592ee),
	.w6(32'hbac1e150),
	.w7(32'h3afa3d5b),
	.w8(32'h3ae142a7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3830c015),
	.w1(32'h3b0524fd),
	.w2(32'h3a82c6c6),
	.w3(32'h385719e3),
	.w4(32'h3a7683bd),
	.w5(32'hbad3741f),
	.w6(32'hb7b9f58e),
	.w7(32'h3aa57211),
	.w8(32'h3a3f8932),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39017aa4),
	.w1(32'h39b35843),
	.w2(32'hba0ebce8),
	.w3(32'hba33e598),
	.w4(32'hb9956367),
	.w5(32'hbaf48e66),
	.w6(32'h39269dd6),
	.w7(32'h39910843),
	.w8(32'h3ae7ec27),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab45781),
	.w1(32'hbac1e871),
	.w2(32'hbae63371),
	.w3(32'h3a679ccb),
	.w4(32'hba149b6d),
	.w5(32'hbb0e066b),
	.w6(32'h39f5d21f),
	.w7(32'hb7b43fb8),
	.w8(32'hba768081),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf419df),
	.w1(32'hbaa5c661),
	.w2(32'h3931ad60),
	.w3(32'hba0fc966),
	.w4(32'h399c4da5),
	.w5(32'hbad92de3),
	.w6(32'hba5452be),
	.w7(32'hb9cb6f1c),
	.w8(32'hbae5680f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dd2eaf),
	.w1(32'h3a35aaa9),
	.w2(32'h38d25fff),
	.w3(32'hb837b361),
	.w4(32'hba276eb7),
	.w5(32'hbabc17c4),
	.w6(32'h391d8487),
	.w7(32'hba8e8d1b),
	.w8(32'hbae43a2e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3fe2a),
	.w1(32'hbaa0c922),
	.w2(32'hba817c19),
	.w3(32'hbb9a5da8),
	.w4(32'h3af7607d),
	.w5(32'h39909382),
	.w6(32'hbad6adaf),
	.w7(32'h3ac3c19d),
	.w8(32'h3a16a72e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfb108),
	.w1(32'hbb52589a),
	.w2(32'hbaea75ec),
	.w3(32'hba0267f8),
	.w4(32'hba42e0fe),
	.w5(32'hba00962a),
	.w6(32'h3a439af5),
	.w7(32'h3ad65914),
	.w8(32'h3a8dcca4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a148bae),
	.w1(32'h39cecd49),
	.w2(32'hb918cc43),
	.w3(32'h3ab289e9),
	.w4(32'h3b7a5bf8),
	.w5(32'h3b9f87af),
	.w6(32'h3abd73b4),
	.w7(32'h3b5d8952),
	.w8(32'h3b89680d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bd979),
	.w1(32'hbb5b5aeb),
	.w2(32'hbb8d6971),
	.w3(32'h3b3ae926),
	.w4(32'h388af58a),
	.w5(32'hbafbf6d5),
	.w6(32'h3b04cd6a),
	.w7(32'h3a579c33),
	.w8(32'hbaf3a81f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5e5a0),
	.w1(32'hba444579),
	.w2(32'h3a06f1d9),
	.w3(32'h3a62b07e),
	.w4(32'h3a8c7571),
	.w5(32'h39bb9052),
	.w6(32'h395987bc),
	.w7(32'hba2309b7),
	.w8(32'hba805b87),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60e31f),
	.w1(32'hbaf98a4f),
	.w2(32'hbb787147),
	.w3(32'h3a98f7b1),
	.w4(32'hbad561e6),
	.w5(32'hbb1f6242),
	.w6(32'h3a8a2a61),
	.w7(32'hbae22a6a),
	.w8(32'hbab2b781),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2670cd),
	.w1(32'hba616836),
	.w2(32'hbaee23e8),
	.w3(32'hbad933c9),
	.w4(32'hb86c98c9),
	.w5(32'hba9359b2),
	.w6(32'hb9b72068),
	.w7(32'h3a14fcf9),
	.w8(32'hba2704d2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e9a2d),
	.w1(32'h3993a4bf),
	.w2(32'h3a7a13d5),
	.w3(32'hb9eb719e),
	.w4(32'h38425000),
	.w5(32'h39da549e),
	.w6(32'h3979fab1),
	.w7(32'h3a4b8d14),
	.w8(32'h3ac08312),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4f0f6),
	.w1(32'h392f45b3),
	.w2(32'h3992774b),
	.w3(32'h3ab6412b),
	.w4(32'h3798fcf7),
	.w5(32'hbab8fdbb),
	.w6(32'h3ab23b83),
	.w7(32'h38e0df48),
	.w8(32'hbaa30927),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16976d),
	.w1(32'h39b438ed),
	.w2(32'h3abca41c),
	.w3(32'hbaf5ef3c),
	.w4(32'h3a1ebb0f),
	.w5(32'h3ac44cfc),
	.w6(32'hb7a0d837),
	.w7(32'h3917f265),
	.w8(32'h3a17f35d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10a6cd),
	.w1(32'h3a1ab5c6),
	.w2(32'hb98f9a25),
	.w3(32'hb9050e05),
	.w4(32'hb9cea3b8),
	.w5(32'hbb01181c),
	.w6(32'h3989da64),
	.w7(32'hba4ea529),
	.w8(32'hbb0d79cf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ef15),
	.w1(32'hbb0cf3e2),
	.w2(32'h3ad925d9),
	.w3(32'hbb19f017),
	.w4(32'h3a67babf),
	.w5(32'h3b83e859),
	.w6(32'hbb4acfa6),
	.w7(32'hbad4374a),
	.w8(32'h3a9cc628),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47a91a),
	.w1(32'hb9ff8b8a),
	.w2(32'h38e2d83d),
	.w3(32'h3adf7f8d),
	.w4(32'h3a96fbba),
	.w5(32'h39bc8edc),
	.w6(32'hb984ae08),
	.w7(32'h39048afd),
	.w8(32'hb98efe6f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8196ad),
	.w1(32'hbb1318bb),
	.w2(32'hbb3b7f60),
	.w3(32'hbaa0fc02),
	.w4(32'hb993b4f2),
	.w5(32'hbac1cabf),
	.w6(32'hba45999f),
	.w7(32'h3b0e2a95),
	.w8(32'hba751d41),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0c0c),
	.w1(32'hbb3a0494),
	.w2(32'hbb457892),
	.w3(32'hbb929477),
	.w4(32'hbb4109b0),
	.w5(32'hbadc5028),
	.w6(32'hbb4fdc8e),
	.w7(32'hbad21062),
	.w8(32'hbaae7b00),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858234),
	.w1(32'h3b49700c),
	.w2(32'h3b40862f),
	.w3(32'h3a37e4f1),
	.w4(32'h3b19ff32),
	.w5(32'h3b159ee0),
	.w6(32'hbacfc4b1),
	.w7(32'h3a3ebefc),
	.w8(32'h3ad1c29a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b849),
	.w1(32'hb9bfe0ad),
	.w2(32'hba11d64f),
	.w3(32'h3a8acbd8),
	.w4(32'h3b74b173),
	.w5(32'h3a6b9685),
	.w6(32'h3afc72c9),
	.w7(32'h3bb0b129),
	.w8(32'h3a9afa4d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca4ce9),
	.w1(32'h3ae2e3fd),
	.w2(32'h3a0f2dee),
	.w3(32'h3afe2c19),
	.w4(32'h3a7ad106),
	.w5(32'hb9b14d54),
	.w6(32'h3b468ba1),
	.w7(32'hb9a9ed39),
	.w8(32'hbb0976d7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807a97),
	.w1(32'hbbf4f324),
	.w2(32'hbbf9737c),
	.w3(32'hbaa1038b),
	.w4(32'hbaef9df1),
	.w5(32'hbb2ad884),
	.w6(32'h397b1c8b),
	.w7(32'hbb02c3c5),
	.w8(32'hbbaad649),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b448bd),
	.w1(32'h39d33bc2),
	.w2(32'h3aa9ffff),
	.w3(32'h3acc6a01),
	.w4(32'hb9b0a866),
	.w5(32'hbaec76fe),
	.w6(32'h3aa063fc),
	.w7(32'hbaa973ad),
	.w8(32'hba872e1f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00bb8e),
	.w1(32'h3a9a799a),
	.w2(32'h39f68656),
	.w3(32'hba4266d6),
	.w4(32'hb8453f2f),
	.w5(32'hbb249043),
	.w6(32'h399f8d57),
	.w7(32'hba75ed8c),
	.w8(32'h3a7343f8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967a15e),
	.w1(32'h3b190908),
	.w2(32'h3ab33f37),
	.w3(32'h394434aa),
	.w4(32'h3aa7ff5f),
	.w5(32'hbb280bbd),
	.w6(32'h3b41959d),
	.w7(32'h3b161006),
	.w8(32'hbaa61dac),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67c0b5),
	.w1(32'hbb743a67),
	.w2(32'hbbdc2ea5),
	.w3(32'hba9b24e0),
	.w4(32'hba9fedd0),
	.w5(32'hbbba8eed),
	.w6(32'h3b122cb7),
	.w7(32'h3a22c57c),
	.w8(32'hbb4daa67),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641abc),
	.w1(32'hbb51a68c),
	.w2(32'hbafd39ad),
	.w3(32'hba4f1ee1),
	.w4(32'hbb180bcf),
	.w5(32'hbb31930b),
	.w6(32'hba7d989a),
	.w7(32'hbb7ebffa),
	.w8(32'hbb801809),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e0a1d),
	.w1(32'hba01363e),
	.w2(32'h3a44a0e3),
	.w3(32'hbba488bd),
	.w4(32'h3a592d5f),
	.w5(32'hb9d528e8),
	.w6(32'hbb47d08c),
	.w7(32'h3b478058),
	.w8(32'h3a86ca79),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a044),
	.w1(32'hba84c592),
	.w2(32'h3b05d2fb),
	.w3(32'hbbc5dddc),
	.w4(32'h3b67ea4f),
	.w5(32'h39978d00),
	.w6(32'hbbb95499),
	.w7(32'h372d8030),
	.w8(32'hbac70709),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20ae65),
	.w1(32'hbade5a19),
	.w2(32'hbba1aab0),
	.w3(32'h3a838515),
	.w4(32'hba1a28fd),
	.w5(32'hbb72b33b),
	.w6(32'h3a8e0939),
	.w7(32'hba8d8f74),
	.w8(32'hbb0b95c8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba53bad),
	.w1(32'hba697d40),
	.w2(32'h395669f7),
	.w3(32'hbaa2aea9),
	.w4(32'h3bbc568e),
	.w5(32'hba6e949a),
	.w6(32'hb9e17053),
	.w7(32'h3bc8b427),
	.w8(32'h3b09a36f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0d04),
	.w1(32'h3b9ca619),
	.w2(32'h3b3977f4),
	.w3(32'h3a6e29ee),
	.w4(32'h3b62ec3d),
	.w5(32'h3b32b8d0),
	.w6(32'h3af4bc99),
	.w7(32'h3b4b947e),
	.w8(32'h3b8122eb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22b5db),
	.w1(32'hbbc13c17),
	.w2(32'hbb63e7ce),
	.w3(32'hbc0b10d0),
	.w4(32'hb9906d8e),
	.w5(32'hbad84439),
	.w6(32'hbabc06d6),
	.w7(32'h3b678434),
	.w8(32'hba3857e2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bca15d),
	.w1(32'hb9ef49dc),
	.w2(32'h3a960eaa),
	.w3(32'h3a9455ac),
	.w4(32'h3a5f8294),
	.w5(32'h3a83ed9f),
	.w6(32'h399b97c3),
	.w7(32'h3b3cf70b),
	.w8(32'h3b1af99a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e234b),
	.w1(32'h3a91f6e4),
	.w2(32'h3a792353),
	.w3(32'h3a762265),
	.w4(32'h39c69cf0),
	.w5(32'hb9463d43),
	.w6(32'h3a25c122),
	.w7(32'h3a31f02b),
	.w8(32'h39c8f05d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b92ba9),
	.w1(32'hba823dbf),
	.w2(32'hb9803aa4),
	.w3(32'hb7e3763d),
	.w4(32'hbaa86e1c),
	.w5(32'h3a091a2c),
	.w6(32'hb99c3f0d),
	.w7(32'hba9d5e75),
	.w8(32'h3a7b078b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5652a),
	.w1(32'h3a90d839),
	.w2(32'hb91106d2),
	.w3(32'h3acca4bc),
	.w4(32'h3afb3d65),
	.w5(32'h3a77120a),
	.w6(32'h3ab7c54b),
	.w7(32'h3b8ef21c),
	.w8(32'h3b1913d6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af87053),
	.w1(32'h3aa34b10),
	.w2(32'hbb3b9d5d),
	.w3(32'h3b5face4),
	.w4(32'h3b5a83fd),
	.w5(32'h3a9cbc5c),
	.w6(32'h3b235198),
	.w7(32'h3b50e4f3),
	.w8(32'h3a9ba088),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05b75c),
	.w1(32'hbad3b172),
	.w2(32'hbb2fc341),
	.w3(32'h3ae6633d),
	.w4(32'hb939d34a),
	.w5(32'hbab98be5),
	.w6(32'h3adc4a65),
	.w7(32'h39b66fff),
	.w8(32'hba137072),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35cb4c),
	.w1(32'hba7482aa),
	.w2(32'hb70d33ae),
	.w3(32'hba64cd12),
	.w4(32'hba5b4850),
	.w5(32'hba6211ff),
	.w6(32'hba6889b8),
	.w7(32'hbac19b68),
	.w8(32'hbb345475),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e8ecb),
	.w1(32'h3b2a4410),
	.w2(32'h3b950e84),
	.w3(32'hba3c1606),
	.w4(32'h3b662c12),
	.w5(32'h38213030),
	.w6(32'h3965006c),
	.w7(32'h3b8275cc),
	.w8(32'h3b06b0d6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f3f06),
	.w1(32'hbaade171),
	.w2(32'h39adf86d),
	.w3(32'h37513360),
	.w4(32'hba0abc78),
	.w5(32'hbad0ac70),
	.w6(32'h39cc0c9b),
	.w7(32'h3acd7102),
	.w8(32'h3af7b49a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34b4df),
	.w1(32'hb9110071),
	.w2(32'hbac1fadb),
	.w3(32'hbab94470),
	.w4(32'h3a6c832e),
	.w5(32'hb99ba21d),
	.w6(32'h37171b23),
	.w7(32'h3b0d05b0),
	.w8(32'h3ab9d277),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90f9ab),
	.w1(32'h3a889a69),
	.w2(32'h3a5d2340),
	.w3(32'h39def38a),
	.w4(32'h39740b8a),
	.w5(32'h39a7fd51),
	.w6(32'h385eeaa1),
	.w7(32'h3a0d187c),
	.w8(32'h3a736cfd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a630c6),
	.w1(32'h3a2bcd02),
	.w2(32'h3a787457),
	.w3(32'h3a6373cd),
	.w4(32'h3994261c),
	.w5(32'h3ada3962),
	.w6(32'h39860c85),
	.w7(32'h39e56e42),
	.w8(32'h3a25f4ed),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b66a4),
	.w1(32'h3a7d3ae8),
	.w2(32'h3b01239b),
	.w3(32'h3ade5ca2),
	.w4(32'h397d92af),
	.w5(32'h3a8b5096),
	.w6(32'h3a79b7f1),
	.w7(32'h3af4574e),
	.w8(32'h3a9b862f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8078e9),
	.w1(32'h39288e75),
	.w2(32'h3a727547),
	.w3(32'h3b02e2fe),
	.w4(32'h3a83a340),
	.w5(32'h3a37e8d3),
	.w6(32'h3ab0fecc),
	.w7(32'h3a1442f8),
	.w8(32'hb89698c0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8b2f6),
	.w1(32'hb9a90b21),
	.w2(32'hb9cc1f3d),
	.w3(32'h3a9de2d0),
	.w4(32'h3aee2d3a),
	.w5(32'hba169805),
	.w6(32'h3a6f923d),
	.w7(32'h3b3ee6f4),
	.w8(32'h3b509f6d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2983ea),
	.w1(32'hba2158d0),
	.w2(32'hba1af04c),
	.w3(32'h3aa850ed),
	.w4(32'h3a1e8e50),
	.w5(32'hb940f557),
	.w6(32'h3b1ca09e),
	.w7(32'h3933ab14),
	.w8(32'hb9b39858),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0401b),
	.w1(32'hba288fb6),
	.w2(32'h3a3667e6),
	.w3(32'hbb08c203),
	.w4(32'hba322a05),
	.w5(32'hba392ee4),
	.w6(32'hba0fd5b3),
	.w7(32'h3aa4ffd4),
	.w8(32'h3acfb17f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e89f0),
	.w1(32'h3b2bcb55),
	.w2(32'h3b28eacb),
	.w3(32'hba00182f),
	.w4(32'h39a5d576),
	.w5(32'hbb266505),
	.w6(32'hbb33d269),
	.w7(32'hbaaa0521),
	.w8(32'hbb04a1c2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91524ed),
	.w1(32'h3a462009),
	.w2(32'h36cf7e76),
	.w3(32'hb78f2b1c),
	.w4(32'hba6eefb4),
	.w5(32'hbb13d51b),
	.w6(32'h3a836523),
	.w7(32'hba348c89),
	.w8(32'hbb1afdd1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3300d1),
	.w1(32'hb95efa33),
	.w2(32'h39394ede),
	.w3(32'hba735cd5),
	.w4(32'h39b31ede),
	.w5(32'h3aee9330),
	.w6(32'h39b0b239),
	.w7(32'h3a821d8a),
	.w8(32'h3a8ea23a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39311659),
	.w1(32'h396ad290),
	.w2(32'hb839ec08),
	.w3(32'h3a89dfef),
	.w4(32'h3987c775),
	.w5(32'hbb078d12),
	.w6(32'h3a1e6151),
	.w7(32'h39cdcbc6),
	.w8(32'h38806cae),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66fc9e),
	.w1(32'h3af7687d),
	.w2(32'h3ae4db29),
	.w3(32'hb680ced9),
	.w4(32'h3aa860d6),
	.w5(32'h3b1b6ae6),
	.w6(32'hba8af7ef),
	.w7(32'h3ac863ed),
	.w8(32'h3b17fe8b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88a80a),
	.w1(32'h3a366f39),
	.w2(32'hbaa824e5),
	.w3(32'h3b4c3e98),
	.w4(32'h390b080d),
	.w5(32'hbb829950),
	.w6(32'h3b5b0838),
	.w7(32'h3b5a602c),
	.w8(32'hbb2918cd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba915bd4),
	.w1(32'hbb393162),
	.w2(32'hbb8174af),
	.w3(32'hbaa02e4e),
	.w4(32'hbaddba97),
	.w5(32'hbb059446),
	.w6(32'hba5cde20),
	.w7(32'h3a81a218),
	.w8(32'h39960767),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92046a3),
	.w1(32'hb7c4bd9e),
	.w2(32'h38e5540b),
	.w3(32'h38fa28f2),
	.w4(32'h39f0ccd4),
	.w5(32'hba644d69),
	.w6(32'hba28d1cc),
	.w7(32'h3a30f776),
	.w8(32'hb87d7aad),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d27609),
	.w1(32'hba31f2e0),
	.w2(32'hb9a522b5),
	.w3(32'h39e82347),
	.w4(32'h3b0aba57),
	.w5(32'h3af07e04),
	.w6(32'hba431a7d),
	.w7(32'h3ae5b417),
	.w8(32'h39d40f8c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f96e7),
	.w1(32'hbaa53ae1),
	.w2(32'hb98a2a28),
	.w3(32'h3a8ec711),
	.w4(32'hba9d46d9),
	.w5(32'hbb218c55),
	.w6(32'h3a7fd7b2),
	.w7(32'hba3ff8dd),
	.w8(32'h3aa5619d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdc487),
	.w1(32'hb99d4383),
	.w2(32'hbaad530c),
	.w3(32'h39f19ffd),
	.w4(32'hba7e6941),
	.w5(32'hba3cef9e),
	.w6(32'hb85ec39d),
	.w7(32'h391f17bf),
	.w8(32'hb91ab959),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab23324),
	.w1(32'hbb2d304f),
	.w2(32'hbb351e15),
	.w3(32'h3956b9ed),
	.w4(32'hbababc6f),
	.w5(32'hb87d2ce7),
	.w6(32'hb9096232),
	.w7(32'hbaec4fa0),
	.w8(32'hbb40cb63),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1b07d),
	.w1(32'hbaea5a67),
	.w2(32'hbb526468),
	.w3(32'hba1de43f),
	.w4(32'h3ad91430),
	.w5(32'hbb309685),
	.w6(32'hb9e03655),
	.w7(32'h3a5ba6a6),
	.w8(32'hbafdbf37),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994604),
	.w1(32'hb9ad15fe),
	.w2(32'hba81bffe),
	.w3(32'hb9158255),
	.w4(32'h3a86c06c),
	.w5(32'hba310a81),
	.w6(32'hba151f35),
	.w7(32'hb92f1a9b),
	.w8(32'hba9fa4b4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8ebb5),
	.w1(32'hba328781),
	.w2(32'hbb07bdda),
	.w3(32'hbacde628),
	.w4(32'hbaad3289),
	.w5(32'hbb9fe575),
	.w6(32'hba747c24),
	.w7(32'hba8c1c36),
	.w8(32'hbafc4785),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacb905),
	.w1(32'hbb2e9609),
	.w2(32'hbb2ca227),
	.w3(32'hbb2ca4a3),
	.w4(32'h399fb35e),
	.w5(32'hbaf12067),
	.w6(32'h395cdc26),
	.w7(32'h3b00a3d9),
	.w8(32'hbaae748e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97de9e),
	.w1(32'h3a8215d0),
	.w2(32'h3ae557fe),
	.w3(32'hba84ca71),
	.w4(32'h3adc7904),
	.w5(32'h3ae3a233),
	.w6(32'hbafe86c3),
	.w7(32'h3a3c710c),
	.w8(32'h3aa9d642),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71ea4f),
	.w1(32'hba6ccc12),
	.w2(32'hbadb781b),
	.w3(32'h3a1941f1),
	.w4(32'h3a185d47),
	.w5(32'hb9e72c25),
	.w6(32'h3a3ec2c6),
	.w7(32'h3afccd78),
	.w8(32'h397fe7c9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce8cc),
	.w1(32'h3a22176b),
	.w2(32'h3a8930d2),
	.w3(32'hba90cedf),
	.w4(32'h3a5626f1),
	.w5(32'hbb19d061),
	.w6(32'h39e0855f),
	.w7(32'h3af9b264),
	.w8(32'h39ac2c10),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73767e),
	.w1(32'h39a81c7f),
	.w2(32'hb90c0c2f),
	.w3(32'h3b0067dc),
	.w4(32'hb85801f8),
	.w5(32'h3ae69b8f),
	.w6(32'hba3cc041),
	.w7(32'hbab5dfa3),
	.w8(32'h392dd318),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d7ac5),
	.w1(32'hbab919c9),
	.w2(32'hb97f11ec),
	.w3(32'h39b2e27b),
	.w4(32'h38fe256a),
	.w5(32'h3abf0610),
	.w6(32'hb928e0fc),
	.w7(32'h3a670bbc),
	.w8(32'h3985eeb1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3929a4de),
	.w1(32'hb9c10f10),
	.w2(32'hb8fec679),
	.w3(32'h3aa22d3a),
	.w4(32'h363fb98c),
	.w5(32'hba151b7b),
	.w6(32'h3a9baa92),
	.w7(32'h3a0817d8),
	.w8(32'h39e28fd6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a7a11),
	.w1(32'h3986daaf),
	.w2(32'h379c0568),
	.w3(32'hb9c6a681),
	.w4(32'h3a27e9cb),
	.w5(32'h3970910f),
	.w6(32'hb9e9b4eb),
	.w7(32'h39c7d48d),
	.w8(32'h3543b8f5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab17e0d),
	.w1(32'h361a56d4),
	.w2(32'h3a9221d4),
	.w3(32'h3998fd55),
	.w4(32'hb9ad0d15),
	.w5(32'h3892d130),
	.w6(32'h3a377046),
	.w7(32'h3a9fb19f),
	.w8(32'h3af600a3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f8540),
	.w1(32'h3a1e6108),
	.w2(32'h3a92e04c),
	.w3(32'h386cd97a),
	.w4(32'h3a6b84b2),
	.w5(32'hb97a183f),
	.w6(32'hba8bfbe7),
	.w7(32'hba218556),
	.w8(32'hba83f26b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01afba),
	.w1(32'hba6f5672),
	.w2(32'hbabc4add),
	.w3(32'hba86637e),
	.w4(32'h3aad2f3f),
	.w5(32'hba7e07d6),
	.w6(32'h3b045c44),
	.w7(32'h3b3f2421),
	.w8(32'hb905630b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394886d9),
	.w1(32'h3a74a0af),
	.w2(32'h39a166b5),
	.w3(32'hba3520f8),
	.w4(32'hb9c40851),
	.w5(32'hb9c622a1),
	.w6(32'hb9372a0e),
	.w7(32'h38684d16),
	.w8(32'hbaa1f112),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a6da7),
	.w1(32'hbb245c9b),
	.w2(32'hbb45fd6f),
	.w3(32'hba68f5a1),
	.w4(32'hbb269ba0),
	.w5(32'h38da6fe2),
	.w6(32'h3ae4bd7d),
	.w7(32'hba672013),
	.w8(32'hbab97375),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b019c5b),
	.w1(32'hba8780dc),
	.w2(32'hbb0635a0),
	.w3(32'h3b133e39),
	.w4(32'hba4f36db),
	.w5(32'hbb192765),
	.w6(32'h38e97228),
	.w7(32'hbadaf0a8),
	.w8(32'hbb82e28f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e866),
	.w1(32'hbad460ad),
	.w2(32'hbb6bfe1b),
	.w3(32'h38095ab5),
	.w4(32'h3a7f1ff3),
	.w5(32'hbb327740),
	.w6(32'hbb073b06),
	.w7(32'h3b25c76c),
	.w8(32'hba212ae7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98a613),
	.w1(32'h3aa96fea),
	.w2(32'hbb4d5c49),
	.w3(32'h3ae9e730),
	.w4(32'h3a61e47e),
	.w5(32'hb91e6d8d),
	.w6(32'h3b31d607),
	.w7(32'hb862aa38),
	.w8(32'h3af900cb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72f346),
	.w1(32'hba7f262d),
	.w2(32'hb773e56d),
	.w3(32'hba8658d4),
	.w4(32'hbab104fe),
	.w5(32'h39aa6901),
	.w6(32'hba1f611f),
	.w7(32'hbaea6b06),
	.w8(32'hba86f010),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea921),
	.w1(32'h39731620),
	.w2(32'h3b24208b),
	.w3(32'h3b294086),
	.w4(32'h3b050432),
	.w5(32'h3b0a2445),
	.w6(32'h3b794bed),
	.w7(32'h3b41867a),
	.w8(32'h3b2d898f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadda365),
	.w1(32'hbae1fac9),
	.w2(32'hba25daa9),
	.w3(32'hba903ba0),
	.w4(32'hba971ca4),
	.w5(32'hbae98d9c),
	.w6(32'h3912d462),
	.w7(32'h39b98dec),
	.w8(32'h3a8009dc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb775136),
	.w1(32'hbb053752),
	.w2(32'h3a96b8a2),
	.w3(32'hbaacfd1b),
	.w4(32'hba357cff),
	.w5(32'hba17c90a),
	.w6(32'hbace52a5),
	.w7(32'hbb507bde),
	.w8(32'hbb33c816),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c661),
	.w1(32'h3b12ca2a),
	.w2(32'h3b13c9e3),
	.w3(32'h3af97f30),
	.w4(32'h3aa04fe0),
	.w5(32'h3b239c0e),
	.w6(32'hb9a444fd),
	.w7(32'hb888ce60),
	.w8(32'h39b19d10),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4796d2),
	.w1(32'hba944b0f),
	.w2(32'hb9e7b56e),
	.w3(32'hbaaa0c91),
	.w4(32'h3a03435e),
	.w5(32'h3a7f47ca),
	.w6(32'hba6835a0),
	.w7(32'h3a636333),
	.w8(32'h398b5032),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47ba5a),
	.w1(32'hba94b482),
	.w2(32'hb9f7e05c),
	.w3(32'h3a57c8b6),
	.w4(32'h3aa56a76),
	.w5(32'hba1f6486),
	.w6(32'hb999f179),
	.w7(32'h3a48d148),
	.w8(32'h3a19f1b4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fbb17),
	.w1(32'hbb175ec8),
	.w2(32'hba3d1a28),
	.w3(32'h3957cd39),
	.w4(32'hb903ff4e),
	.w5(32'hb89e5764),
	.w6(32'h3a866556),
	.w7(32'h39e79881),
	.w8(32'h39b3b8cc),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ee18b),
	.w1(32'hb9fbdd4f),
	.w2(32'h3a481ae9),
	.w3(32'h389de8b0),
	.w4(32'hb97e1bc8),
	.w5(32'hbb1e29f7),
	.w6(32'hb9f45cba),
	.w7(32'hb9e34284),
	.w8(32'hba73b7d3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84e282),
	.w1(32'h3a2db964),
	.w2(32'h3a32d36b),
	.w3(32'h3a11c472),
	.w4(32'h394431d1),
	.w5(32'h3accfd6d),
	.w6(32'hb98e5e33),
	.w7(32'h3b00586f),
	.w8(32'h3ad3f5f1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b6b39),
	.w1(32'h373d8e2e),
	.w2(32'h3a2f3011),
	.w3(32'h3b00615f),
	.w4(32'h39c0669e),
	.w5(32'hb940be2b),
	.w6(32'h3a98badd),
	.w7(32'h3a1b3994),
	.w8(32'h3a815bff),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5cc98),
	.w1(32'h3b74ca33),
	.w2(32'h3adbc8e4),
	.w3(32'h3b9d1a22),
	.w4(32'h3b20e1ed),
	.w5(32'h39c2349e),
	.w6(32'h3bb340b5),
	.w7(32'h3ab0f0ab),
	.w8(32'hba299807),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97dc2a),
	.w1(32'hba034a85),
	.w2(32'h37acc08b),
	.w3(32'hb9636aaf),
	.w4(32'h3aea24c3),
	.w5(32'h3aa9f1c1),
	.w6(32'h3914320e),
	.w7(32'h3a5bebe9),
	.w8(32'h3a908239),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acba670),
	.w1(32'hb9eb4ea4),
	.w2(32'h390eaed0),
	.w3(32'h3b033d4e),
	.w4(32'hba969c6c),
	.w5(32'hba30efc8),
	.w6(32'h3a9117f0),
	.w7(32'hbacdb0dc),
	.w8(32'hb970937f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe0ff6),
	.w1(32'hbb113806),
	.w2(32'hba4f9992),
	.w3(32'h3a7556f6),
	.w4(32'h3acc0f13),
	.w5(32'h3a9cec29),
	.w6(32'h39c4b578),
	.w7(32'h3a8c10ab),
	.w8(32'h3b213ee8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3374a0),
	.w1(32'h39aca91e),
	.w2(32'hbae8e434),
	.w3(32'hbb2a1dc1),
	.w4(32'h3a25af98),
	.w5(32'h3a238a00),
	.w6(32'hbb668def),
	.w7(32'h3b05bca0),
	.w8(32'h39e440d5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e0fda),
	.w1(32'h3ad9f8b8),
	.w2(32'h3ac49c13),
	.w3(32'h3b5eebb6),
	.w4(32'h3a98b2e0),
	.w5(32'hba9501d5),
	.w6(32'h3b6738a2),
	.w7(32'h3ab5a261),
	.w8(32'hb8c8de8b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906d7c3),
	.w1(32'hba2b37f8),
	.w2(32'hbb8e04c0),
	.w3(32'hba44504f),
	.w4(32'h39c325e9),
	.w5(32'hbba56ca0),
	.w6(32'h3b210212),
	.w7(32'h3b42740e),
	.w8(32'h38caf3ab),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dc998),
	.w1(32'h3a7e6373),
	.w2(32'h39e0e78c),
	.w3(32'hb78a03f8),
	.w4(32'hba41e6d5),
	.w5(32'hb7623adc),
	.w6(32'hbaf59741),
	.w7(32'hba5b2228),
	.w8(32'hb8cd65d5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b6e9),
	.w1(32'hb9b87af0),
	.w2(32'hbb670df3),
	.w3(32'h3ac7f9ce),
	.w4(32'h3a6fc63b),
	.w5(32'hbb4da04e),
	.w6(32'h3b3dd583),
	.w7(32'h3b2eacb2),
	.w8(32'h38946b54),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750928),
	.w1(32'hbb427a90),
	.w2(32'hbb88d4d5),
	.w3(32'hbaf9c2e5),
	.w4(32'hba14283a),
	.w5(32'hbafbd5e7),
	.w6(32'hba9307ba),
	.w7(32'hb9571680),
	.w8(32'hba9966a4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3fcb9),
	.w1(32'hbb4a6306),
	.w2(32'hbb7cfb16),
	.w3(32'hbb4b4f74),
	.w4(32'hb96949cd),
	.w5(32'hbb42ca54),
	.w6(32'hbaa64c3c),
	.w7(32'h3b0eb4c8),
	.w8(32'hbafcd192),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108587),
	.w1(32'hb97a51cd),
	.w2(32'h3acf168c),
	.w3(32'h3ab5f900),
	.w4(32'h3a6bf7cd),
	.w5(32'h39ac951a),
	.w6(32'h3a0fd630),
	.w7(32'h3a80d6d8),
	.w8(32'h3ab701d6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab18315),
	.w1(32'hba1e3dff),
	.w2(32'hbaccdfe3),
	.w3(32'h38b72b0d),
	.w4(32'hba4b8637),
	.w5(32'hba9cd0f0),
	.w6(32'h3a3c505c),
	.w7(32'h389804da),
	.w8(32'hba7ca1fc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2882ea),
	.w1(32'h3944be7f),
	.w2(32'hb7da3bbf),
	.w3(32'hba99d565),
	.w4(32'h3a2eb98a),
	.w5(32'h38e42466),
	.w6(32'h397673b4),
	.w7(32'h3a6e64df),
	.w8(32'h3a915560),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3a894),
	.w1(32'h3a6f06e5),
	.w2(32'hb99a4784),
	.w3(32'h3a07d2b6),
	.w4(32'h3a55cd10),
	.w5(32'hb9e5b268),
	.w6(32'h3ad527c1),
	.w7(32'h3b24b86f),
	.w8(32'h39db6085),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf8ee9),
	.w1(32'hbad62216),
	.w2(32'hb819bf4c),
	.w3(32'h3a2c8aaf),
	.w4(32'hba0d646b),
	.w5(32'h3a401256),
	.w6(32'h39be41b1),
	.w7(32'hbad07c46),
	.w8(32'hba5acd8a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c61382),
	.w1(32'h39807f60),
	.w2(32'hbb0af7f0),
	.w3(32'h39c89a66),
	.w4(32'h399b2f44),
	.w5(32'hbadd8e66),
	.w6(32'hba341da8),
	.w7(32'hba6703b1),
	.w8(32'hba9ceba2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad411c),
	.w1(32'hba4d906f),
	.w2(32'hba510b6e),
	.w3(32'hba50cb7a),
	.w4(32'h39c52ed9),
	.w5(32'hb9996155),
	.w6(32'hb8796add),
	.w7(32'hb90f4254),
	.w8(32'hb98940b1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c7cc8),
	.w1(32'hbaa7fdc5),
	.w2(32'hb936ca71),
	.w3(32'hba778ca5),
	.w4(32'h3ae7df0c),
	.w5(32'h3a7d13bb),
	.w6(32'hba8d7d06),
	.w7(32'h3ac8d9d2),
	.w8(32'h3a8457cc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ecdb5d),
	.w1(32'hb84624a5),
	.w2(32'h3a14fa78),
	.w3(32'h39b104ad),
	.w4(32'h3a2a0370),
	.w5(32'h3a1c856c),
	.w6(32'hb9a5b78c),
	.w7(32'h3a23aa91),
	.w8(32'hb95f9085),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf59d34),
	.w1(32'hba95d3f4),
	.w2(32'hba48a78f),
	.w3(32'hba6b6e3c),
	.w4(32'hb7f85f88),
	.w5(32'h3a518e96),
	.w6(32'hba7f63fc),
	.w7(32'h39457f0f),
	.w8(32'hb9265bfb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d9c8),
	.w1(32'hb9b861d5),
	.w2(32'h3b302f74),
	.w3(32'hbafe0208),
	.w4(32'h396c1ca1),
	.w5(32'h3b1d36a1),
	.w6(32'hba3f99ae),
	.w7(32'h3a80f94a),
	.w8(32'h3a2637a7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b171186),
	.w1(32'h3a0993d0),
	.w2(32'hbab6bc8a),
	.w3(32'h3a95054f),
	.w4(32'h3904bf3d),
	.w5(32'hba12a20e),
	.w6(32'h3a928baf),
	.w7(32'hb9a64728),
	.w8(32'hbabe4973),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb884a79),
	.w1(32'hbb8f0445),
	.w2(32'hbc0a275a),
	.w3(32'h3b44d599),
	.w4(32'h3a9d6d54),
	.w5(32'hbbdad70d),
	.w6(32'h3bf33e7f),
	.w7(32'h3c0af465),
	.w8(32'h3b081627),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b7b29),
	.w1(32'hbb50c38a),
	.w2(32'hbb17a959),
	.w3(32'h38d90d5a),
	.w4(32'hbb0fd72e),
	.w5(32'h3a76cac7),
	.w6(32'hbaad10da),
	.w7(32'hbb316c5d),
	.w8(32'hbadb0290),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fce89),
	.w1(32'h3a416ea2),
	.w2(32'h3a9cf7dd),
	.w3(32'hba673b23),
	.w4(32'h3a1a94b8),
	.w5(32'hb92bc2e9),
	.w6(32'h3a357744),
	.w7(32'h39b382e0),
	.w8(32'hb994fd62),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cdff99),
	.w1(32'hba2bede9),
	.w2(32'hba2237ed),
	.w3(32'h3a54c64a),
	.w4(32'hbaa5e672),
	.w5(32'hbb24fcb7),
	.w6(32'h3a81b3ad),
	.w7(32'h398dd426),
	.w8(32'h3a980532),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf2fdb),
	.w1(32'h38dcf0ec),
	.w2(32'hba6f9c67),
	.w3(32'hba0a1017),
	.w4(32'hba1e0a01),
	.w5(32'hba161ce7),
	.w6(32'hb9db0ae5),
	.w7(32'h38995b57),
	.w8(32'hb9ff6154),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9387d2f),
	.w1(32'h39f74fc4),
	.w2(32'hb8c32f34),
	.w3(32'h39d4bda0),
	.w4(32'hb902407f),
	.w5(32'hba326af1),
	.w6(32'h38ff6bfc),
	.w7(32'hb9426880),
	.w8(32'hb941e857),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07856f),
	.w1(32'h3adc815b),
	.w2(32'h3b0eab04),
	.w3(32'hba278e84),
	.w4(32'h3a42862f),
	.w5(32'hba46f4e3),
	.w6(32'hb95817fd),
	.w7(32'h3ad7c9cc),
	.w8(32'hb9795216),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fc5d6),
	.w1(32'hbabf57c7),
	.w2(32'hbaa6a27e),
	.w3(32'hbb18c691),
	.w4(32'hbab58989),
	.w5(32'hbad250d9),
	.w6(32'hba6d14f8),
	.w7(32'hbabf3c1e),
	.w8(32'hbb0d6dd4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bf1c55),
	.w1(32'h3a5415b5),
	.w2(32'h3b21e134),
	.w3(32'h3a4e6f02),
	.w4(32'h3b0fdaa4),
	.w5(32'h3a0fa6b3),
	.w6(32'h3b034be2),
	.w7(32'h3b8ed778),
	.w8(32'h3b449037),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6045c),
	.w1(32'hba959cd8),
	.w2(32'h3aba8952),
	.w3(32'h3975ad81),
	.w4(32'hba4b2b68),
	.w5(32'h3a4ef6c3),
	.w6(32'h3ac4264f),
	.w7(32'hba59c68c),
	.w8(32'h3aa035b7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0c23b),
	.w1(32'h3b9545eb),
	.w2(32'hbbe0b995),
	.w3(32'h3b7a3591),
	.w4(32'h3b9a58b6),
	.w5(32'hbc35db05),
	.w6(32'h3b7f5b24),
	.w7(32'h3bdcd759),
	.w8(32'hbc499ac6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63de51),
	.w1(32'hbbd3eb05),
	.w2(32'hba6c2411),
	.w3(32'hbc3764cb),
	.w4(32'hbb69eeef),
	.w5(32'hbbd5a33d),
	.w6(32'hbbd935af),
	.w7(32'hba29a60b),
	.w8(32'hbbe11b1c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24e1ad),
	.w1(32'h3b47e2fb),
	.w2(32'h3bdc1e84),
	.w3(32'hbc3c6256),
	.w4(32'h3b6f15ff),
	.w5(32'h3af283af),
	.w6(32'hbbe141db),
	.w7(32'hba8fa175),
	.w8(32'h3b0c5745),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d87c),
	.w1(32'hbaa0cae3),
	.w2(32'h3ab7d5f5),
	.w3(32'hbb0c8823),
	.w4(32'h3b359ee6),
	.w5(32'hbb494481),
	.w6(32'hbaac1388),
	.w7(32'hbac1107c),
	.w8(32'hbab30341),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15dc20),
	.w1(32'h36e25102),
	.w2(32'hbb318936),
	.w3(32'h3c262868),
	.w4(32'hb9382cb6),
	.w5(32'hbad7d8c7),
	.w6(32'h3b0ed59b),
	.w7(32'h3afbe399),
	.w8(32'hbb059975),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b955),
	.w1(32'h3b6929a0),
	.w2(32'h3ba2dcb3),
	.w3(32'hb9c027c0),
	.w4(32'h3bc407aa),
	.w5(32'hbc1afe96),
	.w6(32'hbba90d25),
	.w7(32'h3c0432ce),
	.w8(32'h3b1e78a2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdc107),
	.w1(32'hbb8c75ea),
	.w2(32'hbb2ce924),
	.w3(32'hbb2bfdf0),
	.w4(32'hbb72ab2d),
	.w5(32'hbbb9e0f5),
	.w6(32'h3c26ef8d),
	.w7(32'hbbcc91c7),
	.w8(32'hbbc1b10e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cf06d),
	.w1(32'hba1afb97),
	.w2(32'hbc6d20a3),
	.w3(32'h3ab0e7ce),
	.w4(32'h3b9b4488),
	.w5(32'hbc32b18c),
	.w6(32'hbb3485df),
	.w7(32'hbb313a36),
	.w8(32'hbc68488a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee66c2),
	.w1(32'h3b42adaa),
	.w2(32'hbbea40d4),
	.w3(32'hbb55a2a5),
	.w4(32'hbaca4be4),
	.w5(32'hbc95d225),
	.w6(32'hbbd3e700),
	.w7(32'hbb19d38f),
	.w8(32'hbbeb4781),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec3687),
	.w1(32'hbb8437cd),
	.w2(32'hbb949ed1),
	.w3(32'hbc05b2e6),
	.w4(32'hbba5d6c2),
	.w5(32'hbb5f4124),
	.w6(32'hbc526ea6),
	.w7(32'hbbc2afea),
	.w8(32'hbb551676),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eb923),
	.w1(32'hbb3580b2),
	.w2(32'hbc8567fd),
	.w3(32'hbad5b13a),
	.w4(32'hbaa6ce63),
	.w5(32'hbcb52c80),
	.w6(32'h3b0c6afb),
	.w7(32'hbb40a4a7),
	.w8(32'hbc9f4a1a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0cd6c),
	.w1(32'hbc2cfed2),
	.w2(32'hba954f01),
	.w3(32'hbb60f0ee),
	.w4(32'hbbdc2748),
	.w5(32'h3bd2576a),
	.w6(32'hbc2611e4),
	.w7(32'hbbb8c02e),
	.w8(32'h3c020d51),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafdcf4),
	.w1(32'h3bb76f5e),
	.w2(32'hba99d0cb),
	.w3(32'h3b12949c),
	.w4(32'h3b66d17e),
	.w5(32'hbb0a6df6),
	.w6(32'hb99fb828),
	.w7(32'h3b819c21),
	.w8(32'hbb949d6c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbf0d9),
	.w1(32'hbb0456d8),
	.w2(32'h3b6d83b6),
	.w3(32'h3ae8803c),
	.w4(32'hbb88a140),
	.w5(32'h3acac46b),
	.w6(32'hbb30799b),
	.w7(32'hbc075bae),
	.w8(32'hbbc367e7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7a0f6),
	.w1(32'h3aa2037c),
	.w2(32'h3c4ce74e),
	.w3(32'hbaeb7226),
	.w4(32'h3c2aac60),
	.w5(32'h3c185b22),
	.w6(32'hbb8bf79e),
	.w7(32'h3c2d59b9),
	.w8(32'h3bc4e77e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e6d5c),
	.w1(32'hbad95e47),
	.w2(32'hbbd8e256),
	.w3(32'hba8fd15c),
	.w4(32'h3a8cafbe),
	.w5(32'hbba6f8cb),
	.w6(32'h3be1385f),
	.w7(32'h3a28de42),
	.w8(32'hbbd69159),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01fbcb),
	.w1(32'hbaa22ea9),
	.w2(32'hbb57b5fe),
	.w3(32'h3b5e3618),
	.w4(32'h3a89e6e8),
	.w5(32'hbbfc3d6c),
	.w6(32'h3a07f7c8),
	.w7(32'hbc0fe8f8),
	.w8(32'hbbc2c91e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae793e),
	.w1(32'h3bfb5a9e),
	.w2(32'h3c62a896),
	.w3(32'h3be47601),
	.w4(32'h3c2d8f45),
	.w5(32'h3c5d4556),
	.w6(32'h3c44d55d),
	.w7(32'h3b8e9e75),
	.w8(32'h3bbe4341),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96a1a2),
	.w1(32'h3b347164),
	.w2(32'hbb053191),
	.w3(32'h3b1247b0),
	.w4(32'h3b9aa677),
	.w5(32'hbc382436),
	.w6(32'h3b9ab9f1),
	.w7(32'h3a95075b),
	.w8(32'hbb6320b5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ac2a),
	.w1(32'h398596d3),
	.w2(32'hbb786b26),
	.w3(32'hbbc9d2d1),
	.w4(32'hbbefaf9f),
	.w5(32'hbb67cb08),
	.w6(32'hb9b6dc01),
	.w7(32'hbbacfe66),
	.w8(32'hbc11c102),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968cf7c),
	.w1(32'h3ae424cf),
	.w2(32'hbb31e6a1),
	.w3(32'hbc39feaf),
	.w4(32'hbaef1829),
	.w5(32'hbbc08da8),
	.w6(32'hbbe6680e),
	.w7(32'hba25e51f),
	.w8(32'hbc3bcaf7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf127e1),
	.w1(32'h3b503dfb),
	.w2(32'h3b03e188),
	.w3(32'hbbffb093),
	.w4(32'hba2d675f),
	.w5(32'h3bd6749f),
	.w6(32'hbba59d56),
	.w7(32'h3bb4def2),
	.w8(32'h3baf9139),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29fec1),
	.w1(32'hbaf78a50),
	.w2(32'h3ac936c8),
	.w3(32'hbbf93065),
	.w4(32'h3ad1a6b0),
	.w5(32'hbb1d2278),
	.w6(32'hbc01f90a),
	.w7(32'h3a864974),
	.w8(32'hbb14161e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9109f7),
	.w1(32'hbb4ebe98),
	.w2(32'h3c0dc55e),
	.w3(32'hbc0410bf),
	.w4(32'h3a8e1b22),
	.w5(32'h3c068b3c),
	.w6(32'hbb4baa81),
	.w7(32'hbb554576),
	.w8(32'h3b94613e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a068310),
	.w1(32'hbc058f1d),
	.w2(32'hbb6d1c54),
	.w3(32'h3bb67694),
	.w4(32'hbb83886d),
	.w5(32'h3c1bd1f7),
	.w6(32'h3bc6e9e8),
	.w7(32'hbb82f09d),
	.w8(32'h3b82f61a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23ed05),
	.w1(32'hbb7b8f3c),
	.w2(32'h3b58e286),
	.w3(32'h3bb83dc3),
	.w4(32'h3a91f03b),
	.w5(32'hbc577f93),
	.w6(32'h3b76de81),
	.w7(32'hbbb78388),
	.w8(32'hbc1ae269),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f8a3),
	.w1(32'h3ac71d52),
	.w2(32'h3c22ae70),
	.w3(32'hbb10de5a),
	.w4(32'hba87e1ac),
	.w5(32'h3cc98568),
	.w6(32'hbc22f031),
	.w7(32'h3bd17f5b),
	.w8(32'h3c84fa45),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be28660),
	.w1(32'h3a972cf6),
	.w2(32'h3b3c364b),
	.w3(32'h3bd38397),
	.w4(32'hb9dc9a26),
	.w5(32'hbb09034f),
	.w6(32'h3bc6f36d),
	.w7(32'h3999cf67),
	.w8(32'hbbd68414),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba714bce),
	.w1(32'h3bd0b30a),
	.w2(32'h3b34cc38),
	.w3(32'h3741d225),
	.w4(32'h3bdd80b5),
	.w5(32'h3b5644c6),
	.w6(32'hb9103d27),
	.w7(32'h3bcac7ac),
	.w8(32'h3929aa50),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2150da),
	.w1(32'hba9b43d2),
	.w2(32'hbb6a918a),
	.w3(32'h3af1aa85),
	.w4(32'hbba926e1),
	.w5(32'hbb6a613c),
	.w6(32'h3a4c5ddf),
	.w7(32'hbc2e3bfa),
	.w8(32'hbbce8354),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee58ee),
	.w1(32'hbb0e91cd),
	.w2(32'hbc223ecf),
	.w3(32'hbbc1751b),
	.w4(32'hbba28158),
	.w5(32'hbc24698c),
	.w6(32'hbbefa1f3),
	.w7(32'h3b05ea84),
	.w8(32'hbabc3ec0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cddcf),
	.w1(32'hbb645923),
	.w2(32'h3a23a3e7),
	.w3(32'hbb897b3c),
	.w4(32'hbaf8d8a7),
	.w5(32'hbba3d9e2),
	.w6(32'hbb9bf44a),
	.w7(32'hbb530d66),
	.w8(32'hbba6dbf7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3cbb9),
	.w1(32'hbba33b52),
	.w2(32'hbad360a7),
	.w3(32'hbbb63cf5),
	.w4(32'hbba5a0fe),
	.w5(32'hba2cebe0),
	.w6(32'hbb76a228),
	.w7(32'hbac62a62),
	.w8(32'hbb9f7521),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bab5a),
	.w1(32'hbb1140f8),
	.w2(32'h3b76fd68),
	.w3(32'hbbcecf2c),
	.w4(32'hbbc0df91),
	.w5(32'h3a75ec46),
	.w6(32'hbb586ebf),
	.w7(32'hbbf4e8c0),
	.w8(32'h3a7417b6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dd565),
	.w1(32'h3b0a3fc8),
	.w2(32'h3aa13788),
	.w3(32'hbaa2ae76),
	.w4(32'hb96d6daa),
	.w5(32'h39aad840),
	.w6(32'hbb830276),
	.w7(32'hba56552d),
	.w8(32'hbae4212e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658567),
	.w1(32'hbb23fcbb),
	.w2(32'hbbac55af),
	.w3(32'hb743cb9f),
	.w4(32'hbb3fbdcc),
	.w5(32'hbc13e903),
	.w6(32'hb9b9881f),
	.w7(32'hbba3232c),
	.w8(32'hbc0c1a99),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0ddb),
	.w1(32'h39ffdac5),
	.w2(32'hbb6a1012),
	.w3(32'hbba21648),
	.w4(32'h3b50595a),
	.w5(32'hbb819716),
	.w6(32'h3a29918a),
	.w7(32'hba1d73bd),
	.w8(32'hbbf4c6e8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa630a),
	.w1(32'h38ecddd5),
	.w2(32'hbb3c6ea6),
	.w3(32'h3a9033ca),
	.w4(32'hbb08703c),
	.w5(32'hbb585ed1),
	.w6(32'hba5d6bf1),
	.w7(32'hbaa50713),
	.w8(32'hbb84bccc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe8c7),
	.w1(32'hbbba6b54),
	.w2(32'hbb2f77c2),
	.w3(32'hbb4043cf),
	.w4(32'h3a02a6f3),
	.w5(32'hbbacbcc5),
	.w6(32'hbb7e7f2f),
	.w7(32'h3b563646),
	.w8(32'hbbfc9285),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ff9b5),
	.w1(32'hbb156fa6),
	.w2(32'hbb89d330),
	.w3(32'hbc104b1a),
	.w4(32'hbaef11ce),
	.w5(32'hbc3eb1bd),
	.w6(32'hbc258da1),
	.w7(32'hbb9e9a48),
	.w8(32'hbb587783),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3676),
	.w1(32'h3ac44631),
	.w2(32'hb977b148),
	.w3(32'hbbe77ac4),
	.w4(32'h3b7a14d4),
	.w5(32'hbbecf567),
	.w6(32'hbb096d99),
	.w7(32'h3b34bd46),
	.w8(32'hbba2b4e1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba85482),
	.w1(32'h3af13e97),
	.w2(32'hbba53022),
	.w3(32'hbb349bdc),
	.w4(32'hbb781bd7),
	.w5(32'hbbe15469),
	.w6(32'hbb965a8d),
	.w7(32'hbab471cb),
	.w8(32'h3b8634d4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac87a6f),
	.w1(32'hbb6d8e71),
	.w2(32'hbc42ddb6),
	.w3(32'h3bdc50fd),
	.w4(32'h3a5d1047),
	.w5(32'hbbf6a2b2),
	.w6(32'h3bff3a9c),
	.w7(32'hbbc70086),
	.w8(32'hbc12361d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe8dcc),
	.w1(32'hbb2da26e),
	.w2(32'hbc543b1c),
	.w3(32'hbb404fe1),
	.w4(32'h3b8b7402),
	.w5(32'hbb6a4e10),
	.w6(32'h3a528510),
	.w7(32'h3c146115),
	.w8(32'hbae83c6d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ae33),
	.w1(32'hbb2b4707),
	.w2(32'h3b7888b9),
	.w3(32'hbb7cc378),
	.w4(32'hbba25bd5),
	.w5(32'h3bd17a75),
	.w6(32'hbb20d6ac),
	.w7(32'hbaabd64b),
	.w8(32'hbae06516),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ee9e7),
	.w1(32'h3b844fea),
	.w2(32'h3af5284f),
	.w3(32'h39bb441a),
	.w4(32'h3c1a5b1d),
	.w5(32'h3c1a3e7b),
	.w6(32'hbbd856a5),
	.w7(32'h3bf63c83),
	.w8(32'h3b0cfe82),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9da7b),
	.w1(32'h3ad3e780),
	.w2(32'h3a06bdd2),
	.w3(32'hbc117b94),
	.w4(32'h3ba2391f),
	.w5(32'h3b13265e),
	.w6(32'hbc24563b),
	.w7(32'h3bc3ea37),
	.w8(32'hbade687d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed2c1),
	.w1(32'h3bd95f7a),
	.w2(32'h3c136ac2),
	.w3(32'hbaa7dac0),
	.w4(32'h3c393a80),
	.w5(32'h3c5accf9),
	.w6(32'hbac69cf2),
	.w7(32'h3c28a049),
	.w8(32'h3c08b9f4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9f61),
	.w1(32'h3aae4b4e),
	.w2(32'hb9696877),
	.w3(32'h398ae6f6),
	.w4(32'h3b00c2da),
	.w5(32'h3c0e0f98),
	.w6(32'hbab6cff7),
	.w7(32'hbacdf7c3),
	.w8(32'h3acaed34),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81d65f),
	.w1(32'hbb8d414f),
	.w2(32'h3b26e1e8),
	.w3(32'h3bafd1df),
	.w4(32'hbb830962),
	.w5(32'hbbe50e5f),
	.w6(32'hbbc1c07c),
	.w7(32'hbb19b2cf),
	.w8(32'hbb8d9f05),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4fe6c),
	.w1(32'hb9c076e4),
	.w2(32'hbb58591b),
	.w3(32'h3af9b741),
	.w4(32'h39cfd8de),
	.w5(32'h379c8b7c),
	.w6(32'hbb2384ed),
	.w7(32'hbb76e229),
	.w8(32'hbbdab87d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2daf5),
	.w1(32'hb89d1e0d),
	.w2(32'h3b415ed5),
	.w3(32'h3bdb533d),
	.w4(32'hbb045dc7),
	.w5(32'h3bdfb8a1),
	.w6(32'h3b8df3e3),
	.w7(32'hbae4005f),
	.w8(32'h3bb08246),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa40065),
	.w1(32'h3ba88085),
	.w2(32'hbbea5ebc),
	.w3(32'h3b0797c4),
	.w4(32'h39fdf7b9),
	.w5(32'hbc884cba),
	.w6(32'hb8eb9c91),
	.w7(32'hbb5368b2),
	.w8(32'hbc9247e0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69d567),
	.w1(32'hbb485b15),
	.w2(32'hbac20b7e),
	.w3(32'hbca0aea4),
	.w4(32'h3abd3870),
	.w5(32'hbb0f5722),
	.w6(32'hbc6f4a52),
	.w7(32'h3b01599d),
	.w8(32'hbb852daa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8061d1),
	.w1(32'hbb530a83),
	.w2(32'hbc3f3df4),
	.w3(32'hbb7592b4),
	.w4(32'hb9267038),
	.w5(32'hbc2db6c6),
	.w6(32'hbb22ec39),
	.w7(32'h3ad4ef44),
	.w8(32'hbc6b4a79),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc078338),
	.w1(32'h39ac27bf),
	.w2(32'hbac3a74f),
	.w3(32'hbbf5c40d),
	.w4(32'h3bcb3b54),
	.w5(32'hbc2b9b08),
	.w6(32'hbbb7e2c8),
	.w7(32'h3b00abca),
	.w8(32'hbb29c89f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87e2a8),
	.w1(32'hbb1c28d0),
	.w2(32'hbbfba87a),
	.w3(32'hbb675a1f),
	.w4(32'hbb8369d0),
	.w5(32'hbbd90703),
	.w6(32'hbbf713ff),
	.w7(32'hbbdc153c),
	.w8(32'hbb871443),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb035855),
	.w1(32'h390d4e42),
	.w2(32'hbc394609),
	.w3(32'hbac8f792),
	.w4(32'hbb111bc7),
	.w5(32'hbc5920e1),
	.w6(32'h3a81e4b0),
	.w7(32'hbbb18e82),
	.w8(32'hbc67966a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9581de),
	.w1(32'hbc058d0a),
	.w2(32'hbb70834b),
	.w3(32'hbca0b4c1),
	.w4(32'h3b0fee3f),
	.w5(32'h3a8f0d4f),
	.w6(32'hbc72291a),
	.w7(32'h3bb845c6),
	.w8(32'hba246474),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule