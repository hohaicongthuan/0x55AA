module layer_10_featuremap_32(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19f4ac),
	.w1(32'hbb379896),
	.w2(32'h3ad7b2d2),
	.w3(32'hbb94dfee),
	.w4(32'hba979099),
	.w5(32'h3b96ecd2),
	.w6(32'h3b0824f6),
	.w7(32'h3ba3cc13),
	.w8(32'h3bb1dd94),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba767dce),
	.w1(32'h3a1e5ed9),
	.w2(32'h3ba85cac),
	.w3(32'h3bd92719),
	.w4(32'h3ba43f1d),
	.w5(32'h3b85170e),
	.w6(32'h3b661001),
	.w7(32'h3b071f06),
	.w8(32'h3c17112a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e1426),
	.w1(32'h3b9696d4),
	.w2(32'h38a8588b),
	.w3(32'h3be579f7),
	.w4(32'h3b3f2b58),
	.w5(32'hbb7caf17),
	.w6(32'h3bb3626b),
	.w7(32'h3bad9731),
	.w8(32'hb98680f7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02cff0),
	.w1(32'h3ba0cd6d),
	.w2(32'h3b990ec7),
	.w3(32'h3956c192),
	.w4(32'hb9a1f615),
	.w5(32'h3b9b6d99),
	.w6(32'h3805fc86),
	.w7(32'h39a612bc),
	.w8(32'h3c16b0b6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a299ab7),
	.w1(32'h3bc48167),
	.w2(32'hbb2587a4),
	.w3(32'h3baa5ada),
	.w4(32'h3bfca8a3),
	.w5(32'h3af36af4),
	.w6(32'h3bf3a1e2),
	.w7(32'h390eebb8),
	.w8(32'h3b5d0654),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1a368),
	.w1(32'h3be295f6),
	.w2(32'hbbba3ce3),
	.w3(32'h3b66dc42),
	.w4(32'h3b63878b),
	.w5(32'h3c7fd59c),
	.w6(32'h3c28fffd),
	.w7(32'h3b944ff6),
	.w8(32'h3c4f2562),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bede7ea),
	.w1(32'h3b7e8dd1),
	.w2(32'hbaf19d31),
	.w3(32'h3d4e6e3f),
	.w4(32'h3d222aaa),
	.w5(32'h3a9e9140),
	.w6(32'h3d410ba6),
	.w7(32'h3d0d133a),
	.w8(32'h3b454758),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e256),
	.w1(32'hbb820b4c),
	.w2(32'h3abc4ea7),
	.w3(32'hbba38980),
	.w4(32'hbb106eec),
	.w5(32'h3ba21e01),
	.w6(32'h39f3d1cf),
	.w7(32'h3aae0e2c),
	.w8(32'hbae0e8e6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe0112),
	.w1(32'h3b0ecf8c),
	.w2(32'h3abf90ec),
	.w3(32'h3ab03722),
	.w4(32'h3b2f309e),
	.w5(32'hbae25b76),
	.w6(32'hbaa2ca15),
	.w7(32'h3b39ba46),
	.w8(32'h39b39f79),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002a77),
	.w1(32'hbb12ffcc),
	.w2(32'hbbf7c68d),
	.w3(32'h394763d5),
	.w4(32'h39937631),
	.w5(32'hbbdc07f0),
	.w6(32'h3a414f57),
	.w7(32'h3a8a27b0),
	.w8(32'hbc1019ee),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973c16),
	.w1(32'hbb8adc22),
	.w2(32'h389591b4),
	.w3(32'h3b88f4c8),
	.w4(32'h3ad3a1fc),
	.w5(32'hbbc024fd),
	.w6(32'h39e96bed),
	.w7(32'hbad074fa),
	.w8(32'h393c3235),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d99464),
	.w1(32'h39e425a8),
	.w2(32'hbc4116e7),
	.w3(32'hbb325475),
	.w4(32'hbb9e8f93),
	.w5(32'hbc62dffb),
	.w6(32'h3b0e0b52),
	.w7(32'hbbb63803),
	.w8(32'hbc30cb2f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b5cde),
	.w1(32'hbc8ce701),
	.w2(32'h3aa3ad67),
	.w3(32'hbc822937),
	.w4(32'hbc97d973),
	.w5(32'h3b8f04c8),
	.w6(32'hbc651a30),
	.w7(32'hbc8b3611),
	.w8(32'h3bb80d70),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bc918),
	.w1(32'h3b12fc84),
	.w2(32'h3b0ed97e),
	.w3(32'hba0ae678),
	.w4(32'h3be5e56b),
	.w5(32'h3b0563f5),
	.w6(32'h3b81125a),
	.w7(32'h3bb76625),
	.w8(32'h3b9a2969),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3d42),
	.w1(32'h3a67c54a),
	.w2(32'hb817f37a),
	.w3(32'hbb914180),
	.w4(32'hbba9e739),
	.w5(32'h3b12156a),
	.w6(32'hbaa0bc95),
	.w7(32'h3b27c8c3),
	.w8(32'h3aaa3563),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082e00),
	.w1(32'hbbeef58e),
	.w2(32'hba1b4f70),
	.w3(32'hbb621be3),
	.w4(32'hbbba3824),
	.w5(32'h3bd7d25d),
	.w6(32'h3a797361),
	.w7(32'hbb80d992),
	.w8(32'h3b888e7c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9b21),
	.w1(32'h3b9fc38f),
	.w2(32'hbad8f6d2),
	.w3(32'h3cd63851),
	.w4(32'h3ca22acc),
	.w5(32'h3a8aa477),
	.w6(32'h3cb004f9),
	.w7(32'h3c78111c),
	.w8(32'h3b814d3b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9473338),
	.w1(32'h3aa00ab2),
	.w2(32'h3a19d0ed),
	.w3(32'h3ac7779f),
	.w4(32'h3b4f184f),
	.w5(32'h3b9a1f6e),
	.w6(32'h3ba363ba),
	.w7(32'h3b579ea6),
	.w8(32'h3b062eba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa355),
	.w1(32'h3b2c75fe),
	.w2(32'hba30b28a),
	.w3(32'h3abc76b3),
	.w4(32'h3b0c66bf),
	.w5(32'hbb23e082),
	.w6(32'h3bf4c188),
	.w7(32'h3aed4f0f),
	.w8(32'h3b9ff878),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5de939),
	.w1(32'h3b822c6a),
	.w2(32'hba147d22),
	.w3(32'hbb37c301),
	.w4(32'hbb5e25d2),
	.w5(32'h3b1edb89),
	.w6(32'h392a0d2f),
	.w7(32'hb9b878ad),
	.w8(32'h3adb2de0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38529),
	.w1(32'h39dcc1bb),
	.w2(32'hbb824f74),
	.w3(32'h3b9a218f),
	.w4(32'hb8474090),
	.w5(32'hbb88a9af),
	.w6(32'h3b9e084a),
	.w7(32'hbb16fef7),
	.w8(32'hbb7ff421),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ede54),
	.w1(32'hbaf4d342),
	.w2(32'h3a813f26),
	.w3(32'hbb8c3776),
	.w4(32'hbb8a1146),
	.w5(32'hba372513),
	.w6(32'hbaac35e0),
	.w7(32'hbb476a9a),
	.w8(32'hb8ba4cfb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81cf5b),
	.w1(32'hbb2f070f),
	.w2(32'h3c9caa3d),
	.w3(32'hbbc2e771),
	.w4(32'hbae3b320),
	.w5(32'h3c6c5e21),
	.w6(32'hbb5e75f1),
	.w7(32'hb5d16076),
	.w8(32'h3c961177),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66cb5e),
	.w1(32'h3c81bfaf),
	.w2(32'hb9858708),
	.w3(32'h3bd45d03),
	.w4(32'h3c3c35ff),
	.w5(32'h3bb5281a),
	.w6(32'h3c2b52a2),
	.w7(32'h3c412a71),
	.w8(32'hb90d9d8d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc8acd),
	.w1(32'hb73d76eb),
	.w2(32'hb98ddc82),
	.w3(32'h3b89679d),
	.w4(32'hbb05eae9),
	.w5(32'hb9532b9f),
	.w6(32'h3bef629e),
	.w7(32'h3a871825),
	.w8(32'h3ae3c414),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fc02b),
	.w1(32'h3ac9c8f9),
	.w2(32'hb9cb2c54),
	.w3(32'hbb2d2ae6),
	.w4(32'hbb632524),
	.w5(32'hb9eafdb6),
	.w6(32'h3b246448),
	.w7(32'hbb99d2ac),
	.w8(32'h3af90a5d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb244bb3),
	.w1(32'h3ab67f57),
	.w2(32'hb777adb9),
	.w3(32'hbafba0fe),
	.w4(32'hbad0c765),
	.w5(32'hb768b8cc),
	.w6(32'h3b2e4a56),
	.w7(32'hbaf74719),
	.w8(32'hb6f12aaf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a0300),
	.w1(32'hb87d3e5b),
	.w2(32'hb901ed04),
	.w3(32'hb8bdef6f),
	.w4(32'hb8c1efb3),
	.w5(32'hb9143de6),
	.w6(32'hb90e7a33),
	.w7(32'hb8b9b08b),
	.w8(32'hb93ccb0b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848ea03),
	.w1(32'h39320662),
	.w2(32'h399a7848),
	.w3(32'hba2ce9b2),
	.w4(32'hb95cf33b),
	.w5(32'h38398cbb),
	.w6(32'hb9f21c33),
	.w7(32'hb9454579),
	.w8(32'hb81470f0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d40fa),
	.w1(32'h38cbc348),
	.w2(32'h39595e68),
	.w3(32'h39889367),
	.w4(32'h3696d832),
	.w5(32'h3943dbaa),
	.w6(32'h39601c6b),
	.w7(32'h390caf66),
	.w8(32'h393dd124),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a58cec),
	.w1(32'hb7252436),
	.w2(32'hb78d7aab),
	.w3(32'hb708a592),
	.w4(32'hb762782f),
	.w5(32'hb7bb0afe),
	.w6(32'h34f9a9d8),
	.w7(32'hb7419e9e),
	.w8(32'hb7bcef68),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f10ad6),
	.w1(32'hb7f7c303),
	.w2(32'hb7f6d7db),
	.w3(32'h38049547),
	.w4(32'hb81ba080),
	.w5(32'hb888b786),
	.w6(32'h36bd95ce),
	.w7(32'hb77b59d7),
	.w8(32'hb85a77a7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78c7570),
	.w1(32'hb8de9aa7),
	.w2(32'hb908c099),
	.w3(32'hb84a3c4e),
	.w4(32'hb978199f),
	.w5(32'hb93828a7),
	.w6(32'h38e0d101),
	.w7(32'hb8a59f19),
	.w8(32'hb916f0b4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39674317),
	.w1(32'h38b72c81),
	.w2(32'h38e867f4),
	.w3(32'h393aac77),
	.w4(32'h38ff1d4d),
	.w5(32'h393cf4a3),
	.w6(32'h35d3de1f),
	.w7(32'h38622379),
	.w8(32'h391df05f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71226c2),
	.w1(32'hb790d53a),
	.w2(32'hb71c7417),
	.w3(32'hb7285028),
	.w4(32'hb702df2a),
	.w5(32'hb6c131b3),
	.w6(32'hb6fdc051),
	.w7(32'hb67cef92),
	.w8(32'hb6cbcb05),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c6b16b),
	.w1(32'hb70aa03a),
	.w2(32'hb7e39c0a),
	.w3(32'h37f22d54),
	.w4(32'hb727159b),
	.w5(32'hb868a95f),
	.w6(32'h3807315b),
	.w7(32'h370f6f43),
	.w8(32'hb830447c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7410d3),
	.w1(32'hb93f6286),
	.w2(32'hb90886aa),
	.w3(32'h3a5a93fd),
	.w4(32'hb81680e3),
	.w5(32'hb85c3430),
	.w6(32'h39e25510),
	.w7(32'hb8c5be1b),
	.w8(32'h38b01594),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c182ca),
	.w1(32'hb9097e58),
	.w2(32'hba07ac72),
	.w3(32'hb9fca862),
	.w4(32'hba168875),
	.w5(32'hba1b5b2b),
	.w6(32'h3984365e),
	.w7(32'hb7bfd070),
	.w8(32'hb9d82959),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aee29a),
	.w1(32'hb8203b90),
	.w2(32'hb842080a),
	.w3(32'hb988d771),
	.w4(32'hb8a2b417),
	.w5(32'h38613966),
	.w6(32'hba09c910),
	.w7(32'hb9d7eff1),
	.w8(32'hb9a27f31),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3792aa0f),
	.w1(32'h378150be),
	.w2(32'h37b968bb),
	.w3(32'h3798f247),
	.w4(32'h37abab12),
	.w5(32'h381b3356),
	.w6(32'h370a0581),
	.w7(32'h37492acb),
	.w8(32'h37a8b97f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908f1ae),
	.w1(32'h38e25879),
	.w2(32'h3930d3da),
	.w3(32'h3897737a),
	.w4(32'h38a0c9f1),
	.w5(32'h3953311e),
	.w6(32'h38fd12f8),
	.w7(32'h385c4fe3),
	.w8(32'h396fc94d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8504d90),
	.w1(32'hb85c906c),
	.w2(32'hb84426ce),
	.w3(32'hb820424a),
	.w4(32'hb80e5952),
	.w5(32'hb7ddb72b),
	.w6(32'hb8b5d570),
	.w7(32'hb8c7b328),
	.w8(32'hb816c1a6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb704ccee),
	.w1(32'hb9187847),
	.w2(32'hb88873f3),
	.w3(32'h37afaaae),
	.w4(32'hb928990d),
	.w5(32'hb8d3bc3c),
	.w6(32'h3766e4df),
	.w7(32'hb903ee32),
	.w8(32'hb8d530e7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f89d06),
	.w1(32'h389b8ec1),
	.w2(32'h39a949bd),
	.w3(32'hba2df114),
	.w4(32'hb9d987cf),
	.w5(32'h3a22bd29),
	.w6(32'hba124dd6),
	.w7(32'hb9f2f1e3),
	.w8(32'h394045b3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d6481),
	.w1(32'hb89103c4),
	.w2(32'h391dc616),
	.w3(32'h3921668e),
	.w4(32'hb8b7e260),
	.w5(32'h38d67585),
	.w6(32'h38afd250),
	.w7(32'hb8672862),
	.w8(32'h388b2697),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991075b),
	.w1(32'h3916b42e),
	.w2(32'h39bd2e49),
	.w3(32'h395108c5),
	.w4(32'h39313948),
	.w5(32'h39fbb6bf),
	.w6(32'hb9348825),
	.w7(32'hb80f2800),
	.w8(32'h3983636d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a280),
	.w1(32'h3a32c9e0),
	.w2(32'h3a3d21f3),
	.w3(32'h3a3477c9),
	.w4(32'h3a1c0a98),
	.w5(32'h3a2c92b7),
	.w6(32'h39baf604),
	.w7(32'h39f40e76),
	.w8(32'h3a43c83e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c13a17),
	.w1(32'h399e7876),
	.w2(32'h39d9b136),
	.w3(32'h3940c931),
	.w4(32'h3916d02f),
	.w5(32'h39b06c7f),
	.w6(32'h37ca55f1),
	.w7(32'h380e2d9f),
	.w8(32'h38da5c3f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a18aac),
	.w1(32'h373bcd84),
	.w2(32'h38e7c70d),
	.w3(32'hb94df551),
	.w4(32'h38b35edb),
	.w5(32'h3985f842),
	.w6(32'hb99bb82f),
	.w7(32'hb8bdea5e),
	.w8(32'h3911f304),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910abd1),
	.w1(32'h38c9cf65),
	.w2(32'h391e454e),
	.w3(32'h38f5e0b7),
	.w4(32'h397537ee),
	.w5(32'h3988e795),
	.w6(32'hb95ff0b6),
	.w7(32'hb8b4fa78),
	.w8(32'h38aa2a6e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91de77a),
	.w1(32'h38ad01c3),
	.w2(32'h3998d59e),
	.w3(32'hb962a0ad),
	.w4(32'hb8bda257),
	.w5(32'h393e463b),
	.w6(32'hb98bee3d),
	.w7(32'hb83bb3b6),
	.w8(32'h38565c43),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c4785f),
	.w1(32'hb83ddc0a),
	.w2(32'hb7c1aa21),
	.w3(32'hb8032a53),
	.w4(32'hb8191108),
	.w5(32'h36f7f44f),
	.w6(32'hb749a07b),
	.w7(32'hb78734ff),
	.w8(32'h37216f9a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38740757),
	.w1(32'h3830567b),
	.w2(32'h38b19d85),
	.w3(32'h38703d5f),
	.w4(32'h388a0ee4),
	.w5(32'h38f28f61),
	.w6(32'hb82df6cc),
	.w7(32'hb780d280),
	.w8(32'h36c4fdc2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882ea93),
	.w1(32'h38a2a795),
	.w2(32'h39555547),
	.w3(32'h38a63f46),
	.w4(32'h3892945a),
	.w5(32'h3909a3ee),
	.w6(32'hb8fe8d04),
	.w7(32'hb8dededa),
	.w8(32'hb73c6110),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f4d5e6),
	.w1(32'h38003242),
	.w2(32'h389ce0ac),
	.w3(32'hb898174c),
	.w4(32'h36589d9a),
	.w5(32'h385fd987),
	.w6(32'hb8b52303),
	.w7(32'hb7cd98f4),
	.w8(32'h374ef779),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369ba6b8),
	.w1(32'h36b875c2),
	.w2(32'h35dbed2c),
	.w3(32'hb680d553),
	.w4(32'hb64d89e5),
	.w5(32'hb56f873a),
	.w6(32'hb6886bb2),
	.w7(32'hb589c451),
	.w8(32'hb60673f7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356f8c3f),
	.w1(32'hb5b49565),
	.w2(32'hb65ca0ba),
	.w3(32'h361afb1a),
	.w4(32'h34dfa416),
	.w5(32'hb6da6d86),
	.w6(32'h36cf5833),
	.w7(32'h3689e622),
	.w8(32'hb56cbebf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a29fa),
	.w1(32'hb6871a94),
	.w2(32'h373c2645),
	.w3(32'hb7bc5376),
	.w4(32'hb6d7ac66),
	.w5(32'h379b634f),
	.w6(32'hb753cdea),
	.w7(32'hb73b923d),
	.w8(32'h37068077),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823f708),
	.w1(32'hb91dc8be),
	.w2(32'hb8f91397),
	.w3(32'h381a83ba),
	.w4(32'hb90f74d0),
	.w5(32'hb9090969),
	.w6(32'h38dc30d6),
	.w7(32'hb8103dfa),
	.w8(32'hb8e13145),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8067a),
	.w1(32'hb88ea54b),
	.w2(32'h38c44fec),
	.w3(32'hb905f928),
	.w4(32'hb90182d6),
	.w5(32'hb7b7ea75),
	.w6(32'hb75e0264),
	.w7(32'hb83111f3),
	.w8(32'h37aed18c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38040872),
	.w1(32'h388df66e),
	.w2(32'h38cb1c1f),
	.w3(32'hb7c59824),
	.w4(32'h37ae0bd0),
	.w5(32'h381f5560),
	.w6(32'hb75cff91),
	.w7(32'h376071e1),
	.w8(32'h370fd780),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36472cf8),
	.w1(32'hb80e69cf),
	.w2(32'h37d5523a),
	.w3(32'hb7552875),
	.w4(32'hb889101e),
	.w5(32'hb787d48e),
	.w6(32'hb879da46),
	.w7(32'hb892dc45),
	.w8(32'hb7f18c5d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3821b6f2),
	.w1(32'h3794412f),
	.w2(32'h36c0897b),
	.w3(32'h37062056),
	.w4(32'h36fffaf7),
	.w5(32'h365a727c),
	.w6(32'hb74d4050),
	.w7(32'hb69f8e07),
	.w8(32'hb60f50ac),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362ecfe4),
	.w1(32'h36743827),
	.w2(32'hb611e600),
	.w3(32'h36b4c3c0),
	.w4(32'h36d60632),
	.w5(32'h35a498fc),
	.w6(32'h368e1de1),
	.w7(32'h36bb2971),
	.w8(32'h3659962f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f2d563),
	.w1(32'hb73cc562),
	.w2(32'hb833fd2e),
	.w3(32'hb6891eb7),
	.w4(32'h378490b1),
	.w5(32'hb7db551f),
	.w6(32'hb791e6bd),
	.w7(32'hb83027e0),
	.w8(32'hb87276a9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6920f12),
	.w1(32'hb5eb90e9),
	.w2(32'hb700224a),
	.w3(32'hb42d0765),
	.w4(32'h35b9c754),
	.w5(32'hb62001c7),
	.w6(32'h37060a03),
	.w7(32'h3713d4cd),
	.w8(32'h366f96c7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e3286),
	.w1(32'hb8bfcaed),
	.w2(32'hb89c0d04),
	.w3(32'hb843404b),
	.w4(32'hb9008765),
	.w5(32'hb88bd0b7),
	.w6(32'hb828b738),
	.w7(32'hb90d0e57),
	.w8(32'hb9162edd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb756ddee),
	.w1(32'hb8a5f7f4),
	.w2(32'h37dc429b),
	.w3(32'h380e87bc),
	.w4(32'hb8a53546),
	.w5(32'h376307d5),
	.w6(32'hb902c902),
	.w7(32'hb9193e61),
	.w8(32'hb8a1b113),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dfabe4),
	.w1(32'hb73bb43c),
	.w2(32'h3943baee),
	.w3(32'hb901cd5f),
	.w4(32'hb82e6c08),
	.w5(32'h39359934),
	.w6(32'hb9e51428),
	.w7(32'hb9921022),
	.w8(32'hb7184443),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a13b6),
	.w1(32'h38b81eb3),
	.w2(32'h39e43b21),
	.w3(32'h39316f47),
	.w4(32'h39a38925),
	.w5(32'h3a064441),
	.w6(32'hb9bd59b3),
	.w7(32'h3841ea84),
	.w8(32'h395d9544),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3622b293),
	.w1(32'hb5fe7580),
	.w2(32'hb6f5e3b5),
	.w3(32'h360fdca2),
	.w4(32'h32f5dacd),
	.w5(32'hb6eb9004),
	.w6(32'h36843a56),
	.w7(32'h36ed1904),
	.w8(32'hb61b6f3b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60513c5),
	.w1(32'h35a04c91),
	.w2(32'hb6dda1bf),
	.w3(32'h3481d443),
	.w4(32'h3594098b),
	.w5(32'hb70b21c4),
	.w6(32'h364a74a4),
	.w7(32'h36d204b1),
	.w8(32'h358102cc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74b1d25),
	.w1(32'hb770f9bc),
	.w2(32'hb7e576da),
	.w3(32'hb75acd88),
	.w4(32'hb70d0940),
	.w5(32'hb76bf997),
	.w6(32'h3685517e),
	.w7(32'h3721f076),
	.w8(32'hb64478a4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3889efb7),
	.w1(32'hb713ba94),
	.w2(32'h3790847c),
	.w3(32'hb76f9ee6),
	.w4(32'hb781ee67),
	.w5(32'h37fd4958),
	.w6(32'h37e0c562),
	.w7(32'h3837b26f),
	.w8(32'h3904d6b8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37568cd9),
	.w1(32'h37ab45c8),
	.w2(32'h368e3d2e),
	.w3(32'hb7be9ec1),
	.w4(32'h37cf3b4f),
	.w5(32'h372707e2),
	.w6(32'hb83c3c34),
	.w7(32'hb6a2923d),
	.w8(32'h36868d37),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3870c1cf),
	.w1(32'h37a6a502),
	.w2(32'h3833937c),
	.w3(32'h3852edea),
	.w4(32'h3762ebb3),
	.w5(32'hb7af4a71),
	.w6(32'h3814ec1d),
	.w7(32'h385672c4),
	.w8(32'hb86c7129),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a30167),
	.w1(32'h3752e25f),
	.w2(32'hb70653c6),
	.w3(32'hb8298260),
	.w4(32'hb85157c3),
	.w5(32'hb8c0cce7),
	.w6(32'h38c8af63),
	.w7(32'h385a04f9),
	.w8(32'hb8df494d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6083c6b),
	.w1(32'hb7bf0bc7),
	.w2(32'h388e84fd),
	.w3(32'hb780467f),
	.w4(32'hb821becf),
	.w5(32'h38aea5b6),
	.w6(32'hb8e82e6b),
	.w7(32'hb8b98363),
	.w8(32'h377fef92),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb769ecfd),
	.w1(32'h3789bc4b),
	.w2(32'h3941d7e1),
	.w3(32'hb88ba975),
	.w4(32'hb8068c3b),
	.w5(32'h391a58aa),
	.w6(32'hb89969d8),
	.w7(32'hb72db9bd),
	.w8(32'h3917077e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38040141),
	.w1(32'hb7590501),
	.w2(32'h378fff72),
	.w3(32'h383bdb30),
	.w4(32'hb797370d),
	.w5(32'h37ea59be),
	.w6(32'h37984aa9),
	.w7(32'hb71867bb),
	.w8(32'h363b7b53),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3819b847),
	.w1(32'hb7c5ffb8),
	.w2(32'h393bb827),
	.w3(32'h366e8e0f),
	.w4(32'hb8dae38f),
	.w5(32'h38e84d3c),
	.w6(32'h38e8299c),
	.w7(32'h378cfb52),
	.w8(32'h38ce2718),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a2297c),
	.w1(32'hb84669c8),
	.w2(32'hb85de053),
	.w3(32'h384d35b8),
	.w4(32'hb847b953),
	.w5(32'hb8997694),
	.w6(32'h38a72860),
	.w7(32'hb53bc6f0),
	.w8(32'hb89eb8fe),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5884267),
	.w1(32'hb630587a),
	.w2(32'hb6382246),
	.w3(32'hb5b78922),
	.w4(32'hb601d0a2),
	.w5(32'hb68174a0),
	.w6(32'hb5d3810e),
	.w7(32'hb6111679),
	.w8(32'hb6a7a192),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361da36b),
	.w1(32'hb57eb5c0),
	.w2(32'hb5cf1b21),
	.w3(32'hb451dbf3),
	.w4(32'h35b7e81c),
	.w5(32'hb507dfec),
	.w6(32'hb65b294f),
	.w7(32'h3660169b),
	.w8(32'h355af10f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eddf6a),
	.w1(32'hb6837ecf),
	.w2(32'hb72d8e9e),
	.w3(32'hb5a25952),
	.w4(32'hb54628e9),
	.w5(32'hb6c42c9c),
	.w6(32'hb725cc5f),
	.w7(32'hb695648c),
	.w8(32'hb6464925),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37188443),
	.w1(32'h37840c07),
	.w2(32'h37440f30),
	.w3(32'h37299231),
	.w4(32'h375e159a),
	.w5(32'h373ce5d4),
	.w6(32'h36fa203d),
	.w7(32'h370dc072),
	.w8(32'h3735abbb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a79ec1),
	.w1(32'hb604a421),
	.w2(32'h3869164f),
	.w3(32'h37a66a3d),
	.w4(32'h37120e38),
	.w5(32'h38308c79),
	.w6(32'h38e78d13),
	.w7(32'h389fa72e),
	.w8(32'h38c0544c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb2b6ee59),
	.w1(32'hb71c98ca),
	.w2(32'hb7473815),
	.w3(32'hb6c064e9),
	.w4(32'hb7017801),
	.w5(32'hb6ef17e2),
	.w6(32'hb7b72279),
	.w7(32'hb79d864a),
	.w8(32'hb7dc73c6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb750107b),
	.w1(32'h36cb8c0f),
	.w2(32'h379b14dc),
	.w3(32'h38317e6e),
	.w4(32'h3861e739),
	.w5(32'h3860b225),
	.w6(32'h355d3903),
	.w7(32'h37d6437d),
	.w8(32'h35a5e019),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7342fd6),
	.w1(32'hb72795ba),
	.w2(32'hb720cc7a),
	.w3(32'hb8ee1352),
	.w4(32'hb8c89cd9),
	.w5(32'hb88ca589),
	.w6(32'hb887c21d),
	.w7(32'hb893e2c4),
	.w8(32'hb8941b56),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1c808),
	.w1(32'h38726a31),
	.w2(32'h38dddbda),
	.w3(32'hb7e13200),
	.w4(32'h389f3446),
	.w5(32'h38b8400a),
	.w6(32'hb92616d8),
	.w7(32'hb707f30d),
	.w8(32'h37a76006),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f98eb),
	.w1(32'hb8afdf68),
	.w2(32'h3745b410),
	.w3(32'h392d238e),
	.w4(32'hb86bfeba),
	.w5(32'h38be6409),
	.w6(32'h3903fc41),
	.w7(32'h37452323),
	.w8(32'h37e29b4e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eea8f7),
	.w1(32'hb948b744),
	.w2(32'hb91b92c1),
	.w3(32'hb8deec70),
	.w4(32'hb96a4680),
	.w5(32'hb95f3178),
	.w6(32'hb8ad7735),
	.w7(32'hb935df3c),
	.w8(32'hb94831b1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905430f),
	.w1(32'h39059968),
	.w2(32'h3981bfdd),
	.w3(32'h3910b0c3),
	.w4(32'h390d74c7),
	.w5(32'h39c4d1f3),
	.w6(32'hb95e5273),
	.w7(32'hb937d98d),
	.w8(32'h38ea3eac),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e989b7),
	.w1(32'h38e449ff),
	.w2(32'h36ec64cc),
	.w3(32'h3895d37b),
	.w4(32'h393c4dcb),
	.w5(32'h389eb9bd),
	.w6(32'hb8a7b2c9),
	.w7(32'h3809b06f),
	.w8(32'h374a6906),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a32981),
	.w1(32'hb8323472),
	.w2(32'hb82fbb0f),
	.w3(32'h38bce92f),
	.w4(32'hb839931c),
	.w5(32'hb88768c5),
	.w6(32'hb8859f23),
	.w7(32'hb8d3b7fa),
	.w8(32'hb85ba6b2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ef4ab),
	.w1(32'hb975ae4e),
	.w2(32'hb9d7f48f),
	.w3(32'hb9a220a7),
	.w4(32'hb8fd23e5),
	.w5(32'hb9667460),
	.w6(32'hb9b86fe7),
	.w7(32'hb9628f74),
	.w8(32'hb9d9a6da),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e440e6),
	.w1(32'hb737e9e2),
	.w2(32'h3812ddfa),
	.w3(32'h39893687),
	.w4(32'h38539aeb),
	.w5(32'h3899e562),
	.w6(32'hba275a45),
	.w7(32'hb9a721bd),
	.w8(32'hb948ba22),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d7adf1),
	.w1(32'hb9306fe4),
	.w2(32'hb9a79c1d),
	.w3(32'h3a181347),
	.w4(32'h3a08faf5),
	.w5(32'h38d97442),
	.w6(32'hb9e993f2),
	.w7(32'hba1a10de),
	.w8(32'hb9a333b6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926c9fc),
	.w1(32'h379946e9),
	.w2(32'h387fdce1),
	.w3(32'h38c12eb5),
	.w4(32'hb767e8df),
	.w5(32'hb8c6928c),
	.w6(32'h3863cc94),
	.w7(32'h371293b5),
	.w8(32'hb873dfcc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379dd76a),
	.w1(32'h36fed97e),
	.w2(32'h3a312c5b),
	.w3(32'h3a9f5d14),
	.w4(32'h3a27346d),
	.w5(32'h3ab4fc64),
	.w6(32'h39ecfd09),
	.w7(32'hb8c36a88),
	.w8(32'h3a236f45),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47183c),
	.w1(32'h3990ca3e),
	.w2(32'h390eb507),
	.w3(32'h3986557a),
	.w4(32'h355dee24),
	.w5(32'h3868f078),
	.w6(32'hba2280bf),
	.w7(32'hb971f3d4),
	.w8(32'hb94ab190),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f34f9),
	.w1(32'hb615509e),
	.w2(32'h39c67e48),
	.w3(32'h3792642a),
	.w4(32'hb91a8ce4),
	.w5(32'h39e31c40),
	.w6(32'h39464197),
	.w7(32'hb899a593),
	.w8(32'h392e5d49),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39218c62),
	.w1(32'h3784a477),
	.w2(32'h381eb59a),
	.w3(32'hb9cb5333),
	.w4(32'h392d2d89),
	.w5(32'hb7e4a63f),
	.w6(32'hba0e8be7),
	.w7(32'hb9a0cded),
	.w8(32'hb9b46e9e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987810b),
	.w1(32'h3960f3b2),
	.w2(32'h3921f245),
	.w3(32'h39527369),
	.w4(32'h3894bed6),
	.w5(32'h3974c567),
	.w6(32'h3948062d),
	.w7(32'h39b43848),
	.w8(32'h393492d9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed7d0b),
	.w1(32'h38bbaff9),
	.w2(32'hb907d08e),
	.w3(32'hb8e62333),
	.w4(32'h382f501d),
	.w5(32'hb973def6),
	.w6(32'hb8aed951),
	.w7(32'h36feacfa),
	.w8(32'hb90f428e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3715a1c7),
	.w1(32'hb6ae6291),
	.w2(32'h37ca77f8),
	.w3(32'h36a00605),
	.w4(32'hb7c3dbfb),
	.w5(32'hb78bbce3),
	.w6(32'hb7190cb7),
	.w7(32'hb7508a4e),
	.w8(32'hb780b47d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7681403),
	.w1(32'hb79abb55),
	.w2(32'h37058521),
	.w3(32'h3890be45),
	.w4(32'h371d2cc1),
	.w5(32'h3865fc04),
	.w6(32'hb818357e),
	.w7(32'hb8720b10),
	.w8(32'h367908a1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805c6c5),
	.w1(32'hb8ee5443),
	.w2(32'h39ab2036),
	.w3(32'h380786d9),
	.w4(32'hb95c887f),
	.w5(32'h39cdc19c),
	.w6(32'hb9d9f14e),
	.w7(32'hb9ece138),
	.w8(32'hb8de5b76),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385ebc70),
	.w1(32'hb80b7a14),
	.w2(32'h38f408b2),
	.w3(32'hb9285ee1),
	.w4(32'hb731270c),
	.w5(32'h3921c2ac),
	.w6(32'hba298ae6),
	.w7(32'hba05f50e),
	.w8(32'hb8cb2ae4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c92850),
	.w1(32'h380d44b3),
	.w2(32'h3934778f),
	.w3(32'h3986a414),
	.w4(32'h39533e01),
	.w5(32'h3998d26a),
	.w6(32'h362bc20c),
	.w7(32'h388a2179),
	.w8(32'h382b03ae),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb777f098),
	.w1(32'h3806db96),
	.w2(32'h395faefb),
	.w3(32'h379b3e15),
	.w4(32'h38a950c0),
	.w5(32'h39a0e6e7),
	.w6(32'h393a877c),
	.w7(32'h38a31bd8),
	.w8(32'h3983be7f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eb994e),
	.w1(32'hb8e0eb42),
	.w2(32'hb820ff26),
	.w3(32'hb904f30d),
	.w4(32'hb955ebe7),
	.w5(32'hb9094e6c),
	.w6(32'h3834dc4b),
	.w7(32'hb84d6bb8),
	.w8(32'hb8f3dd90),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e0f9c3),
	.w1(32'hb8f8388e),
	.w2(32'h398e3595),
	.w3(32'h399e5cf8),
	.w4(32'h380dda89),
	.w5(32'h392e377f),
	.w6(32'h39c516d7),
	.w7(32'h3906b78b),
	.w8(32'h39b30d41),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886de63),
	.w1(32'h38a93bca),
	.w2(32'h392dd209),
	.w3(32'h38b85403),
	.w4(32'h38bd0159),
	.w5(32'h3980433a),
	.w6(32'hb6409cac),
	.w7(32'h3774b936),
	.w8(32'h3911435b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d41a21),
	.w1(32'h37db712c),
	.w2(32'hb6fc5379),
	.w3(32'h37bd2f0a),
	.w4(32'hb529a79b),
	.w5(32'hb7c206af),
	.w6(32'h3818827c),
	.w7(32'h38566b44),
	.w8(32'h37963679),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61e8a2a),
	.w1(32'h355c6c91),
	.w2(32'hb6a0738f),
	.w3(32'hb6740d8b),
	.w4(32'hb6812c88),
	.w5(32'hb6ae0772),
	.w6(32'h356f37ca),
	.w7(32'h36933f2b),
	.w8(32'hb421d211),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68781ad),
	.w1(32'hb5f9c206),
	.w2(32'hb6b66482),
	.w3(32'h3562c035),
	.w4(32'h35ca546e),
	.w5(32'hb63ce4ba),
	.w6(32'h35d78c51),
	.w7(32'h3526b47d),
	.w8(32'h35cf0d0a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3759392b),
	.w1(32'h372d8a04),
	.w2(32'hb598097a),
	.w3(32'hb4af9acc),
	.w4(32'hb6940692),
	.w5(32'hb7bc9bad),
	.w6(32'h37d18e91),
	.w7(32'h378debd4),
	.w8(32'hb78f9e1e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37680fba),
	.w1(32'hb8d246f2),
	.w2(32'hb88ce453),
	.w3(32'hb7f9c49a),
	.w4(32'hb905570f),
	.w5(32'hb8e44b9d),
	.w6(32'hb883db02),
	.w7(32'hb8e0ec3e),
	.w8(32'hb93bc370),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38985b4c),
	.w1(32'hb812935b),
	.w2(32'h36eec478),
	.w3(32'h381ef6e8),
	.w4(32'hb8881c7d),
	.w5(32'hb6aafa9b),
	.w6(32'h38ae279e),
	.w7(32'h37acab4c),
	.w8(32'h37a02606),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a469ac),
	.w1(32'h388e6c2b),
	.w2(32'h3834e4f1),
	.w3(32'h389c49bf),
	.w4(32'h38609f46),
	.w5(32'h38128dd7),
	.w6(32'h37c2a703),
	.w7(32'h38addaa6),
	.w8(32'h37cbb65a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1e5d9),
	.w1(32'hb75a75b3),
	.w2(32'h37b0c7fc),
	.w3(32'h34003c3e),
	.w4(32'hb628753c),
	.w5(32'h383e49b3),
	.w6(32'hb7a57306),
	.w7(32'h377d792e),
	.w8(32'h38698ad1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6baab9e),
	.w1(32'hb65621d0),
	.w2(32'hb6926a1d),
	.w3(32'hb65b94e9),
	.w4(32'hb52fbf72),
	.w5(32'hb5f809b9),
	.w6(32'h35cb4739),
	.w7(32'h36074d42),
	.w8(32'h351c70da),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372202f0),
	.w1(32'h36f52eed),
	.w2(32'h3730df72),
	.w3(32'h37a73a76),
	.w4(32'hb4a4d855),
	.w5(32'h371d37a1),
	.w6(32'hb76b0ca4),
	.w7(32'hb73020e0),
	.w8(32'h3719c6c2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76cf36d),
	.w1(32'hb6863412),
	.w2(32'h3763af43),
	.w3(32'hb662198e),
	.w4(32'hb654cd05),
	.w5(32'h35dd6134),
	.w6(32'hb757b7a8),
	.w7(32'hb7868172),
	.w8(32'h3742b1be),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a34d9f),
	.w1(32'h37dc9095),
	.w2(32'h37bf81fe),
	.w3(32'h36698785),
	.w4(32'h37a9c3e4),
	.w5(32'h38387aea),
	.w6(32'hb84cabb5),
	.w7(32'hb74defcb),
	.w8(32'h376c4096),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39092d06),
	.w1(32'h379730dd),
	.w2(32'h366d4f33),
	.w3(32'h38e7af13),
	.w4(32'h3807744d),
	.w5(32'hb892d4bb),
	.w6(32'h387cc97b),
	.w7(32'h38295746),
	.w8(32'h38840b54),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8144dca),
	.w1(32'hb8477133),
	.w2(32'hb7924173),
	.w3(32'h37ee872e),
	.w4(32'hb6a67896),
	.w5(32'hb67f5d61),
	.w6(32'hb89ef6b7),
	.w7(32'hb8fb6da3),
	.w8(32'hb7ee11f1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c866f2),
	.w1(32'h34905cfa),
	.w2(32'h35138721),
	.w3(32'h3706dfb8),
	.w4(32'h3520232a),
	.w5(32'hb67619bd),
	.w6(32'h36b89a94),
	.w7(32'h343d2ed1),
	.w8(32'hb714e2eb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8eed0),
	.w1(32'h3919d4b4),
	.w2(32'h388e3c9e),
	.w3(32'h3849b788),
	.w4(32'h37d6f5a4),
	.w5(32'h383f08b9),
	.w6(32'h38f2d087),
	.w7(32'h38abde0e),
	.w8(32'h3849f39c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76100d1),
	.w1(32'hb6fb1ac7),
	.w2(32'hb7245680),
	.w3(32'hb6dc4986),
	.w4(32'h358c380c),
	.w5(32'h36be6b71),
	.w6(32'hb7637676),
	.w7(32'hb4906e9f),
	.w8(32'h36ac6638),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383443fb),
	.w1(32'hb78303d4),
	.w2(32'h3884c681),
	.w3(32'hb7acc118),
	.w4(32'hb7e949a7),
	.w5(32'h38827a38),
	.w6(32'hb90a47e8),
	.w7(32'hb8ab8346),
	.w8(32'h37d3e96e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f2a57f),
	.w1(32'hb7a3b8d2),
	.w2(32'hb885f722),
	.w3(32'hb7fbdcae),
	.w4(32'hb71a537c),
	.w5(32'hb7f3442e),
	.w6(32'hb605223d),
	.w7(32'hb78ac777),
	.w8(32'hb83c7c30),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a42411),
	.w1(32'h36e3d11b),
	.w2(32'h38d93dce),
	.w3(32'h38366558),
	.w4(32'hb6fab9c6),
	.w5(32'h3684b5d0),
	.w6(32'hb666be8c),
	.w7(32'hb8c18f7e),
	.w8(32'hb8b31fca),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f26615),
	.w1(32'hb719e4c1),
	.w2(32'h389dbc4a),
	.w3(32'h382193d0),
	.w4(32'hb63fe964),
	.w5(32'h38bd8180),
	.w6(32'hb766cbfc),
	.w7(32'hb67b9b5a),
	.w8(32'h381f5b21),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d4c099),
	.w1(32'h38168cb9),
	.w2(32'h3836d7f2),
	.w3(32'h38bcdf80),
	.w4(32'h38757162),
	.w5(32'h38b6df4e),
	.w6(32'hb88242f7),
	.w7(32'hb8c646f7),
	.w8(32'hb829ab3f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb4e3d),
	.w1(32'h3803c54c),
	.w2(32'h377cd4bf),
	.w3(32'hb6948fdc),
	.w4(32'h37617f99),
	.w5(32'hb8bc70bf),
	.w6(32'h388b8208),
	.w7(32'h378bd02b),
	.w8(32'hb90b778b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f45c5),
	.w1(32'h37c1c37b),
	.w2(32'h381f2cb5),
	.w3(32'h38cd7e17),
	.w4(32'h38c8ff03),
	.w5(32'h382d41da),
	.w6(32'h38c68dcf),
	.w7(32'h38fb4020),
	.w8(32'h386af82a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390908f5),
	.w1(32'h37ffc1ae),
	.w2(32'h37eee8c6),
	.w3(32'h3924d277),
	.w4(32'h389ca8ec),
	.w5(32'h38f71cfe),
	.w6(32'h38d1f122),
	.w7(32'h38aa858a),
	.w8(32'hb6cdf742),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3782e69a),
	.w1(32'hb7f87c2b),
	.w2(32'h382de143),
	.w3(32'h37b52f2b),
	.w4(32'hb7acbc1d),
	.w5(32'h3885bac4),
	.w6(32'hb6672cb3),
	.w7(32'hb7d07ef1),
	.w8(32'h37a85812),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38841d84),
	.w1(32'h38b35dc7),
	.w2(32'h392044b2),
	.w3(32'h3914de85),
	.w4(32'h392efe0b),
	.w5(32'h399895a4),
	.w6(32'h38231b72),
	.w7(32'h38db33b6),
	.w8(32'h396e6a6f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380453ef),
	.w1(32'h38135f7e),
	.w2(32'h37b4f35c),
	.w3(32'h381a9694),
	.w4(32'h37f58ced),
	.w5(32'h379d2ebb),
	.w6(32'h382206f1),
	.w7(32'hb5982c1f),
	.w8(32'h36801d1f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4880f1d),
	.w1(32'hb60ed604),
	.w2(32'hb5ab51b5),
	.w3(32'h362f6720),
	.w4(32'hb648f65c),
	.w5(32'hb644d7c0),
	.w6(32'h36534738),
	.w7(32'hb5a80820),
	.w8(32'hb66d32c1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34d036a5),
	.w1(32'h35dc45fa),
	.w2(32'h35c07849),
	.w3(32'h35a4a46b),
	.w4(32'h35922c8f),
	.w5(32'h3684dc73),
	.w6(32'h34fd45aa),
	.w7(32'h35ae4818),
	.w8(32'h35e47634),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb650c57a),
	.w1(32'hb7e1f70e),
	.w2(32'hb7cc3bc2),
	.w3(32'h368d67d5),
	.w4(32'hb7d5471e),
	.w5(32'hb750a92b),
	.w6(32'hb657e02e),
	.w7(32'hb786acd0),
	.w8(32'hb732d55f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38421418),
	.w1(32'h38bdfeb4),
	.w2(32'h38efe97b),
	.w3(32'h3721170c),
	.w4(32'h38adbb00),
	.w5(32'h391634a5),
	.w6(32'hb7be1d97),
	.w7(32'h389339ae),
	.w8(32'h3900bb98),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ee0c98),
	.w1(32'hb7851d3d),
	.w2(32'h3880bb68),
	.w3(32'h370a0c52),
	.w4(32'hb805857f),
	.w5(32'h386e47d6),
	.w6(32'h35156d68),
	.w7(32'hb54cf900),
	.w8(32'h376270fb),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3717426e),
	.w1(32'hb49e1fba),
	.w2(32'h36817d39),
	.w3(32'h37207478),
	.w4(32'h36024ae7),
	.w5(32'h368b29ce),
	.w6(32'h36709d77),
	.w7(32'hb3b300ae),
	.w8(32'h369daaad),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad1911),
	.w1(32'hb8187e9f),
	.w2(32'h368a302c),
	.w3(32'h385d16a1),
	.w4(32'hb76986fd),
	.w5(32'h386ebc7f),
	.w6(32'h36609503),
	.w7(32'hb8a811a9),
	.w8(32'h38303c4e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39344e3b),
	.w1(32'h39c1b8c9),
	.w2(32'h394f1e71),
	.w3(32'hb8f2c07c),
	.w4(32'h398cf72b),
	.w5(32'h396975ac),
	.w6(32'hb98798f2),
	.w7(32'hb8a40127),
	.w8(32'h383c08ad),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2c891),
	.w1(32'h3985feb7),
	.w2(32'h3a10a730),
	.w3(32'h3988a889),
	.w4(32'h39951548),
	.w5(32'h3a2cb92e),
	.w6(32'h39bb09b9),
	.w7(32'h39d0c6dc),
	.w8(32'h3a0212fb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787dd99),
	.w1(32'h38417f65),
	.w2(32'h3884ee57),
	.w3(32'hb79d4bce),
	.w4(32'h387cd7e6),
	.w5(32'h3907cd8b),
	.w6(32'hb8df3532),
	.w7(32'hb67eb430),
	.w8(32'h388937aa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e29318),
	.w1(32'hb8797373),
	.w2(32'hb93584ec),
	.w3(32'hb86b2bbe),
	.w4(32'h3887dc5d),
	.w5(32'h389fd17e),
	.w6(32'hb909c8d5),
	.w7(32'hb8cd8d8e),
	.w8(32'hb8f5d1ec),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba460dd7),
	.w1(32'hba147fda),
	.w2(32'h3aab5379),
	.w3(32'hb997c836),
	.w4(32'hb9d10b48),
	.w5(32'h3aaee002),
	.w6(32'hba56c858),
	.w7(32'hba0cfa78),
	.w8(32'h3a4add86),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c727f),
	.w1(32'h3b1cc792),
	.w2(32'h3b5637c5),
	.w3(32'h3ae13f11),
	.w4(32'h3aa54276),
	.w5(32'hbb449070),
	.w6(32'h3aafc49b),
	.w7(32'h3a96361d),
	.w8(32'hbbe004a8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913be1d),
	.w1(32'h3b9f23ed),
	.w2(32'hbb8dd17a),
	.w3(32'h3b07b67d),
	.w4(32'h3ae3a7db),
	.w5(32'hbc459c17),
	.w6(32'hbbeef508),
	.w7(32'hbbfe0618),
	.w8(32'hbc20df86),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9071ce),
	.w1(32'h3a98e77d),
	.w2(32'hbad15805),
	.w3(32'h3b207956),
	.w4(32'hbbd8a131),
	.w5(32'h3ada6c28),
	.w6(32'h3b6f595e),
	.w7(32'hbbb8d21c),
	.w8(32'h3b136bc1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8926ab),
	.w1(32'hbac8715d),
	.w2(32'h3b87a2b5),
	.w3(32'hba2583a4),
	.w4(32'h3a59cb2e),
	.w5(32'h3ba2169d),
	.w6(32'hb94aff75),
	.w7(32'hb9d39eab),
	.w8(32'h3b0c0912),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe07c4c),
	.w1(32'hbbb81f21),
	.w2(32'hba6b9454),
	.w3(32'hbbd71862),
	.w4(32'hbc3e153f),
	.w5(32'h3b3b2a08),
	.w6(32'hbc7d0fb9),
	.w7(32'hbb04f19e),
	.w8(32'h3b636a74),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb155abb),
	.w1(32'hbb829d63),
	.w2(32'hbb37ac03),
	.w3(32'hbc2bf7b1),
	.w4(32'hbb182cc0),
	.w5(32'hba57c578),
	.w6(32'hbc0d43ff),
	.w7(32'h3c196db2),
	.w8(32'hb9a1b982),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53d8ed),
	.w1(32'hb9b74de2),
	.w2(32'hbbe9a67c),
	.w3(32'hba4f4316),
	.w4(32'hbb2f0207),
	.w5(32'hbc3b31c9),
	.w6(32'hba72159e),
	.w7(32'hb9b30aa0),
	.w8(32'hbc1669cd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7bfe3),
	.w1(32'hba33121e),
	.w2(32'h3b11b143),
	.w3(32'hba97401d),
	.w4(32'h3bb2fd41),
	.w5(32'h3a2d92aa),
	.w6(32'hbb257d67),
	.w7(32'h3a40baa7),
	.w8(32'hbab0df5d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ae7dc),
	.w1(32'h3ae5dfad),
	.w2(32'hbbe267d9),
	.w3(32'h3aab009c),
	.w4(32'hbb19b98b),
	.w5(32'hbc024eb2),
	.w6(32'h39c3d359),
	.w7(32'hbaf5cf6a),
	.w8(32'hbc08c096),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64be62),
	.w1(32'h3c2fb97d),
	.w2(32'h3b44a31b),
	.w3(32'h3bc2111b),
	.w4(32'h3c6dd024),
	.w5(32'h3ba69fb4),
	.w6(32'h3be58a7b),
	.w7(32'h3be7bf9e),
	.w8(32'hb9a30281),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bfece),
	.w1(32'h3b791fa1),
	.w2(32'h3c18d2ed),
	.w3(32'h3b96e81c),
	.w4(32'h3af61c82),
	.w5(32'h3c6da617),
	.w6(32'h3b1c1346),
	.w7(32'hba975ca1),
	.w8(32'h3b9aaecf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a161),
	.w1(32'hbac13bd7),
	.w2(32'hbad5c0a7),
	.w3(32'hb9a74237),
	.w4(32'hbbb2e428),
	.w5(32'hbb84b15c),
	.w6(32'hbb7682ce),
	.w7(32'h3a7174b4),
	.w8(32'h390a009a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f4196),
	.w1(32'h3b926442),
	.w2(32'h3a028b77),
	.w3(32'h3c9acaa9),
	.w4(32'h3b44d522),
	.w5(32'h3a8a04b4),
	.w6(32'h3c20bd7c),
	.w7(32'hbb34598b),
	.w8(32'h3b87cb97),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df711),
	.w1(32'hba0c7937),
	.w2(32'h391f36a6),
	.w3(32'hbbb5e993),
	.w4(32'hbb712975),
	.w5(32'h3b1e2eca),
	.w6(32'hb89eb6df),
	.w7(32'h3a3cc14c),
	.w8(32'h3bd2f625),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dd026),
	.w1(32'h3b50de79),
	.w2(32'hba80cb32),
	.w3(32'hb9adbf89),
	.w4(32'h3a1815af),
	.w5(32'hbc71ee76),
	.w6(32'h3be3eb7f),
	.w7(32'h3a95b906),
	.w8(32'hbc3bf6c3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c0db),
	.w1(32'hbc01ed56),
	.w2(32'h3ab01e65),
	.w3(32'hbcb1a7b8),
	.w4(32'h3bbe0353),
	.w5(32'h3a5befc0),
	.w6(32'hbca3fc22),
	.w7(32'h3bcc7574),
	.w8(32'hba561b8c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09e3bc),
	.w1(32'h3b19b2c5),
	.w2(32'h3a752822),
	.w3(32'hba41b3ac),
	.w4(32'hb9ea8160),
	.w5(32'h3c27383d),
	.w6(32'h3afbf55d),
	.w7(32'h3b3ed5bc),
	.w8(32'h3c7a935f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc20bf4),
	.w1(32'hbb872899),
	.w2(32'h3c182fe9),
	.w3(32'h3cbd54a3),
	.w4(32'hbc48d8c8),
	.w5(32'h3c50e065),
	.w6(32'h3c887c77),
	.w7(32'hbc863175),
	.w8(32'h3c37760e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc191839),
	.w1(32'hbc2c0f0f),
	.w2(32'hbc42d7ea),
	.w3(32'hbb5d3c81),
	.w4(32'h3c61fd72),
	.w5(32'hbc545447),
	.w6(32'hb9614f87),
	.w7(32'h3bff80c0),
	.w8(32'hbc8e1d97),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8197cc),
	.w1(32'h3aa96b67),
	.w2(32'h3bf50b3c),
	.w3(32'hbc62285d),
	.w4(32'h3c025782),
	.w5(32'h3bf1b114),
	.w6(32'hbc01ca70),
	.w7(32'h3c1b2b4c),
	.w8(32'hbb357eb2),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75bfde),
	.w1(32'hbc1d9277),
	.w2(32'h3b8bcb98),
	.w3(32'hbc8fd689),
	.w4(32'h398c1efb),
	.w5(32'h3b3a8702),
	.w6(32'hbc02070d),
	.w7(32'h3a63fe1d),
	.w8(32'h3ac02ab7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be12b19),
	.w1(32'h3b4e8401),
	.w2(32'h3a232e53),
	.w3(32'h3bd3f318),
	.w4(32'h3ba6c4b7),
	.w5(32'h3ab41b1a),
	.w6(32'h3bbe2923),
	.w7(32'h3b8fd75f),
	.w8(32'h3b13fe00),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e7c37),
	.w1(32'h3b6304b0),
	.w2(32'h3b4c94ef),
	.w3(32'hbc2e209f),
	.w4(32'h3a977ece),
	.w5(32'hbb85df2f),
	.w6(32'hbc82c809),
	.w7(32'hbb999a65),
	.w8(32'hbb8899de),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099287),
	.w1(32'hbb5ab8e8),
	.w2(32'h3b38de3b),
	.w3(32'h3b5c0505),
	.w4(32'hbb4ad93d),
	.w5(32'h3b831d4b),
	.w6(32'h3c1ef658),
	.w7(32'hbba30068),
	.w8(32'h3c6a6a02),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b676a61),
	.w1(32'hbc2bf801),
	.w2(32'h3bfeb3dc),
	.w3(32'h3bfe2591),
	.w4(32'hbca1e5d1),
	.w5(32'hba9f705a),
	.w6(32'h3b3a507b),
	.w7(32'hbb35f75d),
	.w8(32'hba54206f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb70d67),
	.w1(32'h3bdd39f5),
	.w2(32'h3a4e1218),
	.w3(32'h3c8e9001),
	.w4(32'h3888f997),
	.w5(32'h3b778e7b),
	.w6(32'h3c58b582),
	.w7(32'hbc043721),
	.w8(32'hbb0c338a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb969d7),
	.w1(32'hbbf6e139),
	.w2(32'hbc28a3cb),
	.w3(32'hbbd22ff5),
	.w4(32'hbc2d192d),
	.w5(32'hbc8218b4),
	.w6(32'hbbc1ac43),
	.w7(32'hbb1b9f33),
	.w8(32'hbb99f1dc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf69a),
	.w1(32'h3b89338c),
	.w2(32'hbb936541),
	.w3(32'h3c3df7af),
	.w4(32'h3b96b551),
	.w5(32'h3c0db684),
	.w6(32'h3bc61d35),
	.w7(32'h3b20f338),
	.w8(32'h3c8193d1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5ba6),
	.w1(32'hbac47c71),
	.w2(32'h3ad193a6),
	.w3(32'h3bf594f8),
	.w4(32'hbc944df5),
	.w5(32'hbc6d5bd7),
	.w6(32'h3b45e4c3),
	.w7(32'hbc8f0d97),
	.w8(32'hbc46bc98),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f482d7),
	.w1(32'h3a3ae60d),
	.w2(32'h3c001f4f),
	.w3(32'h3c3e0aca),
	.w4(32'h3acd3ef2),
	.w5(32'h3b9709c5),
	.w6(32'h3c5e7b00),
	.w7(32'hbbd3551c),
	.w8(32'h3c02f8eb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b1a4e),
	.w1(32'h3c5d7fb2),
	.w2(32'hba5f2153),
	.w3(32'h3b4c2309),
	.w4(32'h3c10143b),
	.w5(32'hba8ef4b8),
	.w6(32'hba4ac9cc),
	.w7(32'h3b739078),
	.w8(32'hb9cf2265),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0080aa),
	.w1(32'hbbf4ee87),
	.w2(32'h3b1ce83f),
	.w3(32'hbaa5c6de),
	.w4(32'hbc13cc04),
	.w5(32'h3ba4d7aa),
	.w6(32'hb97b85b5),
	.w7(32'hbc2c5cc9),
	.w8(32'h3befa2ed),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae03cee),
	.w1(32'hba9fa0d5),
	.w2(32'h3afbc059),
	.w3(32'hbb3d45b9),
	.w4(32'hb9ed75e0),
	.w5(32'hba13f710),
	.w6(32'hbb8d8c9f),
	.w7(32'hbba41318),
	.w8(32'h3b996881),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc340796),
	.w1(32'hbbaa45f9),
	.w2(32'hba69a196),
	.w3(32'hbc831e86),
	.w4(32'hbb3d1857),
	.w5(32'hbb41d97e),
	.w6(32'hbc7b3fce),
	.w7(32'hba2b0da9),
	.w8(32'hbc0f43de),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83bff1),
	.w1(32'h3b061a63),
	.w2(32'h3c2edfd8),
	.w3(32'hbcb1988e),
	.w4(32'hb9bfa3a8),
	.w5(32'h3ac0c01b),
	.w6(32'hbbcc64c8),
	.w7(32'hbac7fa00),
	.w8(32'h3bc8dcbf),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82424c),
	.w1(32'h3bafe655),
	.w2(32'h3a589d5c),
	.w3(32'hbc0f1c76),
	.w4(32'h3c37faf2),
	.w5(32'hbb91cc97),
	.w6(32'h3b806555),
	.w7(32'h3c3c87c8),
	.w8(32'h3af136c3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e59f0),
	.w1(32'h3bb20576),
	.w2(32'h3c0bdc01),
	.w3(32'hba8b4ca0),
	.w4(32'hbacdc52f),
	.w5(32'h3c3c0007),
	.w6(32'h3b3da5cf),
	.w7(32'h3b96e93f),
	.w8(32'h3c0ee6e6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adde5b3),
	.w1(32'hbc1a1f12),
	.w2(32'h3b34a3d5),
	.w3(32'hbc1418ca),
	.w4(32'hbc9ba348),
	.w5(32'h3b8905dc),
	.w6(32'hbc9ce6cb),
	.w7(32'hbcb4e221),
	.w8(32'h3bcb1c07),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af45851),
	.w1(32'hbb4448b2),
	.w2(32'hba7560d9),
	.w3(32'h3ad8caef),
	.w4(32'hbb8816bb),
	.w5(32'h3a6072ee),
	.w6(32'h3b8ab416),
	.w7(32'hbb1ba478),
	.w8(32'hb9a93368),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad34d09),
	.w1(32'hb970a7ef),
	.w2(32'hbbf1d14c),
	.w3(32'h3a65be2b),
	.w4(32'hbb1a6134),
	.w5(32'hbc4179c4),
	.w6(32'h3b5dec85),
	.w7(32'h3ace38a5),
	.w8(32'hbc7cce97),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ca263),
	.w1(32'h3c6c35ff),
	.w2(32'h3be1d58f),
	.w3(32'h3c58d24f),
	.w4(32'h3c2d2ae4),
	.w5(32'h3ba3b6d9),
	.w6(32'h3c0fccbd),
	.w7(32'h3b29c904),
	.w8(32'h3bfefc41),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ad100),
	.w1(32'hbbe49164),
	.w2(32'h3ae92f1a),
	.w3(32'h3b8099b1),
	.w4(32'hbc860863),
	.w5(32'h3b49d9fc),
	.w6(32'h3addf6ef),
	.w7(32'hbca6f506),
	.w8(32'h3bb8ab69),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40a920),
	.w1(32'h3a11a884),
	.w2(32'h3baa1d24),
	.w3(32'h3a87e8df),
	.w4(32'h3b1fdf87),
	.w5(32'h39db4e5c),
	.w6(32'h3b4964ee),
	.w7(32'h3ba984ec),
	.w8(32'hba74ad05),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa71da),
	.w1(32'h3bca875c),
	.w2(32'hb811bd87),
	.w3(32'h3a19131f),
	.w4(32'h38d52a8d),
	.w5(32'hbbf5a772),
	.w6(32'h3b47c60e),
	.w7(32'h3b3b672f),
	.w8(32'hbbb76358),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf57b64),
	.w1(32'h3b94070b),
	.w2(32'hbc9118ef),
	.w3(32'h397a8110),
	.w4(32'h3aa5655a),
	.w5(32'hbc9745b8),
	.w6(32'h3b88c77a),
	.w7(32'hbb3bb846),
	.w8(32'hbc550cdd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3a9a2),
	.w1(32'hbaae54c7),
	.w2(32'h3c4ef831),
	.w3(32'hbc4febef),
	.w4(32'h3c1244d6),
	.w5(32'h3cd012ba),
	.w6(32'hbb683adc),
	.w7(32'h3bec0ab2),
	.w8(32'h3c68be75),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab24fe5),
	.w1(32'hbc4cdd53),
	.w2(32'h3b5c9dc1),
	.w3(32'hbb596460),
	.w4(32'hbcc7eb49),
	.w5(32'h3ac30060),
	.w6(32'hbc29eb34),
	.w7(32'hbca81795),
	.w8(32'h39962053),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb0cd),
	.w1(32'h396ae016),
	.w2(32'hbb52f2cf),
	.w3(32'hba8b2f33),
	.w4(32'hbb194ae8),
	.w5(32'h3af74f9b),
	.w6(32'h3a2af653),
	.w7(32'hba77c020),
	.w8(32'h3a87ee54),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf65e),
	.w1(32'h3b7a8347),
	.w2(32'h3c2f03e3),
	.w3(32'h3b48a91b),
	.w4(32'h3b4e0961),
	.w5(32'h3cdddca9),
	.w6(32'h3b80c9e7),
	.w7(32'h3b7cd59e),
	.w8(32'h3cc6b98a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21a4c3),
	.w1(32'hbc971131),
	.w2(32'h3c33000b),
	.w3(32'h3c319990),
	.w4(32'hbcc34b89),
	.w5(32'h3ca73715),
	.w6(32'h3b87083c),
	.w7(32'hbcb24b6e),
	.w8(32'h3cc771b6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf0163),
	.w1(32'hbcbd452d),
	.w2(32'hbb59d8a5),
	.w3(32'h3a07b342),
	.w4(32'hbceb2901),
	.w5(32'hbc65fae6),
	.w6(32'hbb7e1744),
	.w7(32'hbc72055d),
	.w8(32'hbc821eba),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a9317),
	.w1(32'hbaf927b6),
	.w2(32'h3b0af668),
	.w3(32'hb718157c),
	.w4(32'h3c55486f),
	.w5(32'h3b33d887),
	.w6(32'hbacd177b),
	.w7(32'h3bc594e0),
	.w8(32'h3af83d2b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4caf91),
	.w1(32'h3b130a3f),
	.w2(32'h3a28e198),
	.w3(32'hb9d10964),
	.w4(32'h3aac28c5),
	.w5(32'hbb537440),
	.w6(32'h39a0e129),
	.w7(32'h3a9b8c38),
	.w8(32'hbb8477c6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48ca32),
	.w1(32'h3a5db4a0),
	.w2(32'h3b5023b9),
	.w3(32'h3a9dc5ea),
	.w4(32'hb737f2ca),
	.w5(32'h3b911b4a),
	.w6(32'h3b9fe7a0),
	.w7(32'hbaf14cf0),
	.w8(32'h3b7aab1a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d56e),
	.w1(32'h3a465712),
	.w2(32'h3be7f04a),
	.w3(32'h39e77dfd),
	.w4(32'hbaa28961),
	.w5(32'hbc32b2e1),
	.w6(32'h3aeb61d2),
	.w7(32'hb89cb7fb),
	.w8(32'hbc8fb18e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21d891),
	.w1(32'h3c9fcff5),
	.w2(32'hbb5629ad),
	.w3(32'hbc95af10),
	.w4(32'h3ca655dd),
	.w5(32'hbbb902b0),
	.w6(32'hbc07fc64),
	.w7(32'h3c967485),
	.w8(32'hbc1b4821),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b96ed),
	.w1(32'hbb00fd4b),
	.w2(32'hbc99c360),
	.w3(32'hbcc602db),
	.w4(32'h3b2f60d6),
	.w5(32'hbc9ad9b9),
	.w6(32'hbcab18d8),
	.w7(32'h3b48e51e),
	.w8(32'hbc1ec9fc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18cef1),
	.w1(32'hbb72a14f),
	.w2(32'hbba244cd),
	.w3(32'hbc83e6a7),
	.w4(32'h3a2fe688),
	.w5(32'hbbafdb69),
	.w6(32'hbc05c9f2),
	.w7(32'h3c02b74e),
	.w8(32'hba9a5be6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc12939),
	.w1(32'h3b4bc9cb),
	.w2(32'h3bb08a88),
	.w3(32'h3b9f2363),
	.w4(32'hbb2c3ecd),
	.w5(32'h3a949662),
	.w6(32'h3bfb4e0a),
	.w7(32'hbbd0542b),
	.w8(32'h3b16183a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9333b9a),
	.w1(32'hbaf17311),
	.w2(32'h3b383ce6),
	.w3(32'hbba1a6ab),
	.w4(32'hbbec9a44),
	.w5(32'h3b94dce3),
	.w6(32'hbb25d9bf),
	.w7(32'hbbec755d),
	.w8(32'h3bc1b302),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacd220),
	.w1(32'hb9b636a4),
	.w2(32'h3b7b1eb1),
	.w3(32'h3b380914),
	.w4(32'h3b1135e8),
	.w5(32'hbad38735),
	.w6(32'h3bd1d3f0),
	.w7(32'h3b66ceda),
	.w8(32'h3b708bcc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd63de),
	.w1(32'hbae9e893),
	.w2(32'hba29c830),
	.w3(32'h3c3937be),
	.w4(32'hbbcb8a3b),
	.w5(32'h3b91af7b),
	.w6(32'h3c6f1332),
	.w7(32'hbb32d695),
	.w8(32'h3b9ee505),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae57d4b),
	.w1(32'hbbdc91ba),
	.w2(32'hba3194ce),
	.w3(32'h3bc5adca),
	.w4(32'hbb4bffd8),
	.w5(32'h3b8688f0),
	.w6(32'h3c2dfcc9),
	.w7(32'hbaec2a1a),
	.w8(32'h3bd2cb79),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac548d8),
	.w1(32'hba5e2ce9),
	.w2(32'h3b394c7d),
	.w3(32'h394b9791),
	.w4(32'hba8ea35d),
	.w5(32'h3bab18bc),
	.w6(32'h3a162a29),
	.w7(32'h3b24f2f8),
	.w8(32'h3ba37bbd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92d8c),
	.w1(32'hbb9443ac),
	.w2(32'h3bce3604),
	.w3(32'hbc14bcfc),
	.w4(32'hbb15c26d),
	.w5(32'h3bb0444b),
	.w6(32'hbbeaec9c),
	.w7(32'hba980ce1),
	.w8(32'h3b91878c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2e1dd),
	.w1(32'h3b6ba448),
	.w2(32'h3b71f7cb),
	.w3(32'h3bb82225),
	.w4(32'hb995eb06),
	.w5(32'h3b2e6bc1),
	.w6(32'h3b72dcec),
	.w7(32'hbb3fc687),
	.w8(32'h3adb5e1c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b6557),
	.w1(32'h3b0741d3),
	.w2(32'h3bd83276),
	.w3(32'hbab7b557),
	.w4(32'h3a547dc9),
	.w5(32'h3c47e3ad),
	.w6(32'hbac4e09f),
	.w7(32'h3a87130c),
	.w8(32'h3c353e86),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a80be),
	.w1(32'hbb41e4d4),
	.w2(32'h3bdfc4e7),
	.w3(32'h3bd6fb42),
	.w4(32'hbc7eca81),
	.w5(32'h3bf9ee98),
	.w6(32'h3ba34d25),
	.w7(32'hbc468b49),
	.w8(32'h3b67b9f4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf2f76),
	.w1(32'hbc639e0e),
	.w2(32'hbae0faa7),
	.w3(32'hbc1d04f0),
	.w4(32'hbc577f06),
	.w5(32'hbba30de0),
	.w6(32'hbc64c3de),
	.w7(32'hbaca9831),
	.w8(32'hbba6cac1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadff33),
	.w1(32'h3bb8a5b8),
	.w2(32'hbbd2935e),
	.w3(32'h3ac7d460),
	.w4(32'h3b676d42),
	.w5(32'hbc433f66),
	.w6(32'h3ae18949),
	.w7(32'h3a2f125a),
	.w8(32'hbbedb824),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce50c2e),
	.w1(32'hbb901da6),
	.w2(32'h3b20592a),
	.w3(32'hbcb9da05),
	.w4(32'h3c72f7a0),
	.w5(32'h3c024df6),
	.w6(32'hbc163e3d),
	.w7(32'h3c563cfc),
	.w8(32'h3c0d0a03),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf887fc),
	.w1(32'hbbd576bc),
	.w2(32'h3b79814b),
	.w3(32'h3c11cb5f),
	.w4(32'hbc57788c),
	.w5(32'h3bb3524e),
	.w6(32'h3bd1cf68),
	.w7(32'hba8e903a),
	.w8(32'h3b89df52),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb02c),
	.w1(32'h3b9e7d4b),
	.w2(32'h39135b18),
	.w3(32'hbad5ec07),
	.w4(32'hba5772be),
	.w5(32'hbc61c438),
	.w6(32'hbb676e9d),
	.w7(32'hbbd4bdbc),
	.w8(32'hbbeaa242),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd23df0),
	.w1(32'hbb59d91a),
	.w2(32'h3b3acd51),
	.w3(32'hbcab6280),
	.w4(32'hbbd22d48),
	.w5(32'h3a7cd102),
	.w6(32'hbc8e8296),
	.w7(32'h3b8f3e2a),
	.w8(32'hbbb2ccfe),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb890b854),
	.w1(32'hbbe76035),
	.w2(32'h3a9ad476),
	.w3(32'hbc9ca2fd),
	.w4(32'hbc5e7573),
	.w5(32'h3a2ad866),
	.w6(32'hbc9ffcaa),
	.w7(32'hbbf83c70),
	.w8(32'h3c0387f6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc53c9),
	.w1(32'hbacb201f),
	.w2(32'h3a9e8a29),
	.w3(32'h3c183ed6),
	.w4(32'hbb69c61a),
	.w5(32'hbaf73575),
	.w6(32'h3c161f5c),
	.w7(32'hba34b3db),
	.w8(32'hbb78d430),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb445bd1),
	.w1(32'hbb6363a0),
	.w2(32'hb7f06fab),
	.w3(32'hbc24cb92),
	.w4(32'hbbc0fdcc),
	.w5(32'hbc115fee),
	.w6(32'hbbd945a8),
	.w7(32'h3abc9cb7),
	.w8(32'hbbed99dc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb9db2),
	.w1(32'h3c680f38),
	.w2(32'hbbb2a2ab),
	.w3(32'h3c2abeff),
	.w4(32'h3bf1c20a),
	.w5(32'hbbdee359),
	.w6(32'h3ae820c3),
	.w7(32'hb8e4739e),
	.w8(32'hbad160b2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac043ae),
	.w1(32'h3bfbc8e7),
	.w2(32'hbb36d664),
	.w3(32'h3ba82f1f),
	.w4(32'hba534bb1),
	.w5(32'hbc1c9459),
	.w6(32'h3acff378),
	.w7(32'hbbe0bee8),
	.w8(32'hbbed2771),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21f68d),
	.w1(32'h3c255742),
	.w2(32'h3a498736),
	.w3(32'h3ac45170),
	.w4(32'h3ba36791),
	.w5(32'hbb12bad6),
	.w6(32'h3b332546),
	.w7(32'hbb30f59a),
	.w8(32'hba087d4f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8deb45),
	.w1(32'h3ace3314),
	.w2(32'hbc4e0f41),
	.w3(32'hbb071d60),
	.w4(32'h393d5f01),
	.w5(32'hbcdf4799),
	.w6(32'h3a080437),
	.w7(32'hbb9ecd1b),
	.w8(32'hbc7c5a6e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a212),
	.w1(32'h3a3ad626),
	.w2(32'h3afe7849),
	.w3(32'hbb7f45b9),
	.w4(32'hbb9cff5f),
	.w5(32'h3b15ecb0),
	.w6(32'h3b1afdfe),
	.w7(32'hbb9f7ac6),
	.w8(32'hbb0d4ff3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3be5f),
	.w1(32'hbbb8c79f),
	.w2(32'hba0fefd8),
	.w3(32'hbc97522a),
	.w4(32'h3a81c315),
	.w5(32'hbc42f194),
	.w6(32'hbc880e97),
	.w7(32'h3b73962a),
	.w8(32'hbc0da7d6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6986db),
	.w1(32'h3a881430),
	.w2(32'h3acd8ad1),
	.w3(32'hbc7d6de5),
	.w4(32'h3c623f81),
	.w5(32'hbc1f545b),
	.w6(32'hbbdbd0b2),
	.w7(32'h3c3920dc),
	.w8(32'hbbe5293f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48382f),
	.w1(32'h3c5263bb),
	.w2(32'h3b4350e1),
	.w3(32'h3c4a35eb),
	.w4(32'h3c596edf),
	.w5(32'hbbfc025a),
	.w6(32'h3c60e4e7),
	.w7(32'h3b648623),
	.w8(32'hbc1b4f71),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b422eff),
	.w1(32'h3c804129),
	.w2(32'h3b87cba2),
	.w3(32'h3b0d6934),
	.w4(32'h3ca332f8),
	.w5(32'hbbc65e3d),
	.w6(32'h3a885c33),
	.w7(32'h3c5f428b),
	.w8(32'hbc3ca0c1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc420bdc),
	.w1(32'h3b2ce6c0),
	.w2(32'hbba86be5),
	.w3(32'hbcd13f75),
	.w4(32'h3c0ae3ae),
	.w5(32'hbb310990),
	.w6(32'hbc9b4726),
	.w7(32'h3c75367b),
	.w8(32'h3c159b9c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaad4c),
	.w1(32'h3b0f2b30),
	.w2(32'hbaca6f58),
	.w3(32'h3b49808c),
	.w4(32'hbb46323a),
	.w5(32'h3b12838d),
	.w6(32'h3ba62b5b),
	.w7(32'hbbc56cbc),
	.w8(32'h3a216fa4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b5b0),
	.w1(32'h3b1ad67e),
	.w2(32'hbb87d847),
	.w3(32'h39e8e7f5),
	.w4(32'h39ee52a8),
	.w5(32'hbb067a7e),
	.w6(32'hbb3eb2f0),
	.w7(32'hba859274),
	.w8(32'h3b050045),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8c9da),
	.w1(32'h3b3d1a04),
	.w2(32'h3b0b66d9),
	.w3(32'h3ad48429),
	.w4(32'h3bee6cd7),
	.w5(32'hb9fea8f7),
	.w6(32'h3b94a215),
	.w7(32'h3c277c07),
	.w8(32'h3b4241fa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9aea7),
	.w1(32'h390e6c07),
	.w2(32'h3c1b65d9),
	.w3(32'hbb171d40),
	.w4(32'hbb9a7b68),
	.w5(32'h3c429127),
	.w6(32'h3ac08192),
	.w7(32'h3b21c08d),
	.w8(32'h3c5d06b8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae51fef),
	.w1(32'hbc64052c),
	.w2(32'h3b2b2fdc),
	.w3(32'hbabd22b0),
	.w4(32'hbc500011),
	.w5(32'hba8c75d8),
	.w6(32'hbb2b0347),
	.w7(32'hbba40152),
	.w8(32'hbb5b5842),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e110),
	.w1(32'hbb8db6f9),
	.w2(32'h39ef80e0),
	.w3(32'hbca31808),
	.w4(32'hbbcdc2c6),
	.w5(32'h3b4668c4),
	.w6(32'hbca28bf1),
	.w7(32'hbb946e3f),
	.w8(32'h3baec6e6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fee46),
	.w1(32'hb9e13108),
	.w2(32'h3aabfed1),
	.w3(32'hbbfc09e5),
	.w4(32'h3b525ce4),
	.w5(32'h3b163585),
	.w6(32'hbbaaafaf),
	.w7(32'h3beb8431),
	.w8(32'h3b28d305),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc0f42),
	.w1(32'hbb19f01a),
	.w2(32'hbb592566),
	.w3(32'h3b2043e5),
	.w4(32'hba2bd16e),
	.w5(32'hbaffb7d7),
	.w6(32'h3ba0dc2f),
	.w7(32'h3b0f3bf9),
	.w8(32'hb9dd517e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4475a0),
	.w1(32'h3b24fe4e),
	.w2(32'hbab7accd),
	.w3(32'h3ad2017c),
	.w4(32'h3b85c126),
	.w5(32'hbbc6d790),
	.w6(32'h3ae9f700),
	.w7(32'h3b996c5e),
	.w8(32'hbb27f7bc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d5e96),
	.w1(32'hb9f9affa),
	.w2(32'h3a650f92),
	.w3(32'hbc4e5ee4),
	.w4(32'h3bc204d3),
	.w5(32'hbba60c97),
	.w6(32'hbbdd2ba1),
	.w7(32'h3c3fc44c),
	.w8(32'hbbd3f11a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c588b),
	.w1(32'h3a20c826),
	.w2(32'hbbcc5f8c),
	.w3(32'hbb7dbdde),
	.w4(32'hbb8239d2),
	.w5(32'hbc24b95c),
	.w6(32'hbbc9b264),
	.w7(32'hbba53012),
	.w8(32'hbc1aa5de),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4f9fc),
	.w1(32'h3c2ea9f5),
	.w2(32'hbc85a9d4),
	.w3(32'h3c21d926),
	.w4(32'h3bf11cb3),
	.w5(32'hbcb5cc0d),
	.w6(32'h3c052ab0),
	.w7(32'h3b0c87c0),
	.w8(32'hbcb6d2f8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade4487),
	.w1(32'h3c5bb9dd),
	.w2(32'hbbf7d47d),
	.w3(32'h3bd9c6a0),
	.w4(32'h3c842cad),
	.w5(32'hbc90fcfa),
	.w6(32'h3c00411f),
	.w7(32'h399cc7f8),
	.w8(32'hbcaa4f3b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c445fe5),
	.w1(32'h3c7e1a0a),
	.w2(32'h3b94f091),
	.w3(32'h3c46f47e),
	.w4(32'h3c4047e1),
	.w5(32'hbc0dfb6d),
	.w6(32'h3c253305),
	.w7(32'h3b05b1c3),
	.w8(32'hbc85822f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule