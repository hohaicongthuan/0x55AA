module layer_10_featuremap_62(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b076b89),
	.w1(32'hbc2b7830),
	.w2(32'h3c70ef89),
	.w3(32'h3b22612a),
	.w4(32'hbc4a821f),
	.w5(32'h3c071369),
	.w6(32'hba96f363),
	.w7(32'hbb4a014e),
	.w8(32'hba8aa77f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c018163),
	.w1(32'hba51b1d6),
	.w2(32'h3bf1da15),
	.w3(32'h3c765766),
	.w4(32'h3ba666c2),
	.w5(32'h3c509009),
	.w6(32'h3c769a88),
	.w7(32'h3c34338e),
	.w8(32'h3c528644),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b047f),
	.w1(32'hbb129f1a),
	.w2(32'h3a2a9b0b),
	.w3(32'h3b8e8bd8),
	.w4(32'hbc115646),
	.w5(32'hbb1ddc00),
	.w6(32'h3c166bf5),
	.w7(32'hbb34beb1),
	.w8(32'hba90ca0c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7be42),
	.w1(32'hbb5e169b),
	.w2(32'hbc09b2ff),
	.w3(32'h38ffc7e9),
	.w4(32'h3ba15728),
	.w5(32'hbc10176a),
	.w6(32'hbb69426c),
	.w7(32'h3b1c335e),
	.w8(32'hba245dfa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870f2a),
	.w1(32'hbc23dd8a),
	.w2(32'h3b738627),
	.w3(32'hbb88d535),
	.w4(32'hb9888f9d),
	.w5(32'h3b2b38a8),
	.w6(32'hbb0f69d6),
	.w7(32'hbc778d09),
	.w8(32'h3b608089),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc78d20),
	.w1(32'hbb217b02),
	.w2(32'hbb16d199),
	.w3(32'h38a285ff),
	.w4(32'hbb2d1447),
	.w5(32'hbb00aa7f),
	.w6(32'hbaf1e527),
	.w7(32'hbc1d5ed6),
	.w8(32'hbb7c6bd4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cefc4),
	.w1(32'hb98c94f7),
	.w2(32'h39e6ef34),
	.w3(32'hbb8f913d),
	.w4(32'hba8d4738),
	.w5(32'h39fca159),
	.w6(32'hbbe7c5ef),
	.w7(32'hbb8537f3),
	.w8(32'hbc1b1256),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafed3b),
	.w1(32'hbbd9da91),
	.w2(32'h3c73d0f9),
	.w3(32'h3af0fff3),
	.w4(32'h3b539fe9),
	.w5(32'h3c023bee),
	.w6(32'hbc008afd),
	.w7(32'h3b09ae46),
	.w8(32'h3b0ce4f4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bc115),
	.w1(32'hbb8ee2e5),
	.w2(32'h3aba3056),
	.w3(32'h3c7899a7),
	.w4(32'h3be428ec),
	.w5(32'h3934bf1e),
	.w6(32'h3bb3cbd1),
	.w7(32'h3c3d9804),
	.w8(32'hbae94fb2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2381db),
	.w1(32'h3c1c6aef),
	.w2(32'h3c502f83),
	.w3(32'h3bc3335b),
	.w4(32'h3ac7e806),
	.w5(32'h3bf2532c),
	.w6(32'h3b94b865),
	.w7(32'h3aef6d4f),
	.w8(32'h3b922004),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228acf),
	.w1(32'h3b858ac1),
	.w2(32'hbaea926f),
	.w3(32'h3aac0e59),
	.w4(32'h3b0e072b),
	.w5(32'h3a893717),
	.w6(32'h39e60c2b),
	.w7(32'h3b026421),
	.w8(32'h3b4abfb0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f5d51),
	.w1(32'hbb3de679),
	.w2(32'h3babb8cc),
	.w3(32'h3ba8e2f9),
	.w4(32'hbbe36add),
	.w5(32'h3b8b652e),
	.w6(32'h3b506055),
	.w7(32'h3b257aa6),
	.w8(32'h3b41a222),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c323520),
	.w1(32'h3c0eb62d),
	.w2(32'h3c12e7db),
	.w3(32'h3bcec48a),
	.w4(32'h3b75019b),
	.w5(32'h3a712016),
	.w6(32'h3bb85c38),
	.w7(32'h3a88863a),
	.w8(32'h3987b3df),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85f66),
	.w1(32'hbb9a0295),
	.w2(32'h3b5f4633),
	.w3(32'hbb8cbd6e),
	.w4(32'hba79406a),
	.w5(32'hbba37fec),
	.w6(32'hbb8a0a0d),
	.w7(32'hbb0701a8),
	.w8(32'hba9c1aec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94d317),
	.w1(32'hbc61007a),
	.w2(32'hbaff9bd2),
	.w3(32'hbb6af515),
	.w4(32'hbac1e922),
	.w5(32'hbb370591),
	.w6(32'hba8d039f),
	.w7(32'hbbbb1492),
	.w8(32'hbbc38d0f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff63f2),
	.w1(32'h3b2a1c94),
	.w2(32'h3c0a4a9e),
	.w3(32'hbc111e95),
	.w4(32'hbbd679e9),
	.w5(32'h3b3dc5a7),
	.w6(32'hbb17b11f),
	.w7(32'hb9684f5a),
	.w8(32'h3885e236),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00b10),
	.w1(32'h3b840f5b),
	.w2(32'h3b1e0a17),
	.w3(32'hba3b86de),
	.w4(32'h3a8f3852),
	.w5(32'hb9667036),
	.w6(32'hbb3573a2),
	.w7(32'hba7c7853),
	.w8(32'h379fb585),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c246be6),
	.w1(32'hba45e4bb),
	.w2(32'h3c539daa),
	.w3(32'h3b89adca),
	.w4(32'hbb712a8c),
	.w5(32'h3be9f603),
	.w6(32'h3bf55bf4),
	.w7(32'hbb91693e),
	.w8(32'h3c20dc3e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f60791),
	.w1(32'hbae30705),
	.w2(32'h3caa5d5f),
	.w3(32'hbb866767),
	.w4(32'hbb1b1625),
	.w5(32'h3c49dc11),
	.w6(32'hbb0cc9b4),
	.w7(32'hbc07ca66),
	.w8(32'h3bba825d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7daa15),
	.w1(32'h3b5a48ec),
	.w2(32'hbb6eea0f),
	.w3(32'h3bbab426),
	.w4(32'h3c0a8d93),
	.w5(32'hbbb5c18c),
	.w6(32'h3aae358a),
	.w7(32'h3c02354b),
	.w8(32'hbbac2359),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3af01),
	.w1(32'hbc02d7e3),
	.w2(32'h3bcdd3e8),
	.w3(32'hbb9e3d1c),
	.w4(32'hbbb88f6c),
	.w5(32'h3b2fd1e0),
	.w6(32'hbb9f89d9),
	.w7(32'hbad80046),
	.w8(32'hba06065b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba953cc2),
	.w1(32'h3aa89e9a),
	.w2(32'hba33c2ba),
	.w3(32'h3983ef3e),
	.w4(32'hbbb4dc93),
	.w5(32'h3b4caa3e),
	.w6(32'hbb3504d3),
	.w7(32'hbb77e6cd),
	.w8(32'h3b95e5bd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c862e30),
	.w1(32'h3c2876fd),
	.w2(32'h3c101e20),
	.w3(32'h3c8d86d8),
	.w4(32'hbbb01ad3),
	.w5(32'h3c12d13a),
	.w6(32'h3cd9e335),
	.w7(32'h3c114a62),
	.w8(32'h3c5201d2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be66809),
	.w1(32'h3920caaf),
	.w2(32'h3b812d0b),
	.w3(32'h3b43429b),
	.w4(32'hbb92cbfa),
	.w5(32'h3a874734),
	.w6(32'h3b77c5c3),
	.w7(32'hbb0c6f07),
	.w8(32'hbb80b7ae),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b357813),
	.w1(32'hb97ae2a3),
	.w2(32'hbae9a0c1),
	.w3(32'h3ae0ca17),
	.w4(32'hbb83b2d5),
	.w5(32'hbbc67a72),
	.w6(32'h3a6490b0),
	.w7(32'hbc620e22),
	.w8(32'hbbe44d5e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51efca),
	.w1(32'hbc7e828b),
	.w2(32'hba497258),
	.w3(32'h3b9ba071),
	.w4(32'hb9920d2e),
	.w5(32'hbb8791db),
	.w6(32'hbaaaa96f),
	.w7(32'hbb1806f9),
	.w8(32'hbbd20f54),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba598c13),
	.w1(32'hbbe028ef),
	.w2(32'hb9b3576c),
	.w3(32'hb6f6bdaf),
	.w4(32'hbbbbb0bd),
	.w5(32'hba964e07),
	.w6(32'hbbc6f40a),
	.w7(32'hbb7e5098),
	.w8(32'hb9b31ba5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b244020),
	.w1(32'hbb27f253),
	.w2(32'h3ab802cd),
	.w3(32'h3a8c0d16),
	.w4(32'h37fb5d20),
	.w5(32'hbb90d93b),
	.w6(32'hbb1d5399),
	.w7(32'h3a082a51),
	.w8(32'hbc0d5cae),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfa736),
	.w1(32'h3bade2bf),
	.w2(32'hbcf54b97),
	.w3(32'hbb34621c),
	.w4(32'h3ba4478d),
	.w5(32'hbc585b6b),
	.w6(32'hba2a601d),
	.w7(32'h3bbe77c4),
	.w8(32'hbc24a7b3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6061df),
	.w1(32'hb8efb99f),
	.w2(32'h3b6dc295),
	.w3(32'h3d16021f),
	.w4(32'h3b8ebb95),
	.w5(32'hba3cdcfc),
	.w6(32'h3c6deb8d),
	.w7(32'hbc5dab4d),
	.w8(32'hba46a965),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcdec2),
	.w1(32'h3a8e3b35),
	.w2(32'hbc023b70),
	.w3(32'h3bc8de63),
	.w4(32'h3ad08b7f),
	.w5(32'hbc1e40be),
	.w6(32'h3b74586f),
	.w7(32'h3ad0d592),
	.w8(32'hbb3f46e6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8793e),
	.w1(32'hba6589e1),
	.w2(32'hbc0c9b84),
	.w3(32'h3cb2836a),
	.w4(32'hbbe3b140),
	.w5(32'hbb8bb8c1),
	.w6(32'h3c770161),
	.w7(32'hbc03aaa1),
	.w8(32'h3aeed3b9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c302b91),
	.w1(32'h3c04939c),
	.w2(32'h3c4aab65),
	.w3(32'h3cae6f10),
	.w4(32'h3bdff145),
	.w5(32'h3b44c2b0),
	.w6(32'h3c993250),
	.w7(32'hbb99e4ce),
	.w8(32'hba68d366),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ddda7),
	.w1(32'hbb33fd9e),
	.w2(32'hbb45cc38),
	.w3(32'hbbc73723),
	.w4(32'hbbafa451),
	.w5(32'h3b1e636f),
	.w6(32'hbc14cb83),
	.w7(32'hbbf04ffd),
	.w8(32'h3bb3e260),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f2497),
	.w1(32'h398a901d),
	.w2(32'h3906f59e),
	.w3(32'h3c452562),
	.w4(32'hbc911f1f),
	.w5(32'h3b3bc199),
	.w6(32'hbbf593a1),
	.w7(32'h3b2cff2d),
	.w8(32'h3b30a776),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55ff19),
	.w1(32'hbb410a5b),
	.w2(32'hbb53313b),
	.w3(32'hbaacb75e),
	.w4(32'hbb2f0238),
	.w5(32'h3cbc2070),
	.w6(32'h3b0bff33),
	.w7(32'hba5d6da2),
	.w8(32'h3bc03aa0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d29f20e),
	.w1(32'hbc374570),
	.w2(32'h3bda8e16),
	.w3(32'h3d117209),
	.w4(32'hbcb9df8e),
	.w5(32'hbaa5d0d0),
	.w6(32'h3c4f55d6),
	.w7(32'hbbf606a8),
	.w8(32'h3ba91d98),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c749d5e),
	.w1(32'h3ae9cc58),
	.w2(32'hbcc73a54),
	.w3(32'h3c591878),
	.w4(32'h3b652fb4),
	.w5(32'hbc1e56c1),
	.w6(32'h3c3e4b63),
	.w7(32'hbaa01730),
	.w8(32'hbc8649eb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8257e),
	.w1(32'h3c5073c5),
	.w2(32'hbbcfb5ec),
	.w3(32'h3baa2466),
	.w4(32'hbbd09f8e),
	.w5(32'hbc055ed5),
	.w6(32'h3a854fae),
	.w7(32'h3a1f6a9f),
	.w8(32'hbaebce23),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf888a6),
	.w1(32'h3b1d998a),
	.w2(32'hbb8950f1),
	.w3(32'hbb8910eb),
	.w4(32'h3b268b15),
	.w5(32'hbbfe839f),
	.w6(32'h3b250219),
	.w7(32'hbbc94eb8),
	.w8(32'hbbc73187),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb32516),
	.w1(32'hbc7345e8),
	.w2(32'hbb3866dd),
	.w3(32'hbbab36a7),
	.w4(32'hbc5f5354),
	.w5(32'hbb5600f5),
	.w6(32'hbb22f938),
	.w7(32'hbb9adcf2),
	.w8(32'hbba5ed58),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc322bb4),
	.w1(32'h3b7f0225),
	.w2(32'hbc0390c8),
	.w3(32'hbc474a77),
	.w4(32'hb919ced6),
	.w5(32'h3b8b22cc),
	.w6(32'hbbf1e47b),
	.w7(32'hbac88765),
	.w8(32'hbb7dff29),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f6721),
	.w1(32'h3c7b88ff),
	.w2(32'hbbb35319),
	.w3(32'h3ccc318e),
	.w4(32'h3b8f5fd4),
	.w5(32'hbb9549b6),
	.w6(32'h3c85d3a7),
	.w7(32'hbb83e86d),
	.w8(32'hbb95e644),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdbce8),
	.w1(32'h3b7c5f77),
	.w2(32'hba6e091f),
	.w3(32'h3c0b4554),
	.w4(32'h37fbaafa),
	.w5(32'hbc309e6a),
	.w6(32'h3c58b739),
	.w7(32'h3bc603a3),
	.w8(32'h3bd46fce),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81eac4),
	.w1(32'h3be1b439),
	.w2(32'hbc581760),
	.w3(32'h3beff613),
	.w4(32'h3c3ff008),
	.w5(32'hbc380fa2),
	.w6(32'h3c29a64a),
	.w7(32'hbc591f80),
	.w8(32'hbc75b352),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1d81d),
	.w1(32'h3c576fb4),
	.w2(32'h3c8689dc),
	.w3(32'h3d4355a4),
	.w4(32'h3c017359),
	.w5(32'h3b8de267),
	.w6(32'h3d01906e),
	.w7(32'hbc69bf07),
	.w8(32'h3baec3fa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082cda),
	.w1(32'hbb53bbb2),
	.w2(32'h3c9239c4),
	.w3(32'hbb58bdbd),
	.w4(32'h3c87944d),
	.w5(32'h3c38704e),
	.w6(32'h3b2529fb),
	.w7(32'h3b8967ae),
	.w8(32'hbb9df8ac),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b751d81),
	.w1(32'hbc786311),
	.w2(32'h3c3d6261),
	.w3(32'h3a162086),
	.w4(32'hbc993663),
	.w5(32'h3c278688),
	.w6(32'hbad6f436),
	.w7(32'hbc0ba8df),
	.w8(32'h3c8f813d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e9ea7),
	.w1(32'h3bd319ae),
	.w2(32'hba1e280d),
	.w3(32'h3bb554f7),
	.w4(32'h3b7d6dbf),
	.w5(32'h3b894649),
	.w6(32'h3bc4acb3),
	.w7(32'h3b391f6d),
	.w8(32'hbaedd729),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbcf4d),
	.w1(32'h3b37cff6),
	.w2(32'h3a72abdb),
	.w3(32'h3c482bc8),
	.w4(32'h3b1ff07f),
	.w5(32'h3c19baea),
	.w6(32'h3c0f7bb8),
	.w7(32'hbb54030f),
	.w8(32'hbb4f2496),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30aa29),
	.w1(32'hbb873837),
	.w2(32'hbb8d7802),
	.w3(32'hbc3a9bfd),
	.w4(32'hbc570e8d),
	.w5(32'hbc57333a),
	.w6(32'hbca84844),
	.w7(32'h39bce2cc),
	.w8(32'hbc3b918e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b15ad),
	.w1(32'hbb170c57),
	.w2(32'h3c5c7357),
	.w3(32'hbc67975e),
	.w4(32'h3b71798d),
	.w5(32'h3c5e5ae8),
	.w6(32'h3a1f964a),
	.w7(32'hbafd7dd6),
	.w8(32'hbbfa34f9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4bf88),
	.w1(32'hb9a18df5),
	.w2(32'h3b612e9b),
	.w3(32'hbc5753cf),
	.w4(32'h3bc068eb),
	.w5(32'hbb20b078),
	.w6(32'hbbdddf67),
	.w7(32'h3c366d08),
	.w8(32'hbb642237),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38b692),
	.w1(32'hbaf861a7),
	.w2(32'h3abb2c91),
	.w3(32'hba5c54ff),
	.w4(32'hbc472948),
	.w5(32'hbb5714bd),
	.w6(32'hb985fdd3),
	.w7(32'hb996584c),
	.w8(32'h3c92c4b4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ef82d),
	.w1(32'h3b9de6d8),
	.w2(32'hbb0b383b),
	.w3(32'h3c510746),
	.w4(32'hbb90d0b4),
	.w5(32'hbc708d92),
	.w6(32'h3af41f50),
	.w7(32'hbaf0701a),
	.w8(32'hbc2baec6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4011e2),
	.w1(32'hbb2ba5ea),
	.w2(32'hbc01e6dd),
	.w3(32'h3bdc2897),
	.w4(32'hbaaeb5b0),
	.w5(32'h3b52c746),
	.w6(32'hb97e3832),
	.w7(32'hbc2831bd),
	.w8(32'h3baa30ce),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3753f6),
	.w1(32'hbb076f3a),
	.w2(32'hbb3c32da),
	.w3(32'h3c1026e2),
	.w4(32'h3c6f8c29),
	.w5(32'hbc1e7ecc),
	.w6(32'h3b633ddf),
	.w7(32'hba4856d7),
	.w8(32'hbbb23921),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e906),
	.w1(32'h3a18bbc4),
	.w2(32'h3ace401d),
	.w3(32'hbb1b86c3),
	.w4(32'hbb788b77),
	.w5(32'h3a388ff1),
	.w6(32'hb9d1d393),
	.w7(32'hbba81b4e),
	.w8(32'h3ba9e068),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6cfc1),
	.w1(32'h3b221f22),
	.w2(32'hbba92397),
	.w3(32'hbb2237aa),
	.w4(32'h3aee0027),
	.w5(32'hbbdf2eb9),
	.w6(32'h383d13fb),
	.w7(32'h3bc7f1ea),
	.w8(32'hbb592cc1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb127a29),
	.w1(32'hbb9afd0d),
	.w2(32'h3abc978e),
	.w3(32'hbb72a689),
	.w4(32'h391a39a7),
	.w5(32'hbac4d3b1),
	.w6(32'hbb505db5),
	.w7(32'hbb3f4792),
	.w8(32'h3a384a34),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2bc4),
	.w1(32'h3bbc6beb),
	.w2(32'hbb328d89),
	.w3(32'h3c49edf7),
	.w4(32'h3b484ec3),
	.w5(32'hbb435488),
	.w6(32'h3c7bddee),
	.w7(32'hbb3166c7),
	.w8(32'h3acbc4bf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc633857),
	.w1(32'h3bc957a0),
	.w2(32'hbbc77a24),
	.w3(32'h3b497aef),
	.w4(32'h3babd6d2),
	.w5(32'hbc6cd3c2),
	.w6(32'h3a68f8e2),
	.w7(32'hba9120e0),
	.w8(32'h3be031ce),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e6481),
	.w1(32'h3aa0afff),
	.w2(32'h3b9542dd),
	.w3(32'hbc42fceb),
	.w4(32'h3b2695e6),
	.w5(32'h3bee6f6e),
	.w6(32'hba3c76d4),
	.w7(32'h3b77ab68),
	.w8(32'h3b3d0300),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb91cb8),
	.w1(32'hbb727558),
	.w2(32'hbbdaa85f),
	.w3(32'h3b4f54fd),
	.w4(32'hbb3e6ec7),
	.w5(32'hbb5d7e08),
	.w6(32'hbafe5bb7),
	.w7(32'hbb3d75d4),
	.w8(32'hbb4c6fa8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44608b),
	.w1(32'hbb05e1de),
	.w2(32'h3b3e0dd9),
	.w3(32'h3cb7a7c2),
	.w4(32'hbbe21d89),
	.w5(32'h39c2ed14),
	.w6(32'h3c732aa4),
	.w7(32'hbbb0404d),
	.w8(32'hbb627795),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5cea7),
	.w1(32'h3b1260fc),
	.w2(32'h3ba4f17c),
	.w3(32'hb9758e0f),
	.w4(32'hbb82d5bc),
	.w5(32'hba2c74c8),
	.w6(32'hbb272f68),
	.w7(32'hbb1aaa20),
	.w8(32'hbab79ccc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a6d3d),
	.w1(32'h3bc58940),
	.w2(32'h3c86c392),
	.w3(32'hbc7f6503),
	.w4(32'hbc0600ef),
	.w5(32'h3c6174e8),
	.w6(32'hbbe59fee),
	.w7(32'h3b32a8ac),
	.w8(32'h3be078d2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8610f4),
	.w1(32'hbac4e065),
	.w2(32'h3c514ae8),
	.w3(32'hbb6e01b5),
	.w4(32'hba157a64),
	.w5(32'h3c248693),
	.w6(32'hbc0c5110),
	.w7(32'hbb084b43),
	.w8(32'hbaa94473),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c579e3d),
	.w1(32'hbab96df4),
	.w2(32'h3c0442d7),
	.w3(32'h3b894e05),
	.w4(32'hba98f2f6),
	.w5(32'h3bb0d3a7),
	.w6(32'h3b082d43),
	.w7(32'h3b5816e0),
	.w8(32'h3c11ad44),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff9a60),
	.w1(32'hbbcb9961),
	.w2(32'h3bfd2658),
	.w3(32'h3bf7d518),
	.w4(32'hbb9406d2),
	.w5(32'hbb4d2ecd),
	.w6(32'h3bde2d53),
	.w7(32'hbbd49837),
	.w8(32'hbc3a1419),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6e888),
	.w1(32'h3bafeef4),
	.w2(32'h3b64a58f),
	.w3(32'hb92a0751),
	.w4(32'hbaf35125),
	.w5(32'h3a7953df),
	.w6(32'h3b1e7570),
	.w7(32'hbb33b921),
	.w8(32'hbbf805f1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4f130),
	.w1(32'hba6b5c8e),
	.w2(32'h3bce6220),
	.w3(32'hbaf556fe),
	.w4(32'hbbdcfb28),
	.w5(32'h3b7bd34d),
	.w6(32'hbb36de36),
	.w7(32'hba84458e),
	.w8(32'h3b03ac11),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba377e),
	.w1(32'hbc2313ce),
	.w2(32'hbcd027f6),
	.w3(32'hbc91b9de),
	.w4(32'hbb3f5d31),
	.w5(32'hbd20b796),
	.w6(32'hbc351560),
	.w7(32'hbac538b1),
	.w8(32'hbcb48b76),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf5cfc),
	.w1(32'h3bfb0a4e),
	.w2(32'hbbc4265e),
	.w3(32'h3d06db0d),
	.w4(32'hbc0c27fc),
	.w5(32'hbbaf9ac2),
	.w6(32'h3c79a8f9),
	.w7(32'hbb71c5b1),
	.w8(32'hba77674a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d43b1),
	.w1(32'hb832509f),
	.w2(32'h3a6ce903),
	.w3(32'h3c19e1ad),
	.w4(32'h3b73507d),
	.w5(32'hba6acf5b),
	.w6(32'h3c0ebaed),
	.w7(32'hbad44268),
	.w8(32'hbbcb444c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68b293),
	.w1(32'hbbb3f461),
	.w2(32'h3b955313),
	.w3(32'hbba0c677),
	.w4(32'hbc30be00),
	.w5(32'h3b16fa8f),
	.w6(32'hbb9f3961),
	.w7(32'hbbe01867),
	.w8(32'hbab55d1d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8781d3),
	.w1(32'hbc12273d),
	.w2(32'h3b10d068),
	.w3(32'h3c0fc904),
	.w4(32'hbc795847),
	.w5(32'hbb28f898),
	.w6(32'h3c3c8787),
	.w7(32'h3c150758),
	.w8(32'h3b8de57d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf34af2),
	.w1(32'hbc87c3b6),
	.w2(32'hbc23844c),
	.w3(32'h3c6ae16f),
	.w4(32'hbc6720f1),
	.w5(32'hbc4c8fc3),
	.w6(32'h3bbd783f),
	.w7(32'hba4c3aa7),
	.w8(32'hbc659ec0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b57fb),
	.w1(32'h3bb38c35),
	.w2(32'h3b5f7d16),
	.w3(32'h3b9c5b91),
	.w4(32'h3c21107e),
	.w5(32'hb93c7127),
	.w6(32'hbb2edcdc),
	.w7(32'h390bae3d),
	.w8(32'h399456cf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ebdc5),
	.w1(32'hbb1a843d),
	.w2(32'h3c769b85),
	.w3(32'hba1a3fed),
	.w4(32'hbc0f45c4),
	.w5(32'h3a295928),
	.w6(32'hb9bf01b6),
	.w7(32'hbb5a4fe6),
	.w8(32'hbbce07d1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdab9f),
	.w1(32'hbb50e4c6),
	.w2(32'h3c014da9),
	.w3(32'h3b2b5a91),
	.w4(32'h3bab6ce2),
	.w5(32'h3a97eb0a),
	.w6(32'h388fb1ec),
	.w7(32'hbaa15f0e),
	.w8(32'hbb361ba0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbee3e3),
	.w1(32'hbb29d04e),
	.w2(32'h3ce7cb85),
	.w3(32'hb9a2e421),
	.w4(32'hbbc5fe7c),
	.w5(32'h3d5390d7),
	.w6(32'h3a59f4d0),
	.w7(32'hbb66a0f5),
	.w8(32'h3d3c998c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf48e82),
	.w1(32'hbc84ce95),
	.w2(32'hbb981fd4),
	.w3(32'h3ced248e),
	.w4(32'hbbe14160),
	.w5(32'hbb92c674),
	.w6(32'h3c118595),
	.w7(32'h3c453f84),
	.w8(32'hbb90e066),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e4f1f),
	.w1(32'hbbb2be99),
	.w2(32'h3bebb7be),
	.w3(32'hbbe58826),
	.w4(32'hbbd73f09),
	.w5(32'hba96c245),
	.w6(32'hbc0f8095),
	.w7(32'hbc12b1ad),
	.w8(32'h3b0d9110),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5dac5),
	.w1(32'hbbb0d50f),
	.w2(32'h3b9ddd1e),
	.w3(32'hbcae8ee6),
	.w4(32'hbb0046ea),
	.w5(32'h3ba3e0db),
	.w6(32'hbc01b07d),
	.w7(32'hb8e9b074),
	.w8(32'hbc0a3f42),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4e2f2),
	.w1(32'h3c028a86),
	.w2(32'h3ac52781),
	.w3(32'hbca85cc8),
	.w4(32'h3c27ab45),
	.w5(32'hbb7726f9),
	.w6(32'hbc29d4c4),
	.w7(32'hbb43749c),
	.w8(32'hbbf3b7c2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34c99e),
	.w1(32'h3b4e95fd),
	.w2(32'hbb0bf2ce),
	.w3(32'h3b62f79d),
	.w4(32'hbae0ed70),
	.w5(32'hbb791987),
	.w6(32'h3a0d138e),
	.w7(32'hb991cd84),
	.w8(32'hbb948ab4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8780d),
	.w1(32'h3ab61181),
	.w2(32'h3be0cd64),
	.w3(32'hbae27ac0),
	.w4(32'hba73051f),
	.w5(32'h3c28eedc),
	.w6(32'hbb5a544e),
	.w7(32'h3aab7879),
	.w8(32'hbba90ccd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb051d1c),
	.w1(32'hbb4c6dec),
	.w2(32'h3c306d16),
	.w3(32'hbc84ecc4),
	.w4(32'h3bb53774),
	.w5(32'hbb2d09d0),
	.w6(32'hbbae5350),
	.w7(32'h3bbb78fb),
	.w8(32'h3b7b7ff7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c426a8d),
	.w1(32'h3bd481db),
	.w2(32'h3ba72be1),
	.w3(32'h39fa78ad),
	.w4(32'hba1e7a7b),
	.w5(32'h3b9b5121),
	.w6(32'h399b5f3d),
	.w7(32'hbb4db03b),
	.w8(32'h3c39ee9e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74bfbf),
	.w1(32'h3b95931a),
	.w2(32'h3bf4ddbb),
	.w3(32'h3bcef6b0),
	.w4(32'h3ba353d0),
	.w5(32'hbb6efcb2),
	.w6(32'h3b9e3caf),
	.w7(32'h3b062b89),
	.w8(32'h3b82028a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24ad53),
	.w1(32'h3c36edef),
	.w2(32'hba86d771),
	.w3(32'hbc023679),
	.w4(32'hbc1f5a92),
	.w5(32'hbb704d91),
	.w6(32'h3b7928cd),
	.w7(32'hba761bf4),
	.w8(32'hbabc3ca6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c171d),
	.w1(32'hbbda0231),
	.w2(32'hbbecf69b),
	.w3(32'hbb53bbac),
	.w4(32'hbbb69c8a),
	.w5(32'hbbccc922),
	.w6(32'hbb783916),
	.w7(32'hbbb0431f),
	.w8(32'hbba5593a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696be1),
	.w1(32'h3a9909f0),
	.w2(32'h3c89aa3d),
	.w3(32'h3bd93322),
	.w4(32'hbae4db6c),
	.w5(32'h3c2ca0c1),
	.w6(32'h3c234d95),
	.w7(32'h3bb79d9f),
	.w8(32'h3acd6d35),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5021),
	.w1(32'hbad0a07d),
	.w2(32'h3c773d60),
	.w3(32'hbbdb3d62),
	.w4(32'hbaee99ae),
	.w5(32'hbc0f0bb5),
	.w6(32'h3bf81c38),
	.w7(32'h3ba69839),
	.w8(32'hba9dd64a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab9397),
	.w1(32'h3c3ece5b),
	.w2(32'hbc99afd0),
	.w3(32'h3ccde7f3),
	.w4(32'hbb7bad45),
	.w5(32'hbc5d96d2),
	.w6(32'h3cdb0bca),
	.w7(32'hbcaa4291),
	.w8(32'hbc52e5c9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dfe58),
	.w1(32'hbb8a44c2),
	.w2(32'hbc4d685b),
	.w3(32'hbc2de305),
	.w4(32'hbc2ec8a0),
	.w5(32'hbc198aef),
	.w6(32'hbc0fcfa7),
	.w7(32'hbbfca104),
	.w8(32'h3aef2e55),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3090bd),
	.w1(32'h3c2eee07),
	.w2(32'h3ca79ec6),
	.w3(32'h3c521e41),
	.w4(32'h3c6e9f91),
	.w5(32'h3be23ca4),
	.w6(32'h3c52a02c),
	.w7(32'h3c4b625f),
	.w8(32'hbb0b6441),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c324044),
	.w1(32'hbb5a6b5f),
	.w2(32'h3c4e802d),
	.w3(32'h3b49f7a4),
	.w4(32'hbc553f8e),
	.w5(32'h3b63876f),
	.w6(32'hbb2356a3),
	.w7(32'hbb471c60),
	.w8(32'hb85f4884),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb726951c),
	.w1(32'hbb2c9b77),
	.w2(32'hbc7e422c),
	.w3(32'hb9c3f535),
	.w4(32'hbbf7113a),
	.w5(32'hbc4bd2a8),
	.w6(32'h3b9351f2),
	.w7(32'hbc063675),
	.w8(32'hbb0801c7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d093434),
	.w1(32'hbb8289af),
	.w2(32'hbcdd379e),
	.w3(32'h3d251bbc),
	.w4(32'hbc8917af),
	.w5(32'hbc7eae05),
	.w6(32'h3ca848bf),
	.w7(32'hbc5fb43a),
	.w8(32'hbc794723),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb8c22),
	.w1(32'hba202492),
	.w2(32'h3bb43882),
	.w3(32'h3cf238c5),
	.w4(32'hbc8cc527),
	.w5(32'h3aee4d7f),
	.w6(32'h3c31aa7a),
	.w7(32'hbcd5b22a),
	.w8(32'hbbcffe06),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83813c),
	.w1(32'h3c21e21d),
	.w2(32'h3bc20f97),
	.w3(32'h3bc17d87),
	.w4(32'h3a5377b6),
	.w5(32'hbaf1a9ba),
	.w6(32'h3bfb75ec),
	.w7(32'h39d32afa),
	.w8(32'h3bbd97a1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf93bf8),
	.w1(32'hbb3e3a91),
	.w2(32'hbc01780f),
	.w3(32'hbbcbb986),
	.w4(32'h3b7e0435),
	.w5(32'hbc282e7d),
	.w6(32'hb93bac19),
	.w7(32'hbb848a14),
	.w8(32'hbc8a9963),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc148075),
	.w1(32'h3b295758),
	.w2(32'h3c5187e1),
	.w3(32'hb8d45e03),
	.w4(32'h3b017308),
	.w5(32'h3a3ab52e),
	.w6(32'hbc5944a7),
	.w7(32'h3ab4f8a2),
	.w8(32'hbb801868),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91517c4),
	.w1(32'hba838383),
	.w2(32'h3b45c26a),
	.w3(32'hbbac4bfd),
	.w4(32'hba463aa4),
	.w5(32'hbab2aaea),
	.w6(32'h3a0962a3),
	.w7(32'h3aa10dc9),
	.w8(32'hbc4a1172),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86907d),
	.w1(32'h3a60c7f3),
	.w2(32'hbb87ed1c),
	.w3(32'hbb63edeb),
	.w4(32'hba8a9742),
	.w5(32'hbbc00aac),
	.w6(32'hb5c32a54),
	.w7(32'h3b37c350),
	.w8(32'hbc056968),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a0342),
	.w1(32'h3be770a0),
	.w2(32'h3affc5df),
	.w3(32'h3afe94aa),
	.w4(32'h3ba2eb7f),
	.w5(32'hbc535252),
	.w6(32'hbafb0a74),
	.w7(32'h3ac0238e),
	.w8(32'h3b5f03ca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56ee4),
	.w1(32'h3bfb5886),
	.w2(32'hbc0fb8c6),
	.w3(32'hbba9b951),
	.w4(32'h3bf8b303),
	.w5(32'hbc368f86),
	.w6(32'hbb1e9a97),
	.w7(32'h3c3db042),
	.w8(32'hbb15774b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e5a4d),
	.w1(32'hbb550d92),
	.w2(32'hbcb18d79),
	.w3(32'h3cb870be),
	.w4(32'hbbfec2ec),
	.w5(32'hbc59d10f),
	.w6(32'h3c1224cc),
	.w7(32'hbc5311a8),
	.w8(32'hbbb7aa06),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd822f),
	.w1(32'h3c9c1374),
	.w2(32'hbbaeda36),
	.w3(32'h3c112023),
	.w4(32'h3c865410),
	.w5(32'h3ab32ac0),
	.w6(32'h3c5f9e7a),
	.w7(32'h3bd22d31),
	.w8(32'h3b230559),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa8810),
	.w1(32'hb9844515),
	.w2(32'hbafe07f2),
	.w3(32'hb9f5a692),
	.w4(32'h3b640383),
	.w5(32'h3ca41c47),
	.w6(32'h3b4be874),
	.w7(32'h3b2645a9),
	.w8(32'h3cabed24),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb73af1),
	.w1(32'hbcc28d20),
	.w2(32'hbc455623),
	.w3(32'h3cbd9785),
	.w4(32'hbcc68549),
	.w5(32'hbc23604e),
	.w6(32'h3bd18d8a),
	.w7(32'hbbebef7f),
	.w8(32'h3a8b35c8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4facf0),
	.w1(32'h3c68a5bd),
	.w2(32'hb90fc3b8),
	.w3(32'h3c88c538),
	.w4(32'h3b8dbcd0),
	.w5(32'hbbf4da72),
	.w6(32'h3c43cdf4),
	.w7(32'h3bdf9b12),
	.w8(32'hbbad6f02),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80f05),
	.w1(32'h3a4b6730),
	.w2(32'h3ba1b8ca),
	.w3(32'h3c04be80),
	.w4(32'hbb4622cf),
	.w5(32'h3abb0257),
	.w6(32'h3b80e9d7),
	.w7(32'h3a25a00a),
	.w8(32'hba8850da),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaec7d),
	.w1(32'h3929ad69),
	.w2(32'hbad80743),
	.w3(32'hba5b8949),
	.w4(32'hbb00afe8),
	.w5(32'hbae75f0c),
	.w6(32'hbb87b362),
	.w7(32'hbaf6053b),
	.w8(32'hbb685072),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25fde1),
	.w1(32'h3bd443a6),
	.w2(32'h39bd4184),
	.w3(32'h390c31a2),
	.w4(32'h3b355c8f),
	.w5(32'hbb550528),
	.w6(32'h3976c8e3),
	.w7(32'h3b311e2c),
	.w8(32'hbaec28ed),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac13c83),
	.w1(32'hbb69fc3a),
	.w2(32'hbb11b1f6),
	.w3(32'hbb436b9f),
	.w4(32'hbb5a5b67),
	.w5(32'h3b36678a),
	.w6(32'hbb00dd37),
	.w7(32'hbb40bc6a),
	.w8(32'h3bb48435),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a0330),
	.w1(32'hbbce6c34),
	.w2(32'hbc37d735),
	.w3(32'h3c866290),
	.w4(32'hbbc267e3),
	.w5(32'hbc209b55),
	.w6(32'h3bebb9eb),
	.w7(32'hbb80e125),
	.w8(32'hbc06670e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd7aa72),
	.w1(32'hbb0eeffe),
	.w2(32'hbc11dceb),
	.w3(32'h3cbdb04e),
	.w4(32'hbc375ce7),
	.w5(32'hbc583c27),
	.w6(32'h3c3865f2),
	.w7(32'hbcb9c79e),
	.w8(32'hbbd43328),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc746479),
	.w1(32'h3aa132ad),
	.w2(32'hbb1031b7),
	.w3(32'hbc40c8e6),
	.w4(32'h3bb7e732),
	.w5(32'hbb75fee0),
	.w6(32'h3ba5fac6),
	.w7(32'hbb8b23e9),
	.w8(32'hba60189f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac47a48),
	.w1(32'hbae67978),
	.w2(32'h3b9df972),
	.w3(32'hbabe828c),
	.w4(32'hbb1df372),
	.w5(32'h3bc4ad97),
	.w6(32'h3a2377ca),
	.w7(32'hb9a14450),
	.w8(32'h3be2fb9d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7af36),
	.w1(32'h3a48ea63),
	.w2(32'h3b13514c),
	.w3(32'h3be333d3),
	.w4(32'h3b9330aa),
	.w5(32'h3be1034a),
	.w6(32'h3bbb359e),
	.w7(32'h3b0a29fc),
	.w8(32'h3c065f4c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd656c6),
	.w1(32'hbc9a8099),
	.w2(32'hbb91502f),
	.w3(32'h3c10c183),
	.w4(32'hbc4e9416),
	.w5(32'hbc10de65),
	.w6(32'hb9de1cb1),
	.w7(32'hbc8b1133),
	.w8(32'hbbb9fd1b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05764b),
	.w1(32'h3b51d099),
	.w2(32'h3c66b7d7),
	.w3(32'hbb1af575),
	.w4(32'h3af3f2b8),
	.w5(32'h3baf2786),
	.w6(32'h3a5defe9),
	.w7(32'hbac34402),
	.w8(32'hbb1ed7c8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5522fa),
	.w1(32'hbb99b29c),
	.w2(32'hbb81ead0),
	.w3(32'hbc9cea09),
	.w4(32'h39f27492),
	.w5(32'h3bfec995),
	.w6(32'hbc94b517),
	.w7(32'hbbdb92e9),
	.w8(32'hbb4a3eba),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88bf7e),
	.w1(32'hbc0d5888),
	.w2(32'h3a1baefa),
	.w3(32'hbc982bad),
	.w4(32'h3a34f129),
	.w5(32'h3b42aca7),
	.w6(32'hbc7eb92c),
	.w7(32'h3b4c4486),
	.w8(32'h3b40fd70),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85adb9),
	.w1(32'hbb9211ad),
	.w2(32'h3c01778c),
	.w3(32'hbc854a28),
	.w4(32'h3b6fcb8f),
	.w5(32'hbab05a99),
	.w6(32'hbc2cd2f7),
	.w7(32'hbbab0c5f),
	.w8(32'h3bd50273),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfc32c),
	.w1(32'hbb94115e),
	.w2(32'h3c2599e5),
	.w3(32'h3aa9e0e8),
	.w4(32'hbc340191),
	.w5(32'h3b9aed7d),
	.w6(32'hbb4e0a3e),
	.w7(32'hbba5a72b),
	.w8(32'hba33c877),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82d174),
	.w1(32'hbbfe7b0c),
	.w2(32'hbcbd0443),
	.w3(32'hbc4e5d79),
	.w4(32'hbaeb0bda),
	.w5(32'hbcd27ddb),
	.w6(32'hbc1427a1),
	.w7(32'h3b7b7376),
	.w8(32'hbc004e8d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083c0a),
	.w1(32'hbc1ec980),
	.w2(32'hbc6af765),
	.w3(32'h3c9871f9),
	.w4(32'hbc94b8f3),
	.w5(32'hbc4dfda7),
	.w6(32'h3c134288),
	.w7(32'hbc6a3834),
	.w8(32'hbc037501),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacff7d7),
	.w1(32'h3c43c3a2),
	.w2(32'h3c7e10d4),
	.w3(32'h3a8b36c9),
	.w4(32'hbac314df),
	.w5(32'hbb188156),
	.w6(32'h3bab36e6),
	.w7(32'h3b0d5c77),
	.w8(32'hbb154dbe),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31bc4e),
	.w1(32'hbc21d050),
	.w2(32'h3c0bd2c8),
	.w3(32'hbac402e6),
	.w4(32'h3ba4898e),
	.w5(32'h3cb91430),
	.w6(32'h3c377582),
	.w7(32'h3ba9f9ba),
	.w8(32'h3ccff480),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f9fe6),
	.w1(32'h3c255db2),
	.w2(32'hbb4e5f4b),
	.w3(32'h3d3acc7a),
	.w4(32'h3c5795f5),
	.w5(32'hbb94ec0f),
	.w6(32'h3d14e0d0),
	.w7(32'hbc220d81),
	.w8(32'hbaad9295),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c512),
	.w1(32'h3ad6d4df),
	.w2(32'h3c95d0d0),
	.w3(32'h3c11b084),
	.w4(32'hbaed770a),
	.w5(32'h3c02695d),
	.w6(32'h3c7e2dd0),
	.w7(32'h3b388c0b),
	.w8(32'h3c0bde3f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30f1cb),
	.w1(32'hbb932a26),
	.w2(32'hbba09f44),
	.w3(32'hbbc2c817),
	.w4(32'h388b3681),
	.w5(32'hbb86f29f),
	.w6(32'hb8b5a416),
	.w7(32'hba47e603),
	.w8(32'hbc6c85bc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03ae84),
	.w1(32'h3c1a569c),
	.w2(32'h3b68d8ec),
	.w3(32'h3b631c86),
	.w4(32'h3a6f1da6),
	.w5(32'hbb984ef1),
	.w6(32'hba93d0d9),
	.w7(32'h3b677146),
	.w8(32'hbb8c7784),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b455cf9),
	.w1(32'hba7f392a),
	.w2(32'h3c77d94f),
	.w3(32'hbc9ba1aa),
	.w4(32'hbc888b0f),
	.w5(32'h3c1e5631),
	.w6(32'hbc1a12a9),
	.w7(32'hbbfe791c),
	.w8(32'h3c52f169),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43ab06),
	.w1(32'hbb2219f0),
	.w2(32'hbbc9a0c5),
	.w3(32'h3aa2ba09),
	.w4(32'hbafdc801),
	.w5(32'hbb575e28),
	.w6(32'h3af082eb),
	.w7(32'hba8f3374),
	.w8(32'hbbc30d8e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1af12c),
	.w1(32'h3c003e1d),
	.w2(32'h3b48e72d),
	.w3(32'h3c11054b),
	.w4(32'h3bdc3f2d),
	.w5(32'h3b2cf512),
	.w6(32'h3c33896f),
	.w7(32'hbb17363f),
	.w8(32'h3bcd3a6d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5396ec),
	.w1(32'h3afc7ddf),
	.w2(32'hba620edb),
	.w3(32'h3b62a27d),
	.w4(32'h38aab53c),
	.w5(32'h3bab4094),
	.w6(32'h3b7096af),
	.w7(32'h3b559e4c),
	.w8(32'hbb1ca4c2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9754aa),
	.w1(32'hbbc1a5cd),
	.w2(32'h3ac0dd4b),
	.w3(32'h3b9e363f),
	.w4(32'h39dcd9c1),
	.w5(32'hbc79fe17),
	.w6(32'h3c4875f9),
	.w7(32'hbaca1b72),
	.w8(32'hbbead533),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f484a),
	.w1(32'hbc9f8a12),
	.w2(32'h3b2dfb1e),
	.w3(32'h3be1bc98),
	.w4(32'hbc865424),
	.w5(32'hb8d7a2a3),
	.w6(32'h39d7817b),
	.w7(32'h3b7595fc),
	.w8(32'hbba7503d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9822170),
	.w1(32'h39032369),
	.w2(32'h3ad7d96c),
	.w3(32'hbb2f4d13),
	.w4(32'hbbb71ad0),
	.w5(32'hb961ae4b),
	.w6(32'hbbcbb71e),
	.w7(32'hbb9b553d),
	.w8(32'hb9d1b04a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f4efa),
	.w1(32'hba95fbe8),
	.w2(32'hbad62f3a),
	.w3(32'hbaaeb3ae),
	.w4(32'hba27e379),
	.w5(32'hbb9578ec),
	.w6(32'hba5b239e),
	.w7(32'h39fbd7a7),
	.w8(32'hbb303485),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baafcf3),
	.w1(32'h3c4f3a6b),
	.w2(32'h39db9f66),
	.w3(32'hbb8d1abb),
	.w4(32'h3bd7add4),
	.w5(32'hba84ec19),
	.w6(32'h3ac8d60d),
	.w7(32'h3c09746e),
	.w8(32'h3a03c887),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aedd8),
	.w1(32'h3b58a4f9),
	.w2(32'hbc73fe2d),
	.w3(32'h3b88efd7),
	.w4(32'h3997fd91),
	.w5(32'hbc857b6f),
	.w6(32'h3c07e305),
	.w7(32'h38ecdf3b),
	.w8(32'hbadf5eeb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f7e67),
	.w1(32'h3bd5405d),
	.w2(32'h3c7179c3),
	.w3(32'hbaaebeb0),
	.w4(32'hbb0dc57e),
	.w5(32'h3b7565dc),
	.w6(32'hbab444e4),
	.w7(32'hbb45fdec),
	.w8(32'h3c02c04f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0062),
	.w1(32'hbaab0185),
	.w2(32'hbc3788f5),
	.w3(32'hbb92c302),
	.w4(32'h3b374dc6),
	.w5(32'hbc8c8fd1),
	.w6(32'h3b665186),
	.w7(32'h3b97932a),
	.w8(32'hbb5f0860),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17785b),
	.w1(32'h3baf025d),
	.w2(32'h3b221fe3),
	.w3(32'hbb080f6d),
	.w4(32'h3c397f31),
	.w5(32'hbb940812),
	.w6(32'h390182f6),
	.w7(32'h3c5bd265),
	.w8(32'hbb90f95e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb3cea),
	.w1(32'h3a85c123),
	.w2(32'h3ae5aff6),
	.w3(32'h398673a7),
	.w4(32'hbb22ac28),
	.w5(32'hb8ce4b1c),
	.w6(32'hbb8e0122),
	.w7(32'hbc169b27),
	.w8(32'h3822fb42),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c2478),
	.w1(32'hba410c78),
	.w2(32'h3c43255f),
	.w3(32'h3ae44e1c),
	.w4(32'hbbd5c4d0),
	.w5(32'h3c3e6d41),
	.w6(32'h3b616c45),
	.w7(32'hbbff8065),
	.w8(32'h3bb6a7ff),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce67ef),
	.w1(32'hbb58513a),
	.w2(32'hbb32563a),
	.w3(32'h3ab24af3),
	.w4(32'hbbc36255),
	.w5(32'h3c2ade9e),
	.w6(32'h3a852fbf),
	.w7(32'hbbf93a3b),
	.w8(32'h3bceb435),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1828e),
	.w1(32'h3cf13ecb),
	.w2(32'h3c03fea9),
	.w3(32'h3d189f7e),
	.w4(32'h3c3cdb62),
	.w5(32'h3b402cd8),
	.w6(32'h3cbd5e2f),
	.w7(32'h3b9690c3),
	.w8(32'hbb26464f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4ca82),
	.w1(32'hbc1154cc),
	.w2(32'hbb0aab8b),
	.w3(32'hbbb6ef8d),
	.w4(32'hbc2cc756),
	.w5(32'hbb4af0f7),
	.w6(32'hbb264a92),
	.w7(32'h3b394356),
	.w8(32'h39ba4176),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b883cdd),
	.w1(32'hba323d8b),
	.w2(32'h3c323b6f),
	.w3(32'h3bda26ac),
	.w4(32'hbb00b99b),
	.w5(32'h3b393f16),
	.w6(32'h3b94f8b1),
	.w7(32'hba7ae337),
	.w8(32'hbb7c2b4d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86aaae),
	.w1(32'h3c626713),
	.w2(32'h3c3ebfb1),
	.w3(32'h3c23427f),
	.w4(32'h3b2e1e7d),
	.w5(32'hbba46eb0),
	.w6(32'h3b983db3),
	.w7(32'hbb153b82),
	.w8(32'hbad40118),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5834c1),
	.w1(32'h3ae1cc5a),
	.w2(32'hbbabaf36),
	.w3(32'h3c6699cb),
	.w4(32'h3c8c152a),
	.w5(32'hbbc766de),
	.w6(32'hbc145d21),
	.w7(32'hbb96f290),
	.w8(32'hbad54876),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae33a97),
	.w1(32'hbb1b56ea),
	.w2(32'hbb40655d),
	.w3(32'hbb9f680e),
	.w4(32'hbb81c4cf),
	.w5(32'hbba3b768),
	.w6(32'hba6f2141),
	.w7(32'h3b03ad35),
	.w8(32'hba07e221),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d9435),
	.w1(32'h3c4045af),
	.w2(32'h3b279cdc),
	.w3(32'hbb3f19d8),
	.w4(32'h3c6465c2),
	.w5(32'h3bc764a3),
	.w6(32'hbc60212a),
	.w7(32'hbb09bd2e),
	.w8(32'h3ab9eb9f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b594d30),
	.w1(32'h3b8c2f12),
	.w2(32'h3c2b1e47),
	.w3(32'h3c11adb2),
	.w4(32'h3b9494ac),
	.w5(32'h3b90b146),
	.w6(32'h3be06dfe),
	.w7(32'h3c148f2f),
	.w8(32'h3c1cf190),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9daef6),
	.w1(32'hba12b5b7),
	.w2(32'h3c0c18e2),
	.w3(32'hbae32140),
	.w4(32'hbbace822),
	.w5(32'h3c02826a),
	.w6(32'hbba579ca),
	.w7(32'hbbf69b6b),
	.w8(32'hbba56b24),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd537),
	.w1(32'hbc366f28),
	.w2(32'hbacdee4c),
	.w3(32'h3c1a242f),
	.w4(32'h3b77b4ea),
	.w5(32'hbb335655),
	.w6(32'h3bd04b67),
	.w7(32'h3c7b7d55),
	.w8(32'hbaff4782),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75e03),
	.w1(32'hbbad6fd7),
	.w2(32'h3ca1c381),
	.w3(32'h3ac35613),
	.w4(32'hbb172d19),
	.w5(32'h3c1d5942),
	.w6(32'h3b4c66ec),
	.w7(32'h3942b460),
	.w8(32'hb918556c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf4915),
	.w1(32'h3c449ce5),
	.w2(32'h3b86dbf7),
	.w3(32'h3d217de1),
	.w4(32'h3cfa361c),
	.w5(32'hbb9ffbf3),
	.w6(32'h3c94b8b0),
	.w7(32'h3d2abee1),
	.w8(32'h3ab951c7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93e995),
	.w1(32'hbb3a3172),
	.w2(32'hbb909ace),
	.w3(32'hbb5f43cc),
	.w4(32'hbbccb15c),
	.w5(32'hbba5d9e5),
	.w6(32'hbb461a45),
	.w7(32'hb9dfcada),
	.w8(32'h3bf40182),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc49175),
	.w1(32'hbc049829),
	.w2(32'h3b22bedc),
	.w3(32'hbca838c5),
	.w4(32'hbc957af5),
	.w5(32'h3ac02471),
	.w6(32'h3be22068),
	.w7(32'h3b91cd50),
	.w8(32'hbbb5bc7b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f02e0),
	.w1(32'h3c22d9aa),
	.w2(32'h3a8becbc),
	.w3(32'h3b4c2aa0),
	.w4(32'h3c4b152d),
	.w5(32'h39d5f853),
	.w6(32'hbb99b717),
	.w7(32'hbc30432b),
	.w8(32'hb99c6267),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e1c2),
	.w1(32'h3b9d7021),
	.w2(32'hbb4ad7fa),
	.w3(32'h3b433995),
	.w4(32'hbae78648),
	.w5(32'hb9e23fee),
	.w6(32'h3b3d889a),
	.w7(32'h3b6e0880),
	.w8(32'h3c49c8a2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb983e5),
	.w1(32'hbc79fd27),
	.w2(32'hba54d6e7),
	.w3(32'hbc204646),
	.w4(32'hbc36e773),
	.w5(32'h3bb3fb13),
	.w6(32'h3c69660f),
	.w7(32'h3c90d724),
	.w8(32'hbbf684fa),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb04b8e),
	.w1(32'hbb9d4e91),
	.w2(32'h3b380552),
	.w3(32'hbb6e5d71),
	.w4(32'hbbb24037),
	.w5(32'hbb25e9cb),
	.w6(32'hbc5669cd),
	.w7(32'hbc7c7f0e),
	.w8(32'hbc098aee),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c553c),
	.w1(32'h3b80b388),
	.w2(32'hbb27115e),
	.w3(32'h3af12807),
	.w4(32'h398baa24),
	.w5(32'h3c069592),
	.w6(32'hbaf395f5),
	.w7(32'hb86745ef),
	.w8(32'h3c446f10),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc436f4),
	.w1(32'h3c280ad7),
	.w2(32'h3ce9a1b3),
	.w3(32'h3b90304e),
	.w4(32'hbbb58804),
	.w5(32'h3b819e0f),
	.w6(32'h3c356f46),
	.w7(32'hbc7ef725),
	.w8(32'hbca77289),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbe578),
	.w1(32'h3c1da282),
	.w2(32'hba97f08a),
	.w3(32'h3c0c1398),
	.w4(32'hba4db94e),
	.w5(32'hbc6655bf),
	.w6(32'hbcac8395),
	.w7(32'hbc8c3e38),
	.w8(32'h3ba57c8b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f6da4),
	.w1(32'h3c00a7a7),
	.w2(32'h3c9c7837),
	.w3(32'hbb83f7fd),
	.w4(32'h3a7e21a6),
	.w5(32'h3bafb14b),
	.w6(32'h3c2196f8),
	.w7(32'h3c204197),
	.w8(32'h3be293ec),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c376db1),
	.w1(32'h3b5370ee),
	.w2(32'hb99a4b95),
	.w3(32'h3c39ae50),
	.w4(32'h3bb340b2),
	.w5(32'hbb4c41a8),
	.w6(32'h3add5dde),
	.w7(32'h3c4a98b0),
	.w8(32'hbc089043),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14adb9),
	.w1(32'hb97e81b8),
	.w2(32'h3add1c19),
	.w3(32'hba862f2f),
	.w4(32'hbb6de48b),
	.w5(32'h3b8e3094),
	.w6(32'hbac20de9),
	.w7(32'hba4580ad),
	.w8(32'h3c4558bc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff4668),
	.w1(32'h3a8bc086),
	.w2(32'h3c858f10),
	.w3(32'hbc640af8),
	.w4(32'h3b7d885b),
	.w5(32'h3cb1fa89),
	.w6(32'h3c34a101),
	.w7(32'h3c887da8),
	.w8(32'hbc652793),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cfd36),
	.w1(32'h3893a674),
	.w2(32'h3b3a4a57),
	.w3(32'h3cccfeb1),
	.w4(32'h3c3ac0dd),
	.w5(32'h3c218fb9),
	.w6(32'h3a0ce30e),
	.w7(32'h3bc7bfc5),
	.w8(32'hbc795470),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a962fe2),
	.w1(32'h3bf4c663),
	.w2(32'h3c89ce1d),
	.w3(32'h3be13689),
	.w4(32'hbb9b70cc),
	.w5(32'h3c96a270),
	.w6(32'hbc5ce5bf),
	.w7(32'hbc848df9),
	.w8(32'hbc04b715),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9472cf),
	.w1(32'hb69ef31d),
	.w2(32'h3b523fdf),
	.w3(32'h3cf8ea4f),
	.w4(32'h3b9880a2),
	.w5(32'hbbdec9c2),
	.w6(32'h3c1eba8f),
	.w7(32'h3bc62ce7),
	.w8(32'h3a9e7ca6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b450f53),
	.w1(32'h3c1b9b6b),
	.w2(32'hbb1ffefc),
	.w3(32'hbb32084c),
	.w4(32'hbbc87a20),
	.w5(32'hbb5c3025),
	.w6(32'hbc1a02b1),
	.w7(32'hba4fcde7),
	.w8(32'hb898206c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d83bb),
	.w1(32'h3a561ab7),
	.w2(32'h3b9155aa),
	.w3(32'h3b8eb8ac),
	.w4(32'h3bf8b697),
	.w5(32'h3c135b7b),
	.w6(32'hb8a67646),
	.w7(32'h3c3a504d),
	.w8(32'h3c0ec214),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12823e),
	.w1(32'h3c631cb1),
	.w2(32'h3b6542a3),
	.w3(32'h3cf2d3a3),
	.w4(32'h3cdae343),
	.w5(32'hbb684594),
	.w6(32'h3cf16147),
	.w7(32'h3d04d4ab),
	.w8(32'hbb6d294b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b5019),
	.w1(32'h3c9ba7cd),
	.w2(32'h3c09b946),
	.w3(32'h3b90ceb5),
	.w4(32'h3bd42eb5),
	.w5(32'h3a882cb8),
	.w6(32'h3adb7c7c),
	.w7(32'hbbc5333a),
	.w8(32'h3b1cc124),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7295d5),
	.w1(32'h3baad26f),
	.w2(32'hbb7f1fc3),
	.w3(32'h3b6a35af),
	.w4(32'hbc22c412),
	.w5(32'hbc3873cc),
	.w6(32'h3a58fcdc),
	.w7(32'hbbcba896),
	.w8(32'h3b665198),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1621d6),
	.w1(32'h3bae527f),
	.w2(32'h3b5c384f),
	.w3(32'h3b908513),
	.w4(32'h3a8a9763),
	.w5(32'hbc4ab94d),
	.w6(32'h3bf6802b),
	.w7(32'h3c1f3808),
	.w8(32'hbc028f0f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8571d3),
	.w1(32'h3c350963),
	.w2(32'h3c92dd8f),
	.w3(32'hbb51a88f),
	.w4(32'hbc525f73),
	.w5(32'hba9917a3),
	.w6(32'h3b14090a),
	.w7(32'hbc15e267),
	.w8(32'hbb348fbc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3211a3),
	.w1(32'h3bb44416),
	.w2(32'h3bbac7cf),
	.w3(32'hbc8afda0),
	.w4(32'hbbc37529),
	.w5(32'hbba06a06),
	.w6(32'hbbb7498f),
	.w7(32'h3ac1956f),
	.w8(32'hbb90c945),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec65d5),
	.w1(32'hbaf333c1),
	.w2(32'h3ca40d44),
	.w3(32'hbbbb7912),
	.w4(32'hb9883a92),
	.w5(32'hb9cd6d75),
	.w6(32'hbbb47a22),
	.w7(32'h3a99669e),
	.w8(32'hbbb4156a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab3cd6),
	.w1(32'h3c660c17),
	.w2(32'hbbd91dac),
	.w3(32'h3a7955e9),
	.w4(32'hb93e3ff4),
	.w5(32'hbc24ed1a),
	.w6(32'hbc3c4f16),
	.w7(32'hbbf8ca1d),
	.w8(32'hbacd9527),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fafa6),
	.w1(32'hbb644042),
	.w2(32'hbb308621),
	.w3(32'hbbd2f4aa),
	.w4(32'hbc3e7b4c),
	.w5(32'hbc70d521),
	.w6(32'h3b64829d),
	.w7(32'h3aefcfb8),
	.w8(32'hbb85ba28),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14745d),
	.w1(32'h3c259cd1),
	.w2(32'h3b800b69),
	.w3(32'hbc285915),
	.w4(32'h3bae53f9),
	.w5(32'h3ae136e4),
	.w6(32'hbc90e440),
	.w7(32'h3b397fc5),
	.w8(32'hbb5d0f4c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bd0dd),
	.w1(32'hbab04544),
	.w2(32'h3c135e41),
	.w3(32'hbb758729),
	.w4(32'hbbb70515),
	.w5(32'h3bd0cbc8),
	.w6(32'hbb4b839c),
	.w7(32'hbbf44cfa),
	.w8(32'h3b5f9e1d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4192e9),
	.w1(32'h3c15a8ce),
	.w2(32'hbb0380cc),
	.w3(32'h3bb462c7),
	.w4(32'h3a97bae2),
	.w5(32'h3c9a3fd3),
	.w6(32'hb8b2db55),
	.w7(32'h3a8c88c7),
	.w8(32'h3d0f603b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bc398),
	.w1(32'hbcd42cae),
	.w2(32'h3c4b287a),
	.w3(32'h3c417100),
	.w4(32'h3a256730),
	.w5(32'h3832215b),
	.w6(32'h3d3f8edf),
	.w7(32'h3c9b00ff),
	.w8(32'hbc80d6ef),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46926c),
	.w1(32'h3b751446),
	.w2(32'hbafbb2ef),
	.w3(32'h3c447c88),
	.w4(32'h3b6df6cd),
	.w5(32'hb88da572),
	.w6(32'hbc406eaf),
	.w7(32'hbc1f77e9),
	.w8(32'hb94a9111),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2f1df),
	.w1(32'hb8db6275),
	.w2(32'h3c247dfc),
	.w3(32'h3af6d990),
	.w4(32'hbaf7436b),
	.w5(32'h3c14605e),
	.w6(32'h3b2c0382),
	.w7(32'hbb1bf035),
	.w8(32'h3c6990bf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7e67e),
	.w1(32'hbb38da3d),
	.w2(32'hba504fa3),
	.w3(32'hbabf3c1a),
	.w4(32'hbbc654a8),
	.w5(32'h3a9a44b4),
	.w6(32'h3bb2dea6),
	.w7(32'hbb4e8f0a),
	.w8(32'h3b8e3c93),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012117),
	.w1(32'h3a409a5d),
	.w2(32'hbca906ff),
	.w3(32'hbba4fa12),
	.w4(32'hb8e92c30),
	.w5(32'hbc0116af),
	.w6(32'hbba51b7f),
	.w7(32'hba0213d8),
	.w8(32'h3c8f0978),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d2723),
	.w1(32'hbc5ce805),
	.w2(32'h3c94bbea),
	.w3(32'hbc7f7548),
	.w4(32'hb94ef800),
	.w5(32'h3b5aa27c),
	.w6(32'h3cee0ef3),
	.w7(32'h3cfd3b30),
	.w8(32'hbc9e5032),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d055160),
	.w1(32'h3ceb5277),
	.w2(32'hba851608),
	.w3(32'hba4b17ab),
	.w4(32'h3c867264),
	.w5(32'hbbb8662b),
	.w6(32'hbd164ae6),
	.w7(32'hbcbf25ad),
	.w8(32'hbbe5ae4e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8c712),
	.w1(32'hba97da0e),
	.w2(32'h3a6c1b32),
	.w3(32'h3bc3ae65),
	.w4(32'h3b004cc3),
	.w5(32'hbc2984ab),
	.w6(32'h3c270411),
	.w7(32'h3b366cb0),
	.w8(32'hbbcbac25),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a559c),
	.w1(32'h3b1de347),
	.w2(32'h3c016f41),
	.w3(32'h39cef782),
	.w4(32'hbb19a1c5),
	.w5(32'hbc7666eb),
	.w6(32'h3b61729a),
	.w7(32'h3a1f1df9),
	.w8(32'hbce33454),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccda239),
	.w1(32'h3c9349a6),
	.w2(32'hb8ed72fc),
	.w3(32'h3c481a53),
	.w4(32'h3c86b05c),
	.w5(32'hbc503417),
	.w6(32'hbcabf675),
	.w7(32'hbbfd9648),
	.w8(32'hbc987842),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca34264),
	.w1(32'h3c6651a7),
	.w2(32'h3bb3c02f),
	.w3(32'hb9da3763),
	.w4(32'h3c5edf60),
	.w5(32'hbbd2458e),
	.w6(32'hbcc4ce38),
	.w7(32'hbb9ee516),
	.w8(32'h3b9e92ae),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0927ff),
	.w1(32'hbaf3eccb),
	.w2(32'hba78cf5d),
	.w3(32'h3b139fd0),
	.w4(32'hbafffe5f),
	.w5(32'hbb46bd34),
	.w6(32'h3c5b975b),
	.w7(32'h3bdb55bd),
	.w8(32'h388493b9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a40c),
	.w1(32'h3adba398),
	.w2(32'h3b9c9ad0),
	.w3(32'h3bd70519),
	.w4(32'h38c5cbef),
	.w5(32'h3b858bea),
	.w6(32'h3b824ec2),
	.w7(32'hbaf881d8),
	.w8(32'h3b0c13dc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c0965),
	.w1(32'h3a7fe3ba),
	.w2(32'h3b433af2),
	.w3(32'h3bc303c8),
	.w4(32'hba9dd208),
	.w5(32'hbb84e312),
	.w6(32'h3a1b145e),
	.w7(32'hb9c6fd95),
	.w8(32'h3b766087),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaccd0),
	.w1(32'hbab6cf88),
	.w2(32'h3c072f39),
	.w3(32'hbb9511ef),
	.w4(32'hbba4d670),
	.w5(32'h3a0b7a50),
	.w6(32'hba838697),
	.w7(32'hba9ffc0d),
	.w8(32'hbb76ca8e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcacb08c),
	.w1(32'hbcdf9d0f),
	.w2(32'hbc18f7a5),
	.w3(32'h3adc7487),
	.w4(32'hbac24f10),
	.w5(32'hbc3aed43),
	.w6(32'h3cf296dd),
	.w7(32'h3cda0091),
	.w8(32'hbb9ec538),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b31be),
	.w1(32'hbb7903e1),
	.w2(32'h3a1e98ba),
	.w3(32'h3b3fd88f),
	.w4(32'h3b432d89),
	.w5(32'hbc329a37),
	.w6(32'h3ac0f876),
	.w7(32'h3bfcb2c6),
	.w8(32'hbad46dec),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fe289),
	.w1(32'h3c7863ed),
	.w2(32'h3b2d9f26),
	.w3(32'hbbd08808),
	.w4(32'h3aa466be),
	.w5(32'h3c8a0197),
	.w6(32'h3c6b5d72),
	.w7(32'h3bdd707f),
	.w8(32'h3c72fe5d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cbfef),
	.w1(32'hbb998ae6),
	.w2(32'h3bd30f16),
	.w3(32'h3c6b0f06),
	.w4(32'hbc1502c9),
	.w5(32'h3b9360db),
	.w6(32'h3ccc13dd),
	.w7(32'hbbea522a),
	.w8(32'h3a8588e6),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bc07e),
	.w1(32'hba3271d4),
	.w2(32'h3b2a810b),
	.w3(32'hbb9e2d38),
	.w4(32'hbbdb1f44),
	.w5(32'h3a143a98),
	.w6(32'hbab126f4),
	.w7(32'h392c4cf4),
	.w8(32'h3b451a8c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca528e),
	.w1(32'hbb88388f),
	.w2(32'h3c76b39d),
	.w3(32'hba29be0c),
	.w4(32'hbb8948b0),
	.w5(32'h3cb704bd),
	.w6(32'hbb928ef8),
	.w7(32'hbb5890ad),
	.w8(32'hb99fbb3b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c866942),
	.w1(32'hbbbc2c86),
	.w2(32'hbc0426d5),
	.w3(32'h3d036382),
	.w4(32'h3c2f34a7),
	.w5(32'hbbae9eb0),
	.w6(32'h3c028d34),
	.w7(32'h3b7d6a11),
	.w8(32'h3c34d9f6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76c8be),
	.w1(32'hbcc1325e),
	.w2(32'h3c0a8ae4),
	.w3(32'h3bbb0251),
	.w4(32'hbc23e46f),
	.w5(32'h3ad2e743),
	.w6(32'h3c8d6f62),
	.w7(32'h3ba0aa6a),
	.w8(32'hbbcdedcc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d6732),
	.w1(32'h3bb8acda),
	.w2(32'h3cbdcdc8),
	.w3(32'h3bd3577f),
	.w4(32'hba0843d4),
	.w5(32'h3b84feb7),
	.w6(32'hb9bc094c),
	.w7(32'hbb9dc54a),
	.w8(32'h3b691e01),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd54661),
	.w1(32'h3c9a9fe6),
	.w2(32'hbb70f11b),
	.w3(32'h3ab22a23),
	.w4(32'hbb601a51),
	.w5(32'hbac4ddcd),
	.w6(32'hbb3b43ca),
	.w7(32'hbb507770),
	.w8(32'h3abc9592),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fef9),
	.w1(32'hbc07346d),
	.w2(32'hbb94d919),
	.w3(32'hb98621c0),
	.w4(32'hbb112d44),
	.w5(32'hbbf0bc30),
	.w6(32'hbb8736ce),
	.w7(32'hbb89f67b),
	.w8(32'hbc340590),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc116),
	.w1(32'h3bcbcc5f),
	.w2(32'h3b8b84cf),
	.w3(32'h3b18852a),
	.w4(32'h3b2e653c),
	.w5(32'hbbbf67d6),
	.w6(32'hb9b6f47b),
	.w7(32'hb96f1d76),
	.w8(32'hbc83d6e2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95cad2),
	.w1(32'h3c2ba881),
	.w2(32'h3b7ab4bf),
	.w3(32'h3c622141),
	.w4(32'h3c476c03),
	.w5(32'hbb18495e),
	.w6(32'hbc786872),
	.w7(32'hb7b75536),
	.w8(32'h3b4af03b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d368),
	.w1(32'hba3d3d05),
	.w2(32'hbb8ac702),
	.w3(32'hbcdd9168),
	.w4(32'hbc4b9c5b),
	.w5(32'hbc211c68),
	.w6(32'hbb62f876),
	.w7(32'hbb8ff0bb),
	.w8(32'h38037ab6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb243f5),
	.w1(32'h39f42869),
	.w2(32'h3cf3f697),
	.w3(32'h3a973e98),
	.w4(32'h3bbabb64),
	.w5(32'hbb0b2e19),
	.w6(32'h3a8b9264),
	.w7(32'hba16f3cb),
	.w8(32'hbc6c06ff),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b39b2),
	.w1(32'h3aea126a),
	.w2(32'h3c15d9b0),
	.w3(32'hbc01d430),
	.w4(32'hba808b36),
	.w5(32'h3a7f1753),
	.w6(32'hbcb1322e),
	.w7(32'hbbac0934),
	.w8(32'hbc452784),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5101e3),
	.w1(32'h3b6c7978),
	.w2(32'h3c19fa9b),
	.w3(32'h3bfbec09),
	.w4(32'h3bef35cf),
	.w5(32'h3b3c875d),
	.w6(32'hbc21abbf),
	.w7(32'h3b7e865a),
	.w8(32'hba37e1d2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fca8e),
	.w1(32'h3c0f9b04),
	.w2(32'hbb56b535),
	.w3(32'h3c0cc01a),
	.w4(32'h3a9af40c),
	.w5(32'h3b3b0d07),
	.w6(32'h3b7bc4ca),
	.w7(32'hbaab0178),
	.w8(32'h3c800a95),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa74f04),
	.w1(32'h3acefe48),
	.w2(32'hbbd5077f),
	.w3(32'hbb0dfb3d),
	.w4(32'hbc0d13e2),
	.w5(32'hbc63ca23),
	.w6(32'hbae96f6e),
	.w7(32'hbbc911e6),
	.w8(32'h3c0202e0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9db834),
	.w1(32'h3a7a30af),
	.w2(32'hbc3499ae),
	.w3(32'hbc68c024),
	.w4(32'h3ad1d26e),
	.w5(32'hb996bb7f),
	.w6(32'hbbc9ef49),
	.w7(32'h3acb08e9),
	.w8(32'h3b4e7dad),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fdc26),
	.w1(32'hbb88fc03),
	.w2(32'hbb407c90),
	.w3(32'h3ae9c0b5),
	.w4(32'hbbbf243c),
	.w5(32'hba2bd3c0),
	.w6(32'h3c09b883),
	.w7(32'h3ba22740),
	.w8(32'h3b3e0de4),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9598e),
	.w1(32'h3a8d59af),
	.w2(32'hba6591ee),
	.w3(32'hbbb88331),
	.w4(32'hbc0afaa3),
	.w5(32'h3b98c7e8),
	.w6(32'hbc289912),
	.w7(32'hbbc47887),
	.w8(32'h3c27eaaa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3da4a5),
	.w1(32'hbb81b2b3),
	.w2(32'h390f3ffd),
	.w3(32'h3bc76f0d),
	.w4(32'hbb2827b3),
	.w5(32'h3bad0f78),
	.w6(32'h3c059640),
	.w7(32'h3ac72e46),
	.w8(32'h3b1a44cf),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27d487),
	.w1(32'hbb63a87e),
	.w2(32'h3bd499b0),
	.w3(32'hbac38828),
	.w4(32'hbc1d67a7),
	.w5(32'h3c697659),
	.w6(32'hbb8c0b72),
	.w7(32'hba449265),
	.w8(32'h3c6f8062),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90257c6),
	.w1(32'h39037541),
	.w2(32'hb9a42881),
	.w3(32'h3c00b487),
	.w4(32'hbb5d6670),
	.w5(32'hbb991247),
	.w6(32'h3b657266),
	.w7(32'hbaef5a66),
	.w8(32'hbb090d51),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70425d),
	.w1(32'h3b1a8dca),
	.w2(32'h3a932858),
	.w3(32'h3a6c5190),
	.w4(32'h3bb38cba),
	.w5(32'hbc2e9018),
	.w6(32'h3aa4d666),
	.w7(32'h3b71553b),
	.w8(32'h3baf6eb5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d5dbe),
	.w1(32'h3c15869c),
	.w2(32'hbc0eead3),
	.w3(32'hbba3552c),
	.w4(32'h3beffa64),
	.w5(32'hbb4111fa),
	.w6(32'h3c6f1a2d),
	.w7(32'hbb0f24af),
	.w8(32'h3b139cb5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc85c6),
	.w1(32'hb7b2fe3b),
	.w2(32'h3c8c7e8a),
	.w3(32'h3c35eaab),
	.w4(32'h3c02f64d),
	.w5(32'h3ada7866),
	.w6(32'hbbdc0bd4),
	.w7(32'hbb1e1245),
	.w8(32'hbc25ea4c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95f9c3),
	.w1(32'h3b4525b3),
	.w2(32'hbbfa55fd),
	.w3(32'hbbe117d2),
	.w4(32'hbb34ca47),
	.w5(32'hbb3e83d4),
	.w6(32'hbc633d10),
	.w7(32'hbc3082a2),
	.w8(32'hbae3a054),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5eadc),
	.w1(32'h3ac96d73),
	.w2(32'h3c8a9408),
	.w3(32'hbbc62b44),
	.w4(32'hbc6f7a00),
	.w5(32'h3c3cd47a),
	.w6(32'h3b8f4706),
	.w7(32'hb9fe9483),
	.w8(32'h3ba73776),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc096956),
	.w1(32'hbc4fc2c5),
	.w2(32'h3c8d18a9),
	.w3(32'hba4621e4),
	.w4(32'hbb8414e9),
	.w5(32'h3b79b877),
	.w6(32'h3c030b8a),
	.w7(32'h3c0abfd4),
	.w8(32'hbc0eb482),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfd6db),
	.w1(32'h3bc73827),
	.w2(32'h3c2f1933),
	.w3(32'hbbbf61b6),
	.w4(32'h3a260ab0),
	.w5(32'h3c32fffd),
	.w6(32'hbc49b94f),
	.w7(32'hbc418487),
	.w8(32'h3ba927bf),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b0bd2),
	.w1(32'h3c401274),
	.w2(32'hbaf3069a),
	.w3(32'h3c443f88),
	.w4(32'h3cb3efe2),
	.w5(32'hbaa3f314),
	.w6(32'h3be2afff),
	.w7(32'h3c38f639),
	.w8(32'h39bb9fcc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a6cec),
	.w1(32'h3b0ab37c),
	.w2(32'h3c8f5841),
	.w3(32'h3b296f4c),
	.w4(32'h3b823b8b),
	.w5(32'hb990823d),
	.w6(32'h394049fa),
	.w7(32'h3bad96a1),
	.w8(32'hbb80a5bd),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c512d96),
	.w1(32'h3c0ff74a),
	.w2(32'hbb3ef97a),
	.w3(32'h3bc0547d),
	.w4(32'h3b3879fa),
	.w5(32'hbb76326a),
	.w6(32'hbb9f8c48),
	.w7(32'hb8ae5ed2),
	.w8(32'h3ade2469),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59ecf5),
	.w1(32'h3c11662e),
	.w2(32'hbbd597f9),
	.w3(32'h3afc14ff),
	.w4(32'h3b6c0f47),
	.w5(32'hbc3b3af0),
	.w6(32'h39e299c4),
	.w7(32'h3bb1c3b9),
	.w8(32'hbc47e27f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d213c),
	.w1(32'h3b7ed130),
	.w2(32'h3aa28edf),
	.w3(32'h3b469112),
	.w4(32'h3c0c4d98),
	.w5(32'h3b9fc59f),
	.w6(32'hbbd9bf68),
	.w7(32'hbc223644),
	.w8(32'h3ca0eafa),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf62160),
	.w1(32'hbb024520),
	.w2(32'h3c5cb2c5),
	.w3(32'h3b20372d),
	.w4(32'h3bd93dbb),
	.w5(32'h3c61dced),
	.w6(32'hbbec910e),
	.w7(32'h3b2d2374),
	.w8(32'hbbb288eb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbfb302),
	.w1(32'h3bf314a4),
	.w2(32'hba1b07fc),
	.w3(32'h3b36bcfb),
	.w4(32'h3b87bf9d),
	.w5(32'h3a22f9e5),
	.w6(32'hbc0cb52a),
	.w7(32'hbc0362ca),
	.w8(32'h3acab936),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ecd89),
	.w1(32'hbb8f3a5a),
	.w2(32'hba903c59),
	.w3(32'hba869b42),
	.w4(32'hbb8057d2),
	.w5(32'hbb25c41e),
	.w6(32'hb98e1524),
	.w7(32'h3a99ecc0),
	.w8(32'h3b09a6cf),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1d5d6),
	.w1(32'hbbcac2c8),
	.w2(32'h3bb79923),
	.w3(32'hbb63a43e),
	.w4(32'hbb20bb3f),
	.w5(32'h3a106b4b),
	.w6(32'h3b2b921f),
	.w7(32'h3b93bf4b),
	.w8(32'hbbdf89c2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0614b6),
	.w1(32'h3977a8b8),
	.w2(32'h3b13937d),
	.w3(32'h3c887d0d),
	.w4(32'h3b8e808f),
	.w5(32'hb8ee631d),
	.w6(32'hbba96200),
	.w7(32'h3ba897a5),
	.w8(32'hba3a53bd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad17fc0),
	.w1(32'h3af8c8a4),
	.w2(32'h3b07036d),
	.w3(32'hbb0bf31f),
	.w4(32'hbb105ac8),
	.w5(32'h3b81d13e),
	.w6(32'hbb1cf91a),
	.w7(32'hba24381c),
	.w8(32'hbb73a8ed),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef96bb),
	.w1(32'h3ae98539),
	.w2(32'h3b6b168a),
	.w3(32'h3bd3f2db),
	.w4(32'hbbd2c0bf),
	.w5(32'h3bebc14a),
	.w6(32'h3be2b393),
	.w7(32'h3b6c89c7),
	.w8(32'h3cf8ff94),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd12660a),
	.w1(32'hbcb35eb7),
	.w2(32'hbcda7cb1),
	.w3(32'h3ba3c4b4),
	.w4(32'hbbacb5c9),
	.w5(32'h3b2438f4),
	.w6(32'h3d182a60),
	.w7(32'h3cc08c94),
	.w8(32'h3d1e3294),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4f0edf),
	.w1(32'hbcc1868e),
	.w2(32'h3b3c9809),
	.w3(32'hba355d0f),
	.w4(32'hbc430eb3),
	.w5(32'h3ac3ff3c),
	.w6(32'h3d46267e),
	.w7(32'h3cc0fad1),
	.w8(32'hba7cd500),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule