module layer_10_featuremap_19(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990ed9),
	.w1(32'h3a8554e1),
	.w2(32'hbb5eccf9),
	.w3(32'hbc03abce),
	.w4(32'hbb25aa5a),
	.w5(32'hbbfd9ea7),
	.w6(32'hbbf153ae),
	.w7(32'hbb561d96),
	.w8(32'hbc14ec6e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8329dae),
	.w1(32'hbbafdf57),
	.w2(32'hb9872e3c),
	.w3(32'hbaf78166),
	.w4(32'h39e867e2),
	.w5(32'hbb98d764),
	.w6(32'hbb4fa48c),
	.w7(32'hbc080d20),
	.w8(32'hbb84ca9a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae025),
	.w1(32'h3bdcd739),
	.w2(32'hbbf4510d),
	.w3(32'h3b4a6069),
	.w4(32'h3b342f8a),
	.w5(32'hbbb0d882),
	.w6(32'hbc06b2db),
	.w7(32'hbb9e4a92),
	.w8(32'h3bc3f03c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc264c82),
	.w1(32'hbc62a58b),
	.w2(32'hbc228cda),
	.w3(32'hbc2dd799),
	.w4(32'hbc280f32),
	.w5(32'hba2e224f),
	.w6(32'hba5d38c3),
	.w7(32'hbab0c4c8),
	.w8(32'hbba77eac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac27450),
	.w1(32'hbbe4bed5),
	.w2(32'hbc4dfc4b),
	.w3(32'hbb9ca566),
	.w4(32'hbbccff8e),
	.w5(32'hbbf5e85d),
	.w6(32'h3b85d76b),
	.w7(32'h3c115e26),
	.w8(32'hbb1c6529),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1de08),
	.w1(32'hbac33276),
	.w2(32'h3d87b9ae),
	.w3(32'hbc14d466),
	.w4(32'hba8dbf57),
	.w5(32'h3d15738a),
	.w6(32'hbbe3fbdc),
	.w7(32'hbbb36174),
	.w8(32'hbcb95fd2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db65054),
	.w1(32'h3d89812b),
	.w2(32'hbc36d4a6),
	.w3(32'hbc7f65b0),
	.w4(32'h3b6c0e5b),
	.w5(32'hbc9877e3),
	.w6(32'hbe03e3e6),
	.w7(32'hbd8c95c6),
	.w8(32'h3b5cf60c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94d723),
	.w1(32'hbc4c5354),
	.w2(32'h3b280d45),
	.w3(32'hbd185373),
	.w4(32'hbc9ba0fb),
	.w5(32'h3c7a95d3),
	.w6(32'hbb0a7ed0),
	.w7(32'h3c386a95),
	.w8(32'h3be1ec92),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b185fec),
	.w1(32'hbb61dd92),
	.w2(32'hba95c5cf),
	.w3(32'h3a82eed5),
	.w4(32'hbbaabfa7),
	.w5(32'hba42f3cf),
	.w6(32'h3b4af44f),
	.w7(32'h3acc7c60),
	.w8(32'hb9dd7994),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b7646),
	.w1(32'hbbb89651),
	.w2(32'hbc93fb76),
	.w3(32'h3b87f95c),
	.w4(32'hbb7440af),
	.w5(32'hba19c83b),
	.w6(32'h3c4f6fce),
	.w7(32'hbb176813),
	.w8(32'h3c6e635d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd379a2d),
	.w1(32'hbd27a184),
	.w2(32'hbb831690),
	.w3(32'h3c4cccfd),
	.w4(32'hbc198f07),
	.w5(32'hbbb79568),
	.w6(32'h3d87ea69),
	.w7(32'h3ca9abbf),
	.w8(32'hbaac6100),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d4a2),
	.w1(32'hba2d095d),
	.w2(32'h3cf5a743),
	.w3(32'hbc54e94d),
	.w4(32'hbc1b1df5),
	.w5(32'h3bfeefa0),
	.w6(32'hbc26e1d3),
	.w7(32'hbc24896c),
	.w8(32'hbaf3adfe),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2be92f),
	.w1(32'h3d25df03),
	.w2(32'h39eacdb8),
	.w3(32'hba1a1fac),
	.w4(32'h3c41f3d1),
	.w5(32'hb8b4107a),
	.w6(32'hbd01941f),
	.w7(32'hbc71aa39),
	.w8(32'hba8e8b26),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9256b),
	.w1(32'hbb10e1d9),
	.w2(32'hbb516393),
	.w3(32'hbbd8cffe),
	.w4(32'hbb381947),
	.w5(32'h3b1731c1),
	.w6(32'hbbc62de8),
	.w7(32'hb9775178),
	.w8(32'hbacf3c59),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a9a51),
	.w1(32'h3aa01946),
	.w2(32'hbaab9300),
	.w3(32'hbad0c006),
	.w4(32'h3bc29562),
	.w5(32'hbbd2c31d),
	.w6(32'hbb8384f2),
	.w7(32'hbae14c92),
	.w8(32'hba83ed71),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cfa31),
	.w1(32'h3b0112fa),
	.w2(32'h3bee3339),
	.w3(32'hbc8a8443),
	.w4(32'hbc2da072),
	.w5(32'h3c0e8d83),
	.w6(32'hbc2893bc),
	.w7(32'hbb9a7f15),
	.w8(32'h3c27a0d5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc854f27),
	.w1(32'hbca985c7),
	.w2(32'hbaf5918e),
	.w3(32'h3bc13c18),
	.w4(32'hbc5a91af),
	.w5(32'h3addd78d),
	.w6(32'h3cfa168a),
	.w7(32'h393d8c28),
	.w8(32'h3ba81b6c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa50d83),
	.w1(32'h3a2a42a3),
	.w2(32'h3b094112),
	.w3(32'hbc0b05ea),
	.w4(32'hbb8cae35),
	.w5(32'h3b1235e7),
	.w6(32'h3bd1fe1d),
	.w7(32'h3c0f9ad9),
	.w8(32'hba95df92),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff282),
	.w1(32'hb92f5ef3),
	.w2(32'h3c624313),
	.w3(32'hbb1b5e83),
	.w4(32'hbb08ef24),
	.w5(32'h3c1ff15e),
	.w6(32'hbc174eb6),
	.w7(32'hbb6ae9d0),
	.w8(32'h3bfbfff4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468967),
	.w1(32'h3c16e74d),
	.w2(32'hbc17929e),
	.w3(32'h3c4d1078),
	.w4(32'h3c1e6f46),
	.w5(32'hbbf66b7c),
	.w6(32'hbb846f24),
	.w7(32'h3b971d71),
	.w8(32'hba39addd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ce95),
	.w1(32'hbb4b3189),
	.w2(32'hbac1263f),
	.w3(32'hbb8a27a1),
	.w4(32'hb9f9e41b),
	.w5(32'hbb851f3b),
	.w6(32'h3b586bbc),
	.w7(32'h39133928),
	.w8(32'h3b277cb7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba456fd3),
	.w1(32'hbbb5f95e),
	.w2(32'h3c4087c7),
	.w3(32'h3b26f0e8),
	.w4(32'hbabb7f9f),
	.w5(32'h3bf0eb1b),
	.w6(32'h3b8095df),
	.w7(32'hb647d613),
	.w8(32'hba4ebef5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17b5bb),
	.w1(32'h3cb97b49),
	.w2(32'hbc93195a),
	.w3(32'hbbf32f3f),
	.w4(32'h3b1f1f12),
	.w5(32'hbc71b249),
	.w6(32'hbcb5dd4a),
	.w7(32'hbbff3313),
	.w8(32'h3c0a6f2f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3382c4),
	.w1(32'hbcea26d5),
	.w2(32'h3a8da368),
	.w3(32'h3c16453a),
	.w4(32'hbc0b7353),
	.w5(32'h392eb3cf),
	.w6(32'h3d809bc8),
	.w7(32'h3c917012),
	.w8(32'hbb64a18d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71f738),
	.w1(32'hbb3ea8b5),
	.w2(32'hba656150),
	.w3(32'hbab38851),
	.w4(32'hbb67c250),
	.w5(32'h3ba8221b),
	.w6(32'hbba9dfe5),
	.w7(32'hbbd565d0),
	.w8(32'h3c5252dc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e2d3b8),
	.w1(32'h3a70798c),
	.w2(32'h3b3f4ab1),
	.w3(32'h3bef116c),
	.w4(32'h3b7990fd),
	.w5(32'hbb9e27b1),
	.w6(32'h3c3bc62b),
	.w7(32'h3b83f104),
	.w8(32'hbbc5ab14),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacde148),
	.w1(32'hbbefa96a),
	.w2(32'hb9b32989),
	.w3(32'hbb7c1b82),
	.w4(32'hbb9b5e79),
	.w5(32'h3ba7619e),
	.w6(32'h38550bcf),
	.w7(32'h3b3cc8c2),
	.w8(32'h3a87e265),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb29b1a),
	.w1(32'h3b221e66),
	.w2(32'hbc561285),
	.w3(32'h3cc83aa9),
	.w4(32'h3c1f5e1f),
	.w5(32'hbc376738),
	.w6(32'h3c5c0697),
	.w7(32'h3b61cb93),
	.w8(32'hbbbba9b2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2876cf),
	.w1(32'hbb9f806a),
	.w2(32'h3b2e02f4),
	.w3(32'hbc1a9fb2),
	.w4(32'h3b03c209),
	.w5(32'hbaf8a813),
	.w6(32'hbb3712ae),
	.w7(32'h3aeffe00),
	.w8(32'h3b923454),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f5f2),
	.w1(32'h3b7d7d28),
	.w2(32'hbc165cfe),
	.w3(32'h396c0872),
	.w4(32'hbb6cb177),
	.w5(32'h3bae3f31),
	.w6(32'h3bd11732),
	.w7(32'hbb2cc443),
	.w8(32'hbbd29243),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939eea),
	.w1(32'hbb637fb0),
	.w2(32'hb9c5f545),
	.w3(32'h3ce2933c),
	.w4(32'h3c89305f),
	.w5(32'h3a54fc7f),
	.w6(32'h3c50bdd5),
	.w7(32'h3b316290),
	.w8(32'hbb29e3ff),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33cb90),
	.w1(32'h3754f806),
	.w2(32'hbb657905),
	.w3(32'h3ae564a3),
	.w4(32'h3b86334b),
	.w5(32'hbae81a5f),
	.w6(32'hbad117dd),
	.w7(32'hb861b22d),
	.w8(32'hba616dae),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab17d5c),
	.w1(32'hb9aa87ed),
	.w2(32'hbb3dc8a1),
	.w3(32'hbb331a7a),
	.w4(32'hba307ab4),
	.w5(32'h3c228f76),
	.w6(32'hbb45238c),
	.w7(32'hbb197d63),
	.w8(32'hbb96c3cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c191997),
	.w1(32'hba415af9),
	.w2(32'h3b1c2e9a),
	.w3(32'h3cbb12d1),
	.w4(32'h3c42c5da),
	.w5(32'h3b028077),
	.w6(32'h3c08e757),
	.w7(32'hba907b91),
	.w8(32'h3b3acdf5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927ed5f),
	.w1(32'h39563093),
	.w2(32'hbb62d0c9),
	.w3(32'h3b38898f),
	.w4(32'h3ad9afa2),
	.w5(32'hbc409543),
	.w6(32'h3b1502e5),
	.w7(32'h3be5597c),
	.w8(32'hbbbf9637),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76ecdf),
	.w1(32'hbc0dca89),
	.w2(32'hbb9fd469),
	.w3(32'hbd067b69),
	.w4(32'hbcb6a5a0),
	.w5(32'hbbf73cc6),
	.w6(32'hbccdc21a),
	.w7(32'hbc7deeb6),
	.w8(32'hbb108cfa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbde3af),
	.w1(32'h3af75f98),
	.w2(32'hbb977182),
	.w3(32'hbc1cf7a1),
	.w4(32'h3b02702b),
	.w5(32'h3a74262a),
	.w6(32'hbbb498cd),
	.w7(32'hbad8b3ae),
	.w8(32'hbc464594),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3909),
	.w1(32'hbc9cea75),
	.w2(32'hbb5c3c0f),
	.w3(32'h3c143d9b),
	.w4(32'hbbc87e1b),
	.w5(32'hbbc8cb29),
	.w6(32'hbad63d4b),
	.w7(32'hbc8dcd0d),
	.w8(32'hbbc8b3dc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8878006),
	.w1(32'hbb9b904b),
	.w2(32'hbbfb98fa),
	.w3(32'h3b59f497),
	.w4(32'hba5bb557),
	.w5(32'h3b0f554d),
	.w6(32'h392f80d2),
	.w7(32'hbb99edca),
	.w8(32'hba89bc15),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa612d9),
	.w1(32'hbba2edb4),
	.w2(32'h3bd788e3),
	.w3(32'h3c2159fb),
	.w4(32'h39afecfc),
	.w5(32'h3b3a5e32),
	.w6(32'h3c0e9c4e),
	.w7(32'hbb45d305),
	.w8(32'h3b1ecfc6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b016bb0),
	.w1(32'h3b425426),
	.w2(32'hbb106666),
	.w3(32'hbb02841d),
	.w4(32'h3b2bfc68),
	.w5(32'hb97dc2d8),
	.w6(32'h3a32efc2),
	.w7(32'h3afb78ab),
	.w8(32'hbac9d280),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38edfb3a),
	.w1(32'hbb21fefb),
	.w2(32'h3b67db12),
	.w3(32'h3ba31c7e),
	.w4(32'h3ac9b4d1),
	.w5(32'hbae581f4),
	.w6(32'h3ac1c179),
	.w7(32'h3b2d3aed),
	.w8(32'hbb0fd89c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059424),
	.w1(32'h3adaf01f),
	.w2(32'h3b94b531),
	.w3(32'hb9174fee),
	.w4(32'hbb72985c),
	.w5(32'h3b2412e4),
	.w6(32'hb9353138),
	.w7(32'hbb07160b),
	.w8(32'h3c1b8f86),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8579d1),
	.w1(32'h3c4410a2),
	.w2(32'h3b821a4b),
	.w3(32'h3b024029),
	.w4(32'h3c24a2a3),
	.w5(32'h3c02f17a),
	.w6(32'h3c07b6a1),
	.w7(32'h3c8968f5),
	.w8(32'h3bc88945),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99cb22),
	.w1(32'h3ad92a12),
	.w2(32'h3b93883f),
	.w3(32'h3bdf98e7),
	.w4(32'h3bea9872),
	.w5(32'h3b88beec),
	.w6(32'h3b8aaaee),
	.w7(32'h3b90c58e),
	.w8(32'h3b84474e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b552),
	.w1(32'hb9f42bda),
	.w2(32'h3a0ab6e8),
	.w3(32'h3a18a32a),
	.w4(32'h3b2aeed7),
	.w5(32'h3b9355c4),
	.w6(32'h3b1500cd),
	.w7(32'h3989108f),
	.w8(32'h3b74d34e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4057d7),
	.w1(32'h3a8285ec),
	.w2(32'h3b582847),
	.w3(32'h3b7b417e),
	.w4(32'h3b9cbf17),
	.w5(32'hba0fc6f1),
	.w6(32'h3b173670),
	.w7(32'h3ae3a2fa),
	.w8(32'hb9a20aad),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e4c6a),
	.w1(32'h3bbe2bfb),
	.w2(32'h3c63878e),
	.w3(32'hbaaa7cab),
	.w4(32'h3b5483eb),
	.w5(32'hbb87d0d3),
	.w6(32'hbb82f714),
	.w7(32'h3bcf1b94),
	.w8(32'h3c5081c3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa38ed),
	.w1(32'h3ae408a7),
	.w2(32'h3bb1ab55),
	.w3(32'hbd04e49b),
	.w4(32'hbca85463),
	.w5(32'h3b92a691),
	.w6(32'hbc79f563),
	.w7(32'hbb8c9eea),
	.w8(32'h3b4bb9cf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbe8f1),
	.w1(32'h3b442f3f),
	.w2(32'hba01c571),
	.w3(32'h3b5003dd),
	.w4(32'h3b33acff),
	.w5(32'h3994c1f5),
	.w6(32'h3b6e6d81),
	.w7(32'h3bcc9a9f),
	.w8(32'h3b076135),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39686474),
	.w1(32'hba854bb0),
	.w2(32'h3a8d31f7),
	.w3(32'hbb4201c1),
	.w4(32'h3ac45069),
	.w5(32'hbbe98faa),
	.w6(32'h3a868129),
	.w7(32'hba93d406),
	.w8(32'hbb5cf794),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd34e5),
	.w1(32'hbb22cb64),
	.w2(32'h3b2fedb8),
	.w3(32'hbb06cb14),
	.w4(32'hbb892e38),
	.w5(32'h3b3c2548),
	.w6(32'hbbc0d346),
	.w7(32'hbba704cd),
	.w8(32'h3b42c2ec),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b692d),
	.w1(32'h3a3a8b7c),
	.w2(32'h39f8809a),
	.w3(32'h3ae19e46),
	.w4(32'hbb85ef9c),
	.w5(32'h3b6e6f3c),
	.w6(32'h3a341e4b),
	.w7(32'hbae6a52a),
	.w8(32'h3ba1385b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6eeb4),
	.w1(32'hb9214f0c),
	.w2(32'h3b4904fb),
	.w3(32'hba31d933),
	.w4(32'h3a8ef7db),
	.w5(32'h3b0c551d),
	.w6(32'hba561b16),
	.w7(32'h3a3c9711),
	.w8(32'h3b617916),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37b0c8),
	.w1(32'h3a555f6b),
	.w2(32'hbb3bd900),
	.w3(32'hbb2c5a1e),
	.w4(32'hb83568c2),
	.w5(32'hbb4c0c0b),
	.w6(32'h3aa37520),
	.w7(32'hb95d3e07),
	.w8(32'h3b193e2d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c63f0),
	.w1(32'h3ae268d5),
	.w2(32'h3a8fcde0),
	.w3(32'h3b38fb1c),
	.w4(32'h3b15a6ce),
	.w5(32'h3ad9be2c),
	.w6(32'h3b0bb407),
	.w7(32'h3b61b405),
	.w8(32'h3bb377f5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6aee),
	.w1(32'h3af72f64),
	.w2(32'hbc2f29ad),
	.w3(32'h3b50176f),
	.w4(32'h3b933dd1),
	.w5(32'hbba9d7ee),
	.w6(32'h3a46d0a2),
	.w7(32'h3ba9c1c1),
	.w8(32'hbbd266a5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08decf),
	.w1(32'hbc463aa7),
	.w2(32'h3aad7e52),
	.w3(32'hbb155728),
	.w4(32'hbc1a4131),
	.w5(32'h3b4550dd),
	.w6(32'hbb29e49e),
	.w7(32'hbc0a511d),
	.w8(32'h3b767eb2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30979e),
	.w1(32'hbaf65039),
	.w2(32'hbc22d0c7),
	.w3(32'h3c3c49b2),
	.w4(32'h3be9c8dd),
	.w5(32'hbc0b854c),
	.w6(32'h3c645697),
	.w7(32'h3c405835),
	.w8(32'hbc1def22),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb76879),
	.w1(32'hbbd4af63),
	.w2(32'hbc49c876),
	.w3(32'hbbd51423),
	.w4(32'hbb946634),
	.w5(32'hbc01b9be),
	.w6(32'hbbf4eb65),
	.w7(32'hbbe74efb),
	.w8(32'hbc049e4d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0df0c4),
	.w1(32'hbbde0997),
	.w2(32'hb9ba278c),
	.w3(32'hba4a9f33),
	.w4(32'h3ab76f3e),
	.w5(32'hbac87518),
	.w6(32'hbb330a7c),
	.w7(32'h3a5ce5db),
	.w8(32'h3b0eb2d5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba0f11),
	.w1(32'h3c037b91),
	.w2(32'hba0d02b0),
	.w3(32'h3a7567f5),
	.w4(32'h3c020b85),
	.w5(32'h3ba6517b),
	.w6(32'hbb0fa946),
	.w7(32'hb8db18d3),
	.w8(32'h3b2dbcaf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefa2f8),
	.w1(32'hbac51d0b),
	.w2(32'hb97676ac),
	.w3(32'hbb5d61f7),
	.w4(32'hba8fb1ed),
	.w5(32'h3b6c466d),
	.w6(32'hbba28448),
	.w7(32'hbaa0f9bd),
	.w8(32'hbb55f566),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7e69a),
	.w1(32'hbb4679dd),
	.w2(32'h3a769966),
	.w3(32'h3b2fb2bf),
	.w4(32'h3b2cd0eb),
	.w5(32'h3b5f7427),
	.w6(32'hba1bd019),
	.w7(32'hb9d4d7dc),
	.w8(32'hba8293a0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b69fc),
	.w1(32'h3b87f759),
	.w2(32'hbb44e566),
	.w3(32'h3b0976af),
	.w4(32'h3b253361),
	.w5(32'hbaf473e7),
	.w6(32'h3ad37058),
	.w7(32'hb91a29f5),
	.w8(32'hbb9eece3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45823b),
	.w1(32'h3b0fbbca),
	.w2(32'h3c705f77),
	.w3(32'h3a0f11dc),
	.w4(32'h3b095413),
	.w5(32'h3cf92a77),
	.w6(32'hbb39b63a),
	.w7(32'hba6060c1),
	.w8(32'h3cbf3e27),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d092fd1),
	.w1(32'h3d0b04e3),
	.w2(32'h3bacd5bd),
	.w3(32'h3d8208b9),
	.w4(32'h3d5cde15),
	.w5(32'h3b4a34cf),
	.w6(32'h3d36741a),
	.w7(32'h3d262165),
	.w8(32'h3acbe11c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26cecf),
	.w1(32'h39f9b75c),
	.w2(32'h3a086d5a),
	.w3(32'hbb621e15),
	.w4(32'hbb7e568e),
	.w5(32'h3abdad9c),
	.w6(32'hba858c38),
	.w7(32'hbb2e5827),
	.w8(32'h3848fe53),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be463),
	.w1(32'hba49fd4b),
	.w2(32'h3a81ca6f),
	.w3(32'hbbf1dd83),
	.w4(32'hbb475365),
	.w5(32'h3b334483),
	.w6(32'hbbc074b0),
	.w7(32'hbb21c95c),
	.w8(32'h3ba43b5c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3810d5),
	.w1(32'hbabcfd04),
	.w2(32'hbc04a353),
	.w3(32'h3c0ca0d4),
	.w4(32'h3b7c877c),
	.w5(32'hbc17caed),
	.w6(32'h3c2487f0),
	.w7(32'h3b479376),
	.w8(32'hbc04fdeb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51be7),
	.w1(32'hbb0be8a5),
	.w2(32'h3960ed5b),
	.w3(32'hbb8e0908),
	.w4(32'h3af24626),
	.w5(32'h3b44b258),
	.w6(32'hbbb0416f),
	.w7(32'h3b21ef96),
	.w8(32'h3b4ac19e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba583332),
	.w1(32'h3b1f5e36),
	.w2(32'hbaeec9ed),
	.w3(32'h3b0266ba),
	.w4(32'h3b6ecc4f),
	.w5(32'hbb02e364),
	.w6(32'h3aaff3a5),
	.w7(32'h3a88ca1b),
	.w8(32'hba017a01),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba996482),
	.w1(32'hbae0c934),
	.w2(32'hbbe84e0b),
	.w3(32'hb868c40f),
	.w4(32'hbb3840ca),
	.w5(32'hbaee2c3c),
	.w6(32'hbb4c880b),
	.w7(32'hb9210408),
	.w8(32'hbb857c79),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0daee),
	.w1(32'hbb8f920a),
	.w2(32'h3c0d002c),
	.w3(32'hbb265bc3),
	.w4(32'hbb523579),
	.w5(32'h3ac304e3),
	.w6(32'hbb964664),
	.w7(32'hbb9adb5a),
	.w8(32'h3c14f7e8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d20a5),
	.w1(32'h39385be2),
	.w2(32'h3a37708c),
	.w3(32'hbc5f988b),
	.w4(32'hbc109a35),
	.w5(32'h3a3d3d55),
	.w6(32'hbb93ba4c),
	.w7(32'hba8af715),
	.w8(32'h3ac69236),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa44d0),
	.w1(32'hba29dcc2),
	.w2(32'h3a96789a),
	.w3(32'hbbbc5044),
	.w4(32'hbb370311),
	.w5(32'hbb24568f),
	.w6(32'hbbec0d4f),
	.w7(32'hbbbe23f9),
	.w8(32'h3a9dca92),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d1d0f),
	.w1(32'hb971c119),
	.w2(32'h3bb10b04),
	.w3(32'hbb0b05a0),
	.w4(32'hbb58ec21),
	.w5(32'h3ab15fae),
	.w6(32'hbb61bc1a),
	.w7(32'hba706365),
	.w8(32'h3a37d12e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecca6f),
	.w1(32'h3a290aee),
	.w2(32'h3c0ccca0),
	.w3(32'hbb06659a),
	.w4(32'h3a220c03),
	.w5(32'h3c3d69d3),
	.w6(32'hbb9847ed),
	.w7(32'h3a0bb0be),
	.w8(32'h3bf9c232),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49d055),
	.w1(32'h3b9f0fe4),
	.w2(32'h3b855108),
	.w3(32'h3c012587),
	.w4(32'h3bcefc5e),
	.w5(32'h3b848e14),
	.w6(32'h3bfd7d4b),
	.w7(32'h3bf66cc8),
	.w8(32'h3bb8be6b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831898),
	.w1(32'h3bb14f9d),
	.w2(32'h3b871edc),
	.w3(32'h3c84ccd1),
	.w4(32'h3c2d7f7f),
	.w5(32'h3b6646e1),
	.w6(32'h3bdce837),
	.w7(32'h3bc1df7c),
	.w8(32'h3b29f1d2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a70609),
	.w1(32'hb918fa34),
	.w2(32'h3c3c3a22),
	.w3(32'h3b30df89),
	.w4(32'h3b266049),
	.w5(32'h3d1cd0ff),
	.w6(32'h3b1d854f),
	.w7(32'h3ab35970),
	.w8(32'h3cb5471c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d294457),
	.w1(32'h3cbb7f7a),
	.w2(32'h3bc35d4e),
	.w3(32'h3db9ca9e),
	.w4(32'h3d842207),
	.w5(32'h3b870d9c),
	.w6(32'h3d851dc3),
	.w7(32'h3d22789b),
	.w8(32'hbae0faba),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c4564),
	.w1(32'h3bdd5a14),
	.w2(32'h392e89e0),
	.w3(32'hbb9a85ef),
	.w4(32'h3c4a6bd2),
	.w5(32'hbb752920),
	.w6(32'hbb4f239d),
	.w7(32'h3bc1405d),
	.w8(32'hbaa073bd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb570f0f),
	.w1(32'h3b24d1ad),
	.w2(32'hbb3a9928),
	.w3(32'hbb9358b8),
	.w4(32'h3b199c9a),
	.w5(32'h3a94891e),
	.w6(32'hbb9f3e8e),
	.w7(32'hbb10ca37),
	.w8(32'hba8524a9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373fe714),
	.w1(32'h397c1da0),
	.w2(32'h3b780876),
	.w3(32'hba55c20d),
	.w4(32'h3b4d03e2),
	.w5(32'hba0c7ac4),
	.w6(32'h3a4d6b40),
	.w7(32'h3b6eddbe),
	.w8(32'hbab4ad81),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1165),
	.w1(32'hbab045a6),
	.w2(32'hb9b3d249),
	.w3(32'hbb9144f7),
	.w4(32'hbabfe7e3),
	.w5(32'h3aea85f3),
	.w6(32'hbba1bd70),
	.w7(32'hbb5a03de),
	.w8(32'h3aa5814b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fc754),
	.w1(32'hba9043af),
	.w2(32'h3b04b9c6),
	.w3(32'h3bc6052a),
	.w4(32'h3a688871),
	.w5(32'h3bc01ddf),
	.w6(32'h3bd3ac51),
	.w7(32'h3b005395),
	.w8(32'h3bb27c8e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f08f0),
	.w1(32'h3b436c10),
	.w2(32'hba6bbf77),
	.w3(32'h3bb19d93),
	.w4(32'h3bb9669a),
	.w5(32'h39ba531f),
	.w6(32'h3bc245a6),
	.w7(32'h3baca06f),
	.w8(32'h3b2fe725),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2ef16),
	.w1(32'hbb464d89),
	.w2(32'hbb58ce0f),
	.w3(32'hbb88da82),
	.w4(32'hba8aa85c),
	.w5(32'hb812d328),
	.w6(32'h38140b63),
	.w7(32'hba325ae1),
	.w8(32'h3bb2f58b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cb402),
	.w1(32'hbad03374),
	.w2(32'hbb97dfd2),
	.w3(32'h3a8b91b3),
	.w4(32'h3b97e09d),
	.w5(32'h3b2e528a),
	.w6(32'h3b0aef72),
	.w7(32'h3b8aeba5),
	.w8(32'hbc047c11),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b16e5),
	.w1(32'h388633da),
	.w2(32'hbb613ab7),
	.w3(32'h3bf8ef5e),
	.w4(32'h3b4c7cd7),
	.w5(32'hba182e60),
	.w6(32'hbc0897e7),
	.w7(32'hbc419e93),
	.w8(32'hbb31b8c8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa9ada),
	.w1(32'h3bd01ff6),
	.w2(32'h3b9c2d7b),
	.w3(32'h3bbaa2f2),
	.w4(32'h3c0d7ec1),
	.w5(32'hb97749e3),
	.w6(32'hb8f43094),
	.w7(32'h3c0626ee),
	.w8(32'h394714ff),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75a4bf),
	.w1(32'hbbcaff21),
	.w2(32'hbc6e8f3c),
	.w3(32'hbb43547f),
	.w4(32'hbb9048aa),
	.w5(32'hbc27dfd9),
	.w6(32'hbb35a793),
	.w7(32'hbbbf1154),
	.w8(32'hbc0f87bf),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc087d3f),
	.w1(32'hbbaa57b3),
	.w2(32'h3b946b7d),
	.w3(32'h3bb5f5d5),
	.w4(32'h3b732195),
	.w5(32'h3afb0ada),
	.w6(32'h3b7f3558),
	.w7(32'h3b9cf6d1),
	.w8(32'h3bd10b46),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52d038),
	.w1(32'hbb3bf51b),
	.w2(32'hbad5e1dc),
	.w3(32'hbb9295a6),
	.w4(32'hbbdfff28),
	.w5(32'hb96b0869),
	.w6(32'hbbaf32e1),
	.w7(32'hbbb428fb),
	.w8(32'hb90f1183),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72d41a),
	.w1(32'hbb919569),
	.w2(32'h3bde0e78),
	.w3(32'hbb982cce),
	.w4(32'hbbb229b1),
	.w5(32'h3be2c48e),
	.w6(32'hbb032d14),
	.w7(32'h39d9c572),
	.w8(32'h3c03e40e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee22fb),
	.w1(32'h3bee4420),
	.w2(32'hbb774e37),
	.w3(32'h3bf6ad6b),
	.w4(32'h3bf1742b),
	.w5(32'h3b9638d4),
	.w6(32'h3bdbdde9),
	.w7(32'h3b96d9e5),
	.w8(32'hba2d0182),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adba4f0),
	.w1(32'h3acc056c),
	.w2(32'h3bc655b6),
	.w3(32'hbac3d69b),
	.w4(32'h3afca591),
	.w5(32'h3c0c3fd2),
	.w6(32'hba9a1de3),
	.w7(32'hb92c99ca),
	.w8(32'h3a9d6ff1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c7f4),
	.w1(32'h3bb103de),
	.w2(32'hbaf62881),
	.w3(32'h3b3fbec4),
	.w4(32'h3b846e7f),
	.w5(32'hb99ee38d),
	.w6(32'hbb1899ad),
	.w7(32'h3990958d),
	.w8(32'h3b2af44f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4b8b4),
	.w1(32'hbc7a8bd0),
	.w2(32'h3c0817a4),
	.w3(32'hbbcfeb9c),
	.w4(32'hbc75d34d),
	.w5(32'hba4aa420),
	.w6(32'hba963d2f),
	.w7(32'hbc0c4e9e),
	.w8(32'h3b404520),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ef87c),
	.w1(32'hbb99c3ae),
	.w2(32'hba09d152),
	.w3(32'hbaa8f33c),
	.w4(32'hbb96884f),
	.w5(32'h3af29088),
	.w6(32'h3825e6c0),
	.w7(32'hbb27de19),
	.w8(32'hbb82c3a3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e6a5d),
	.w1(32'h3b66f38b),
	.w2(32'h39c2db00),
	.w3(32'h3a945ded),
	.w4(32'hbb1d86df),
	.w5(32'h3ba018f8),
	.w6(32'hbaadd32c),
	.w7(32'h3a8686ca),
	.w8(32'h3bc97430),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895535),
	.w1(32'hbb349a41),
	.w2(32'h3ba19e9d),
	.w3(32'hbb1a153d),
	.w4(32'hbb1681dc),
	.w5(32'h3b95c86a),
	.w6(32'hbb91aeb3),
	.w7(32'hbb860ce1),
	.w8(32'h3a495af3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bbf4e),
	.w1(32'hba377c9e),
	.w2(32'h3be4fa29),
	.w3(32'hb6a8c924),
	.w4(32'h3ad5434c),
	.w5(32'h3c09e841),
	.w6(32'hb9f17eda),
	.w7(32'hbb4dbacd),
	.w8(32'h3b6d3c94),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c11f),
	.w1(32'h3bda53e6),
	.w2(32'h3c0de798),
	.w3(32'h3befed1a),
	.w4(32'h3b8a1011),
	.w5(32'h3c28d0ce),
	.w6(32'h3bbf3181),
	.w7(32'h3a9a380d),
	.w8(32'h3c1ed46a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb970e13d),
	.w1(32'hb9bb26d4),
	.w2(32'hba94ffb1),
	.w3(32'hbb0616f5),
	.w4(32'h3999b84b),
	.w5(32'hb8e25baa),
	.w6(32'h3a7d3269),
	.w7(32'hba8900f8),
	.w8(32'hbac20ae5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb174d62),
	.w1(32'h3895549b),
	.w2(32'hbb273a37),
	.w3(32'hbb459be7),
	.w4(32'h39a144f4),
	.w5(32'hbaf101f8),
	.w6(32'hbb01c6cd),
	.w7(32'hba86a6ca),
	.w8(32'h3b627919),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d7e17),
	.w1(32'hbbb13661),
	.w2(32'hbb86b3a7),
	.w3(32'hbbaad587),
	.w4(32'hbbef088b),
	.w5(32'h398a0b33),
	.w6(32'h3a9ae4bd),
	.w7(32'hb983bd2c),
	.w8(32'h3aa0f17f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eaebb),
	.w1(32'h39885c03),
	.w2(32'h3bc229d2),
	.w3(32'h3a3957a2),
	.w4(32'hbb0de3fc),
	.w5(32'h3bb46456),
	.w6(32'h3a0503f2),
	.w7(32'hbab6db19),
	.w8(32'h3afb886d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4aba5f),
	.w1(32'h3b1b4a89),
	.w2(32'h3b8a2ef7),
	.w3(32'h3b26165e),
	.w4(32'h3b0597fe),
	.w5(32'h3bb72d40),
	.w6(32'h3a929ced),
	.w7(32'h3b226b4d),
	.w8(32'h3a2a7b60),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdec975),
	.w1(32'h3b20a8d6),
	.w2(32'h3ae26f14),
	.w3(32'h3b4de63d),
	.w4(32'h3b7b6bdc),
	.w5(32'h3b1e3c92),
	.w6(32'h3bbaf44b),
	.w7(32'h3a05b62a),
	.w8(32'h3b1f04d5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84c2ee),
	.w1(32'hba0d0d96),
	.w2(32'hbbd614e6),
	.w3(32'h3b9671c9),
	.w4(32'h3b27b52c),
	.w5(32'h3a98ce38),
	.w6(32'h3b26a867),
	.w7(32'h3b53433c),
	.w8(32'h3aa13cfc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76174c),
	.w1(32'hbb9457d4),
	.w2(32'hb99f7498),
	.w3(32'hbbd92d92),
	.w4(32'h3b5a715b),
	.w5(32'h3b7af1e4),
	.w6(32'hbb43b8b6),
	.w7(32'h3bfa2c13),
	.w8(32'h3b33c4dc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49d82e),
	.w1(32'h3b2c006c),
	.w2(32'h3b5a964d),
	.w3(32'h3b8b030f),
	.w4(32'h3b186d48),
	.w5(32'h3b1ddadf),
	.w6(32'hbab8df6d),
	.w7(32'h388a0c0e),
	.w8(32'h3b83e329),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10cb20),
	.w1(32'hbac98ace),
	.w2(32'hbb54789b),
	.w3(32'h3b08ea59),
	.w4(32'h3b229d35),
	.w5(32'hbb1944c7),
	.w6(32'h3b3a9b2c),
	.w7(32'h3bee5737),
	.w8(32'h3b4d05ca),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd12776),
	.w1(32'hbc034a17),
	.w2(32'hbc60a088),
	.w3(32'hbb70362e),
	.w4(32'hbb91a53d),
	.w5(32'hbc246d96),
	.w6(32'h3b52a9f8),
	.w7(32'h3a9d722c),
	.w8(32'hbc1959e7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b2a8b),
	.w1(32'hbc3f2ba4),
	.w2(32'hb92ac429),
	.w3(32'hbc0ecb76),
	.w4(32'hbc11aabf),
	.w5(32'h3a520d2d),
	.w6(32'hbb932ca4),
	.w7(32'hbbc03266),
	.w8(32'h3a59cea0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b8a77),
	.w1(32'hbb288a92),
	.w2(32'hba607b70),
	.w3(32'h3a85bf03),
	.w4(32'h3b2cb554),
	.w5(32'hbb6e5bd7),
	.w6(32'h3ac835e3),
	.w7(32'h3b4ad6d9),
	.w8(32'hba82f60a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0af0f),
	.w1(32'hbafa0733),
	.w2(32'h395f48a4),
	.w3(32'hbb65f42d),
	.w4(32'hbb26d94e),
	.w5(32'hbbd26283),
	.w6(32'hba42c3a3),
	.w7(32'h3b7de903),
	.w8(32'hbae18ac1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1c8ab),
	.w1(32'h39170ccc),
	.w2(32'h3b1f59c5),
	.w3(32'hbbdb4f8c),
	.w4(32'hbb0ffaed),
	.w5(32'h3a2a0389),
	.w6(32'h3ace76c6),
	.w7(32'hba775c35),
	.w8(32'h3ab8a2d4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cbe0a),
	.w1(32'hba4a8a87),
	.w2(32'hb9330e5c),
	.w3(32'hbafff655),
	.w4(32'hbb012bd3),
	.w5(32'hbb3108a4),
	.w6(32'h3b621cd5),
	.w7(32'h3a97b551),
	.w8(32'hbb12513f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a4041),
	.w1(32'hbb1e5031),
	.w2(32'hbc0e32bb),
	.w3(32'hbc0748b0),
	.w4(32'hbc0b7362),
	.w5(32'hbc01dd03),
	.w6(32'hbc29cb46),
	.w7(32'hbc07705d),
	.w8(32'hbc345112),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea7185),
	.w1(32'hbc4e3968),
	.w2(32'hbb747383),
	.w3(32'hbb2bab61),
	.w4(32'hbbfabe26),
	.w5(32'hba18462b),
	.w6(32'hbbcbd0ce),
	.w7(32'hbc3dbaf1),
	.w8(32'h3ac7016e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04eb24),
	.w1(32'hba779a72),
	.w2(32'hbbafb39f),
	.w3(32'hb983c419),
	.w4(32'h39ce3b02),
	.w5(32'hbbad37e1),
	.w6(32'h3b274cc7),
	.w7(32'hbb8cb729),
	.w8(32'hb992117a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31ec8),
	.w1(32'h39745b45),
	.w2(32'hbb16d13d),
	.w3(32'hbb73c7a2),
	.w4(32'h3ad77922),
	.w5(32'hbb8c80ef),
	.w6(32'h39fc40a2),
	.w7(32'h3b5ec1ac),
	.w8(32'hba3daaf0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90431a),
	.w1(32'hbab28a72),
	.w2(32'hbb19a7cc),
	.w3(32'h3bb55331),
	.w4(32'h3b8a56e3),
	.w5(32'hbb70dce9),
	.w6(32'h3a698290),
	.w7(32'h3be0d0bb),
	.w8(32'hbb578429),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa5e43),
	.w1(32'hbb37ab8c),
	.w2(32'hba4be361),
	.w3(32'hbbb437f1),
	.w4(32'h3bf4bd42),
	.w5(32'hba869004),
	.w6(32'hbb8ffaca),
	.w7(32'h3b97740c),
	.w8(32'hb9ecec6a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d843e),
	.w1(32'hb9b64fa9),
	.w2(32'hbb8ee098),
	.w3(32'hbbd40927),
	.w4(32'h3ae165fa),
	.w5(32'hba81ff20),
	.w6(32'hbbcaa380),
	.w7(32'h3a897dfb),
	.w8(32'h3bd5e18e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7cbf1),
	.w1(32'hbb877b14),
	.w2(32'h3b065041),
	.w3(32'hbb21b7e0),
	.w4(32'h3ac179ba),
	.w5(32'h3bd96cf0),
	.w6(32'hbbc5e28f),
	.w7(32'hbbd8d669),
	.w8(32'h3bae0e4a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecb09f),
	.w1(32'hbb2dcaf6),
	.w2(32'hbb5d1d89),
	.w3(32'hb937aaf8),
	.w4(32'h3a0b7c87),
	.w5(32'h38870edb),
	.w6(32'hba70002d),
	.w7(32'hb9020879),
	.w8(32'hbae6a1dd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac19dc3),
	.w1(32'hbb654524),
	.w2(32'h3877d8b4),
	.w3(32'h3ba5e11b),
	.w4(32'hba8d683c),
	.w5(32'h3a6b0f17),
	.w6(32'h39ddd9a8),
	.w7(32'h3b221601),
	.w8(32'h3ad6f1f7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388998fa),
	.w1(32'h3a610c21),
	.w2(32'h3bf77134),
	.w3(32'hb8d17c86),
	.w4(32'h3af2675e),
	.w5(32'hbab6cd3c),
	.w6(32'hb9ff988f),
	.w7(32'h3adebcf8),
	.w8(32'hbb514402),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ca75),
	.w1(32'hba1be2ba),
	.w2(32'h3b6a2eb8),
	.w3(32'hbb96d0fb),
	.w4(32'hbb0886f7),
	.w5(32'h3bc94e97),
	.w6(32'hbac7604f),
	.w7(32'hbb71d53f),
	.w8(32'h3b6cac6c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b244a2f),
	.w1(32'hb9c2224f),
	.w2(32'hbc1bd3a1),
	.w3(32'h3b92c5a5),
	.w4(32'h3aa86238),
	.w5(32'hbc429fa7),
	.w6(32'h3b6061be),
	.w7(32'h3ad79a4f),
	.w8(32'hbb454e0d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae614c),
	.w1(32'hbbf72829),
	.w2(32'hbb4dee2b),
	.w3(32'hbca43bf3),
	.w4(32'hbbffd883),
	.w5(32'hbb819673),
	.w6(32'hbc5214ab),
	.w7(32'hbb00f441),
	.w8(32'h3b789a10),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40984f),
	.w1(32'hbc40a6a7),
	.w2(32'hbb1c67f4),
	.w3(32'hbbebc23c),
	.w4(32'hbbc7a39c),
	.w5(32'h3b9b98b1),
	.w6(32'hb9d8dc71),
	.w7(32'hbb1489f2),
	.w8(32'h39ff8b5b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8c6e),
	.w1(32'hbb7de46e),
	.w2(32'hbafaea4b),
	.w3(32'hba14908a),
	.w4(32'hbb099632),
	.w5(32'hbac9e90a),
	.w6(32'hbb8b45f5),
	.w7(32'hbb3aacf5),
	.w8(32'h376f44b6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb510fe9),
	.w1(32'hbb0d6a40),
	.w2(32'hbb23ab09),
	.w3(32'hbb7a0c8f),
	.w4(32'hba7a2cf7),
	.w5(32'h3bada86b),
	.w6(32'hbbb62d4c),
	.w7(32'hba933138),
	.w8(32'hbb0f2a03),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebd3eb),
	.w1(32'hb9f0b84c),
	.w2(32'h3ac0bd76),
	.w3(32'h3cda9ca7),
	.w4(32'h3c80ef10),
	.w5(32'h3a944eff),
	.w6(32'h3c66ea8d),
	.w7(32'h3bc427ff),
	.w8(32'h3b6b18cd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5fec6),
	.w1(32'h3ad149aa),
	.w2(32'hbc545310),
	.w3(32'hbb82f3c8),
	.w4(32'hb7aec132),
	.w5(32'hbc9d77b2),
	.w6(32'hba9290b6),
	.w7(32'h3a265d7f),
	.w8(32'hbc7feb40),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac6701),
	.w1(32'hbc99433c),
	.w2(32'h3a881643),
	.w3(32'hbcf684bb),
	.w4(32'hbce3d797),
	.w5(32'hbb17fd88),
	.w6(32'hbcd3dde9),
	.w7(32'hbcc2764a),
	.w8(32'h3a464489),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4b4f6),
	.w1(32'hbb9646be),
	.w2(32'h3a821aca),
	.w3(32'h3bd0950e),
	.w4(32'hba6a86ea),
	.w5(32'h399ae6cf),
	.w6(32'h3bda9e93),
	.w7(32'h3a67dd63),
	.w8(32'hba2d9a29),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75d167),
	.w1(32'hba4f3f16),
	.w2(32'h3b3dfe1d),
	.w3(32'hbb4883d5),
	.w4(32'hbbaaa4bb),
	.w5(32'h3b8bd495),
	.w6(32'h3a0b78c7),
	.w7(32'h3b08f994),
	.w8(32'h3b44b2f1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab60aea),
	.w1(32'h3a5bb432),
	.w2(32'h3c248883),
	.w3(32'h3a23e628),
	.w4(32'h3ae602b0),
	.w5(32'h3cafdf28),
	.w6(32'h3ad23f9a),
	.w7(32'h3b7fc05b),
	.w8(32'h3c6c385f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc117f7),
	.w1(32'h3c8b6c11),
	.w2(32'h3af87016),
	.w3(32'h3d3fa7a6),
	.w4(32'h3d14d92a),
	.w5(32'h3b234396),
	.w6(32'h3d131592),
	.w7(32'h3cdc63d8),
	.w8(32'h3b5becc8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c5b2b),
	.w1(32'h3b278dec),
	.w2(32'h3a4fe8f9),
	.w3(32'h3b388153),
	.w4(32'h3b8e8526),
	.w5(32'h3b07eef9),
	.w6(32'h3b6bee88),
	.w7(32'h3b5cc939),
	.w8(32'h3aa2eb61),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f42af),
	.w1(32'h3aea94e1),
	.w2(32'h3a91c481),
	.w3(32'h3b26810f),
	.w4(32'h39803e80),
	.w5(32'h3b4947a5),
	.w6(32'h3bac5d68),
	.w7(32'h3b181d56),
	.w8(32'h3b511bd4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb106b91),
	.w1(32'h3bd9b6c8),
	.w2(32'h3a95b0cf),
	.w3(32'hbb6aabcf),
	.w4(32'hbabd01bb),
	.w5(32'h3916891f),
	.w6(32'hbaf0736f),
	.w7(32'h3ad6c618),
	.w8(32'h3ad9c74f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77b14c),
	.w1(32'h39ac4ec7),
	.w2(32'h3a918d39),
	.w3(32'h3a1444bd),
	.w4(32'h39f382d2),
	.w5(32'h3b0faa56),
	.w6(32'h3ad3416e),
	.w7(32'h3b049a91),
	.w8(32'h3a8f6860),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38a5e1),
	.w1(32'h3a2d96dd),
	.w2(32'h3b21e747),
	.w3(32'h3b2b99a6),
	.w4(32'hbaa84b07),
	.w5(32'h3b03c351),
	.w6(32'hbac7718e),
	.w7(32'hba147a16),
	.w8(32'hb8ab0bf7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10f359),
	.w1(32'h3831163e),
	.w2(32'hbba5d791),
	.w3(32'hbbb20ba8),
	.w4(32'hbacd644a),
	.w5(32'hbb09e0e6),
	.w6(32'hbb8309b9),
	.w7(32'hbb061def),
	.w8(32'hbbb401b8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb938cf),
	.w1(32'hbbf030df),
	.w2(32'h3b3e75d0),
	.w3(32'hbba839aa),
	.w4(32'hbbc9930d),
	.w5(32'h3b8fae10),
	.w6(32'hbc3a2827),
	.w7(32'hbc372dbd),
	.w8(32'h378ac502),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b702ce0),
	.w1(32'h3a017ab6),
	.w2(32'hbb76d930),
	.w3(32'h3c17a002),
	.w4(32'h3b1f4b70),
	.w5(32'hbb8bda45),
	.w6(32'h3c0cbc69),
	.w7(32'h3b8e21e5),
	.w8(32'h39a4e727),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21706d),
	.w1(32'hbb570454),
	.w2(32'h3b22a466),
	.w3(32'hbc1335f0),
	.w4(32'hbbcc9b85),
	.w5(32'h3b49600c),
	.w6(32'hbb46e929),
	.w7(32'hbb826efe),
	.w8(32'hba167668),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb112835),
	.w1(32'h393a6dd0),
	.w2(32'hbb04c639),
	.w3(32'hb9fbf3cd),
	.w4(32'hb957e863),
	.w5(32'hbaf29fb0),
	.w6(32'h3b01f3a4),
	.w7(32'hbb3606cd),
	.w8(32'hba28bb60),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab34f1),
	.w1(32'hbaf49e1a),
	.w2(32'hbbaf1306),
	.w3(32'hbaa2641b),
	.w4(32'hba34b632),
	.w5(32'hbc1a1411),
	.w6(32'h3af47147),
	.w7(32'h391e6d88),
	.w8(32'hbb9ccc44),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2df629),
	.w1(32'h3b34a2e6),
	.w2(32'hbbf0223a),
	.w3(32'hbc5be96c),
	.w4(32'h3bdd8eaa),
	.w5(32'hbc7278d8),
	.w6(32'hbb88bae2),
	.w7(32'h3bcdabbd),
	.w8(32'hbc5ab5cc),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a8c8b),
	.w1(32'h3b071f5e),
	.w2(32'hbb820134),
	.w3(32'hbc8d54d7),
	.w4(32'h3b1d57a6),
	.w5(32'hbb547a69),
	.w6(32'hbc218e89),
	.w7(32'h3a00622c),
	.w8(32'hbb391097),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4ff26),
	.w1(32'h39cb6f59),
	.w2(32'h3b69e7c3),
	.w3(32'hbb61f562),
	.w4(32'hbb228c5f),
	.w5(32'h3c3b4352),
	.w6(32'hbbab6e12),
	.w7(32'hbb887f2a),
	.w8(32'h3c1b667f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36ccd),
	.w1(32'h3b9fe580),
	.w2(32'hbc672306),
	.w3(32'h3c013315),
	.w4(32'h3b0b4890),
	.w5(32'hbbd777c3),
	.w6(32'h3bb644dc),
	.w7(32'h3b791ac6),
	.w8(32'h3c069449),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2437e8),
	.w1(32'hbc2f8fd4),
	.w2(32'h3a0a7145),
	.w3(32'hbced2d2e),
	.w4(32'hbcd26dfb),
	.w5(32'h3ba2cb9b),
	.w6(32'hbc087111),
	.w7(32'hbc11ce5c),
	.w8(32'h3b0eb21a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee5e8),
	.w1(32'hb9c77b78),
	.w2(32'hbbeb860b),
	.w3(32'h3bb5f58f),
	.w4(32'h3b779519),
	.w5(32'hbb460004),
	.w6(32'hbb289d9e),
	.w7(32'hbb7e43ab),
	.w8(32'h3b77b2eb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb358d8c),
	.w1(32'hbc124232),
	.w2(32'h3b3330c6),
	.w3(32'hbb525f64),
	.w4(32'hbcee8326),
	.w5(32'h3b2956bf),
	.w6(32'hbc5e65bf),
	.w7(32'hbcbb8bb5),
	.w8(32'h3b81b5b6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b8864),
	.w1(32'hbacd59b1),
	.w2(32'hbadab004),
	.w3(32'hb937ae4f),
	.w4(32'hbadd0e77),
	.w5(32'hbc48dfbe),
	.w6(32'hbaa93030),
	.w7(32'hbb696c0e),
	.w8(32'hbbe1524f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954a87b),
	.w1(32'hbaf48921),
	.w2(32'hbbe9967f),
	.w3(32'hbc16a8dc),
	.w4(32'hbbd4ab79),
	.w5(32'hbc28f05e),
	.w6(32'hbc04be62),
	.w7(32'hbc567cd1),
	.w8(32'hbc534f64),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7f50c),
	.w1(32'h3b421348),
	.w2(32'h3b7c79d5),
	.w3(32'hbb6f0d4c),
	.w4(32'h39d1f1b9),
	.w5(32'h3c654a80),
	.w6(32'hbc286fae),
	.w7(32'hbb99eb20),
	.w8(32'h3a3d4437),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dc936),
	.w1(32'h3baaa3a9),
	.w2(32'hbb2e845c),
	.w3(32'h3c180697),
	.w4(32'h3c350828),
	.w5(32'hbbc7d299),
	.w6(32'h3c48d03b),
	.w7(32'h3c66fe77),
	.w8(32'h3a81a3e2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f1c32),
	.w1(32'h3b11028b),
	.w2(32'hb9d056cd),
	.w3(32'hbcae271c),
	.w4(32'hbc99fb71),
	.w5(32'h3abd8ba5),
	.w6(32'hbc087e63),
	.w7(32'hbc22c498),
	.w8(32'h3ba3a55c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb873de4),
	.w1(32'hbb72f27d),
	.w2(32'hb94a1746),
	.w3(32'hbc1f37cd),
	.w4(32'hbbd7777e),
	.w5(32'h3c8e3e97),
	.w6(32'hbc014c03),
	.w7(32'hbc0ff821),
	.w8(32'h3b82cc8b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a1a1c),
	.w1(32'hbbec390e),
	.w2(32'h3ad561d7),
	.w3(32'h3b54d42a),
	.w4(32'hbc8d3e86),
	.w5(32'h3b00198a),
	.w6(32'h3b989d7f),
	.w7(32'hbc06b375),
	.w8(32'h3c5d206d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902933),
	.w1(32'hbb6c388d),
	.w2(32'h3b84c702),
	.w3(32'h3c03986a),
	.w4(32'h3bcd19db),
	.w5(32'h3a830e69),
	.w6(32'h3c453243),
	.w7(32'h3bb9a41d),
	.w8(32'h3b15d6c4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac79822),
	.w1(32'hbab77068),
	.w2(32'hbae4cbfd),
	.w3(32'hbb8ec1f5),
	.w4(32'hbb5fee63),
	.w5(32'h3b30ef39),
	.w6(32'hbb7779cd),
	.w7(32'hbad4dc36),
	.w8(32'h3b556d12),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a92e9),
	.w1(32'h3afd03a3),
	.w2(32'h3afb5846),
	.w3(32'hbc251b9b),
	.w4(32'h3aa1affa),
	.w5(32'h3c5c98ce),
	.w6(32'hbbfb35b5),
	.w7(32'h3c4a985e),
	.w8(32'h3bac5e75),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840b90),
	.w1(32'hbb7a3458),
	.w2(32'h3c9495fb),
	.w3(32'h3b24f534),
	.w4(32'h3ada590e),
	.w5(32'h3cf08841),
	.w6(32'h3a5fba97),
	.w7(32'h3bfe1177),
	.w8(32'h3cc69022),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14a24f),
	.w1(32'h3bb715bb),
	.w2(32'h3c07b42f),
	.w3(32'h3c313a91),
	.w4(32'hbadf0f80),
	.w5(32'h3ceb9738),
	.w6(32'h3c51158e),
	.w7(32'hbb0312db),
	.w8(32'h3cb7bde4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868c3b),
	.w1(32'hbc974d9e),
	.w2(32'hbb4c3a46),
	.w3(32'h3c03d541),
	.w4(32'hbce33df5),
	.w5(32'hbbc871ca),
	.w6(32'h3c137df5),
	.w7(32'hbca63c06),
	.w8(32'hbbac4dbd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b2b0e),
	.w1(32'h3a31d92f),
	.w2(32'h3c0c5396),
	.w3(32'hbb98d7c7),
	.w4(32'hbaeb4928),
	.w5(32'h3c63d6a4),
	.w6(32'hbb6292a3),
	.w7(32'hba30abc5),
	.w8(32'h3c2b5832),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4874c2),
	.w1(32'h3a3fc6ef),
	.w2(32'hbab7bc30),
	.w3(32'h3c6b5081),
	.w4(32'h3bcf2035),
	.w5(32'h3c39ffe3),
	.w6(32'h3bd59c4b),
	.w7(32'h3b9f4075),
	.w8(32'h3c3f9bda),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b741dab),
	.w1(32'h3b664fa9),
	.w2(32'h3b522ed2),
	.w3(32'h3bfa4915),
	.w4(32'h3b9e507d),
	.w5(32'h3c01ac84),
	.w6(32'h3be5e6e1),
	.w7(32'h3c194b60),
	.w8(32'h3b8609b0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2b639),
	.w1(32'hbc5b2fd0),
	.w2(32'h3ba9a479),
	.w3(32'hbc38c051),
	.w4(32'hbca26b43),
	.w5(32'h3bacd834),
	.w6(32'h3b8b5464),
	.w7(32'hbb11cdc5),
	.w8(32'h3c12e36f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc4435),
	.w1(32'h3b9109af),
	.w2(32'h3abe39b4),
	.w3(32'h3c43e8c2),
	.w4(32'h3c195ece),
	.w5(32'h3c38d69b),
	.w6(32'h3c49ebc8),
	.w7(32'h3c4fccac),
	.w8(32'h3c1ba8ef),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f711ca),
	.w1(32'h3ac07466),
	.w2(32'h3bd154cd),
	.w3(32'h3b96ba0a),
	.w4(32'hbab5b71b),
	.w5(32'h3c3e39ea),
	.w6(32'hba43c7a9),
	.w7(32'hbb243206),
	.w8(32'h3bd31c99),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca50a3c),
	.w1(32'h3bc97c77),
	.w2(32'hbbf6703c),
	.w3(32'h3c22ebe4),
	.w4(32'h3b9db7da),
	.w5(32'hba25f7ff),
	.w6(32'h3c0ccebc),
	.w7(32'h3c59ea76),
	.w8(32'hbba3ef5b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc0869),
	.w1(32'h3bab5b69),
	.w2(32'hba609756),
	.w3(32'hbc59f6f5),
	.w4(32'hbc19fc29),
	.w5(32'h3b4404d4),
	.w6(32'hbc19cc69),
	.w7(32'hbc06f070),
	.w8(32'h3baa4909),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccde7a2),
	.w1(32'hbc46f2c0),
	.w2(32'h3b6a5f89),
	.w3(32'hbce2fa4c),
	.w4(32'hbcb0ab95),
	.w5(32'h3c12443e),
	.w6(32'hbc911418),
	.w7(32'hbc8b6d1c),
	.w8(32'h3c03bc44),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14248c),
	.w1(32'hbb3d6ab3),
	.w2(32'h3b80ac0a),
	.w3(32'hba2152ab),
	.w4(32'hbc3e4a63),
	.w5(32'h3c063596),
	.w6(32'hbb7be467),
	.w7(32'hbc043168),
	.w8(32'h3ad24dfd),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06693d),
	.w1(32'h3c982456),
	.w2(32'h3b59e48c),
	.w3(32'h3b353b1f),
	.w4(32'h3c7230bd),
	.w5(32'h3bdb69e4),
	.w6(32'hbbed7897),
	.w7(32'h3bd73307),
	.w8(32'h3ba81b66),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3b04d),
	.w1(32'h392e4f85),
	.w2(32'h3b816f7c),
	.w3(32'hb6a5f2af),
	.w4(32'hbbbace3c),
	.w5(32'h3a684e68),
	.w6(32'hbbb2433f),
	.w7(32'hbb917f69),
	.w8(32'hbbb60c40),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b6345),
	.w1(32'h3c073756),
	.w2(32'h3bf7f21a),
	.w3(32'h3c47dd65),
	.w4(32'h3c73f778),
	.w5(32'h3c01d5b7),
	.w6(32'h3b974107),
	.w7(32'h3c6f1612),
	.w8(32'h3bdf4bf1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d929),
	.w1(32'hbbb21732),
	.w2(32'hbb8c06f5),
	.w3(32'hbbc94755),
	.w4(32'hbc09b85a),
	.w5(32'h3af7976c),
	.w6(32'hba49021b),
	.w7(32'hbb974025),
	.w8(32'hbb9a90ea),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb6c0),
	.w1(32'hbb1d14f2),
	.w2(32'h39613bc8),
	.w3(32'hbb775786),
	.w4(32'h3bb20788),
	.w5(32'h3bae47bb),
	.w6(32'hbb4d9915),
	.w7(32'hbb6d851b),
	.w8(32'hb99c1d96),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4321),
	.w1(32'h3bb9cc96),
	.w2(32'h3beda56a),
	.w3(32'h3afbf764),
	.w4(32'h39e613e1),
	.w5(32'h3c1a3714),
	.w6(32'hbb9b570b),
	.w7(32'hba541fa7),
	.w8(32'h3bb9dbed),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b858e2b),
	.w1(32'h3a51e85f),
	.w2(32'hbac00a72),
	.w3(32'h3bdaf2ab),
	.w4(32'h3b7012ed),
	.w5(32'hb9f6c4a3),
	.w6(32'h3ba57bee),
	.w7(32'h3b988664),
	.w8(32'h39ffd773),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb465944),
	.w1(32'h3c1e3a45),
	.w2(32'h3b249273),
	.w3(32'hbc16cdde),
	.w4(32'h3b9a6389),
	.w5(32'hbb7b97e4),
	.w6(32'hbc02e0d6),
	.w7(32'h3af01756),
	.w8(32'hbb0d47a9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0933cc),
	.w1(32'h3b80fdb0),
	.w2(32'h3b2b732a),
	.w3(32'hbbd8471b),
	.w4(32'h3bc5b09f),
	.w5(32'h3bee9b1b),
	.w6(32'hbb682fd0),
	.w7(32'h3b845142),
	.w8(32'hbb2adea9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9cd51),
	.w1(32'hbc8d66b2),
	.w2(32'hbb91462c),
	.w3(32'hba3a5e01),
	.w4(32'hbc4554d4),
	.w5(32'h39cbee84),
	.w6(32'hba98483a),
	.w7(32'h3aa2ffa8),
	.w8(32'hbbbba010),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddbdaa),
	.w1(32'hbbd7c12c),
	.w2(32'hba80a960),
	.w3(32'h3c086861),
	.w4(32'hbb4cc0f3),
	.w5(32'hbbbf899b),
	.w6(32'h3ba12eae),
	.w7(32'hbb969566),
	.w8(32'hbb9ac11a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52d934),
	.w1(32'h3c347de1),
	.w2(32'hbbdf64a9),
	.w3(32'hbc075c63),
	.w4(32'h3bf7f158),
	.w5(32'hbc5d113a),
	.w6(32'hbc08ccb2),
	.w7(32'h3c0359b0),
	.w8(32'hbbc8870a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aee62),
	.w1(32'hbb4ba962),
	.w2(32'h3b61a27f),
	.w3(32'hbc9153a6),
	.w4(32'hbb55fafa),
	.w5(32'h3b87300a),
	.w6(32'hbc140f98),
	.w7(32'hbadf2a10),
	.w8(32'h3c28a380),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227640),
	.w1(32'hb9c939b1),
	.w2(32'h3ba35735),
	.w3(32'hbc25c9ad),
	.w4(32'hbc0c8ee2),
	.w5(32'h3c029726),
	.w6(32'hb733252b),
	.w7(32'h3a62ef98),
	.w8(32'h3a290c98),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba676004),
	.w1(32'hbc323b47),
	.w2(32'hbc4c6b96),
	.w3(32'h3ab1bdd3),
	.w4(32'hbcc8e59f),
	.w5(32'hbc87a08a),
	.w6(32'h3ad2f5a2),
	.w7(32'hbcad7251),
	.w8(32'hbc098480),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7a66c),
	.w1(32'hbba84e3e),
	.w2(32'hba5de914),
	.w3(32'hbcf5f794),
	.w4(32'hbc58008d),
	.w5(32'hbbb15910),
	.w6(32'hbcd164ba),
	.w7(32'hbc5b390f),
	.w8(32'hbb94391e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960971e),
	.w1(32'h3b8cbc9d),
	.w2(32'h3bf63acf),
	.w3(32'hbbd8746a),
	.w4(32'h3b2365fc),
	.w5(32'h3d069933),
	.w6(32'hbbd93c00),
	.w7(32'h3971152f),
	.w8(32'h3cd3a949),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72a91d0),
	.w1(32'hbca82445),
	.w2(32'hba0f0fd2),
	.w3(32'h3c6a534f),
	.w4(32'hbc920056),
	.w5(32'h3b5ba381),
	.w6(32'h3c3a8692),
	.w7(32'hbc8bbb94),
	.w8(32'h3bfdd394),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53870),
	.w1(32'h3b1f56a3),
	.w2(32'h3c4f12ec),
	.w3(32'h3c4bb273),
	.w4(32'hbb92757c),
	.w5(32'h3c548288),
	.w6(32'h3bee4fed),
	.w7(32'hbbc560b2),
	.w8(32'h3c58f5f4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b079327),
	.w1(32'h3b6e9c42),
	.w2(32'h3c31af64),
	.w3(32'h3c3400da),
	.w4(32'h3bb2f636),
	.w5(32'h3cba18f3),
	.w6(32'h3c053cd6),
	.w7(32'h39c8d0c1),
	.w8(32'h3c236f9b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc7044),
	.w1(32'hbc53d0b1),
	.w2(32'h3ad200ee),
	.w3(32'h3b2b2e8e),
	.w4(32'hbc8b2cd5),
	.w5(32'hb9083a82),
	.w6(32'h3c369096),
	.w7(32'hbc2992d5),
	.w8(32'h3b7dfd0e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfff2a6),
	.w1(32'h3a45ae1c),
	.w2(32'h3a50d4ba),
	.w3(32'hbc8a155b),
	.w4(32'hbaa94064),
	.w5(32'h3c0ceb48),
	.w6(32'hbc28698a),
	.w7(32'h3b479118),
	.w8(32'h3c12bb2c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbe226),
	.w1(32'h3981962a),
	.w2(32'hba434b69),
	.w3(32'h3c32684c),
	.w4(32'hbaebbefb),
	.w5(32'h399643a5),
	.w6(32'h3be4858d),
	.w7(32'hb7ddd700),
	.w8(32'h39473539),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b4d1b),
	.w1(32'h3b62cac3),
	.w2(32'hbbb4e3af),
	.w3(32'hbb4db5d7),
	.w4(32'h3b929213),
	.w5(32'hbb84f7f7),
	.w6(32'hbb856061),
	.w7(32'h3b8a348b),
	.w8(32'hbc08fdcd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc98410),
	.w1(32'hbcef1ecd),
	.w2(32'h3cb72105),
	.w3(32'hbd09c19f),
	.w4(32'hbd156211),
	.w5(32'h3ca4b510),
	.w6(32'hbd02c808),
	.w7(32'hbcfb983d),
	.w8(32'h3c63c3ca),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddd9fc),
	.w1(32'hbc2e342e),
	.w2(32'h3c55f9f6),
	.w3(32'h3c42eeda),
	.w4(32'hbc06790a),
	.w5(32'h3cad0f19),
	.w6(32'h3ca42a91),
	.w7(32'hbaae9ba9),
	.w8(32'h3c52a932),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9475a),
	.w1(32'h3bf383be),
	.w2(32'hbae78cdd),
	.w3(32'h3c242f1a),
	.w4(32'hb81cbe20),
	.w5(32'hbb26db7e),
	.w6(32'h3bee9829),
	.w7(32'h3b6a655d),
	.w8(32'hbb8b4bc5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd5f473),
	.w1(32'hbd117346),
	.w2(32'hbc6c2d32),
	.w3(32'hbd33867d),
	.w4(32'hbd48278d),
	.w5(32'hbc26a37d),
	.w6(32'hbd22927d),
	.w7(32'hbce23723),
	.w8(32'hbbf8e967),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60ddee),
	.w1(32'hba4276ed),
	.w2(32'h3bab6bb9),
	.w3(32'hbc01c7d9),
	.w4(32'hbb93c38b),
	.w5(32'h3b83317b),
	.w6(32'hbc08b688),
	.w7(32'hbc0994b1),
	.w8(32'h3a9cfa6a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803f5d),
	.w1(32'hbb54ab8d),
	.w2(32'h3bbf2845),
	.w3(32'hbbb40c62),
	.w4(32'hbba5e2ba),
	.w5(32'h3c1eaf33),
	.w6(32'hbbcc1978),
	.w7(32'hbb7fb053),
	.w8(32'h3c576d41),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c95d5),
	.w1(32'h3b98f550),
	.w2(32'h3c08de4f),
	.w3(32'h3c4d2248),
	.w4(32'h3b206c09),
	.w5(32'h3bbe2ffb),
	.w6(32'h3c28df94),
	.w7(32'h3c3544af),
	.w8(32'h3b6f590f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55ed26),
	.w1(32'h3bf4a10b),
	.w2(32'h3a85c111),
	.w3(32'hbbe9fe68),
	.w4(32'hbbf5d123),
	.w5(32'hbaa0df99),
	.w6(32'hbc879399),
	.w7(32'hbc612efb),
	.w8(32'hb6e7e2d1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb40c49),
	.w1(32'h3bdde3c1),
	.w2(32'hba66f6fe),
	.w3(32'hbc1d47d8),
	.w4(32'h3b90a4e4),
	.w5(32'hbca9379f),
	.w6(32'hbc514b83),
	.w7(32'hbb01ce3d),
	.w8(32'hbc7f33f4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca23afb),
	.w1(32'h3d1cb804),
	.w2(32'h3c0fe3e5),
	.w3(32'h3bd6ecec),
	.w4(32'h3d22485b),
	.w5(32'h3b096c78),
	.w6(32'h3b52f3a3),
	.w7(32'h3cde76a6),
	.w8(32'h3b5989f7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc164dad),
	.w1(32'hbc5bb312),
	.w2(32'h3a6d177c),
	.w3(32'hbc47a29c),
	.w4(32'hbc8da98e),
	.w5(32'hbaac8fcf),
	.w6(32'hbbc0934b),
	.w7(32'hbc4d71ee),
	.w8(32'hb927e1dd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1674d),
	.w1(32'h3ba5fa1a),
	.w2(32'hbc04ebc5),
	.w3(32'hb6e36b00),
	.w4(32'h3b702d21),
	.w5(32'h3afd20a2),
	.w6(32'h3b7ac97e),
	.w7(32'h3bda99dd),
	.w8(32'hbac5c51f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0c38e),
	.w1(32'hbbc7621b),
	.w2(32'hbc20eb03),
	.w3(32'hbb46cbad),
	.w4(32'h3b2e74ad),
	.w5(32'hbc9ec29e),
	.w6(32'h3966a050),
	.w7(32'hba89c5ec),
	.w8(32'hbbce1654),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187591),
	.w1(32'hbb39f378),
	.w2(32'h3b48fe62),
	.w3(32'hbc88a94a),
	.w4(32'hbc3d6704),
	.w5(32'h3c9b73b6),
	.w6(32'hbc1ef6d0),
	.w7(32'h3bae4ce0),
	.w8(32'h3b23aab9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0984fd),
	.w1(32'hbc2d6b1e),
	.w2(32'h3be2905b),
	.w3(32'h3c00fc68),
	.w4(32'hbc85d807),
	.w5(32'h3c2d394c),
	.w6(32'hbb4a271d),
	.w7(32'hbc40705b),
	.w8(32'h3c589588),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63811b),
	.w1(32'h3b8ad316),
	.w2(32'h3c404bb5),
	.w3(32'h3c9b5673),
	.w4(32'h3c0bd9e8),
	.w5(32'h3cb2776d),
	.w6(32'h3c099f30),
	.w7(32'h3c18c2f0),
	.w8(32'h3ca04f01),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f0444),
	.w1(32'h3c3932c4),
	.w2(32'hbbaf5b53),
	.w3(32'h3c0d4753),
	.w4(32'h3bd6c2c1),
	.w5(32'hbc3197d7),
	.w6(32'h3bed29f1),
	.w7(32'hbb0f1bec),
	.w8(32'hbc66cc1f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00a5dd),
	.w1(32'h3b7498a8),
	.w2(32'h3bbfbc43),
	.w3(32'h3bf70441),
	.w4(32'h3c04443c),
	.w5(32'h3bfd8973),
	.w6(32'h3bfa67f8),
	.w7(32'h3c375a29),
	.w8(32'h3c4f6cb4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aa065),
	.w1(32'hbb9190a6),
	.w2(32'h3c20f799),
	.w3(32'h3b14f6d5),
	.w4(32'h3bfd7bc9),
	.w5(32'h3c728cad),
	.w6(32'h3c3e79f0),
	.w7(32'h3bcba24c),
	.w8(32'h3c302ab4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b670600),
	.w1(32'h397c5866),
	.w2(32'h3b4af08b),
	.w3(32'h3bce3faf),
	.w4(32'hbb0f6387),
	.w5(32'h3c0ae26c),
	.w6(32'h3be293e7),
	.w7(32'h3b55ba0a),
	.w8(32'h3bf0c9a3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43503b),
	.w1(32'h3b130f3a),
	.w2(32'hb8a3411d),
	.w3(32'h3b5f00d6),
	.w4(32'hba0872d8),
	.w5(32'h39c1656d),
	.w6(32'hbc013cf1),
	.w7(32'hbc332c90),
	.w8(32'h3b033e49),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a367a01),
	.w1(32'hb9857459),
	.w2(32'h3c5961c6),
	.w3(32'h3b029299),
	.w4(32'hbb8d61ed),
	.w5(32'h3c08b3ef),
	.w6(32'hbbd99414),
	.w7(32'hbc2cc6ab),
	.w8(32'h3c017183),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c01e4),
	.w1(32'hbcafe470),
	.w2(32'h3b60d557),
	.w3(32'hbc81624d),
	.w4(32'hbc9fd9e0),
	.w5(32'h3c777837),
	.w6(32'hbba80fa6),
	.w7(32'hbc0caf89),
	.w8(32'h3c716e46),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7533c14),
	.w1(32'hbab95655),
	.w2(32'h3a18738f),
	.w3(32'h3b1251af),
	.w4(32'hbbc206ff),
	.w5(32'h3ba47e4e),
	.w6(32'h3a43c782),
	.w7(32'hbbacfa0e),
	.w8(32'h3bf6c9b9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bc575),
	.w1(32'hbc9823c6),
	.w2(32'h3bc9bf08),
	.w3(32'hbcc5fce9),
	.w4(32'hbcd3340d),
	.w5(32'h3c195971),
	.w6(32'hbc6ba757),
	.w7(32'hbc86b2e9),
	.w8(32'h3b1f03f5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b3f1),
	.w1(32'hbc8e8e27),
	.w2(32'h3bd5f85b),
	.w3(32'hbadb0ce6),
	.w4(32'hbc76c62a),
	.w5(32'h3c4505aa),
	.w6(32'hb93484a1),
	.w7(32'hbc17dd98),
	.w8(32'h3c039dcb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7065c8),
	.w1(32'h3b0bb5a6),
	.w2(32'h3bb008bb),
	.w3(32'h3bc9af68),
	.w4(32'hbc2ea6ca),
	.w5(32'h3c47035b),
	.w6(32'h3bbdf7e8),
	.w7(32'hbc217965),
	.w8(32'h3c7b4d59),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad03b1b),
	.w1(32'hbaf3a011),
	.w2(32'h3b207715),
	.w3(32'h3c275af9),
	.w4(32'h3aea1de1),
	.w5(32'hba2fa24e),
	.w6(32'h3c816078),
	.w7(32'h3bec11ce),
	.w8(32'h3a9ee150),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe21c8c),
	.w1(32'hbbabdd09),
	.w2(32'h3b914e84),
	.w3(32'h3be86b9c),
	.w4(32'hbae9efaf),
	.w5(32'h3b8582c5),
	.w6(32'h3a88c870),
	.w7(32'h3b1ee0c4),
	.w8(32'h3b97c5b5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf81cb),
	.w1(32'hbbd86fa8),
	.w2(32'hbb485cac),
	.w3(32'hbc7cfe97),
	.w4(32'hbc9d7a80),
	.w5(32'h3bb6c22b),
	.w6(32'hbbce4ab7),
	.w7(32'hbc4f55d0),
	.w8(32'h3c06b7dd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030629),
	.w1(32'hbc917d40),
	.w2(32'h3c5262b1),
	.w3(32'h37c7183f),
	.w4(32'hbcb7dbc8),
	.w5(32'h3cbab923),
	.w6(32'hbb8be22d),
	.w7(32'hbc1496fc),
	.w8(32'h3c826ac4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390930dc),
	.w1(32'h3a0661be),
	.w2(32'h3aca0e35),
	.w3(32'h3b8393a1),
	.w4(32'hbbd8b889),
	.w5(32'h38d75831),
	.w6(32'h3c5d3b32),
	.w7(32'h3c3fd741),
	.w8(32'hb9bed11d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46860),
	.w1(32'h3b23bed9),
	.w2(32'h3bd0c405),
	.w3(32'h3ae4a1f0),
	.w4(32'hbc09e222),
	.w5(32'h3b5f8bb5),
	.w6(32'hba9d4f9a),
	.w7(32'hbbe0357a),
	.w8(32'hbb2367d1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad994dc),
	.w1(32'h3b816cf0),
	.w2(32'hbb75a3fe),
	.w3(32'h3be33b04),
	.w4(32'h3c0fbb6c),
	.w5(32'hb6fc9411),
	.w6(32'h3b90cf7e),
	.w7(32'h3c1c2498),
	.w8(32'h3b87c5b2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fdbee),
	.w1(32'h3a59fd6c),
	.w2(32'h3c00b8cc),
	.w3(32'hbb186123),
	.w4(32'h3a9d3b50),
	.w5(32'h3c0420f8),
	.w6(32'h3bc19e08),
	.w7(32'h3b4fac46),
	.w8(32'h3a6ecff5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba05b52),
	.w1(32'h39eac11d),
	.w2(32'h3c8465fd),
	.w3(32'h3bd7f249),
	.w4(32'h3b1d5e55),
	.w5(32'h3ce56440),
	.w6(32'hb975f1fe),
	.w7(32'hbb0506ba),
	.w8(32'h3c2b911e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c268e69),
	.w1(32'h3acf629c),
	.w2(32'h3bf4bd07),
	.w3(32'h3c55ae6c),
	.w4(32'hbb94405e),
	.w5(32'h3bd00926),
	.w6(32'h3bbda221),
	.w7(32'hba99de99),
	.w8(32'h3c261854),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9030a2),
	.w1(32'hbc379b6b),
	.w2(32'hbc2487e7),
	.w3(32'h3c042451),
	.w4(32'hb811a89c),
	.w5(32'hbb1b3e6f),
	.w6(32'h3c30e347),
	.w7(32'h3c0bccef),
	.w8(32'hbba812fc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1772a7),
	.w1(32'hbbeccd08),
	.w2(32'hbb7deb73),
	.w3(32'h3ae99a7c),
	.w4(32'hbbe0cbac),
	.w5(32'hbb95a3ca),
	.w6(32'hbbb6adf5),
	.w7(32'h3a559323),
	.w8(32'hbbbcaba3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5db12a),
	.w1(32'h3a3ef0b1),
	.w2(32'h3b9ece08),
	.w3(32'hbbb201e2),
	.w4(32'h3ad46aa1),
	.w5(32'h3c1cad98),
	.w6(32'hbbc0d005),
	.w7(32'hba33aebe),
	.w8(32'h3c1308db),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d310a),
	.w1(32'hbba7a962),
	.w2(32'h3c552dff),
	.w3(32'h3b86f993),
	.w4(32'hbbb8050a),
	.w5(32'h3d1e475a),
	.w6(32'h3b34bbc8),
	.w7(32'hbb842781),
	.w8(32'h3d0f3433),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b2a7),
	.w1(32'hbb0eccc7),
	.w2(32'hbbeb166e),
	.w3(32'h3d073c3b),
	.w4(32'hbc47dadd),
	.w5(32'hbba6f7ac),
	.w6(32'h3cc78277),
	.w7(32'hbb83ce3f),
	.w8(32'hba8c933a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473978),
	.w1(32'hbba08c64),
	.w2(32'h3c790943),
	.w3(32'hbc07be08),
	.w4(32'h3a082f99),
	.w5(32'h3ce0cf06),
	.w6(32'hbb5691ea),
	.w7(32'h3b1090fc),
	.w8(32'h3c98296d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba715ae),
	.w1(32'h3aa8caac),
	.w2(32'h3c0f1fef),
	.w3(32'h3be7214f),
	.w4(32'hbbc9926b),
	.w5(32'h3b48f27c),
	.w6(32'h3c383db4),
	.w7(32'h3bfb22b3),
	.w8(32'h3c124c5e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b516ec2),
	.w1(32'hbc4a55e8),
	.w2(32'hbb35f723),
	.w3(32'hbbb281f2),
	.w4(32'hbca75c6d),
	.w5(32'hb9d6bd8d),
	.w6(32'hbc0b1fec),
	.w7(32'hbc044407),
	.w8(32'h3b5999f8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b8aa3),
	.w1(32'hbc933fef),
	.w2(32'hbc37de5d),
	.w3(32'hbc9a736d),
	.w4(32'hbcda9cf0),
	.w5(32'h3a318d22),
	.w6(32'hbc7c88f9),
	.w7(32'hbc875814),
	.w8(32'h3a75dd2d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule