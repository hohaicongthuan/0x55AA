module layer_10_featuremap_87(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39470c1c),
	.w1(32'h3b489186),
	.w2(32'h38285b96),
	.w3(32'hba275f8c),
	.w4(32'h389fbcbd),
	.w5(32'h3b047794),
	.w6(32'hbd059e74),
	.w7(32'hbae369c4),
	.w8(32'h3aa910f7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd116629),
	.w1(32'hba1acc81),
	.w2(32'h3be6f7d4),
	.w3(32'hbb935876),
	.w4(32'hbac9177b),
	.w5(32'h3ba21831),
	.w6(32'h3b803310),
	.w7(32'h3b5a6c53),
	.w8(32'h3c259011),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77a8d),
	.w1(32'hbad668a5),
	.w2(32'hbaab3031),
	.w3(32'h3b202afb),
	.w4(32'h3a8993df),
	.w5(32'h3a8dbcb4),
	.w6(32'h3a847dc7),
	.w7(32'hba4c95d7),
	.w8(32'h3a39f2e5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0d9d6),
	.w1(32'h392d3f9d),
	.w2(32'h3a959a34),
	.w3(32'hbb076952),
	.w4(32'h3ab32183),
	.w5(32'hba7564b6),
	.w6(32'hba57025c),
	.w7(32'hbb206629),
	.w8(32'h3ac6dbe5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a3a3f),
	.w1(32'hbb630dcd),
	.w2(32'h395bebfc),
	.w3(32'hbb2ce95c),
	.w4(32'hba32ca37),
	.w5(32'hb7ac5815),
	.w6(32'hbae77416),
	.w7(32'h390b8370),
	.w8(32'hbc414b95),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82fa5a),
	.w1(32'hba1a166a),
	.w2(32'hba18dc6c),
	.w3(32'hba1ce4f2),
	.w4(32'hbb11d448),
	.w5(32'h3a3dbc0e),
	.w6(32'hbc21b6ed),
	.w7(32'hb8be5b80),
	.w8(32'h39fe1169),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf09ea6),
	.w1(32'hbbc16b8e),
	.w2(32'hbc9811eb),
	.w3(32'h3c363271),
	.w4(32'h3c12ef30),
	.w5(32'hbc3aca2b),
	.w6(32'h3bf8de64),
	.w7(32'hbb8928ea),
	.w8(32'hbbcdb11b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931994),
	.w1(32'h3c5d6623),
	.w2(32'hbbbdc75a),
	.w3(32'h3baa54ef),
	.w4(32'h3cab4d50),
	.w5(32'h3c24c63b),
	.w6(32'h3b9b6560),
	.w7(32'hbca39a6b),
	.w8(32'h3b1fecc6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc323505),
	.w1(32'h3c314cd8),
	.w2(32'hbb2cb43c),
	.w3(32'h3b82c06c),
	.w4(32'hb967ffc6),
	.w5(32'h3b00e1c9),
	.w6(32'h3b05ea31),
	.w7(32'hb91ddf4c),
	.w8(32'h393177ac),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2518),
	.w1(32'hbb9177ff),
	.w2(32'hbc0f1386),
	.w3(32'h3be4df1d),
	.w4(32'hbb49548e),
	.w5(32'hbbf31868),
	.w6(32'h3aee36ef),
	.w7(32'hbc0d2878),
	.w8(32'hbbc7acf0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ebf7d),
	.w1(32'hbab745fb),
	.w2(32'h39c6a80b),
	.w3(32'h3b1c3824),
	.w4(32'h3c565025),
	.w5(32'hbd2d02d5),
	.w6(32'h3b8dea7b),
	.w7(32'hb953c029),
	.w8(32'hb989c9e9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd36f3),
	.w1(32'hbbd6888f),
	.w2(32'hbd009c68),
	.w3(32'h3c194e98),
	.w4(32'hbac7ae38),
	.w5(32'hbc9a4974),
	.w6(32'h3c22e889),
	.w7(32'h3a5be52d),
	.w8(32'hbc878fce),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbad675),
	.w1(32'hbb8f102a),
	.w2(32'hbbfc49af),
	.w3(32'h3c1bbe74),
	.w4(32'hb97070d4),
	.w5(32'hbc0782f8),
	.w6(32'h3a03b5e1),
	.w7(32'hbbf6a263),
	.w8(32'hbc8fb6bf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccdc84),
	.w1(32'hbc00d9e1),
	.w2(32'hb9837df8),
	.w3(32'h3b894d6c),
	.w4(32'h3be7d61a),
	.w5(32'h3b859797),
	.w6(32'hba124ef6),
	.w7(32'h3d092b04),
	.w8(32'h3a20b8c3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22568c),
	.w1(32'hbaeb3803),
	.w2(32'h3ac8b528),
	.w3(32'hbb2cc7e6),
	.w4(32'h3a9b876e),
	.w5(32'h3b65bb18),
	.w6(32'h3ba296ab),
	.w7(32'h3bbfd80b),
	.w8(32'h3b813485),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194c30),
	.w1(32'h3b13070a),
	.w2(32'h3c733c8c),
	.w3(32'hbb134b07),
	.w4(32'h3ab0233b),
	.w5(32'h3c0673b7),
	.w6(32'hbb34dd3e),
	.w7(32'hbb25a1b8),
	.w8(32'h3c936aa6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42f47f),
	.w1(32'h3d023f89),
	.w2(32'h3aecef83),
	.w3(32'hba8df3b1),
	.w4(32'h397ef2bd),
	.w5(32'hbc2b6d2c),
	.w6(32'hba287ecc),
	.w7(32'h3a05b3cc),
	.w8(32'h3b37f834),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc62069),
	.w1(32'hbd02e669),
	.w2(32'hbcddc855),
	.w3(32'h3bf34926),
	.w4(32'h3a98fecd),
	.w5(32'hbc4e2f62),
	.w6(32'hbc93fe5e),
	.w7(32'hbd33a2c2),
	.w8(32'hbcd29d29),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b35c5),
	.w1(32'hbc9a11b5),
	.w2(32'hbc00355a),
	.w3(32'h3bcc9dc5),
	.w4(32'hba55c0c5),
	.w5(32'hbb0471ae),
	.w6(32'hbc005eca),
	.w7(32'hbc651524),
	.w8(32'hbc7e6388),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff0dbf),
	.w1(32'hb9f620e2),
	.w2(32'h3b9dba8a),
	.w3(32'h3ae78ac8),
	.w4(32'h3bab1a7c),
	.w5(32'h3aed208b),
	.w6(32'h3a361a8f),
	.w7(32'hbad5a35e),
	.w8(32'hb9a00ef5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b50b),
	.w1(32'hb984a73b),
	.w2(32'h3bab54a2),
	.w3(32'hb98019b9),
	.w4(32'h3b0844a1),
	.w5(32'h3ad60c28),
	.w6(32'hbbe54e8e),
	.w7(32'h3a5ba84f),
	.w8(32'h3b9d9697),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132ece),
	.w1(32'h3a85d5a2),
	.w2(32'h3a90db2e),
	.w3(32'hba0c4159),
	.w4(32'h394104d1),
	.w5(32'h3a8a9cac),
	.w6(32'h3af18eae),
	.w7(32'h3b4f2a81),
	.w8(32'h3b89e904),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc31a6d),
	.w1(32'h3c96bb5e),
	.w2(32'hbc4919d3),
	.w3(32'h3cd5737e),
	.w4(32'h3bc3face),
	.w5(32'hbc5b95a8),
	.w6(32'hbba699ef),
	.w7(32'hbbe2b0db),
	.w8(32'hbd02833f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1f73),
	.w1(32'h3ae3b541),
	.w2(32'hb985faa3),
	.w3(32'h3b9b3e3c),
	.w4(32'h39c42136),
	.w5(32'h38ec38a1),
	.w6(32'h39d1298e),
	.w7(32'hbb6bf735),
	.w8(32'hbb960cb5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0253d4),
	.w1(32'hbb569c38),
	.w2(32'h3c4e8bc4),
	.w3(32'hbbe852a5),
	.w4(32'h3c08b6d0),
	.w5(32'h3c52add6),
	.w6(32'h3b8717d3),
	.w7(32'h3bfa0b8b),
	.w8(32'h3c97f0da),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a039f),
	.w1(32'h3b1c09ea),
	.w2(32'h3ad7c9df),
	.w3(32'hbb7cf859),
	.w4(32'h3bc4e1f2),
	.w5(32'h3b3f6774),
	.w6(32'h3beb7d64),
	.w7(32'h3aa44083),
	.w8(32'h3ab8263b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c58e9),
	.w1(32'h3b0df29e),
	.w2(32'h3b1ee5d2),
	.w3(32'hbb3bac2c),
	.w4(32'hbad61b6e),
	.w5(32'h3a456cd6),
	.w6(32'h3b4cd059),
	.w7(32'h3adb3378),
	.w8(32'h397353d5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d189c),
	.w1(32'hbca6995e),
	.w2(32'hbb3b9289),
	.w3(32'h3c8a6a66),
	.w4(32'hbc9f14a8),
	.w5(32'hbd350270),
	.w6(32'h3c9fb91c),
	.w7(32'h3ca4bd97),
	.w8(32'h3c5f4f13),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5b4e7),
	.w1(32'hbb5d1ccc),
	.w2(32'h3d0adf72),
	.w3(32'hba1c6934),
	.w4(32'h3b2e6aee),
	.w5(32'h3a22f066),
	.w6(32'h3c0af281),
	.w7(32'hbaa04b96),
	.w8(32'h3b51e227),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcf49c),
	.w1(32'hbc1d599c),
	.w2(32'h3b8255e7),
	.w3(32'h36d99940),
	.w4(32'h3c916a0f),
	.w5(32'hbc2992ee),
	.w6(32'h3ca8ad3c),
	.w7(32'h3b32296c),
	.w8(32'h3bceb557),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bfcb5),
	.w1(32'h3b5fbcb8),
	.w2(32'hbb549655),
	.w3(32'hba6fbcac),
	.w4(32'h3accf820),
	.w5(32'hbaa7c8b5),
	.w6(32'hbb95d8ca),
	.w7(32'h3aae63a5),
	.w8(32'h3bccfaaf),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ec08e),
	.w1(32'h3bae98ea),
	.w2(32'hbb4d27c7),
	.w3(32'h3a188901),
	.w4(32'h3bc14716),
	.w5(32'h3b915c40),
	.w6(32'h3b84f89a),
	.w7(32'hbc18c29c),
	.w8(32'hbb674589),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c858a),
	.w1(32'h3bbf04d8),
	.w2(32'hba4dda4c),
	.w3(32'hb976b50f),
	.w4(32'h3b939cf2),
	.w5(32'hbb01e6f7),
	.w6(32'h3ab78c57),
	.w7(32'hba8122d3),
	.w8(32'hbb3c5c38),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144951),
	.w1(32'h3c9cabd0),
	.w2(32'h3af56bd8),
	.w3(32'hbb739e5a),
	.w4(32'h3b53d783),
	.w5(32'h3bd12b9b),
	.w6(32'h394fe9ab),
	.w7(32'h3c1cb068),
	.w8(32'h3be9ea2d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2101bf),
	.w1(32'h3a8ba356),
	.w2(32'h3b45eced),
	.w3(32'h3946f1f8),
	.w4(32'hbb49d5a7),
	.w5(32'hbbb3dcf3),
	.w6(32'h3ae8fef5),
	.w7(32'hbc0063f3),
	.w8(32'hbbd3cc4a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c048d87),
	.w1(32'hba606a4e),
	.w2(32'hbc71bcd2),
	.w3(32'h3be49ddf),
	.w4(32'h3c22594f),
	.w5(32'h3bad0793),
	.w6(32'hba29abc6),
	.w7(32'hba6dedb2),
	.w8(32'hbc3d578f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03601),
	.w1(32'h3cbedd60),
	.w2(32'h3c1f1b24),
	.w3(32'h3cbba075),
	.w4(32'h3d315891),
	.w5(32'hba8d9f15),
	.w6(32'h3cb46f72),
	.w7(32'h3d143872),
	.w8(32'h3bfb594f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863b0a),
	.w1(32'hbc52dd69),
	.w2(32'h3c417c38),
	.w3(32'hbbefcbe6),
	.w4(32'hbbb4928d),
	.w5(32'hbb8dcd9b),
	.w6(32'h3b14e050),
	.w7(32'h3bee0ee0),
	.w8(32'h3caeb3e2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbac35f),
	.w1(32'hbc867907),
	.w2(32'hbc245d23),
	.w3(32'hbb766fc5),
	.w4(32'hbccb67e9),
	.w5(32'hbcafc63c),
	.w6(32'h3bfa31f9),
	.w7(32'hbb976cd1),
	.w8(32'h3c173088),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2770c),
	.w1(32'h398db37a),
	.w2(32'hb920da20),
	.w3(32'h38e2ac4b),
	.w4(32'h3c87798f),
	.w5(32'h3acec7c1),
	.w6(32'h3ca71cd4),
	.w7(32'h3bb9b761),
	.w8(32'h3b6671f3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b15f59),
	.w1(32'hbb2029c2),
	.w2(32'hbb981c41),
	.w3(32'h3b73554c),
	.w4(32'h390458c4),
	.w5(32'hba04fc33),
	.w6(32'hb993dd99),
	.w7(32'hbad3be0c),
	.w8(32'hbae4c71c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f97b),
	.w1(32'hbadca3c7),
	.w2(32'h3a512646),
	.w3(32'hbb905dac),
	.w4(32'hbb6e9a71),
	.w5(32'hb9945a59),
	.w6(32'hbbe9e197),
	.w7(32'hbbe291c0),
	.w8(32'hbb6618b7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7073e1),
	.w1(32'h3b89a9b9),
	.w2(32'h3a2565dd),
	.w3(32'h3a678e57),
	.w4(32'hbc4cb880),
	.w5(32'hbb26b719),
	.w6(32'h3b13d85d),
	.w7(32'h3af4868d),
	.w8(32'h3b492d37),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d49ab),
	.w1(32'hba8d65b7),
	.w2(32'hbb5193b1),
	.w3(32'h3bc01001),
	.w4(32'hbbb3096d),
	.w5(32'hbc0ce883),
	.w6(32'hbc49e634),
	.w7(32'hbcf35627),
	.w8(32'hbcd67c95),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39807093),
	.w1(32'h3c2f2696),
	.w2(32'h3c3cd86d),
	.w3(32'h3b515c2c),
	.w4(32'h3b960c2f),
	.w5(32'h3b01f3eb),
	.w6(32'h3b438180),
	.w7(32'h3b8b5731),
	.w8(32'h3b1c2031),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff7b6b),
	.w1(32'h3adb98cf),
	.w2(32'hbbe5e72e),
	.w3(32'h3bc4f059),
	.w4(32'hbae806d4),
	.w5(32'hbae4003c),
	.w6(32'h3c4897d9),
	.w7(32'h3adad7c8),
	.w8(32'hbc074eb4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9665a0),
	.w1(32'hb9758c8a),
	.w2(32'hbae717cb),
	.w3(32'h3cdc63c0),
	.w4(32'h3ad226dd),
	.w5(32'h3b4e46f9),
	.w6(32'h3a9a5e00),
	.w7(32'h3c207d74),
	.w8(32'h3b1557a6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce2b387),
	.w1(32'h3c2bde3f),
	.w2(32'hbb957315),
	.w3(32'h3ca78c26),
	.w4(32'h3c8fc7c3),
	.w5(32'hbc43cd66),
	.w6(32'hbcc01598),
	.w7(32'hbcfd57b9),
	.w8(32'hbd26312f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db9614),
	.w1(32'h3b479765),
	.w2(32'hbc2d0e4f),
	.w3(32'hbb9157be),
	.w4(32'h3b8c1c8b),
	.w5(32'hb9cae8fc),
	.w6(32'h3aaf0f91),
	.w7(32'hba9913e3),
	.w8(32'hbb6912e8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb968882),
	.w1(32'h3b680936),
	.w2(32'hba5289e8),
	.w3(32'hbba3f964),
	.w4(32'h3b8fa37e),
	.w5(32'hba63d697),
	.w6(32'hba4e7999),
	.w7(32'hba877488),
	.w8(32'hbaf47f8e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a127f21),
	.w1(32'h3b5831ca),
	.w2(32'h38d11f1c),
	.w3(32'h3a3b5ee8),
	.w4(32'h3a6dbfc7),
	.w5(32'hb83c871f),
	.w6(32'hb95ba591),
	.w7(32'h3b02ef67),
	.w8(32'hbaf01f31),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c608),
	.w1(32'h3b623a43),
	.w2(32'hbafe663f),
	.w3(32'h3d12b6fd),
	.w4(32'hbac4a83e),
	.w5(32'h3b106e8d),
	.w6(32'hbc262398),
	.w7(32'hb928c3c9),
	.w8(32'hb840c9ae),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf94729),
	.w1(32'h3bbf114e),
	.w2(32'hbad4ab0c),
	.w3(32'hbab9a696),
	.w4(32'hbbf55941),
	.w5(32'hbac15852),
	.w6(32'h3a7c9c96),
	.w7(32'h3b047d3c),
	.w8(32'hbb2952d1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c203b30),
	.w1(32'h3af9a13a),
	.w2(32'hbc66b932),
	.w3(32'h3c6a6e24),
	.w4(32'h3c385d0d),
	.w5(32'hbc10afcb),
	.w6(32'hbc1001ce),
	.w7(32'hbcae096d),
	.w8(32'hbcec9744),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c2b71),
	.w1(32'h3ab8cd94),
	.w2(32'hba9f6bd7),
	.w3(32'hbb60fd4f),
	.w4(32'h395badce),
	.w5(32'hbb8838c0),
	.w6(32'h3b040146),
	.w7(32'hbc054479),
	.w8(32'hb9eb7570),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0a767),
	.w1(32'hbb6eabb6),
	.w2(32'hb9304f28),
	.w3(32'h3ad9553e),
	.w4(32'hbb826972),
	.w5(32'h3c691727),
	.w6(32'hb9aa5822),
	.w7(32'h3b61641f),
	.w8(32'hb9998f4f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3cded),
	.w1(32'hbb151da4),
	.w2(32'hbb30fbab),
	.w3(32'hbbdc561f),
	.w4(32'hbac34d4e),
	.w5(32'hbae40855),
	.w6(32'h3cb7bef9),
	.w7(32'hbb85473e),
	.w8(32'hbb127913),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b393a5b),
	.w1(32'h3b67ddd2),
	.w2(32'h3b492f93),
	.w3(32'hbbec46bc),
	.w4(32'h3b117871),
	.w5(32'hbb21ce82),
	.w6(32'h39d10052),
	.w7(32'h3a240daf),
	.w8(32'h3bc49b3b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b335f3e),
	.w1(32'hbc0863b1),
	.w2(32'h3b81be4b),
	.w3(32'hbb74433d),
	.w4(32'h3c2e5bce),
	.w5(32'h3bebed89),
	.w6(32'hbae6e9b1),
	.w7(32'hba5c4ee1),
	.w8(32'h3abb08fe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c74f0),
	.w1(32'h3a2813d2),
	.w2(32'hbb1c481e),
	.w3(32'h3b516860),
	.w4(32'hbb1b9f2d),
	.w5(32'hbbd33b42),
	.w6(32'h3b1a4535),
	.w7(32'hbb3b3a99),
	.w8(32'h3b80415c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8675cc),
	.w1(32'h3b10b20a),
	.w2(32'h3b81bf12),
	.w3(32'h3b962cb4),
	.w4(32'h3b22d0a1),
	.w5(32'hba9d3b99),
	.w6(32'hbc8765ec),
	.w7(32'hbc116f3b),
	.w8(32'hbc501927),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855184),
	.w1(32'hbb011a67),
	.w2(32'h3aa7aa50),
	.w3(32'hbb4d4871),
	.w4(32'hbae47b46),
	.w5(32'hbbe31a06),
	.w6(32'hbb4fc940),
	.w7(32'hbb49b844),
	.w8(32'h3b2014f7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ff3e),
	.w1(32'hbb94b860),
	.w2(32'hbb6187dd),
	.w3(32'h3c93a092),
	.w4(32'h3b42b66f),
	.w5(32'h3a921a73),
	.w6(32'hbb461bf5),
	.w7(32'h3b1a13ae),
	.w8(32'h3b45fc15),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62eac6),
	.w1(32'hbb0110cd),
	.w2(32'h3c37f128),
	.w3(32'hbb6879f0),
	.w4(32'h3ad63c46),
	.w5(32'hbc0f47fd),
	.w6(32'h3b210692),
	.w7(32'h3ba50037),
	.w8(32'hbc1818f3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab7f3b),
	.w1(32'h3ad6ca01),
	.w2(32'h3b1004a5),
	.w3(32'hbb99e7dd),
	.w4(32'hbaa16e8d),
	.w5(32'h3b97e9cc),
	.w6(32'hbc2d9bc7),
	.w7(32'h3cdd708f),
	.w8(32'h3b1029ab),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4c995),
	.w1(32'hbb07478f),
	.w2(32'h3a86e4c4),
	.w3(32'h3a423bd2),
	.w4(32'hbb4146ac),
	.w5(32'hb43a7bfd),
	.w6(32'h3c299da1),
	.w7(32'h3d8e9e57),
	.w8(32'h3b46d66c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba969cc8),
	.w1(32'h3b650d3b),
	.w2(32'hbc0ebb3c),
	.w3(32'h3cac81da),
	.w4(32'hbbaa4784),
	.w5(32'hbcefabaf),
	.w6(32'h3cab3f7e),
	.w7(32'h3b129b4c),
	.w8(32'h3c1e36e6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c414049),
	.w1(32'hbc80deed),
	.w2(32'hbcaab2a8),
	.w3(32'h3bee43d9),
	.w4(32'hbb71613e),
	.w5(32'hbc3417bf),
	.w6(32'h3c2b0b95),
	.w7(32'hbc8d5a10),
	.w8(32'hbd294af7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf7cc7),
	.w1(32'hb8624912),
	.w2(32'hbb55eb21),
	.w3(32'h3adc40e8),
	.w4(32'hbb301d89),
	.w5(32'hbb169fe7),
	.w6(32'hbc4f4ec8),
	.w7(32'hbc9d7588),
	.w8(32'hbc98c28f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84fbb2),
	.w1(32'hbc3dbbb6),
	.w2(32'hbb050491),
	.w3(32'hbc44a9b0),
	.w4(32'hbb5c4e2e),
	.w5(32'h3ae976ca),
	.w6(32'hbaf35bdc),
	.w7(32'hba5d6370),
	.w8(32'h3c4fde73),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5621dd),
	.w1(32'hbb3d12c7),
	.w2(32'h3732b450),
	.w3(32'h3ac15b4e),
	.w4(32'hbbbbbfb3),
	.w5(32'h3a33856b),
	.w6(32'hbb48975b),
	.w7(32'h3b811d83),
	.w8(32'h3badbdf5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acf47d),
	.w1(32'h3beea398),
	.w2(32'hbad1ccdb),
	.w3(32'hbb36f7dd),
	.w4(32'h3b02ccfa),
	.w5(32'h3abb9efe),
	.w6(32'h3b0fc1d7),
	.w7(32'hbaf56b22),
	.w8(32'hbb992fad),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc892a),
	.w1(32'h3b13e2ef),
	.w2(32'h3b8ab0d0),
	.w3(32'h3ba442fb),
	.w4(32'h3b8b963c),
	.w5(32'hbbe3278a),
	.w6(32'hb9c38525),
	.w7(32'hbac62d66),
	.w8(32'h3a659c38),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b554de8),
	.w1(32'h3aa486e1),
	.w2(32'hbc87bf80),
	.w3(32'h39f1d845),
	.w4(32'h3b578cb8),
	.w5(32'hbb1a0c1c),
	.w6(32'h3bbec30f),
	.w7(32'hbc12ec0c),
	.w8(32'hbbd44279),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf29863),
	.w1(32'hba787ed5),
	.w2(32'hb85d101d),
	.w3(32'h3b4cbbcc),
	.w4(32'h3b88bfbe),
	.w5(32'hbb606907),
	.w6(32'h3caa133c),
	.w7(32'hbb9683bd),
	.w8(32'hbb9ceb47),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf696),
	.w1(32'h3bc4c257),
	.w2(32'hbc1bb914),
	.w3(32'hba132e2f),
	.w4(32'h3b5801e7),
	.w5(32'hbb70a341),
	.w6(32'h3b5cbafd),
	.w7(32'hbbc3c6c2),
	.w8(32'hb8dd00d8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e583e),
	.w1(32'hbb2a70b4),
	.w2(32'h3977f007),
	.w3(32'h3c2bd7b5),
	.w4(32'h3bbc8e77),
	.w5(32'hbae6df7a),
	.w6(32'h3ba3b76a),
	.w7(32'hbc377b04),
	.w8(32'hbcab9d65),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf07a5),
	.w1(32'hbc2cb793),
	.w2(32'hbb3be814),
	.w3(32'h3c84afa2),
	.w4(32'h3bd77c75),
	.w5(32'h3be966c6),
	.w6(32'h3becede4),
	.w7(32'hbb3b8188),
	.w8(32'h3c5806c9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2b9bc),
	.w1(32'h3b607bde),
	.w2(32'h3b059a7b),
	.w3(32'h3b8ae929),
	.w4(32'h3a493e72),
	.w5(32'hbb7accad),
	.w6(32'h3a87ec59),
	.w7(32'hb9c79218),
	.w8(32'hba18b326),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69c4d5),
	.w1(32'hbb5c0d39),
	.w2(32'hbc0cd14d),
	.w3(32'h3ba5a54b),
	.w4(32'hbadb9406),
	.w5(32'hbcb3b4b3),
	.w6(32'h3c0ba6b7),
	.w7(32'hbb072608),
	.w8(32'h3c12c0a2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2850b),
	.w1(32'h3a231b46),
	.w2(32'hba04c971),
	.w3(32'h3ab84323),
	.w4(32'h3bf0e46c),
	.w5(32'hb9ecd7bd),
	.w6(32'hbc574fa0),
	.w7(32'h3ba4f925),
	.w8(32'hbb310712),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba31ae9),
	.w1(32'h3bd93af4),
	.w2(32'hbae4920e),
	.w3(32'h3c2063af),
	.w4(32'hba470e72),
	.w5(32'hbc20327e),
	.w6(32'hbaf86257),
	.w7(32'hbb865db6),
	.w8(32'hbbbf93e5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35c14c),
	.w1(32'hbaee9efa),
	.w2(32'hbb04f356),
	.w3(32'hbc1edfce),
	.w4(32'hbc108ed2),
	.w5(32'h3b20dd4e),
	.w6(32'h39b2e551),
	.w7(32'hbafbeacb),
	.w8(32'hbbcef61e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f7055),
	.w1(32'hbb32c9f8),
	.w2(32'h3b685d1c),
	.w3(32'hbc12554e),
	.w4(32'h3b30e0a5),
	.w5(32'h3a5da854),
	.w6(32'h3a5cd597),
	.w7(32'hbba4d484),
	.w8(32'h3bac70f9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c4892),
	.w1(32'hbb92c45a),
	.w2(32'h3c790356),
	.w3(32'h3b4cd806),
	.w4(32'h3b3d3f9e),
	.w5(32'hbb21c023),
	.w6(32'hba9666ab),
	.w7(32'h3b30fbae),
	.w8(32'h3b374d6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f6c2),
	.w1(32'hbb6521fa),
	.w2(32'hb99d717c),
	.w3(32'hbc02048a),
	.w4(32'hbb346d93),
	.w5(32'h3ab8fa06),
	.w6(32'h3ac1adbe),
	.w7(32'hbb044eb6),
	.w8(32'h37743a71),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981a054),
	.w1(32'hbc31ff93),
	.w2(32'h3b32596e),
	.w3(32'h3b6c8e08),
	.w4(32'h3c022184),
	.w5(32'h3b1a26ff),
	.w6(32'hba96494a),
	.w7(32'h3bbb4dd7),
	.w8(32'h3ba0b390),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a50673),
	.w1(32'h3b2ca575),
	.w2(32'h3b69173d),
	.w3(32'h3a852ebe),
	.w4(32'hbac8a7be),
	.w5(32'h3caf81d6),
	.w6(32'h3b52ffac),
	.w7(32'hbc311b03),
	.w8(32'h3b41b542),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849712),
	.w1(32'h3a9e4e50),
	.w2(32'h3c1859cc),
	.w3(32'h3b929006),
	.w4(32'hb9fbc899),
	.w5(32'h3a1c9434),
	.w6(32'h3c021412),
	.w7(32'hbabf5239),
	.w8(32'hbabd3aa0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32e038),
	.w1(32'h3af38043),
	.w2(32'hbc004993),
	.w3(32'h3b6409e0),
	.w4(32'hba555672),
	.w5(32'hbc1dc90e),
	.w6(32'hbc193404),
	.w7(32'hbc9f3f40),
	.w8(32'hbcbeaa50),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932824),
	.w1(32'hbbe84e93),
	.w2(32'hbb745446),
	.w3(32'h3a517d10),
	.w4(32'hbc0a9159),
	.w5(32'hbb94ac16),
	.w6(32'hbb6c052b),
	.w7(32'hbc0bb237),
	.w8(32'h3be0ed36),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130f20),
	.w1(32'h3ba5aa70),
	.w2(32'hbc9fe47a),
	.w3(32'h3c86f265),
	.w4(32'h3ab6e7b0),
	.w5(32'hbc85c039),
	.w6(32'h3c80af59),
	.w7(32'h3baa2a8e),
	.w8(32'hbc914c13),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeda078),
	.w1(32'h3b48eb79),
	.w2(32'hba94293f),
	.w3(32'h3c81bdd7),
	.w4(32'hbc281e3d),
	.w5(32'hbc208831),
	.w6(32'h3bf08bd2),
	.w7(32'hbc3fe6e6),
	.w8(32'h3c2abd89),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17a905),
	.w1(32'hbbce25e1),
	.w2(32'h3c53f595),
	.w3(32'h3bce7a88),
	.w4(32'hbaa49814),
	.w5(32'hb9deecfa),
	.w6(32'hbbefe7c1),
	.w7(32'hbc951f94),
	.w8(32'hbc0f2ab5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc943f9e),
	.w1(32'hbbe3c2e6),
	.w2(32'h39f79bf7),
	.w3(32'hba61093e),
	.w4(32'h3a283a07),
	.w5(32'hbbe0b7b0),
	.w6(32'h3bc38a5c),
	.w7(32'h3bec25f3),
	.w8(32'h3b3dadae),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8521c8),
	.w1(32'hbc037a5a),
	.w2(32'hbb08630f),
	.w3(32'hbba101c0),
	.w4(32'hbc05ffd8),
	.w5(32'h39e56e62),
	.w6(32'h3c91731a),
	.w7(32'h3c788e74),
	.w8(32'h3c9f886c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59d6c3),
	.w1(32'hbb0ac342),
	.w2(32'h3b4e7532),
	.w3(32'hbc3bbedd),
	.w4(32'h3b232f74),
	.w5(32'h3a981f3d),
	.w6(32'hbae8a1a5),
	.w7(32'h3a30f344),
	.w8(32'h3a8daa87),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be73ab4),
	.w1(32'h3b065583),
	.w2(32'hbbda6a9e),
	.w3(32'h3c0706bd),
	.w4(32'h3b6c9d5f),
	.w5(32'hbb428a19),
	.w6(32'hbc0d7e33),
	.w7(32'hbc94225b),
	.w8(32'hbc94071f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb259d9),
	.w1(32'h3d0a16ae),
	.w2(32'hbc874dd3),
	.w3(32'h3c3f4c22),
	.w4(32'hbc08374c),
	.w5(32'hbd048f25),
	.w6(32'h3c2b5ae1),
	.w7(32'h3aeaea5a),
	.w8(32'h3c7aeb45),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c16d),
	.w1(32'h3d09fb3d),
	.w2(32'h3cfca7a8),
	.w3(32'h3cc4738d),
	.w4(32'h3d0d3749),
	.w5(32'h3d1e17fb),
	.w6(32'h3ca16c7c),
	.w7(32'h3d14ba3b),
	.w8(32'hbc230e6b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e69c),
	.w1(32'h3ac4a4ea),
	.w2(32'h3b7a8ed1),
	.w3(32'hbb820736),
	.w4(32'h3b230b1b),
	.w5(32'h3c222aea),
	.w6(32'h3c3e42cd),
	.w7(32'h3cc5da02),
	.w8(32'h3cb05d76),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cbdd8),
	.w1(32'h3bdda06e),
	.w2(32'h3cf6509e),
	.w3(32'hbb888f44),
	.w4(32'h3aca49d3),
	.w5(32'h3bbeb0c7),
	.w6(32'h3cf8c988),
	.w7(32'h3b57b39f),
	.w8(32'h3bb1f786),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c099e48),
	.w1(32'h3b882842),
	.w2(32'hbcc6e661),
	.w3(32'h3bfc3478),
	.w4(32'h3c4040ab),
	.w5(32'hbb47cf4d),
	.w6(32'h3c4f23f9),
	.w7(32'h3c84b880),
	.w8(32'hbc3d1824),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fea4d4),
	.w1(32'h3c8b90d0),
	.w2(32'hbb82c4e1),
	.w3(32'h3a325674),
	.w4(32'h3afb25bb),
	.w5(32'h3b7d112c),
	.w6(32'h3b36d486),
	.w7(32'hbae71750),
	.w8(32'hbadb2b50),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a7cce),
	.w1(32'h3cac40c0),
	.w2(32'h3cdfa05b),
	.w3(32'h3cafe919),
	.w4(32'h3ce1a4a0),
	.w5(32'h3cddee44),
	.w6(32'h3c337d18),
	.w7(32'h3b8f8e09),
	.w8(32'h3acfd188),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb091105),
	.w1(32'hbbc156a6),
	.w2(32'hbc66539d),
	.w3(32'hba21182d),
	.w4(32'hbbf8a2fa),
	.w5(32'hbbdb5f23),
	.w6(32'hb8794fa2),
	.w7(32'hbb8c337f),
	.w8(32'hbb381bc4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0660ca),
	.w1(32'h3c1bea5b),
	.w2(32'h3ba62741),
	.w3(32'h3b32b256),
	.w4(32'hb8daa56a),
	.w5(32'h3a868666),
	.w6(32'h39a1cfe8),
	.w7(32'hb98308df),
	.w8(32'h3a72f53e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b57c2),
	.w1(32'hbb637eaf),
	.w2(32'h3a038f3e),
	.w3(32'hbb07457e),
	.w4(32'h3bf23932),
	.w5(32'h3ba7da27),
	.w6(32'h3b30ecf3),
	.w7(32'h3b2cd71c),
	.w8(32'h3b398f90),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12446e),
	.w1(32'h3a71d131),
	.w2(32'hbb99726e),
	.w3(32'hbbcc168d),
	.w4(32'h3a933946),
	.w5(32'hbb6cb858),
	.w6(32'hbb8a3660),
	.w7(32'hbc17b29e),
	.w8(32'hbc90edbd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d91f2),
	.w1(32'h399ec12a),
	.w2(32'h3b24dfdb),
	.w3(32'hbb58a650),
	.w4(32'hbb28e0d3),
	.w5(32'h3c1a0a51),
	.w6(32'h3bf7c36a),
	.w7(32'hbaef4c09),
	.w8(32'h3bb9a234),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1d724),
	.w1(32'hbc948e38),
	.w2(32'hbbf6cb24),
	.w3(32'h3b732e5f),
	.w4(32'hbc87a1d8),
	.w5(32'hbc1182b8),
	.w6(32'h3c56a6c4),
	.w7(32'hbb9ae75c),
	.w8(32'h3bc8ec8b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e37a80),
	.w1(32'hb967a9b5),
	.w2(32'h3ba1b2ef),
	.w3(32'hbbc01dd9),
	.w4(32'hbb0c9eca),
	.w5(32'h3bda37ea),
	.w6(32'h3b6f23d4),
	.w7(32'h39ab63eb),
	.w8(32'h3bbdf7d3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2afae2),
	.w1(32'h3b58ac10),
	.w2(32'h3b676dc6),
	.w3(32'hbbab850a),
	.w4(32'h3b28ffc6),
	.w5(32'h3b2e10f7),
	.w6(32'h3bf4424f),
	.w7(32'h39b61276),
	.w8(32'hbc5fe921),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6905f4),
	.w1(32'hbbb62007),
	.w2(32'h3c12351a),
	.w3(32'h3c34c73b),
	.w4(32'h3cdc07a7),
	.w5(32'h3b55c6b8),
	.w6(32'h3b38d0d0),
	.w7(32'h3bf26779),
	.w8(32'h3b60c30f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03979d),
	.w1(32'hbc554c4d),
	.w2(32'hbc01c679),
	.w3(32'hba05671d),
	.w4(32'h3b6a436c),
	.w5(32'hbbd09648),
	.w6(32'hbb8de04a),
	.w7(32'hbb26db78),
	.w8(32'hbadb9bfd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc9916),
	.w1(32'hbabb9afd),
	.w2(32'hbbcd16d0),
	.w3(32'h3b6398df),
	.w4(32'hb8d57551),
	.w5(32'h3a84dfe4),
	.w6(32'h3c09e6e4),
	.w7(32'h38836394),
	.w8(32'h3d04f52b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe42f19),
	.w1(32'h3a757530),
	.w2(32'h3b2f72d9),
	.w3(32'h3a8c4ac4),
	.w4(32'h3a35ac50),
	.w5(32'hba6ad3bd),
	.w6(32'hbc1e5c8b),
	.w7(32'h3c0af878),
	.w8(32'hbbeec3ba),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a5b3),
	.w1(32'hbba7f9d8),
	.w2(32'hbb831252),
	.w3(32'hbc49216a),
	.w4(32'hbb1899ee),
	.w5(32'hbc47f7ea),
	.w6(32'hbc08e759),
	.w7(32'hbbc94322),
	.w8(32'h3abee046),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accec3e),
	.w1(32'h3b87da48),
	.w2(32'hba3932ab),
	.w3(32'hb9025b3d),
	.w4(32'hbbe9d520),
	.w5(32'h39d9b8d2),
	.w6(32'hbb59d2d9),
	.w7(32'h3bba3913),
	.w8(32'h3a7f5780),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70a4aa),
	.w1(32'h3a35b487),
	.w2(32'hbc5126c1),
	.w3(32'h3c501d44),
	.w4(32'h3a7113f1),
	.w5(32'h3b2e1610),
	.w6(32'h3b070f10),
	.w7(32'hbc58700e),
	.w8(32'hbb84c37d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9da687),
	.w1(32'h3a053a3a),
	.w2(32'hba57c749),
	.w3(32'hbb453a79),
	.w4(32'hbb24cd9b),
	.w5(32'h3ca9855f),
	.w6(32'h3b8b9001),
	.w7(32'h39884d34),
	.w8(32'h3b3c8de2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c091024),
	.w1(32'h3b9aa640),
	.w2(32'hbc2a8cb4),
	.w3(32'h3c006c5e),
	.w4(32'h3c3afa27),
	.w5(32'hbb97c034),
	.w6(32'h3b342f37),
	.w7(32'hbb7cb002),
	.w8(32'hbc2c40c9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1672a2),
	.w1(32'hbc494643),
	.w2(32'h3b9dce1d),
	.w3(32'hbb59043f),
	.w4(32'hbc5f18be),
	.w5(32'h3b963c5a),
	.w6(32'h3c057d75),
	.w7(32'h3c2589ae),
	.w8(32'h3c696708),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab78474),
	.w1(32'h3bff620b),
	.w2(32'h3be1c7c9),
	.w3(32'h37ea99e6),
	.w4(32'hbb516b6a),
	.w5(32'hbb8572eb),
	.w6(32'hbbbde3f6),
	.w7(32'hbb3eadb7),
	.w8(32'h3b9179c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100080),
	.w1(32'hb98a8889),
	.w2(32'hb9fd5d8e),
	.w3(32'hbb9f27ad),
	.w4(32'hba2df269),
	.w5(32'h3b20a6ce),
	.w6(32'hbad95461),
	.w7(32'h39c026f2),
	.w8(32'hb64158f7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c81f6),
	.w1(32'hb65c002b),
	.w2(32'hbb9d6ed6),
	.w3(32'h3b8e1f2b),
	.w4(32'hbae3b9f2),
	.w5(32'h3c1c5369),
	.w6(32'hba68beb0),
	.w7(32'h383b1164),
	.w8(32'h3abeca5c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c042d),
	.w1(32'hbc260a31),
	.w2(32'hbb510c3f),
	.w3(32'hb97bbdf9),
	.w4(32'h3a73fa9b),
	.w5(32'h3bb78e6f),
	.w6(32'hbbc52df2),
	.w7(32'hbbd250d3),
	.w8(32'h39c85738),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0b642),
	.w1(32'hbc0579df),
	.w2(32'hbc8ca47f),
	.w3(32'h3b12a5d9),
	.w4(32'h3bd9b835),
	.w5(32'hb90583d6),
	.w6(32'h3c82719f),
	.w7(32'hbc9e3c22),
	.w8(32'hbd197bd7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399eb6f3),
	.w1(32'hbc22894b),
	.w2(32'hbc37fc72),
	.w3(32'h3c3e7d14),
	.w4(32'hbc439d18),
	.w5(32'hbc2228f2),
	.w6(32'hbb2891b7),
	.w7(32'hbcc0fb7b),
	.w8(32'hbcc26289),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec415f),
	.w1(32'hba9b4722),
	.w2(32'hbbcf508e),
	.w3(32'h3b9e6b9e),
	.w4(32'h39e03c06),
	.w5(32'h3c6f5f32),
	.w6(32'h3ab20da7),
	.w7(32'hbba0f1ed),
	.w8(32'h397b3107),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e5ab5),
	.w1(32'h3c17d06b),
	.w2(32'h3b011c11),
	.w3(32'hbaf318cf),
	.w4(32'hbb9e7660),
	.w5(32'hbc05499c),
	.w6(32'hbb7ae6d3),
	.w7(32'hbc348435),
	.w8(32'hbba97c5e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffb550),
	.w1(32'h3b82ab99),
	.w2(32'hbb60916f),
	.w3(32'h3c3695a6),
	.w4(32'h3b12fd2d),
	.w5(32'h3d2ba69d),
	.w6(32'hbaf82e53),
	.w7(32'h3b2989d5),
	.w8(32'h3b5de958),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86e753),
	.w1(32'hba4f200d),
	.w2(32'h3b6e91b8),
	.w3(32'h3c3f5866),
	.w4(32'hb94b8196),
	.w5(32'h3b135c9a),
	.w6(32'h3c01d5b0),
	.w7(32'hbc247131),
	.w8(32'hbbae0d9b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98a77a),
	.w1(32'hbbbf1eeb),
	.w2(32'h3b715826),
	.w3(32'hbbdd6756),
	.w4(32'hb9b90bb5),
	.w5(32'h3c4d9c07),
	.w6(32'h3bc74e14),
	.w7(32'h3c972442),
	.w8(32'h3bf2c81e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63f4e1),
	.w1(32'hbb97883d),
	.w2(32'hbc80cd14),
	.w3(32'h3c8d0f71),
	.w4(32'h3b808125),
	.w5(32'hbc3cdf2e),
	.w6(32'hbaf82efd),
	.w7(32'hbb6098ce),
	.w8(32'hbc893228),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba676a15),
	.w1(32'hbb1769a3),
	.w2(32'h3c15e199),
	.w3(32'hb928176d),
	.w4(32'hbbc71463),
	.w5(32'h3c23223f),
	.w6(32'h3bdb045a),
	.w7(32'h3b46942f),
	.w8(32'h3c85e666),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c810bce),
	.w1(32'h3acda4ea),
	.w2(32'h3b989a69),
	.w3(32'h3bbdb7af),
	.w4(32'hbb97b74b),
	.w5(32'h3a079f02),
	.w6(32'h3acbd60e),
	.w7(32'h3b0429d0),
	.w8(32'hbbeb8885),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56dd20),
	.w1(32'h3ca1a9b2),
	.w2(32'hbc41798d),
	.w3(32'h3c9f9957),
	.w4(32'h3bd83d4f),
	.w5(32'hbc0d33bd),
	.w6(32'hbc2799a2),
	.w7(32'hbbabf75f),
	.w8(32'hbcb1dc36),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0fc5d),
	.w1(32'h3b251573),
	.w2(32'hbc2b2fb5),
	.w3(32'hbb6afced),
	.w4(32'h3cbb2f7c),
	.w5(32'h3b19711f),
	.w6(32'hbc0a5288),
	.w7(32'hba5a2c34),
	.w8(32'h3b567065),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934667),
	.w1(32'h3c840a81),
	.w2(32'hbaff74ab),
	.w3(32'hbb43f1c2),
	.w4(32'h3c213bf9),
	.w5(32'hbb303c08),
	.w6(32'h3c235740),
	.w7(32'hbb761755),
	.w8(32'h3a058da8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d6b8e),
	.w1(32'hbaf0228b),
	.w2(32'hbb8d030d),
	.w3(32'h3bf2f0e4),
	.w4(32'h3a676c4e),
	.w5(32'h3b29b47e),
	.w6(32'h3afb9f48),
	.w7(32'h3bd4b820),
	.w8(32'hbb956973),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba524f8),
	.w1(32'h3c54c4bc),
	.w2(32'hbc9598fe),
	.w3(32'hbb10edfd),
	.w4(32'hbc58d63e),
	.w5(32'hbc2e2641),
	.w6(32'h3c5b637d),
	.w7(32'hbc8289f7),
	.w8(32'h3b0ecae3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f7ef1),
	.w1(32'h3a4fcb03),
	.w2(32'h39270ecc),
	.w3(32'h379ba07f),
	.w4(32'h3c93024d),
	.w5(32'hbbc84686),
	.w6(32'h3967e0c5),
	.w7(32'hbbb02520),
	.w8(32'hbbe832b5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cb54c),
	.w1(32'h3ba13fe1),
	.w2(32'hbba4c55c),
	.w3(32'hbc015719),
	.w4(32'hba69b8c2),
	.w5(32'h3afb29e7),
	.w6(32'h3cb34dd5),
	.w7(32'hbc3e79b5),
	.w8(32'hb9819e4b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe981aa),
	.w1(32'h3b011408),
	.w2(32'hb98b4c13),
	.w3(32'hb9b08dba),
	.w4(32'h3b0dc8da),
	.w5(32'h3bb98fce),
	.w6(32'h3b1f909d),
	.w7(32'hbbdbd455),
	.w8(32'h398b1dfc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5ee30),
	.w1(32'h3c0691f9),
	.w2(32'hbb5ebf15),
	.w3(32'h3b3917f8),
	.w4(32'h380ea976),
	.w5(32'h3a2cbd56),
	.w6(32'hba931729),
	.w7(32'h3b83af3a),
	.w8(32'hbab1df73),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac12f0d),
	.w1(32'hbbce00ed),
	.w2(32'hbbb2bee7),
	.w3(32'hbc154612),
	.w4(32'hba247961),
	.w5(32'h3a9afd17),
	.w6(32'hba06c411),
	.w7(32'h3bd5b52f),
	.w8(32'h3bce655c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a36ec),
	.w1(32'hbc39c946),
	.w2(32'h3b4c34cc),
	.w3(32'h3bbe7edc),
	.w4(32'hbca3d3b4),
	.w5(32'hbc064af0),
	.w6(32'hbb46b9ba),
	.w7(32'hbc34dce9),
	.w8(32'hbc820d9f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192ffc),
	.w1(32'hbbc15281),
	.w2(32'hbbcc52e7),
	.w3(32'hbb493ee0),
	.w4(32'hbb670fe6),
	.w5(32'hbc129a03),
	.w6(32'hba89019f),
	.w7(32'h3b0dc559),
	.w8(32'hbb4bde0e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4520f),
	.w1(32'hbb1a470c),
	.w2(32'hbba84574),
	.w3(32'h3c618d7c),
	.w4(32'hbc150e43),
	.w5(32'hbc158e3c),
	.w6(32'hbbbfec24),
	.w7(32'hbc37a246),
	.w8(32'hbbfe58ed),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85fc0f),
	.w1(32'hbbb17cb2),
	.w2(32'hbb5f418d),
	.w3(32'h3c373f1f),
	.w4(32'hbbc2231c),
	.w5(32'h3b1b54ae),
	.w6(32'h3b599e20),
	.w7(32'hba297fcb),
	.w8(32'hbc903220),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a0025),
	.w1(32'h39a0da2d),
	.w2(32'hbbbd41ee),
	.w3(32'h3c20328c),
	.w4(32'hbbcc4068),
	.w5(32'h3b8173b9),
	.w6(32'hbb402377),
	.w7(32'h3adbcaf0),
	.w8(32'hbc1d15b3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17c3ed),
	.w1(32'hbd05995b),
	.w2(32'hbc028453),
	.w3(32'hbb848f4c),
	.w4(32'hbcbd3aca),
	.w5(32'hbcd8d301),
	.w6(32'h38abb1a6),
	.w7(32'hbc0d8d00),
	.w8(32'hba6946c8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d302b),
	.w1(32'h3af1c2b6),
	.w2(32'hba20fbbf),
	.w3(32'hb97f7d62),
	.w4(32'h38e7b9f3),
	.w5(32'h3b722294),
	.w6(32'h3ca0ae39),
	.w7(32'hbb604d7b),
	.w8(32'h3baf8285),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7d6e0),
	.w1(32'hba76f092),
	.w2(32'h3a78815c),
	.w3(32'h3c2430f1),
	.w4(32'h3a7ef4a8),
	.w5(32'hbb31cda9),
	.w6(32'hbb8bd7e7),
	.w7(32'h39d640ac),
	.w8(32'hb92fd46b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ea5b),
	.w1(32'hbb8f4407),
	.w2(32'hbbe294aa),
	.w3(32'hbb6c3550),
	.w4(32'hba779af9),
	.w5(32'hbc83e618),
	.w6(32'h3c395502),
	.w7(32'h3ab7b85b),
	.w8(32'h3b50a047),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b92eb),
	.w1(32'h39eb5549),
	.w2(32'h3b73c660),
	.w3(32'hbb904c29),
	.w4(32'hbbaca0e4),
	.w5(32'hbb384627),
	.w6(32'hbbd423b5),
	.w7(32'h3bead080),
	.w8(32'h3bed3784),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb193),
	.w1(32'h3cb2ca9a),
	.w2(32'h397f011a),
	.w3(32'h3a0309ee),
	.w4(32'h3b6e847d),
	.w5(32'h3b0847ac),
	.w6(32'hbb2219b1),
	.w7(32'h3be0e768),
	.w8(32'h3bf280ae),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9026e2),
	.w1(32'hba35b0dd),
	.w2(32'hbab485c2),
	.w3(32'h3ab2da66),
	.w4(32'hba3bec8b),
	.w5(32'hbbc4281c),
	.w6(32'h3b1c7c5d),
	.w7(32'hbb0b8127),
	.w8(32'hbc1d7f92),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b210b90),
	.w1(32'h394593dd),
	.w2(32'hbb50070e),
	.w3(32'hbb484a88),
	.w4(32'h3bce512d),
	.w5(32'h3b931388),
	.w6(32'h392b9791),
	.w7(32'h3be12798),
	.w8(32'h3cd12a35),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b593ceb),
	.w1(32'h3b1f0e26),
	.w2(32'hbbf570b4),
	.w3(32'h3c166415),
	.w4(32'hbbed0ba5),
	.w5(32'hbc6320d8),
	.w6(32'hb9f20613),
	.w7(32'hbc11d890),
	.w8(32'hbc5d12dd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0ebd6),
	.w1(32'hbb54c094),
	.w2(32'hb9830d6e),
	.w3(32'h3b25c75a),
	.w4(32'hbb924ac3),
	.w5(32'hbbf43a8f),
	.w6(32'h3c72defd),
	.w7(32'hbb7cfd76),
	.w8(32'hbc11c8e6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb4101),
	.w1(32'hbc3dff9c),
	.w2(32'hbad82104),
	.w3(32'hbbcb34b5),
	.w4(32'h3c4dc2dc),
	.w5(32'hbb483087),
	.w6(32'h3a448999),
	.w7(32'hbc3e8474),
	.w8(32'hbbcff9f2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d86d4),
	.w1(32'hb9b46467),
	.w2(32'hbb4eb396),
	.w3(32'hb9e99155),
	.w4(32'h3ac287f2),
	.w5(32'h391aea7c),
	.w6(32'hb91ed095),
	.w7(32'hbaab124b),
	.w8(32'h3aa22336),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae33004),
	.w1(32'hbbd89a2f),
	.w2(32'hbbe334cc),
	.w3(32'h3c3163bb),
	.w4(32'h38cc4ecc),
	.w5(32'hbb7aec64),
	.w6(32'h39617072),
	.w7(32'hbc22a502),
	.w8(32'hbcb718a0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d87cd),
	.w1(32'h3bea5808),
	.w2(32'hbb21317b),
	.w3(32'hbbc81fce),
	.w4(32'hba797137),
	.w5(32'hbbb57c1c),
	.w6(32'hbbec085d),
	.w7(32'hba86d050),
	.w8(32'h3ac2d6e8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69ee43),
	.w1(32'h3a9c21b9),
	.w2(32'h3b919243),
	.w3(32'h3b5649f9),
	.w4(32'h390108b1),
	.w5(32'h39c5ae39),
	.w6(32'hbbe57962),
	.w7(32'h3b064f94),
	.w8(32'hba59ec44),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f0b0f),
	.w1(32'h3b8cca3d),
	.w2(32'h3c1fe926),
	.w3(32'hbc2f1f27),
	.w4(32'hba90911e),
	.w5(32'h3b058663),
	.w6(32'hbb8a686f),
	.w7(32'h3b897df8),
	.w8(32'h3c9f43d8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c330b3e),
	.w1(32'hbb23aac4),
	.w2(32'hbc01d088),
	.w3(32'h3c336a8b),
	.w4(32'hbba7f7c5),
	.w5(32'hbc12e7de),
	.w6(32'h3c274643),
	.w7(32'hbc47f112),
	.w8(32'hbce77d00),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecfdd1),
	.w1(32'h3a36fc26),
	.w2(32'h3a9439ee),
	.w3(32'h3b8bc099),
	.w4(32'hb766fdc7),
	.w5(32'hbaafbc49),
	.w6(32'hbb16f0d7),
	.w7(32'h3bebd8d3),
	.w8(32'hbc1a0ec1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eea2c),
	.w1(32'hb6c8ddcc),
	.w2(32'h3b7ba69e),
	.w3(32'h3a10a296),
	.w4(32'hbab38060),
	.w5(32'h3bbbc2ec),
	.w6(32'h3a985e88),
	.w7(32'h3bb7fcac),
	.w8(32'h3c06ffa3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fc504),
	.w1(32'hb99daaae),
	.w2(32'h3ad00822),
	.w3(32'h3b6b8d42),
	.w4(32'hba61d686),
	.w5(32'hbbce67a7),
	.w6(32'h3c0dc597),
	.w7(32'h3bca8fec),
	.w8(32'hba4ee669),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c3efc),
	.w1(32'hbbb85f5b),
	.w2(32'hbc005659),
	.w3(32'hb7ffa699),
	.w4(32'hbc1866c4),
	.w5(32'hbb8bab51),
	.w6(32'hbc6852c8),
	.w7(32'hbc4ec446),
	.w8(32'hbc456717),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc2b56),
	.w1(32'hbb023265),
	.w2(32'hbb2e050f),
	.w3(32'hbacee1f0),
	.w4(32'hbb033323),
	.w5(32'h3bda5016),
	.w6(32'hba316f93),
	.w7(32'h3aa14e42),
	.w8(32'hbb1e9b1b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73e8c1),
	.w1(32'h3b2b2f5b),
	.w2(32'hbbcf5296),
	.w3(32'h3b001c15),
	.w4(32'h3b304284),
	.w5(32'hbb8077a4),
	.w6(32'hbc21c9b3),
	.w7(32'hbbf43316),
	.w8(32'hbc83d152),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d921),
	.w1(32'h39bddcc4),
	.w2(32'hbabf5bfc),
	.w3(32'h3a15b428),
	.w4(32'h3a64f0a4),
	.w5(32'h3b42e2ac),
	.w6(32'h39c72843),
	.w7(32'h3bf98c7e),
	.w8(32'h3c693524),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71be6c),
	.w1(32'hba72a3b7),
	.w2(32'h3b6bfdf3),
	.w3(32'h3b1ad72d),
	.w4(32'hbab04d43),
	.w5(32'h3b79c838),
	.w6(32'h3b8f944c),
	.w7(32'h3b51b4af),
	.w8(32'h3c0017fa),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab52027),
	.w1(32'hba04842e),
	.w2(32'h3b3bb442),
	.w3(32'hbc1829f0),
	.w4(32'h3c4e87c4),
	.w5(32'h3af9320b),
	.w6(32'h3967029d),
	.w7(32'hbbe1e320),
	.w8(32'hbb10dfd3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066502),
	.w1(32'hbb5afb51),
	.w2(32'hba59e7a4),
	.w3(32'h39746436),
	.w4(32'h3a0eb39d),
	.w5(32'h3b5ac09e),
	.w6(32'h3a100d19),
	.w7(32'hb91d9c51),
	.w8(32'hbb723866),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af8c3c),
	.w1(32'h3c8acf2b),
	.w2(32'h3bd032ad),
	.w3(32'h3b7ac342),
	.w4(32'h3b233d4c),
	.w5(32'h3bc91a66),
	.w6(32'h39a39556),
	.w7(32'hb9a23496),
	.w8(32'h3accbba4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb462f1e),
	.w1(32'h36e88518),
	.w2(32'h3b57c238),
	.w3(32'h380abd88),
	.w4(32'hb652a888),
	.w5(32'h3bc8309c),
	.w6(32'hb8bba37a),
	.w7(32'h3bfe7e4f),
	.w8(32'h3b905e0f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949d3c0),
	.w1(32'hbb2de46a),
	.w2(32'h3b77d959),
	.w3(32'hbbb1779c),
	.w4(32'h3b8a4a49),
	.w5(32'h3afc63e2),
	.w6(32'h3b11de94),
	.w7(32'hba57011f),
	.w8(32'h3bad6992),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9530eff),
	.w1(32'h3c2e2eaf),
	.w2(32'h3a6ff52d),
	.w3(32'h3ab42d83),
	.w4(32'hb863f885),
	.w5(32'h3b6921ef),
	.w6(32'hb74fb066),
	.w7(32'hbc00ff28),
	.w8(32'hbabf5311),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aa53f),
	.w1(32'hbbbc83a0),
	.w2(32'hba1b07c0),
	.w3(32'h3887a282),
	.w4(32'hb9cd1c31),
	.w5(32'hbb18e649),
	.w6(32'h3aa6692f),
	.w7(32'hbb98f729),
	.w8(32'hbb97284f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c319e55),
	.w1(32'h3a133d8d),
	.w2(32'hba8041a9),
	.w3(32'hbb85928a),
	.w4(32'h3bf635ff),
	.w5(32'hbb1f7ac0),
	.w6(32'h3b5dc516),
	.w7(32'h3c878ce9),
	.w8(32'h3b994319),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c2057),
	.w1(32'h3c1565bd),
	.w2(32'h3b1082b2),
	.w3(32'h3c08998e),
	.w4(32'h3c527ec7),
	.w5(32'h3c3ce9aa),
	.w6(32'h3be8e73f),
	.w7(32'h3c3a68b7),
	.w8(32'h3a6e2dd8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8d386),
	.w1(32'h3a9d3a57),
	.w2(32'h39f7bbc6),
	.w3(32'h3a2f926d),
	.w4(32'hba43bc98),
	.w5(32'hbae0eaef),
	.w6(32'hba8224ac),
	.w7(32'hbb9260bf),
	.w8(32'h3abf7ec8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a3e7a),
	.w1(32'hbb4dc138),
	.w2(32'hbc0556bb),
	.w3(32'h3c49651b),
	.w4(32'hbb2f3700),
	.w5(32'hbc01ffc4),
	.w6(32'hbc70fb50),
	.w7(32'hbcd5d234),
	.w8(32'hbd13028c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08f734),
	.w1(32'hbbb203e3),
	.w2(32'h3c96aadc),
	.w3(32'h3be41abc),
	.w4(32'hbb63b997),
	.w5(32'hbc4e12e6),
	.w6(32'h3d00603b),
	.w7(32'h3c5f4231),
	.w8(32'h3cb04957),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c285ede),
	.w1(32'h3bd21e4b),
	.w2(32'hbb1d1c24),
	.w3(32'h3ae791d6),
	.w4(32'hb9f2490d),
	.w5(32'hbbce0712),
	.w6(32'h3bff990c),
	.w7(32'h3b2b5e94),
	.w8(32'hbb1b72fd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5163d),
	.w1(32'hbac58be7),
	.w2(32'hbac6aa78),
	.w3(32'hbbaf5346),
	.w4(32'h38b5c339),
	.w5(32'hba166683),
	.w6(32'hba7000b2),
	.w7(32'h3a99b771),
	.w8(32'h3c258e07),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384cc5),
	.w1(32'hbbebf707),
	.w2(32'hbbfc3bc5),
	.w3(32'h39d99172),
	.w4(32'hba8885a4),
	.w5(32'hb9d3bd36),
	.w6(32'hbb41445e),
	.w7(32'hbad9c87f),
	.w8(32'h3918ba1e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940da0f),
	.w1(32'h3b64f958),
	.w2(32'h3b1146c7),
	.w3(32'h3a3d801c),
	.w4(32'h3983d0a0),
	.w5(32'h3a3cd62d),
	.w6(32'hb8954d55),
	.w7(32'h3b38b66c),
	.w8(32'h3b183680),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7671),
	.w1(32'h3bdf53e7),
	.w2(32'hbba35e2e),
	.w3(32'h3bf84c0d),
	.w4(32'h3c0b7dbe),
	.w5(32'hbbc5cf6a),
	.w6(32'h3af828c5),
	.w7(32'h3ac43921),
	.w8(32'hbc86e9d7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe9ce5),
	.w1(32'hbab0e767),
	.w2(32'hbac6c117),
	.w3(32'h3bb26b51),
	.w4(32'h3b3b030f),
	.w5(32'h3ac7ec8e),
	.w6(32'h3acdb928),
	.w7(32'hbb4a6c15),
	.w8(32'hbc5da02d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91514e),
	.w1(32'h3b86fdf3),
	.w2(32'h3bb4e5e4),
	.w3(32'h3b02a0b2),
	.w4(32'h3bd4d707),
	.w5(32'h3c190fcb),
	.w6(32'h3a966a6a),
	.w7(32'h3bd1428f),
	.w8(32'h3bbca0d7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17de73),
	.w1(32'h3b87062b),
	.w2(32'h3c4dd404),
	.w3(32'hbbe11d64),
	.w4(32'hbb4c0c8f),
	.w5(32'hb8efd0cc),
	.w6(32'h3bdc10f9),
	.w7(32'hba3835d8),
	.w8(32'h3bb3efad),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8d456),
	.w1(32'h3a84b109),
	.w2(32'hbc3fc3cf),
	.w3(32'h3b5a973e),
	.w4(32'h3a062e4a),
	.w5(32'hbc17ca70),
	.w6(32'hb9d4550b),
	.w7(32'hbc7e5d35),
	.w8(32'hbc95c489),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a28f),
	.w1(32'h3bd041b5),
	.w2(32'h3b8187e0),
	.w3(32'hbbf71d75),
	.w4(32'hbc64376d),
	.w5(32'hbb3d4038),
	.w6(32'h3b20043d),
	.w7(32'h3ad95296),
	.w8(32'h3bbf5296),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bf616),
	.w1(32'h3cc79c5d),
	.w2(32'h39bc9aa2),
	.w3(32'h3ae403a0),
	.w4(32'h3b1905d6),
	.w5(32'hbb100288),
	.w6(32'hbb190d72),
	.w7(32'hbb457c6f),
	.w8(32'h3bb4ffb3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49162e),
	.w1(32'hba2c630c),
	.w2(32'h3af5ecef),
	.w3(32'h3ce4d064),
	.w4(32'h3a217884),
	.w5(32'h3bc7f8c7),
	.w6(32'hbb336c48),
	.w7(32'h3c0d38f0),
	.w8(32'hba506494),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886c1c2),
	.w1(32'h3b557461),
	.w2(32'h3a5e5c28),
	.w3(32'h3b88e82b),
	.w4(32'hbb39aa63),
	.w5(32'h3b31e313),
	.w6(32'h3a40fe31),
	.w7(32'hba89fb13),
	.w8(32'hbb53aa0a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5e29),
	.w1(32'hba155851),
	.w2(32'hbb8e0523),
	.w3(32'h3ba19c6d),
	.w4(32'hbb435db6),
	.w5(32'hbbad7ffe),
	.w6(32'h3ae710ce),
	.w7(32'hbbf67293),
	.w8(32'hbc7a9bcf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64508a),
	.w1(32'hbb090f79),
	.w2(32'h3916852e),
	.w3(32'hbbf475f4),
	.w4(32'h3a0fd578),
	.w5(32'h39227e9b),
	.w6(32'hb971b3b9),
	.w7(32'hbab44805),
	.w8(32'h3b64fa14),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba598b47),
	.w1(32'hb87e3374),
	.w2(32'h3ad5db42),
	.w3(32'h3a8506e5),
	.w4(32'h3992280e),
	.w5(32'hbaac8956),
	.w6(32'h3bce493d),
	.w7(32'h3b50dc3a),
	.w8(32'h3bb30c2f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2503e8),
	.w1(32'h39415b7c),
	.w2(32'hbb8ff658),
	.w3(32'hba9f6213),
	.w4(32'h3b693f4a),
	.w5(32'hbb293eda),
	.w6(32'hba774709),
	.w7(32'hbc395d2b),
	.w8(32'h3a9579e7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe5c85),
	.w1(32'hbc282c80),
	.w2(32'h3b102f8c),
	.w3(32'hbb141c9a),
	.w4(32'h3bb9a8db),
	.w5(32'h3c328d28),
	.w6(32'hbab131c2),
	.w7(32'h3bda8473),
	.w8(32'h3c103620),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a922cb),
	.w1(32'hba0d2de1),
	.w2(32'h3b316b8c),
	.w3(32'h3badde70),
	.w4(32'hbc50a281),
	.w5(32'h3abb8f6b),
	.w6(32'hbb33c939),
	.w7(32'hbaea94b3),
	.w8(32'hbc4dcd25),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9852303),
	.w1(32'hbaf44fbb),
	.w2(32'hbb8bcc5e),
	.w3(32'hbc15ad34),
	.w4(32'hb956bdd7),
	.w5(32'hbbb58faf),
	.w6(32'hbb212df3),
	.w7(32'hbbac3a6a),
	.w8(32'hbc0b36f4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9450eb),
	.w1(32'hbaec4d5e),
	.w2(32'h3b6daefb),
	.w3(32'hbaa73415),
	.w4(32'hba89d848),
	.w5(32'h3ad5cd99),
	.w6(32'hbbbc8b35),
	.w7(32'hbc53545d),
	.w8(32'h3c8b70be),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba494a),
	.w1(32'hbad6bdfb),
	.w2(32'hb9d41ad0),
	.w3(32'h3c91e862),
	.w4(32'hb9a6312d),
	.w5(32'hbbc7e64c),
	.w6(32'h3a9d0344),
	.w7(32'hbc3e1408),
	.w8(32'h39dd6454),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c507685),
	.w1(32'hbb8ae0f4),
	.w2(32'hbc1db500),
	.w3(32'h3c155c77),
	.w4(32'hbb3e0941),
	.w5(32'hbc8a3de1),
	.w6(32'h3c120bf3),
	.w7(32'hbc375229),
	.w8(32'hbce7d5e3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2e24f),
	.w1(32'h3bd567d9),
	.w2(32'hbcb2ac9b),
	.w3(32'hbbd833a1),
	.w4(32'hbbe8ae4a),
	.w5(32'hbabd72ff),
	.w6(32'hbb4425e8),
	.w7(32'hbc58999d),
	.w8(32'hbc94b7e6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ed7d2),
	.w1(32'h3af964b0),
	.w2(32'h3b190702),
	.w3(32'hba11fcc5),
	.w4(32'h3b9c88f9),
	.w5(32'h3a3ea055),
	.w6(32'hba829031),
	.w7(32'hb9c613ab),
	.w8(32'hbb1dcc1e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dd466),
	.w1(32'h3bee4f5a),
	.w2(32'hbc91c339),
	.w3(32'h3be24640),
	.w4(32'hbbe88498),
	.w5(32'hbc9d8f81),
	.w6(32'h3c7799ac),
	.w7(32'h3c96bf74),
	.w8(32'h3c018181),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce632a),
	.w1(32'hb9acde23),
	.w2(32'hbb2214f5),
	.w3(32'h3b8c00d5),
	.w4(32'hbc45b7b0),
	.w5(32'hb7dc64a4),
	.w6(32'hbafb9ddf),
	.w7(32'hba7147fc),
	.w8(32'hb70cca09),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f9d93),
	.w1(32'hba79f1e5),
	.w2(32'hba3827c3),
	.w3(32'hbb4be00c),
	.w4(32'h3c471585),
	.w5(32'h3c69fccf),
	.w6(32'hb9eb0472),
	.w7(32'hbb196baa),
	.w8(32'hbabd4f2e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2736ee),
	.w1(32'h3c082042),
	.w2(32'hbcf85615),
	.w3(32'h3bbe6085),
	.w4(32'h3ca88a67),
	.w5(32'hbc384413),
	.w6(32'h3ca35ac9),
	.w7(32'h3c44e085),
	.w8(32'hbd165605),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb44c64),
	.w1(32'hbb575516),
	.w2(32'hbbeb2c95),
	.w3(32'h3cd405af),
	.w4(32'h3b6fb4e7),
	.w5(32'hbc23a42b),
	.w6(32'hbc298c9a),
	.w7(32'hbd0c2039),
	.w8(32'hbcaa3f08),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c100d4b),
	.w1(32'h3bb10910),
	.w2(32'h3b7f239b),
	.w3(32'h3c7c1774),
	.w4(32'h3c55ea9d),
	.w5(32'hbc0f13b9),
	.w6(32'hb9d95a40),
	.w7(32'h3b2d8df8),
	.w8(32'hbc6fb311),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0b0fd),
	.w1(32'hbb37d7e5),
	.w2(32'hb940e593),
	.w3(32'hbc6f1ceb),
	.w4(32'hbbd4a592),
	.w5(32'hbacaf54d),
	.w6(32'hba35aced),
	.w7(32'hbb29d1dc),
	.w8(32'h3bfad362),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f1360),
	.w1(32'hbbedef64),
	.w2(32'h3b77afde),
	.w3(32'hbb9b7261),
	.w4(32'hbadec42b),
	.w5(32'h3c6d24da),
	.w6(32'h3bcfc481),
	.w7(32'h3b161c85),
	.w8(32'h3c96fd25),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb7468),
	.w1(32'hbb59ef4a),
	.w2(32'hbaa61235),
	.w3(32'hbb8eaef1),
	.w4(32'h3b24371c),
	.w5(32'h3bc695e9),
	.w6(32'h3a8abcf1),
	.w7(32'hb952403f),
	.w8(32'h39bbddcc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb6108),
	.w1(32'hba5ff261),
	.w2(32'h3ae3a553),
	.w3(32'hbb2e1dcc),
	.w4(32'hbb3727d1),
	.w5(32'h38f90fad),
	.w6(32'h3acb8b34),
	.w7(32'h3b610c74),
	.w8(32'hba60f4f0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb258ab3),
	.w1(32'hbc2ab282),
	.w2(32'hbb43c8f6),
	.w3(32'h3bc7a308),
	.w4(32'hba4bb4d3),
	.w5(32'h39b4f0f5),
	.w6(32'hbb3f5b02),
	.w7(32'hbc880336),
	.w8(32'hba7d450b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ffce),
	.w1(32'hbb208552),
	.w2(32'hbb335b03),
	.w3(32'h3bba89a1),
	.w4(32'hba3d8196),
	.w5(32'h3babc8a6),
	.w6(32'hbaa9675f),
	.w7(32'hbb1cd5cd),
	.w8(32'hb96f722b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39cba8),
	.w1(32'hbbbb0e58),
	.w2(32'hbc58ecc7),
	.w3(32'h3c1f6642),
	.w4(32'hbb97202a),
	.w5(32'hbb62f011),
	.w6(32'hbbbebb3f),
	.w7(32'h3bad6473),
	.w8(32'hbc04e307),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78a63),
	.w1(32'hb962e7af),
	.w2(32'hbbacf824),
	.w3(32'hbbf5e875),
	.w4(32'hbc1e19b6),
	.w5(32'h3c0c26a2),
	.w6(32'h3bf8081a),
	.w7(32'hbc35ca8e),
	.w8(32'hbcc7dfd2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5627dc),
	.w1(32'hb895a41d),
	.w2(32'hbaf025bd),
	.w3(32'hbc26349c),
	.w4(32'hbbd05329),
	.w5(32'h3accdd15),
	.w6(32'h398b6e7a),
	.w7(32'hbc47c170),
	.w8(32'hbb7914ec),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54d4dd),
	.w1(32'hbba9d101),
	.w2(32'h3c8c72a3),
	.w3(32'h3bc43e46),
	.w4(32'hbbebb094),
	.w5(32'hbbf10914),
	.w6(32'hb87c540e),
	.w7(32'h3c4e546e),
	.w8(32'hba9f88b8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b33c7),
	.w1(32'h3bb4b848),
	.w2(32'h3b95ec3c),
	.w3(32'h3c81a822),
	.w4(32'h3c6cc487),
	.w5(32'h3bc15720),
	.w6(32'hba83e6c1),
	.w7(32'hbc483f6d),
	.w8(32'hbd0bd2ec),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df3606),
	.w1(32'hbc5c7fa2),
	.w2(32'hbbcf1eda),
	.w3(32'h3c062092),
	.w4(32'hbbea6a87),
	.w5(32'hbb04cd75),
	.w6(32'hbbcc4d61),
	.w7(32'hbc9302e7),
	.w8(32'hbc90d77c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ddd21),
	.w1(32'h3ab96e8d),
	.w2(32'hbb3c7f87),
	.w3(32'hbae44634),
	.w4(32'hbbdf9f47),
	.w5(32'h3c50f036),
	.w6(32'hbc26d202),
	.w7(32'h3c1eeb52),
	.w8(32'h3b8c48c1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb641fe),
	.w1(32'h3c38ec29),
	.w2(32'hbafb6985),
	.w3(32'h3c1acc03),
	.w4(32'hbc45433b),
	.w5(32'hbbf8242f),
	.w6(32'hb9838647),
	.w7(32'hbb636cc7),
	.w8(32'hbce0388e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054a60),
	.w1(32'h3b4875fb),
	.w2(32'h3cdcc5fc),
	.w3(32'h3bc7b0fe),
	.w4(32'h3b6388d1),
	.w5(32'hbbbf9c0f),
	.w6(32'h3b9b5423),
	.w7(32'h3c987db4),
	.w8(32'hbca9cc9a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed8496),
	.w1(32'h3b66a89d),
	.w2(32'hbbcf27b4),
	.w3(32'h3bcdd650),
	.w4(32'hbb50d384),
	.w5(32'hbbd16d12),
	.w6(32'h3d16a0a2),
	.w7(32'hba81b9ba),
	.w8(32'h3c251278),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6abe6b),
	.w1(32'hbbb63738),
	.w2(32'hba1c8609),
	.w3(32'h3b1d0bd4),
	.w4(32'h37d5d30c),
	.w5(32'h3b377992),
	.w6(32'hbc8c0e1b),
	.w7(32'hba30f8e2),
	.w8(32'hb95f0886),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0aa58),
	.w1(32'hba4cff9d),
	.w2(32'hbab5ca5b),
	.w3(32'hbb746b8d),
	.w4(32'h3bdb6ff4),
	.w5(32'hbb59cbcc),
	.w6(32'hbb81af38),
	.w7(32'hb6358747),
	.w8(32'hbbf45a6a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b008a51),
	.w1(32'h3b9223cc),
	.w2(32'h3baae5db),
	.w3(32'hbc05ee16),
	.w4(32'hbadf5470),
	.w5(32'h3b4f2113),
	.w6(32'hbb9d7213),
	.w7(32'hba85c950),
	.w8(32'h3bc38082),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95da2c),
	.w1(32'hbbc04796),
	.w2(32'hba00d86a),
	.w3(32'h3acca1d3),
	.w4(32'hbb917ccd),
	.w5(32'hbabe7f2a),
	.w6(32'h3c452e2b),
	.w7(32'h3c1b88be),
	.w8(32'hbb9001d4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431e84),
	.w1(32'h3c22620b),
	.w2(32'hba70780b),
	.w3(32'hbb464662),
	.w4(32'h3c829232),
	.w5(32'hbc80cbb7),
	.w6(32'hbc6b3483),
	.w7(32'hbbc44845),
	.w8(32'hbc1c0622),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ee995),
	.w1(32'hbbaa0fb9),
	.w2(32'hbc586407),
	.w3(32'h3ae3d6b3),
	.w4(32'hbc477900),
	.w5(32'hbc808ad1),
	.w6(32'h3c5857b9),
	.w7(32'h3a35b3e9),
	.w8(32'hbc17fed8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea6537),
	.w1(32'hbc045a9a),
	.w2(32'hbbc8b58d),
	.w3(32'hbc0942e9),
	.w4(32'hbace227d),
	.w5(32'hbc1acda8),
	.w6(32'h3abf28ed),
	.w7(32'h3aacacb7),
	.w8(32'h3ab31567),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25c067),
	.w1(32'h3a280f73),
	.w2(32'hbb61c0f9),
	.w3(32'hb9803009),
	.w4(32'h3a43d221),
	.w5(32'hbba27ebb),
	.w6(32'hbb790df3),
	.w7(32'h3c215dec),
	.w8(32'hbc26cc95),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e6e7fd),
	.w1(32'h39f96a32),
	.w2(32'hbbd22ee0),
	.w3(32'h3c1b4f5d),
	.w4(32'h3b79c321),
	.w5(32'hba939c5f),
	.w6(32'h3c02b1f5),
	.w7(32'h3a894c29),
	.w8(32'hbae24aa3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830a20),
	.w1(32'h3883615f),
	.w2(32'h398fb8a7),
	.w3(32'h3c147cd0),
	.w4(32'hbb11496c),
	.w5(32'h3a6d6f5f),
	.w6(32'h39df149c),
	.w7(32'h3c9e81a4),
	.w8(32'hbb37e6ef),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d08ff),
	.w1(32'hbbd862f5),
	.w2(32'h3acae0f6),
	.w3(32'h3a24e96a),
	.w4(32'hbc34dce7),
	.w5(32'h3b9cd083),
	.w6(32'h3b4eb4a8),
	.w7(32'h3b92f243),
	.w8(32'hbc980cf1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f34b),
	.w1(32'h3b91235a),
	.w2(32'h3b9f0eef),
	.w3(32'hbc942939),
	.w4(32'hbb966ed3),
	.w5(32'hbb68c45a),
	.w6(32'hbc28ec89),
	.w7(32'h3c4ad749),
	.w8(32'h3c131c9e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f848a),
	.w1(32'h3bad0b36),
	.w2(32'hbb2a4352),
	.w3(32'hbbce37be),
	.w4(32'hbc2bb91d),
	.w5(32'hbb129735),
	.w6(32'h3b9fe6e7),
	.w7(32'hbb72e7c8),
	.w8(32'h3c4a0898),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a954781),
	.w1(32'hba8bbe31),
	.w2(32'h379466b9),
	.w3(32'h3a11dcf8),
	.w4(32'h3bd92176),
	.w5(32'h3b395d15),
	.w6(32'hbc4e563e),
	.w7(32'h3703e0a6),
	.w8(32'h3b2c8f9f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a83eb),
	.w1(32'hbc1f5284),
	.w2(32'hbaab51b9),
	.w3(32'h3c603fab),
	.w4(32'hbb8426ee),
	.w5(32'hbc7a739c),
	.w6(32'h3c0dc467),
	.w7(32'h3b6e5925),
	.w8(32'h3cd6bfed),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6fbdd),
	.w1(32'hbc1262ad),
	.w2(32'hbb025722),
	.w3(32'h3c5c7c10),
	.w4(32'hbc545940),
	.w5(32'hbb8b6e55),
	.w6(32'hbc533df5),
	.w7(32'hbc1340cb),
	.w8(32'hbb9e5e8a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca561d9),
	.w1(32'hbc034c8c),
	.w2(32'h3c235966),
	.w3(32'hbc8c8572),
	.w4(32'hbb873668),
	.w5(32'h3a7c5e2a),
	.w6(32'h3d12654e),
	.w7(32'hbb56647c),
	.w8(32'hbc9a66a8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0d71f),
	.w1(32'hba2ec980),
	.w2(32'h3c2e9511),
	.w3(32'h3bafb802),
	.w4(32'h3c553830),
	.w5(32'hbb9a17d0),
	.w6(32'h3c820469),
	.w7(32'h3c2ce6e0),
	.w8(32'h3c09a675),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3575ca),
	.w1(32'hba279f01),
	.w2(32'hbab2f723),
	.w3(32'hbbd57ecb),
	.w4(32'hbb094542),
	.w5(32'hbab1e3cd),
	.w6(32'hbb11727c),
	.w7(32'hbb88be77),
	.w8(32'h3abc4498),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd38a),
	.w1(32'h3b9fe5f2),
	.w2(32'h3b9917e1),
	.w3(32'h3cab3dbb),
	.w4(32'h3b5cbe2e),
	.w5(32'hba364a3f),
	.w6(32'hbc10a4cd),
	.w7(32'hbb770b4a),
	.w8(32'hbb31c006),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule