module layer_10_featuremap_91(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b82393),
	.w1(32'hbab4fc7e),
	.w2(32'hbaba0e96),
	.w3(32'hbabd9882),
	.w4(32'h3b9e728b),
	.w5(32'hbb825958),
	.w6(32'hbbf82abb),
	.w7(32'h3bab20aa),
	.w8(32'h3aa7f1bc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcda320),
	.w1(32'hbb4730ea),
	.w2(32'h3ae9c47c),
	.w3(32'h389e9109),
	.w4(32'hba87d515),
	.w5(32'hba753eda),
	.w6(32'h394ea882),
	.w7(32'h3b27730a),
	.w8(32'hb9b5fead),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8dc89),
	.w1(32'hbb4e1566),
	.w2(32'h3bed4abe),
	.w3(32'hbb1ac313),
	.w4(32'h3ba9b239),
	.w5(32'hbb2a5ed6),
	.w6(32'hbc6ca522),
	.w7(32'h3a3d08f1),
	.w8(32'h3a8f05c3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180e4e),
	.w1(32'h3b807d1e),
	.w2(32'h3b362a6a),
	.w3(32'hb8f034ea),
	.w4(32'h3b75725b),
	.w5(32'hba000fc4),
	.w6(32'h3ae5ce47),
	.w7(32'h3b1cd16c),
	.w8(32'hbb1e0fb5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52e5c3),
	.w1(32'h3a7e28b1),
	.w2(32'h3b4f0584),
	.w3(32'hb90e907d),
	.w4(32'hbab1c5a9),
	.w5(32'hbaa45f6f),
	.w6(32'h3bab0a13),
	.w7(32'hba7b2c47),
	.w8(32'h3c1180bf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2383ee),
	.w1(32'hbb71d674),
	.w2(32'hbb633ed8),
	.w3(32'hbaa5ce5f),
	.w4(32'h3b66e314),
	.w5(32'hbad02ee4),
	.w6(32'h3a9ed6fb),
	.w7(32'hbb4c1779),
	.w8(32'h3ab31086),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c53ddb),
	.w1(32'hb988baa1),
	.w2(32'hbb2faa0f),
	.w3(32'h3b3d17e0),
	.w4(32'hbc87f566),
	.w5(32'h3d2a4b08),
	.w6(32'h3a575979),
	.w7(32'hbb440113),
	.w8(32'h3b05e1d7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc5b78),
	.w1(32'h3aac5606),
	.w2(32'hbbe36f53),
	.w3(32'h3bd890f0),
	.w4(32'hbae20be7),
	.w5(32'hba270136),
	.w6(32'h3b203575),
	.w7(32'hba67dc23),
	.w8(32'h3b43daa1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e37ab),
	.w1(32'h3c83bbeb),
	.w2(32'hb9aa503e),
	.w3(32'hbaf91cfb),
	.w4(32'h3b0a732f),
	.w5(32'hbb575063),
	.w6(32'hbabbf898),
	.w7(32'hb9e3650b),
	.w8(32'h38451746),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f84df),
	.w1(32'h38c8258d),
	.w2(32'hbb41e7a5),
	.w3(32'hba4fa410),
	.w4(32'h39742eb2),
	.w5(32'hbaa5cce2),
	.w6(32'hbb0ed2c1),
	.w7(32'hbcaa53cc),
	.w8(32'hba9066d8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768638),
	.w1(32'hbb58c136),
	.w2(32'hb9cb9d51),
	.w3(32'hbb2583e6),
	.w4(32'hbbf443ae),
	.w5(32'hbb081a0c),
	.w6(32'hbaef856a),
	.w7(32'h39c31d07),
	.w8(32'h39d0791c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba988452),
	.w1(32'h39f0096d),
	.w2(32'h3c8b2778),
	.w3(32'hba18a405),
	.w4(32'h3b9b737c),
	.w5(32'hb9992817),
	.w6(32'h3b1ef696),
	.w7(32'hb87cc5ca),
	.w8(32'hbb9e4989),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af529ba),
	.w1(32'h3a3d2613),
	.w2(32'hba609ebc),
	.w3(32'h3a8720d5),
	.w4(32'hba72473d),
	.w5(32'h3b9bb582),
	.w6(32'h3a74fd56),
	.w7(32'h3af632c1),
	.w8(32'h3aecd211),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c815a47),
	.w1(32'h3b9dbc40),
	.w2(32'hbaea5530),
	.w3(32'h3a289fd0),
	.w4(32'hbc9e31a9),
	.w5(32'hbb53008a),
	.w6(32'hb9b43ed3),
	.w7(32'hb6a337d6),
	.w8(32'hbb335dec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba941),
	.w1(32'hba63f1a9),
	.w2(32'hba5ae7ac),
	.w3(32'hb8fc54ed),
	.w4(32'hb97366c6),
	.w5(32'hbb2db3dc),
	.w6(32'h3b4fb9fe),
	.w7(32'hbb0f590a),
	.w8(32'h3be400d8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6783c70),
	.w1(32'h3aa36cb3),
	.w2(32'h3aa5f1c4),
	.w3(32'h3d22efb1),
	.w4(32'hba5ea018),
	.w5(32'hba948189),
	.w6(32'hbaf5f921),
	.w7(32'hb98f20ca),
	.w8(32'h3be89b8a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83db15b),
	.w1(32'h3c587f81),
	.w2(32'h3b14cb38),
	.w3(32'hba2ea42a),
	.w4(32'hb79ae8b6),
	.w5(32'hbcaaa00d),
	.w6(32'h3a2493c8),
	.w7(32'hba85fb5b),
	.w8(32'h3a92ccd9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb310d6f),
	.w1(32'hbb638b58),
	.w2(32'hbb0b104a),
	.w3(32'hbb538479),
	.w4(32'hbb527d6a),
	.w5(32'hb9031a41),
	.w6(32'hbbd2ea51),
	.w7(32'h3bdc7e26),
	.w8(32'hbb343ebc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e94a),
	.w1(32'h3ba56052),
	.w2(32'h3b5adeaa),
	.w3(32'h3add4d7b),
	.w4(32'h3a955f4a),
	.w5(32'h3bb8ac88),
	.w6(32'h38483148),
	.w7(32'hbbca9e81),
	.w8(32'hba4ed012),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6612ea),
	.w1(32'h3b1a9560),
	.w2(32'hbbd2c557),
	.w3(32'hbb4204dc),
	.w4(32'h3a9b59dc),
	.w5(32'h3aec2f57),
	.w6(32'h3a6764bb),
	.w7(32'h3b31307d),
	.w8(32'hbb4f5b6e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60a5a7),
	.w1(32'hbac1817a),
	.w2(32'hbbe79706),
	.w3(32'h3a8a3059),
	.w4(32'hb88a5297),
	.w5(32'h3a4bd607),
	.w6(32'h3cbc7f03),
	.w7(32'hba3c1695),
	.w8(32'hbb07a887),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b10a7),
	.w1(32'h3a87cc5c),
	.w2(32'h3a876e7d),
	.w3(32'h3a361aba),
	.w4(32'hb9386384),
	.w5(32'hbafa50af),
	.w6(32'h3b47dc00),
	.w7(32'hb932b0a5),
	.w8(32'hba935bbb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b335d22),
	.w1(32'hb9afeae5),
	.w2(32'hbca6360c),
	.w3(32'h3a785449),
	.w4(32'hbae28aeb),
	.w5(32'hbb311efa),
	.w6(32'hbb00605e),
	.w7(32'hba168a3c),
	.w8(32'hbc02b20c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9908ba9),
	.w1(32'hbbd497ac),
	.w2(32'hba91fc63),
	.w3(32'hba28e610),
	.w4(32'h3ab2a2cf),
	.w5(32'h3b64160e),
	.w6(32'hb9e07886),
	.w7(32'hba5b06fe),
	.w8(32'h3a649e69),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae49c7c),
	.w1(32'h3ad96b4b),
	.w2(32'h3b88bba9),
	.w3(32'hbaeceab2),
	.w4(32'h3acb3b95),
	.w5(32'h3af774d5),
	.w6(32'hba0f38d7),
	.w7(32'h3a5c7d35),
	.w8(32'hba060307),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04987f),
	.w1(32'h3aeeb564),
	.w2(32'h3b12d351),
	.w3(32'h3b062836),
	.w4(32'hbc67c998),
	.w5(32'hbab4924a),
	.w6(32'hbbe8d5c7),
	.w7(32'hba856014),
	.w8(32'hba674da1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24d963),
	.w1(32'h3ab81a46),
	.w2(32'hbc0bf8d7),
	.w3(32'h3b8e5136),
	.w4(32'h3b6d984b),
	.w5(32'hba2bd28a),
	.w6(32'hbb9727d2),
	.w7(32'hba9630cc),
	.w8(32'hbb481a8b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb830557),
	.w1(32'h39061655),
	.w2(32'hbc0af845),
	.w3(32'hbb2df1e1),
	.w4(32'h3b87b139),
	.w5(32'hbbf21c93),
	.w6(32'h3bf45101),
	.w7(32'h3d1782be),
	.w8(32'hbaa07185),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb98dd6),
	.w1(32'hbaf86b95),
	.w2(32'h3c45dfde),
	.w3(32'hba156be6),
	.w4(32'h3a9beda8),
	.w5(32'hbbdbce91),
	.w6(32'hb9b0c71d),
	.w7(32'hbb0c2ad2),
	.w8(32'h3b8ce2e0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c159),
	.w1(32'h37c8c333),
	.w2(32'hbac26ccd),
	.w3(32'h3b8343ee),
	.w4(32'h3c911b5a),
	.w5(32'hba16176a),
	.w6(32'hbb287c8f),
	.w7(32'hbba59cb6),
	.w8(32'hbc053ca5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63622),
	.w1(32'hba043f4f),
	.w2(32'h3b113cb9),
	.w3(32'hbab8f450),
	.w4(32'hbb4386fb),
	.w5(32'h3a2c1b34),
	.w6(32'h3b535d7d),
	.w7(32'h393908a6),
	.w8(32'h3c656899),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7af7),
	.w1(32'hbbcb0e40),
	.w2(32'h3aba40a5),
	.w3(32'hbbd48562),
	.w4(32'hbb02123c),
	.w5(32'hbba779fc),
	.w6(32'hbaf372e3),
	.w7(32'h3bfd9969),
	.w8(32'h3b6bf9f2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831f26),
	.w1(32'hbc0d1519),
	.w2(32'hbb51cb73),
	.w3(32'h3b672c29),
	.w4(32'h3ba302b1),
	.w5(32'h3a9a5c6b),
	.w6(32'h3ad59b48),
	.w7(32'hbbb0f46e),
	.w8(32'hb7f1d2d9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0ff95),
	.w1(32'h3c42b3a1),
	.w2(32'h3c18d39b),
	.w3(32'hbb141961),
	.w4(32'hbb3a5c9f),
	.w5(32'hba513251),
	.w6(32'hba52a402),
	.w7(32'hb9f84b4d),
	.w8(32'hbab055cf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac61902),
	.w1(32'hbb7347d3),
	.w2(32'hba1a8ed2),
	.w3(32'h3a2c6029),
	.w4(32'hb869f45c),
	.w5(32'hbbcb1ffe),
	.w6(32'hbb27af3b),
	.w7(32'h3b8481d4),
	.w8(32'hbc39effa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5db1b2),
	.w1(32'hba8c376a),
	.w2(32'h3a10df71),
	.w3(32'h3a552495),
	.w4(32'h3ac020cf),
	.w5(32'hbbcb2104),
	.w6(32'hbc3f08d7),
	.w7(32'h3bce01a2),
	.w8(32'hba31fb27),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865cd0),
	.w1(32'h3bd69aeb),
	.w2(32'hbbebdb41),
	.w3(32'hba6f51ab),
	.w4(32'h3c1d207a),
	.w5(32'hbcb33963),
	.w6(32'hbad79411),
	.w7(32'hbab879a8),
	.w8(32'hbc131bb2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba475391),
	.w1(32'h3a3bc836),
	.w2(32'hbb810925),
	.w3(32'hbaedf07e),
	.w4(32'h3c59759f),
	.w5(32'h3a5e68f8),
	.w6(32'h3b23f38a),
	.w7(32'hbb43870f),
	.w8(32'h3b81bdd8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fb49c),
	.w1(32'hbbb7b2a7),
	.w2(32'hbaf66bd7),
	.w3(32'h3b5f8c2b),
	.w4(32'hbb2c23b9),
	.w5(32'h3b39da6a),
	.w6(32'h3ba5928b),
	.w7(32'h3b481678),
	.w8(32'h3bc363cd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb275a4d),
	.w1(32'h3ac384bb),
	.w2(32'hb96e0ad5),
	.w3(32'hbbb901b5),
	.w4(32'h3c54bde6),
	.w5(32'h3c1a2107),
	.w6(32'h3cf1374d),
	.w7(32'hbc0375a7),
	.w8(32'h3c987661),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3765db2e),
	.w1(32'hbbf22283),
	.w2(32'h3b84bf52),
	.w3(32'h3c93da00),
	.w4(32'h3c20c8ff),
	.w5(32'hba7c8f5e),
	.w6(32'hb9281a59),
	.w7(32'hbbb9c1e8),
	.w8(32'h3b0b7d58),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07f33f),
	.w1(32'h3980b269),
	.w2(32'hbb97f8dd),
	.w3(32'hba93ce0d),
	.w4(32'hbbb60cc7),
	.w5(32'h3b81a1bb),
	.w6(32'h3b165ac3),
	.w7(32'h3adacf92),
	.w8(32'hbc5ea5d1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a9bce),
	.w1(32'h3b87ea73),
	.w2(32'hbc288a62),
	.w3(32'hba82a2c3),
	.w4(32'h3bbdc9ee),
	.w5(32'h3b8bfcac),
	.w6(32'hb8b07cef),
	.w7(32'hba32c9e4),
	.w8(32'h3b85c8a9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be04f7d),
	.w1(32'hbba0e96d),
	.w2(32'h3a5a2f01),
	.w3(32'hbb654237),
	.w4(32'h3b740404),
	.w5(32'hb9a02e3f),
	.w6(32'hbbd27537),
	.w7(32'hbbfe784d),
	.w8(32'hbb736e3b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fb62d),
	.w1(32'hbcc3962f),
	.w2(32'hbaf10af5),
	.w3(32'h3b531b5f),
	.w4(32'h3a6b4abe),
	.w5(32'hbbfbf9aa),
	.w6(32'h3afe8678),
	.w7(32'hbb03e67f),
	.w8(32'h39276f8c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac55a),
	.w1(32'h3b2f2bc5),
	.w2(32'hbb94b246),
	.w3(32'hbb8f1e68),
	.w4(32'hbb14c379),
	.w5(32'h3cd7c25a),
	.w6(32'h3c7af59b),
	.w7(32'h3af3c608),
	.w8(32'hbace0a73),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c69e48),
	.w1(32'hbb6a9d93),
	.w2(32'hb9cc95f8),
	.w3(32'h3cc9bdfc),
	.w4(32'h3a773b98),
	.w5(32'hbc9005f2),
	.w6(32'h38776a5b),
	.w7(32'hba36fa1c),
	.w8(32'h3943a0b7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b993797),
	.w1(32'hbb1a85ca),
	.w2(32'h3b95c4ab),
	.w3(32'h3aeedfee),
	.w4(32'h3c54bb2e),
	.w5(32'h3a039877),
	.w6(32'h3b87c057),
	.w7(32'hbb852962),
	.w8(32'h393c3b35),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107cba),
	.w1(32'h3b4d3339),
	.w2(32'hbc4d0621),
	.w3(32'hbb250ef0),
	.w4(32'hbb3289f7),
	.w5(32'hbb97ee96),
	.w6(32'h3ad29f4d),
	.w7(32'h3b783d2e),
	.w8(32'hbb73e239),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ce901),
	.w1(32'h3a9f83a7),
	.w2(32'hbb337c32),
	.w3(32'hbb2694ea),
	.w4(32'hbb7775b6),
	.w5(32'h3b88a689),
	.w6(32'h3b549333),
	.w7(32'hb891cbb6),
	.w8(32'hbafe57f9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994ec64),
	.w1(32'h3c1c24f0),
	.w2(32'hbaad22c4),
	.w3(32'hbb16103e),
	.w4(32'hb9975290),
	.w5(32'h38b64f2b),
	.w6(32'hbb0537d1),
	.w7(32'hbaecc995),
	.w8(32'h3b2b1f20),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a76ec),
	.w1(32'hbb52665e),
	.w2(32'hbaaba2cf),
	.w3(32'hbc8af58f),
	.w4(32'h3a83e901),
	.w5(32'hbbb7dcee),
	.w6(32'h3bcb6f5c),
	.w7(32'hbb272210),
	.w8(32'h3b763578),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4caba),
	.w1(32'hba29afec),
	.w2(32'hb9d35dbd),
	.w3(32'h3bba0206),
	.w4(32'hba70559d),
	.w5(32'h3b250f2b),
	.w6(32'h3a72daef),
	.w7(32'hbb8d2e3c),
	.w8(32'hbc0da5a3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa211a3),
	.w1(32'hbb89ae3e),
	.w2(32'h3ac413c9),
	.w3(32'h3b267802),
	.w4(32'hbb18a791),
	.w5(32'hbb760208),
	.w6(32'hbaab43a9),
	.w7(32'h3bdf13ab),
	.w8(32'h39ec1fbe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89165b),
	.w1(32'hbb684bb9),
	.w2(32'hbb68e671),
	.w3(32'hbb94521d),
	.w4(32'hba6d49bc),
	.w5(32'hbb272889),
	.w6(32'hbb3294bf),
	.w7(32'h3b27ee5a),
	.w8(32'h3a810ca9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe1c98),
	.w1(32'hbb9c30cc),
	.w2(32'hba542940),
	.w3(32'h3b6f3abc),
	.w4(32'hbc66249c),
	.w5(32'h3923a769),
	.w6(32'h3aa92f15),
	.w7(32'h3c0e6f45),
	.w8(32'hbba787ad),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09142d),
	.w1(32'hbb00349f),
	.w2(32'hbbb62712),
	.w3(32'hbc81c6e4),
	.w4(32'h3aade7e4),
	.w5(32'hbb92af34),
	.w6(32'h3c893d66),
	.w7(32'h3abfebf0),
	.w8(32'hbba05b30),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4024),
	.w1(32'h3b24e473),
	.w2(32'h3c105939),
	.w3(32'hbbc5b57e),
	.w4(32'h39b85465),
	.w5(32'hbc292700),
	.w6(32'hbc2b5c17),
	.w7(32'h39d7ad43),
	.w8(32'hbb17b7a6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48db1a),
	.w1(32'hbc3bae05),
	.w2(32'h3b7dcbe6),
	.w3(32'h3b77907a),
	.w4(32'h39b02e72),
	.w5(32'h3b107ace),
	.w6(32'hbc0ba882),
	.w7(32'hb7ed91bb),
	.w8(32'hbacea5fb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e8a6),
	.w1(32'hba97174a),
	.w2(32'hbbc5a0fd),
	.w3(32'hbbd1a629),
	.w4(32'hbb5e3aa6),
	.w5(32'hba3538bf),
	.w6(32'h39e434f6),
	.w7(32'h39b0ec20),
	.w8(32'h3c1db965),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac53f2a),
	.w1(32'h3acc5f25),
	.w2(32'hbb730e20),
	.w3(32'h3891e46e),
	.w4(32'hbc39bab3),
	.w5(32'hbb579481),
	.w6(32'h3b2361fa),
	.w7(32'h3b0db4a9),
	.w8(32'h3be52bfe),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd7573),
	.w1(32'hbba01476),
	.w2(32'hba212988),
	.w3(32'hbc07d11d),
	.w4(32'h3bcb3c29),
	.w5(32'h3c084982),
	.w6(32'h3b625fb9),
	.w7(32'h3bf45815),
	.w8(32'h3b1ccc1f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c61049),
	.w1(32'hbb20991b),
	.w2(32'hbac08b15),
	.w3(32'hbc454611),
	.w4(32'h3aa855cc),
	.w5(32'hb7b7d242),
	.w6(32'h391ef4e4),
	.w7(32'hbbbd19c9),
	.w8(32'h3c02f732),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ba69),
	.w1(32'hbc7d35a4),
	.w2(32'hba62e5ea),
	.w3(32'hbbc81f97),
	.w4(32'hbbbee4d3),
	.w5(32'h3d5b40e8),
	.w6(32'h3c1f69b8),
	.w7(32'h3a0387d3),
	.w8(32'hbcabdf1e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e8afd),
	.w1(32'h3b9df544),
	.w2(32'h3b7ef27c),
	.w3(32'hbc1bd70a),
	.w4(32'h3a341124),
	.w5(32'h3c8d8e3f),
	.w6(32'h3ac9e99d),
	.w7(32'h3c4ecdda),
	.w8(32'hbba0ea23),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9d738),
	.w1(32'h3bf02a36),
	.w2(32'h3b96fdde),
	.w3(32'hbb992e60),
	.w4(32'h3a8d6f10),
	.w5(32'h36144722),
	.w6(32'hb93abeea),
	.w7(32'h3c18f015),
	.w8(32'hbbd7fafe),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7cf34),
	.w1(32'h3b7cd98d),
	.w2(32'hbc11070b),
	.w3(32'hbb30dc1e),
	.w4(32'h3b92ea06),
	.w5(32'hba8ebde5),
	.w6(32'h38c0de84),
	.w7(32'hbb6049e1),
	.w8(32'hbbb5668b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e5bdd),
	.w1(32'h3d0ffd55),
	.w2(32'hbcd93322),
	.w3(32'h3bbd08bc),
	.w4(32'hbb7a3285),
	.w5(32'hb98b8e76),
	.w6(32'hbaeda027),
	.w7(32'hbaaf22ec),
	.w8(32'hb993889c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ea023),
	.w1(32'h3c47168e),
	.w2(32'hba53b36f),
	.w3(32'h39b3af18),
	.w4(32'hb9c217dd),
	.w5(32'h3c441a5f),
	.w6(32'hbb1d7ec7),
	.w7(32'h3ba1be1c),
	.w8(32'h3badfa8f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc985),
	.w1(32'hbb61c95c),
	.w2(32'hbc3859d8),
	.w3(32'hbc44a33e),
	.w4(32'hba49a4d5),
	.w5(32'h3b811e3e),
	.w6(32'hbb894665),
	.w7(32'h3b99e461),
	.w8(32'h3b5e08a2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbb4be),
	.w1(32'h3c4e15c4),
	.w2(32'hbadf94fd),
	.w3(32'hbc5b541f),
	.w4(32'h3c8a7ad6),
	.w5(32'hbbfded5e),
	.w6(32'h3a03a672),
	.w7(32'h3bb57b98),
	.w8(32'hbc45efcd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410508),
	.w1(32'h3b823f9e),
	.w2(32'h397250b0),
	.w3(32'h3c216c00),
	.w4(32'hbbe6cfd7),
	.w5(32'hbc2b4b44),
	.w6(32'hba66b460),
	.w7(32'hbaff3ff3),
	.w8(32'hbc5c046d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0127a0),
	.w1(32'hbbdc8764),
	.w2(32'hbc01ffd6),
	.w3(32'hba682ce4),
	.w4(32'hbae5a905),
	.w5(32'h3ab3cb20),
	.w6(32'hbb25703c),
	.w7(32'h3b10a7ff),
	.w8(32'hb9c76112),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a3d15),
	.w1(32'hb8976b1c),
	.w2(32'hba9176cd),
	.w3(32'hbb975d59),
	.w4(32'hbb6e974e),
	.w5(32'hbc04e596),
	.w6(32'h3c88e805),
	.w7(32'hbbda3f82),
	.w8(32'hba1f9408),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525569),
	.w1(32'h3b5baeec),
	.w2(32'hb949c796),
	.w3(32'hbb1161cf),
	.w4(32'h3c54c954),
	.w5(32'hbb9730dd),
	.w6(32'hbc4a32ff),
	.w7(32'h3c04bb7f),
	.w8(32'h380ddd9e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b165a76),
	.w1(32'hbc2675e5),
	.w2(32'hbc7af354),
	.w3(32'hbba1f40e),
	.w4(32'hbb1169d0),
	.w5(32'hbb7e05fb),
	.w6(32'hbca35966),
	.w7(32'hbbc701fa),
	.w8(32'hbcc1c2b1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe95c5),
	.w1(32'hbb274b83),
	.w2(32'h3a982512),
	.w3(32'hb87caf49),
	.w4(32'hbb6cc2ff),
	.w5(32'hbbed67e2),
	.w6(32'hbad120e3),
	.w7(32'hb8d3eab6),
	.w8(32'h3b91333a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e85f7),
	.w1(32'h3bc7a94a),
	.w2(32'h3c37cb2d),
	.w3(32'hbcb5b84a),
	.w4(32'hbb11164b),
	.w5(32'hbb506e92),
	.w6(32'hbbbafc49),
	.w7(32'hbcbab6ed),
	.w8(32'h3cbc4a9e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41871),
	.w1(32'h3b0087cc),
	.w2(32'hbaafe658),
	.w3(32'hbab8129d),
	.w4(32'hb98bb676),
	.w5(32'hbb03c0a1),
	.w6(32'hbb4f1736),
	.w7(32'hbbffa40e),
	.w8(32'hbb2fd9c0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c7a32),
	.w1(32'hbb4af264),
	.w2(32'hbd04e413),
	.w3(32'h3abaa8e4),
	.w4(32'h3b75892c),
	.w5(32'h3b18aa9f),
	.w6(32'h3ac2c376),
	.w7(32'hbc087aad),
	.w8(32'hbb206434),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33c819),
	.w1(32'h3af4a2b9),
	.w2(32'h3b21dfcb),
	.w3(32'h3b1e095f),
	.w4(32'hbb3bb64e),
	.w5(32'hbb262c22),
	.w6(32'hb9299dfb),
	.w7(32'h3b9a9bec),
	.w8(32'hbb0cef7e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0221be),
	.w1(32'hbb9fda13),
	.w2(32'hbb8ae372),
	.w3(32'h3bbce14e),
	.w4(32'hba1e8215),
	.w5(32'hbc682e5b),
	.w6(32'hbbc3188e),
	.w7(32'h3a685b6e),
	.w8(32'h3c938087),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa6808),
	.w1(32'hbca9a593),
	.w2(32'h3a979179),
	.w3(32'h3be1debf),
	.w4(32'h39a8e727),
	.w5(32'hbbd63a95),
	.w6(32'h3b1bb737),
	.w7(32'h3c8eb29a),
	.w8(32'h3b79bf3e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79ca09),
	.w1(32'h3a1dfab5),
	.w2(32'hb966a72f),
	.w3(32'h39deae08),
	.w4(32'h3a2cb692),
	.w5(32'hb9d5dcc8),
	.w6(32'h3ae9bc88),
	.w7(32'h3a8f8684),
	.w8(32'hbb48c345),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9eb16),
	.w1(32'h3b2b254d),
	.w2(32'h3d185f79),
	.w3(32'h39dbf235),
	.w4(32'hba2499b8),
	.w5(32'h3a9d86ee),
	.w6(32'hbb49f98a),
	.w7(32'h3910ce6a),
	.w8(32'hbb6cb4fc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0018a0),
	.w1(32'h398122d0),
	.w2(32'h3b6137ef),
	.w3(32'hbb6a2fc6),
	.w4(32'hba287f42),
	.w5(32'h38d43c85),
	.w6(32'h39332e50),
	.w7(32'hbd16ccbe),
	.w8(32'hbb067533),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0b7dc),
	.w1(32'hbd0eacd1),
	.w2(32'h3b1d8460),
	.w3(32'h3b19ce08),
	.w4(32'hba6d28e7),
	.w5(32'hbb3bbb9b),
	.w6(32'h3ac0a625),
	.w7(32'hb9cecfb3),
	.w8(32'hbb0f885f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9b7bb),
	.w1(32'h3b08720b),
	.w2(32'hbae3f456),
	.w3(32'h38b6242b),
	.w4(32'h3b347c7c),
	.w5(32'h3aa5e3d0),
	.w6(32'h3b477702),
	.w7(32'h3aaa32d5),
	.w8(32'hba6c7e6f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabdc58),
	.w1(32'h3abba177),
	.w2(32'hbb0f7d04),
	.w3(32'h3aa7ed75),
	.w4(32'hbac9c73f),
	.w5(32'h3abd7745),
	.w6(32'h3a4644fc),
	.w7(32'hbad4b5b7),
	.w8(32'hbb1ff4e1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fa8f6),
	.w1(32'h3b16dc09),
	.w2(32'hbb925fb8),
	.w3(32'hb9319a5b),
	.w4(32'hbb61bc17),
	.w5(32'hbab782b1),
	.w6(32'h3ad8628a),
	.w7(32'hbb1e89a5),
	.w8(32'hb9c9938a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f8f8e),
	.w1(32'h3abcd8a0),
	.w2(32'hb9db95f9),
	.w3(32'h39148b10),
	.w4(32'hb9eac2bc),
	.w5(32'hbb1490bc),
	.w6(32'hbc5563ec),
	.w7(32'hbc3289f0),
	.w8(32'h391c3e7a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edf6e2),
	.w1(32'h3af2dc7a),
	.w2(32'h3ad52daf),
	.w3(32'h3a7aca09),
	.w4(32'h3b9aa8ab),
	.w5(32'h3bd3ebd7),
	.w6(32'h39efeaa4),
	.w7(32'hbadb38a8),
	.w8(32'hba9af2b5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b85703),
	.w1(32'h3b4a49ff),
	.w2(32'h3bbef51f),
	.w3(32'h3b8f5a59),
	.w4(32'hbb8354dc),
	.w5(32'hbb0175df),
	.w6(32'h3c801ba5),
	.w7(32'hbb935e05),
	.w8(32'h3b8d5d55),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f983d),
	.w1(32'hbc414d59),
	.w2(32'h3c433129),
	.w3(32'h3a859d5b),
	.w4(32'h3ba2d29c),
	.w5(32'hba0e7342),
	.w6(32'hba3068a9),
	.w7(32'h3b1ef8f7),
	.w8(32'hba683a14),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3859ac),
	.w1(32'hbb94092c),
	.w2(32'hb8d9cdfa),
	.w3(32'h3b217d20),
	.w4(32'h3aa2d714),
	.w5(32'hbafbc1b9),
	.w6(32'h39084d45),
	.w7(32'hb884469f),
	.w8(32'hbb82b0fe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc3580),
	.w1(32'h39b6f70f),
	.w2(32'hba7303bd),
	.w3(32'h39fc8c2a),
	.w4(32'h3b40e99f),
	.w5(32'h3c78bc8d),
	.w6(32'h3badb36f),
	.w7(32'h3ba16200),
	.w8(32'hba014ef6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a224987),
	.w1(32'hbd01c654),
	.w2(32'h3b086104),
	.w3(32'hbd429f28),
	.w4(32'h3b11fe56),
	.w5(32'h3a91ef21),
	.w6(32'hba203f86),
	.w7(32'h3a4761a1),
	.w8(32'h37d9bda5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bd10e),
	.w1(32'hb952ccfb),
	.w2(32'hbb091212),
	.w3(32'hb9ca4161),
	.w4(32'h3acc4dfb),
	.w5(32'hbaac638c),
	.w6(32'h3aaf6cad),
	.w7(32'h3aa55efd),
	.w8(32'h3b4b0aab),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e94edf),
	.w1(32'h3d0a99c2),
	.w2(32'hbbac829e),
	.w3(32'hba195194),
	.w4(32'h3b65b9ce),
	.w5(32'h3c0a3ced),
	.w6(32'hb993c2fe),
	.w7(32'h39aa9c62),
	.w8(32'h3d260feb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39327b46),
	.w1(32'h39626c17),
	.w2(32'hb91955cb),
	.w3(32'h3a50cb1f),
	.w4(32'hbaa3e060),
	.w5(32'hba2d45b2),
	.w6(32'h39311daa),
	.w7(32'h3aff5f43),
	.w8(32'h3ad4be91),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fedf6),
	.w1(32'hbb28de86),
	.w2(32'hba78a0f5),
	.w3(32'h3a912e33),
	.w4(32'hbb77b582),
	.w5(32'h39ae9cd9),
	.w6(32'hbae3219e),
	.w7(32'hbaaeb67c),
	.w8(32'hba7faa86),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6f2a7),
	.w1(32'h3ad5c599),
	.w2(32'h3d1363c3),
	.w3(32'h3b4413cb),
	.w4(32'hba75f421),
	.w5(32'h392c6cf3),
	.w6(32'h3cc6a48b),
	.w7(32'hba407cdf),
	.w8(32'hb988ab74),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3713e),
	.w1(32'hbb2f9360),
	.w2(32'hbd24a697),
	.w3(32'hbc422bd3),
	.w4(32'hbaeff1ce),
	.w5(32'h3a556f3e),
	.w6(32'h3af8166f),
	.w7(32'h3af277c5),
	.w8(32'hbc3b826b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb43007),
	.w1(32'h3bef40b6),
	.w2(32'hbcbc7f2d),
	.w3(32'hb7f84e72),
	.w4(32'h3911682d),
	.w5(32'h39654dfd),
	.w6(32'hbaac53c0),
	.w7(32'hba751c04),
	.w8(32'h3b501783),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d406f),
	.w1(32'hbd10bb02),
	.w2(32'hbaadd792),
	.w3(32'h3bbfafeb),
	.w4(32'h3b07da06),
	.w5(32'h3ba168df),
	.w6(32'hb89cb07d),
	.w7(32'h3a439cc5),
	.w8(32'hbb1432d9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5978),
	.w1(32'h3b5a3501),
	.w2(32'hb982b4c1),
	.w3(32'h3b09ece9),
	.w4(32'hb98b0b40),
	.w5(32'h3af70ad2),
	.w6(32'hb8a3c346),
	.w7(32'hbc08bab1),
	.w8(32'h3a29a339),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e90d),
	.w1(32'h3c3d93c1),
	.w2(32'h3b3cdf53),
	.w3(32'h3b060207),
	.w4(32'hb9628b05),
	.w5(32'hb90800af),
	.w6(32'h3ba72b59),
	.w7(32'hbab5222a),
	.w8(32'hb99c667c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec6662),
	.w1(32'hba04beeb),
	.w2(32'h398c121a),
	.w3(32'hb8dd4099),
	.w4(32'h3b12b898),
	.w5(32'hbacc6339),
	.w6(32'h3a0f526f),
	.w7(32'hb9cea23e),
	.w8(32'h3adabd8b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba590188),
	.w1(32'hbaa34f08),
	.w2(32'h3a34e33a),
	.w3(32'hbc4a91f1),
	.w4(32'hb9d04b9c),
	.w5(32'hba301883),
	.w6(32'h3a9b46f4),
	.w7(32'hbb2e0bf2),
	.w8(32'hbb158f5b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46dd6),
	.w1(32'hb9061eca),
	.w2(32'hbb299235),
	.w3(32'hb99898a3),
	.w4(32'h3a1800af),
	.w5(32'h3bf4d3d6),
	.w6(32'hb991aded),
	.w7(32'h37dfefc2),
	.w8(32'h3ac6886b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc9f26),
	.w1(32'h3b8286d3),
	.w2(32'h3b42b722),
	.w3(32'h3ab84712),
	.w4(32'hbb89f528),
	.w5(32'h3bea7e1a),
	.w6(32'h3b60d424),
	.w7(32'h3c09f538),
	.w8(32'h3ab9122a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b170e63),
	.w1(32'hba986169),
	.w2(32'h3b235a66),
	.w3(32'h3b6f57a9),
	.w4(32'hbb4ea904),
	.w5(32'hbafcb515),
	.w6(32'h3ae1eca4),
	.w7(32'h3b6ade81),
	.w8(32'h3ae268be),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8e68),
	.w1(32'hba9cee2a),
	.w2(32'hbacd0267),
	.w3(32'h3b39c6c7),
	.w4(32'hb9b0a544),
	.w5(32'h3abbf097),
	.w6(32'hbaa9e84e),
	.w7(32'hbae182be),
	.w8(32'hbc1ed11d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c3990),
	.w1(32'h38d46761),
	.w2(32'hbb80eb7a),
	.w3(32'h3cc68cd1),
	.w4(32'hbb04a3d6),
	.w5(32'hb9a1f77f),
	.w6(32'h3a19f9a6),
	.w7(32'hbbaef91e),
	.w8(32'hbac3b142),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d41d6),
	.w1(32'hba259697),
	.w2(32'h3a23a015),
	.w3(32'h3a36c753),
	.w4(32'h3ac42c67),
	.w5(32'hbc8065c9),
	.w6(32'h3a82a688),
	.w7(32'h3a386fbf),
	.w8(32'h3a57e1ca),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cb6fb2),
	.w1(32'h3aa24575),
	.w2(32'hbb40b067),
	.w3(32'hbb0ec5b2),
	.w4(32'h3b21d132),
	.w5(32'hbb4e1ea5),
	.w6(32'h3a80c5c7),
	.w7(32'hb9a2e013),
	.w8(32'h38cb82fc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba246a8),
	.w1(32'hb9ca1726),
	.w2(32'h3a57896e),
	.w3(32'h387dfd66),
	.w4(32'hbb706946),
	.w5(32'h39c7c6b2),
	.w6(32'hbb189899),
	.w7(32'h38dcbb60),
	.w8(32'h3b297c4b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b50751),
	.w1(32'h3a28461f),
	.w2(32'hb9bc4be2),
	.w3(32'hbb946297),
	.w4(32'h39268ef1),
	.w5(32'h3b3962af),
	.w6(32'hb8f4af71),
	.w7(32'h3b18cc83),
	.w8(32'h39e5fde4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa36821),
	.w1(32'hbb59dcb9),
	.w2(32'hbc353474),
	.w3(32'hb8bc3270),
	.w4(32'hb93cdc21),
	.w5(32'hba4a35a8),
	.w6(32'hbb3a6f73),
	.w7(32'h3a305fe9),
	.w8(32'hba0d4004),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef75d),
	.w1(32'hbb2abe6b),
	.w2(32'h3ae6675a),
	.w3(32'hba76c11e),
	.w4(32'hb8452033),
	.w5(32'hb74f2e3e),
	.w6(32'h3a2e0b25),
	.w7(32'h39aef9fb),
	.w8(32'hb9d1f8ed),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb569991),
	.w1(32'hba5b0f6c),
	.w2(32'h3b271f11),
	.w3(32'h399b5f6f),
	.w4(32'hb9271fbf),
	.w5(32'h3b1cef3b),
	.w6(32'h3b3b8b60),
	.w7(32'h3c971d15),
	.w8(32'hbb4caf85),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76bc55),
	.w1(32'h3b13018b),
	.w2(32'h3ad956ee),
	.w3(32'hba50504f),
	.w4(32'hbae5360a),
	.w5(32'hbbdf8b52),
	.w6(32'hbb1863f7),
	.w7(32'h3a3c26be),
	.w8(32'h3a0c9113),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a4ef9),
	.w1(32'hbaba534d),
	.w2(32'h39542448),
	.w3(32'h3cadfae4),
	.w4(32'hbaf71bd5),
	.w5(32'hbb533c6c),
	.w6(32'hbb137fcd),
	.w7(32'hbb0b039a),
	.w8(32'hba896192),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87c2f),
	.w1(32'hbbc22472),
	.w2(32'hbb16aaef),
	.w3(32'hb85150be),
	.w4(32'h3adde4e7),
	.w5(32'h3ad414da),
	.w6(32'hba8f92f0),
	.w7(32'hb92697d6),
	.w8(32'hbad0aa6a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba399187),
	.w1(32'hbb1f8bd5),
	.w2(32'hba25cce5),
	.w3(32'hba9d88e1),
	.w4(32'hbaa6db6e),
	.w5(32'hbc5d71a9),
	.w6(32'hbb10c0b1),
	.w7(32'hbcb6ee4d),
	.w8(32'hb9b84dc9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992e5b9),
	.w1(32'hb660634c),
	.w2(32'h380164c1),
	.w3(32'hb9d8e959),
	.w4(32'hbab6fe1b),
	.w5(32'hb9418793),
	.w6(32'h3b4f8b54),
	.w7(32'h380871f8),
	.w8(32'hbb14cfa0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4d12e),
	.w1(32'hbb044300),
	.w2(32'h3a2375bf),
	.w3(32'hbb12bf52),
	.w4(32'hbb44d64a),
	.w5(32'h3d080bb4),
	.w6(32'hba0702c8),
	.w7(32'h3a5f6171),
	.w8(32'hbb1931fd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8f874),
	.w1(32'h3c50d78e),
	.w2(32'hba89dbda),
	.w3(32'hbb8fbbaf),
	.w4(32'hbb2b2140),
	.w5(32'h3ac7e7dd),
	.w6(32'h3b195625),
	.w7(32'h3afde82d),
	.w8(32'h39ed8e93),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2995e),
	.w1(32'h3a9b6585),
	.w2(32'h3a46ca18),
	.w3(32'hbab21d7b),
	.w4(32'hba85dff8),
	.w5(32'hbb2310a1),
	.w6(32'h3a144020),
	.w7(32'h3a8983d5),
	.w8(32'h3c37896b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e140f),
	.w1(32'h38596ac2),
	.w2(32'h3cb15241),
	.w3(32'hbac35de5),
	.w4(32'hb80fdb6a),
	.w5(32'hba27c25f),
	.w6(32'h397678a3),
	.w7(32'h39e016f2),
	.w8(32'hbb19733f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8897196),
	.w1(32'hb88b4c13),
	.w2(32'hb816de72),
	.w3(32'h3cf4aad5),
	.w4(32'hba928d45),
	.w5(32'hbb1730a9),
	.w6(32'hb90a6c13),
	.w7(32'hbc693e4a),
	.w8(32'hba232d7e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f2664),
	.w1(32'hbbef13ec),
	.w2(32'hb9eba191),
	.w3(32'hbc8804b3),
	.w4(32'hbc3f19bd),
	.w5(32'h3b7d7d1b),
	.w6(32'hba386581),
	.w7(32'h390a3b3c),
	.w8(32'hb9cb1336),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea622),
	.w1(32'h3b78e0b3),
	.w2(32'h39305295),
	.w3(32'hbab9a1cc),
	.w4(32'hbb7e81c4),
	.w5(32'hbbca484a),
	.w6(32'hbaacfd0b),
	.w7(32'hbbb9426f),
	.w8(32'hbab9e652),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0880f),
	.w1(32'hbb11dae0),
	.w2(32'hb8e630d1),
	.w3(32'h3b05f9fd),
	.w4(32'h3b0474ac),
	.w5(32'hbaaf100b),
	.w6(32'h3a2fc578),
	.w7(32'hba0e6e47),
	.w8(32'h3a794cbf),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad133e4),
	.w1(32'h3756ae68),
	.w2(32'hbad7717d),
	.w3(32'hbaffc08d),
	.w4(32'h3b5a0cb3),
	.w5(32'h3c286973),
	.w6(32'h3999de71),
	.w7(32'hba74299b),
	.w8(32'hba4f0e2c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7ee5a),
	.w1(32'hb7c35e9c),
	.w2(32'h39a6a328),
	.w3(32'h3b729b52),
	.w4(32'h3a85a6b1),
	.w5(32'hba47d710),
	.w6(32'h3a029739),
	.w7(32'hba54097d),
	.w8(32'h3993dfdd),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba934f21),
	.w1(32'hb9e50174),
	.w2(32'h3b831165),
	.w3(32'hb8f77dcc),
	.w4(32'hbb977888),
	.w5(32'h39ea4b86),
	.w6(32'hba2280bf),
	.w7(32'hbc8ec773),
	.w8(32'hba9dd737),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c3f6),
	.w1(32'hbb4ed2ed),
	.w2(32'hbac9d545),
	.w3(32'h3b291354),
	.w4(32'hbaf8605f),
	.w5(32'hba542f24),
	.w6(32'h398ce9db),
	.w7(32'hbaea5c97),
	.w8(32'hba74d46b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5577fc),
	.w1(32'hbb1aa112),
	.w2(32'hb8f3eef2),
	.w3(32'hba974de5),
	.w4(32'h3a34b1cc),
	.w5(32'hbb158326),
	.w6(32'hbb77e94a),
	.w7(32'h3a8d79ef),
	.w8(32'h3b653f30),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa96954),
	.w1(32'hba91c203),
	.w2(32'h3ac85ae2),
	.w3(32'hb8a77e2c),
	.w4(32'hbb05d618),
	.w5(32'h3aa85aa7),
	.w6(32'h3ba70316),
	.w7(32'h38e9d93b),
	.w8(32'h3b14ad52),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a345e),
	.w1(32'hbac6cd4c),
	.w2(32'hb98dafa2),
	.w3(32'h3af2943b),
	.w4(32'hbb93a44b),
	.w5(32'hba817cd1),
	.w6(32'hba39e96b),
	.w7(32'h3b673374),
	.w8(32'hba15a324),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f693b),
	.w1(32'hbc6328d0),
	.w2(32'h3a712fc0),
	.w3(32'hbb0aff4d),
	.w4(32'h3b59ec05),
	.w5(32'hbac33045),
	.w6(32'h3b6c3f64),
	.w7(32'h3cc2f13f),
	.w8(32'hbb33eea7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08982a),
	.w1(32'hb9eaa807),
	.w2(32'h3a6993dd),
	.w3(32'hbaf1857a),
	.w4(32'hbc3adc53),
	.w5(32'hbb0b5ac0),
	.w6(32'h38dcc062),
	.w7(32'hbad45772),
	.w8(32'hb9ed3c47),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53e26b),
	.w1(32'h3a79d278),
	.w2(32'hba523d2d),
	.w3(32'h39564e6a),
	.w4(32'hbad4ee83),
	.w5(32'h3ab3beda),
	.w6(32'hbc3e2a99),
	.w7(32'hbb7fce56),
	.w8(32'h3b2ec5e7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b7335),
	.w1(32'hbaae7ac9),
	.w2(32'hba8bc731),
	.w3(32'hba28740b),
	.w4(32'hbbf9f650),
	.w5(32'h3987e348),
	.w6(32'hbb178b1e),
	.w7(32'h398cc86b),
	.w8(32'h3a01b0eb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1188),
	.w1(32'h3b30a561),
	.w2(32'h3a5edf68),
	.w3(32'h3b540307),
	.w4(32'hba679afb),
	.w5(32'hb8c219d9),
	.w6(32'h3a21f6c7),
	.w7(32'hbba53c6c),
	.w8(32'h398fa56a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50c584),
	.w1(32'hba853ac5),
	.w2(32'hbab6f41f),
	.w3(32'h3ae1736d),
	.w4(32'h39ec4d34),
	.w5(32'h3a965635),
	.w6(32'h3b844eb1),
	.w7(32'hbb25121e),
	.w8(32'h3a4e97f3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6f377),
	.w1(32'hbaa99809),
	.w2(32'h3ad0038c),
	.w3(32'hbc4a6110),
	.w4(32'hbc26958d),
	.w5(32'hbb431660),
	.w6(32'hbb947fbf),
	.w7(32'hbb046b87),
	.w8(32'hbb0aeb29),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b7cae),
	.w1(32'h3acadbf8),
	.w2(32'h3aae9b7e),
	.w3(32'h3accc4ec),
	.w4(32'hba8b6532),
	.w5(32'hbb2e5aa2),
	.w6(32'h3974317e),
	.w7(32'h38e4945e),
	.w8(32'h3b39b22a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce93532),
	.w1(32'h393f54f6),
	.w2(32'hbb50eb0c),
	.w3(32'h3a2305c8),
	.w4(32'hbafce477),
	.w5(32'h3ad5d93a),
	.w6(32'h3a691e8d),
	.w7(32'hb940d167),
	.w8(32'hbb8ea6c8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4c603),
	.w1(32'h3b2a5173),
	.w2(32'hbacbf21b),
	.w3(32'h3b1a9133),
	.w4(32'h3ae13852),
	.w5(32'hba68e468),
	.w6(32'hbbe38a11),
	.w7(32'h3cbad26a),
	.w8(32'hbb9f187a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c52807),
	.w1(32'h3a341207),
	.w2(32'hbb6f5d7f),
	.w3(32'h3900038f),
	.w4(32'hbb82a01c),
	.w5(32'hbc11a793),
	.w6(32'hbb86d0e8),
	.w7(32'hb97a24cf),
	.w8(32'hbb208471),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43548a),
	.w1(32'hba8e92e9),
	.w2(32'hbbbf0e40),
	.w3(32'hba4c1e05),
	.w4(32'hba1769d5),
	.w5(32'hbae157f8),
	.w6(32'h3b07d3cf),
	.w7(32'hbaa4bff8),
	.w8(32'hba8cb3cb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab6bc1),
	.w1(32'hbb2279d9),
	.w2(32'h39c1a4b4),
	.w3(32'h39ca735f),
	.w4(32'h3a23f53e),
	.w5(32'hb487ea8f),
	.w6(32'hbc40e5b0),
	.w7(32'h3905744a),
	.w8(32'hba2475c8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390585a5),
	.w1(32'hbb0e85f2),
	.w2(32'h39cff5d9),
	.w3(32'hbafef0c7),
	.w4(32'h3ab0605d),
	.w5(32'h389348a4),
	.w6(32'h3b4926e5),
	.w7(32'hbab64fa8),
	.w8(32'hbb0df726),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75f1df),
	.w1(32'hb891bf78),
	.w2(32'h3a49c7ca),
	.w3(32'h3a7db765),
	.w4(32'h3abd25b1),
	.w5(32'h3c3f6614),
	.w6(32'h3d1bab11),
	.w7(32'hbb2f0ac7),
	.w8(32'h3a9d2095),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb3605),
	.w1(32'h3b2c5062),
	.w2(32'h39f66658),
	.w3(32'hbaaf4286),
	.w4(32'hbbc3778e),
	.w5(32'h3abced1a),
	.w6(32'h3ad252de),
	.w7(32'hbb241b5c),
	.w8(32'h3a7f43eb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4ac22),
	.w1(32'h3cb4062e),
	.w2(32'h39d39935),
	.w3(32'h3b490905),
	.w4(32'hbb18a269),
	.w5(32'h3a9a691c),
	.w6(32'hbb127157),
	.w7(32'hbaa589db),
	.w8(32'hbad5cf98),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94172c),
	.w1(32'hbb1a9667),
	.w2(32'hb89ee1d6),
	.w3(32'h3cc7f01e),
	.w4(32'h3a5d6d59),
	.w5(32'h3983a02b),
	.w6(32'hb993afaa),
	.w7(32'h3d05c775),
	.w8(32'hba2f355b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e877f),
	.w1(32'h38545dec),
	.w2(32'h3908c8aa),
	.w3(32'h3960234c),
	.w4(32'hbb2dd3f8),
	.w5(32'hbbc79058),
	.w6(32'hba899161),
	.w7(32'hbc8ac8c2),
	.w8(32'hbc330df1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39988503),
	.w1(32'hbacce8a8),
	.w2(32'hba9bede0),
	.w3(32'hb8810eb7),
	.w4(32'hbb316379),
	.w5(32'h3bb55a98),
	.w6(32'h3b7999bc),
	.w7(32'h3b4d9c9f),
	.w8(32'hbafcec30),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8826bd),
	.w1(32'hbb323615),
	.w2(32'hba072392),
	.w3(32'h3a5eae2c),
	.w4(32'h3a30baf3),
	.w5(32'hbb0916c8),
	.w6(32'hbb693d63),
	.w7(32'h3a9e0b59),
	.w8(32'h3a795c96),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f7b3),
	.w1(32'h3b150d3a),
	.w2(32'h3a69352f),
	.w3(32'h3b049865),
	.w4(32'h3c060653),
	.w5(32'h3a0e7849),
	.w6(32'hba91d41c),
	.w7(32'hbb01667f),
	.w8(32'h3986c55b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b62c79),
	.w1(32'hb91d80cf),
	.w2(32'hb9a84fe4),
	.w3(32'hba0fdd11),
	.w4(32'hb9aba4a1),
	.w5(32'hb980b1f2),
	.w6(32'h3c1eb79a),
	.w7(32'h3ba45ece),
	.w8(32'h39969b88),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8edde0),
	.w1(32'h3ab89f8f),
	.w2(32'h38ed268d),
	.w3(32'hb9308d86),
	.w4(32'hbb0c92fb),
	.w5(32'h371f79da),
	.w6(32'hbaaae885),
	.w7(32'hb8c23d50),
	.w8(32'hbbdf4908),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc536b91),
	.w1(32'hba933a43),
	.w2(32'h3a0b0ef7),
	.w3(32'h3b2557df),
	.w4(32'hbaa1426b),
	.w5(32'hbb89a13d),
	.w6(32'hba71e206),
	.w7(32'hb950f7cb),
	.w8(32'hba9a4195),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1308de),
	.w1(32'hbb066bc5),
	.w2(32'h3aa7c4a1),
	.w3(32'h3a638806),
	.w4(32'hb9e53fdc),
	.w5(32'hbb397775),
	.w6(32'hba87908b),
	.w7(32'hb9dd1500),
	.w8(32'h3a75a2c0),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf1ffb),
	.w1(32'h3ac1a1fe),
	.w2(32'h3b68d1f9),
	.w3(32'h3b1aa36f),
	.w4(32'hbb234469),
	.w5(32'hbac56cc1),
	.w6(32'hbb931f37),
	.w7(32'h3b7204fa),
	.w8(32'hbb8be9bd),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae92702),
	.w1(32'h3a5fd458),
	.w2(32'h3a39e332),
	.w3(32'h3b6edb0f),
	.w4(32'hba63a53c),
	.w5(32'hbab57ff1),
	.w6(32'h3a36585a),
	.w7(32'h3b06e904),
	.w8(32'hbb0ac75b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68ec5),
	.w1(32'hbb306d38),
	.w2(32'hbc09dc73),
	.w3(32'h3c2900a0),
	.w4(32'hb93f8dd9),
	.w5(32'hbc29b210),
	.w6(32'hbb810d51),
	.w7(32'hbadce4fc),
	.w8(32'h3b93a50a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867ac8),
	.w1(32'hba1d1761),
	.w2(32'hbb5b1404),
	.w3(32'h399d1e07),
	.w4(32'hbb8f85cd),
	.w5(32'h3b379965),
	.w6(32'hba875a34),
	.w7(32'h3b2b9f5c),
	.w8(32'h39795a36),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38387),
	.w1(32'h3c23bca2),
	.w2(32'h3b11ea5b),
	.w3(32'hbc32b414),
	.w4(32'hbb572038),
	.w5(32'hbb94e619),
	.w6(32'h3c315fab),
	.w7(32'h3acc3057),
	.w8(32'hbb280f8f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f40a),
	.w1(32'hba1a197c),
	.w2(32'hbb734a46),
	.w3(32'h3bb1feca),
	.w4(32'h3bb2f07a),
	.w5(32'hbb7d5616),
	.w6(32'hb9582ff3),
	.w7(32'hbab83812),
	.w8(32'h3d23f5d7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad02a2d),
	.w1(32'h39db0bdc),
	.w2(32'h3a6d43ad),
	.w3(32'h3c08d209),
	.w4(32'hbb1d64eb),
	.w5(32'hbc3eb396),
	.w6(32'hbbf58833),
	.w7(32'hbbee6b0b),
	.w8(32'hbaf2e15a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b636e9d),
	.w1(32'h3b15991f),
	.w2(32'h3bdcf946),
	.w3(32'h39e79926),
	.w4(32'h3af2afc3),
	.w5(32'hbb25f9b8),
	.w6(32'hba894a39),
	.w7(32'hbb96bb8f),
	.w8(32'hbbd34452),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fda87),
	.w1(32'h3b3e0250),
	.w2(32'hbb07de3c),
	.w3(32'h3b343d72),
	.w4(32'h37b5da39),
	.w5(32'hba67067f),
	.w6(32'hbaf775a3),
	.w7(32'h3b89704e),
	.w8(32'h3a0a60c5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84324d8),
	.w1(32'h39cc667e),
	.w2(32'h3afbb57f),
	.w3(32'hbb79536d),
	.w4(32'h3a185c35),
	.w5(32'h3a91b754),
	.w6(32'hbb8c69ec),
	.w7(32'hbb36551f),
	.w8(32'hbb98c39a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aa3be),
	.w1(32'hbad0cbb4),
	.w2(32'h3b9d7978),
	.w3(32'hbbb06195),
	.w4(32'h3bb54999),
	.w5(32'h3bb1a107),
	.w6(32'h3bdedd70),
	.w7(32'h3b20daed),
	.w8(32'hbb36b138),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab12277),
	.w1(32'hbb97c075),
	.w2(32'hbb64245a),
	.w3(32'hbb0cd0f8),
	.w4(32'h3b44ec7f),
	.w5(32'hbc0b7e20),
	.w6(32'h3a7a961a),
	.w7(32'hba40cc92),
	.w8(32'h37a2fc46),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe09e36),
	.w1(32'hbbb71570),
	.w2(32'hbd415ca3),
	.w3(32'hbc15e5c1),
	.w4(32'h3bac75a8),
	.w5(32'h3c217dc9),
	.w6(32'hbbb5e555),
	.w7(32'hb83e97b6),
	.w8(32'h3b071e20),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c1ad7f),
	.w1(32'h3aa3193b),
	.w2(32'hbbe2da91),
	.w3(32'hbb4816e0),
	.w4(32'h39d2db48),
	.w5(32'hbc1c780d),
	.w6(32'hbbd0cb51),
	.w7(32'hbc4ee1f1),
	.w8(32'h39c68399),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace5316),
	.w1(32'hbb949ebd),
	.w2(32'hbb34b9a2),
	.w3(32'h3bf8f4b7),
	.w4(32'hbae39879),
	.w5(32'hbb9dc042),
	.w6(32'h390fcd7b),
	.w7(32'h3b11abbf),
	.w8(32'hbb0c101e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadd857),
	.w1(32'hbd259e0f),
	.w2(32'h3a9be3f4),
	.w3(32'hbd1a3155),
	.w4(32'h3794b9a4),
	.w5(32'hbb147619),
	.w6(32'h363f72e8),
	.w7(32'h3a980244),
	.w8(32'hba17bd15),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb278b52),
	.w1(32'hbc6943cd),
	.w2(32'h3bc55f9f),
	.w3(32'h3b722b94),
	.w4(32'hbba93c26),
	.w5(32'h3aa1d8ce),
	.w6(32'hbc01e414),
	.w7(32'h3b294803),
	.w8(32'hbb94c094),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44247c),
	.w1(32'hbb9ec0a6),
	.w2(32'hbc40f151),
	.w3(32'h3d884190),
	.w4(32'h3b459dee),
	.w5(32'hba8fd511),
	.w6(32'h3c1065b8),
	.w7(32'h3ac76d4d),
	.w8(32'h3a21bf03),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe57eb2),
	.w1(32'h3b8cf36c),
	.w2(32'hbbb25c8c),
	.w3(32'h3b189a1b),
	.w4(32'h3a841feb),
	.w5(32'hbbdf41d1),
	.w6(32'hbb26db2a),
	.w7(32'hbac4b564),
	.w8(32'hba5aa2ad),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b751c36),
	.w1(32'hbc0de863),
	.w2(32'hbb84a5da),
	.w3(32'hbaf77fef),
	.w4(32'hbb8ceb4c),
	.w5(32'hb8ea0630),
	.w6(32'hb9e35180),
	.w7(32'h3baf6fb3),
	.w8(32'hbba5a790),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ff97d),
	.w1(32'hbc4a32d7),
	.w2(32'hbb78c88b),
	.w3(32'h373fc160),
	.w4(32'h3b192802),
	.w5(32'hbbe328da),
	.w6(32'h399d0dfe),
	.w7(32'hba473a8b),
	.w8(32'hbb939da4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103ccc),
	.w1(32'hbbef15e0),
	.w2(32'hba33a0fa),
	.w3(32'hb9b68563),
	.w4(32'h39d940b0),
	.w5(32'hbacc54ca),
	.w6(32'hbc4f6e53),
	.w7(32'hbb90f597),
	.w8(32'hb95941cd),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd2f8f),
	.w1(32'hbbc9eeed),
	.w2(32'hbb6f65c7),
	.w3(32'hbc022488),
	.w4(32'hbc8a8129),
	.w5(32'hbb854246),
	.w6(32'h3acfb7ba),
	.w7(32'h3c17a731),
	.w8(32'hbb94e561),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb30e),
	.w1(32'hbbc7b2ac),
	.w2(32'hbb77ed7e),
	.w3(32'hbc63acc0),
	.w4(32'hb9a88f2a),
	.w5(32'hba27cdc9),
	.w6(32'hbbd9895b),
	.w7(32'h3b521217),
	.w8(32'hbc1c15fd),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08f67),
	.w1(32'hbc23845d),
	.w2(32'hbba3b8d8),
	.w3(32'h3b4c7f46),
	.w4(32'h3ba678a1),
	.w5(32'hbb096996),
	.w6(32'hbc210826),
	.w7(32'hbb3523b7),
	.w8(32'hbb782417),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676dc7),
	.w1(32'h3ae80228),
	.w2(32'hbb5d719d),
	.w3(32'hbb054edd),
	.w4(32'hbaa6ebab),
	.w5(32'hbbdfacfe),
	.w6(32'hb8988044),
	.w7(32'hbb9debf4),
	.w8(32'hba5eea6f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab52f0),
	.w1(32'h3bf42f4c),
	.w2(32'hbb99fc8b),
	.w3(32'hbab1496f),
	.w4(32'h3c8a447c),
	.w5(32'h3910177b),
	.w6(32'h37f16c71),
	.w7(32'hbb07839b),
	.w8(32'h3aef22cd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fba51),
	.w1(32'h3b5f8e94),
	.w2(32'h3b74a239),
	.w3(32'h3b8ccf5e),
	.w4(32'hbb6305fc),
	.w5(32'h3b41f689),
	.w6(32'hbc806e75),
	.w7(32'h3adc2b0a),
	.w8(32'h3a2f532f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e76c),
	.w1(32'hbb25e1c9),
	.w2(32'hbbb41a95),
	.w3(32'hbbb7072d),
	.w4(32'hbba8e97f),
	.w5(32'h3b843bb2),
	.w6(32'hba893f00),
	.w7(32'h3bbbc8fb),
	.w8(32'h3b931c30),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f427),
	.w1(32'hbb84c5d7),
	.w2(32'h3b558538),
	.w3(32'h3c3d8163),
	.w4(32'hbba88563),
	.w5(32'h3c8f0874),
	.w6(32'hb9e5273c),
	.w7(32'hbbfea9e1),
	.w8(32'h3a4cfac5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57bfee),
	.w1(32'hbb98232f),
	.w2(32'hbb0cd8ee),
	.w3(32'h3b30110a),
	.w4(32'hba8b3ec5),
	.w5(32'h3b9097f6),
	.w6(32'hbbe16fac),
	.w7(32'hbb0305a7),
	.w8(32'h3b0eb4dc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac507c),
	.w1(32'hbbedde41),
	.w2(32'hba489a2c),
	.w3(32'hbc0bdbd0),
	.w4(32'h3c9efcf6),
	.w5(32'h3ac0319f),
	.w6(32'h3c3c3b29),
	.w7(32'h3a069c29),
	.w8(32'h3b87b56e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5977),
	.w1(32'hbc4069f2),
	.w2(32'hbb9544f7),
	.w3(32'h3b0297c6),
	.w4(32'hbabf468c),
	.w5(32'h3a83b893),
	.w6(32'hbbe4d098),
	.w7(32'hbb66b8ca),
	.w8(32'hbb0da88d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5a8cb),
	.w1(32'h3bcfbab6),
	.w2(32'hbb03d7e5),
	.w3(32'h3c97a4e4),
	.w4(32'hbb6cfe10),
	.w5(32'hba8f09b9),
	.w6(32'h3c1d53a7),
	.w7(32'h3a6b1d67),
	.w8(32'h3a9831ed),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbc458),
	.w1(32'hbb6820ca),
	.w2(32'hbb8f66e3),
	.w3(32'h3b44d019),
	.w4(32'h3a300924),
	.w5(32'h3abbbdb1),
	.w6(32'h3a940789),
	.w7(32'h3bf0f376),
	.w8(32'h39b2f8cf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fb612),
	.w1(32'h39f24f13),
	.w2(32'hba5fc3c6),
	.w3(32'h3b318b6d),
	.w4(32'h3b32ca34),
	.w5(32'hbae2a651),
	.w6(32'hbc303f0d),
	.w7(32'h3a9e50fd),
	.w8(32'h3aac7a48),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9843925),
	.w1(32'hbbbed089),
	.w2(32'hbb6f5c81),
	.w3(32'hbbb11240),
	.w4(32'h3b69a16c),
	.w5(32'h3a2cee06),
	.w6(32'hbc08975e),
	.w7(32'h3a6a3781),
	.w8(32'h3a0f4baf),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d95a),
	.w1(32'h3ca3a349),
	.w2(32'hbb253577),
	.w3(32'h3b0c7fe7),
	.w4(32'h3952b268),
	.w5(32'hbb4142e7),
	.w6(32'h389071fe),
	.w7(32'hbaff0c05),
	.w8(32'hbb000862),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1e20),
	.w1(32'h3bd9e47a),
	.w2(32'hba5c2a8b),
	.w3(32'hb9a091ec),
	.w4(32'h3c09a712),
	.w5(32'hbaad5eef),
	.w6(32'hba122760),
	.w7(32'h3cf82905),
	.w8(32'hbbf1b0d2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe84082),
	.w1(32'h3ae9deb2),
	.w2(32'hba24a53d),
	.w3(32'h3be1673b),
	.w4(32'h3b408aea),
	.w5(32'h3c356b19),
	.w6(32'h3b60a5ed),
	.w7(32'h3b7cbae7),
	.w8(32'hbb0973d6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96cec0),
	.w1(32'h3b4d0a7a),
	.w2(32'h3b1911f6),
	.w3(32'h3c98dc9a),
	.w4(32'hbc58589e),
	.w5(32'h3b8831da),
	.w6(32'hbba00343),
	.w7(32'h3b567304),
	.w8(32'hbbbec571),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb780ea1a),
	.w1(32'h3c2bce39),
	.w2(32'h3ba11d0f),
	.w3(32'hbc55c20a),
	.w4(32'h370ba19e),
	.w5(32'h3c4b630f),
	.w6(32'h3b984c0b),
	.w7(32'hbafeb005),
	.w8(32'hbb36fd81),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57df26),
	.w1(32'h3c1ec0d8),
	.w2(32'hbafde7f2),
	.w3(32'hbb12c6da),
	.w4(32'h3a4220c6),
	.w5(32'hbacda364),
	.w6(32'hbb4720fe),
	.w7(32'hbbfe42eb),
	.w8(32'hbbd76d4b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc25a),
	.w1(32'hbb16a2a6),
	.w2(32'hb6662fda),
	.w3(32'hba6ecbfa),
	.w4(32'h3992b747),
	.w5(32'hba897634),
	.w6(32'hbb74c73f),
	.w7(32'h3c0c549a),
	.w8(32'hb97cf03b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134e1c),
	.w1(32'hbb01107b),
	.w2(32'hbb12598c),
	.w3(32'h3b842b5f),
	.w4(32'hbb872287),
	.w5(32'h3b3c1474),
	.w6(32'h3b4df8dd),
	.w7(32'h3b3613f7),
	.w8(32'h3b31547f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394921),
	.w1(32'hb95443be),
	.w2(32'hbbefcd2d),
	.w3(32'hbcfdf9b6),
	.w4(32'hbb8a4f25),
	.w5(32'hbb1d7d15),
	.w6(32'hbb545a13),
	.w7(32'h3c11065d),
	.w8(32'h3bbf322a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a8b65),
	.w1(32'hb99165f6),
	.w2(32'hbb05ef96),
	.w3(32'hbb2fcdea),
	.w4(32'h39d6f148),
	.w5(32'hba4a6155),
	.w6(32'hbc30e0e7),
	.w7(32'h3b3bca44),
	.w8(32'hbb673eed),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9125e9),
	.w1(32'h3bd83b72),
	.w2(32'hbb722f87),
	.w3(32'h3b90b543),
	.w4(32'hba795cfa),
	.w5(32'h3b1373fb),
	.w6(32'hbcca7216),
	.w7(32'h3aa9ef03),
	.w8(32'h3c03e868),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd326424),
	.w1(32'h3a517e36),
	.w2(32'h3ac57bd7),
	.w3(32'h3b6ac7b1),
	.w4(32'hbbe74a40),
	.w5(32'h3b6377db),
	.w6(32'h3b23aefc),
	.w7(32'hb885fab7),
	.w8(32'h3bba7e45),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeb3fb),
	.w1(32'hbab38838),
	.w2(32'hbbd9fe2b),
	.w3(32'hbbbbfd30),
	.w4(32'h3d33832a),
	.w5(32'h3b04b3ff),
	.w6(32'hbb4a0940),
	.w7(32'h3bc066a2),
	.w8(32'h3a2655f2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad88b1c),
	.w1(32'hbadd9007),
	.w2(32'h3bd6144d),
	.w3(32'h3bb14baa),
	.w4(32'h3be31559),
	.w5(32'h3b91a913),
	.w6(32'h3b012747),
	.w7(32'h3b9fc57b),
	.w8(32'hbc50f88a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2577bc),
	.w1(32'hbb7b581e),
	.w2(32'hba9cea28),
	.w3(32'h3b9dd718),
	.w4(32'hbb862f9b),
	.w5(32'h3aa76825),
	.w6(32'h3b2fd22c),
	.w7(32'h3c8cd49c),
	.w8(32'hbb90e834),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af91c03),
	.w1(32'hbcbb6dd0),
	.w2(32'hba9c8050),
	.w3(32'hbac966ab),
	.w4(32'h3bb67f24),
	.w5(32'h3a8edcce),
	.w6(32'hbaf4c53c),
	.w7(32'hbab127cd),
	.w8(32'h3bc0ebff),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1271ba),
	.w1(32'hbad0221d),
	.w2(32'h39893b73),
	.w3(32'h3becadbf),
	.w4(32'h3b80db0e),
	.w5(32'hbb838b13),
	.w6(32'h3a79bc0a),
	.w7(32'hba8ef9a6),
	.w8(32'hbb3ddcc2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb611fde),
	.w1(32'h3a3b722b),
	.w2(32'h39481eaf),
	.w3(32'h3a78e541),
	.w4(32'hb97aa977),
	.w5(32'hbd193a3f),
	.w6(32'h3b72bd8f),
	.w7(32'h3aad8690),
	.w8(32'hbb2f11fe),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1f90e),
	.w1(32'hba8f8d9b),
	.w2(32'hbb2da5bd),
	.w3(32'h39d398d6),
	.w4(32'hbb8bafa5),
	.w5(32'h3a6fce07),
	.w6(32'hba2c8ce5),
	.w7(32'h3b04a120),
	.w8(32'hba2159f4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e960a),
	.w1(32'hbb918a8c),
	.w2(32'hbb806fe1),
	.w3(32'h3a016b73),
	.w4(32'hba4f7cb1),
	.w5(32'h3c15e0e0),
	.w6(32'hba9ee31a),
	.w7(32'h3b899f26),
	.w8(32'h3acccb6b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc57eec),
	.w1(32'hbbd3216a),
	.w2(32'h3b76fcd6),
	.w3(32'h3c4f85df),
	.w4(32'h3ac2c281),
	.w5(32'hbb319784),
	.w6(32'hbb4f09bc),
	.w7(32'hbb3d0f8a),
	.w8(32'h3b81145a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26ca69),
	.w1(32'hbb771f7a),
	.w2(32'hba5c486c),
	.w3(32'h3b437896),
	.w4(32'h3a8150de),
	.w5(32'h3aba5e6e),
	.w6(32'h3b9699a6),
	.w7(32'hb9ceecd7),
	.w8(32'h3c2fdfef),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f6783),
	.w1(32'h3b831cad),
	.w2(32'hbcab7793),
	.w3(32'hbb4c86d1),
	.w4(32'hbb0b71a0),
	.w5(32'h3b403efc),
	.w6(32'hba4df980),
	.w7(32'hbb996206),
	.w8(32'h3be90a79),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ea5a),
	.w1(32'hbab4e39e),
	.w2(32'hbb139e82),
	.w3(32'hba875cde),
	.w4(32'h3bef4d98),
	.w5(32'h38d01810),
	.w6(32'hbb4c2d7a),
	.w7(32'hba441a97),
	.w8(32'hba155435),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b325cbd),
	.w1(32'hbba71a87),
	.w2(32'hb8c4b413),
	.w3(32'hbba878b8),
	.w4(32'hbaeca300),
	.w5(32'h39b5759d),
	.w6(32'h3b995ce1),
	.w7(32'h3c0ce6a2),
	.w8(32'hbbfc4ed1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02eac6),
	.w1(32'hbab7aad3),
	.w2(32'h395a4854),
	.w3(32'hba2e417b),
	.w4(32'hbbf6f241),
	.w5(32'hbca4c589),
	.w6(32'h3b2918a3),
	.w7(32'hbb532652),
	.w8(32'hbb8d4613),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b80d5b),
	.w1(32'hbc07d2c9),
	.w2(32'hbb857c03),
	.w3(32'hbb092e64),
	.w4(32'hba3b4751),
	.w5(32'hbb354536),
	.w6(32'h3ba20968),
	.w7(32'h3bb0a622),
	.w8(32'hba7a15e5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5a4f),
	.w1(32'hbb14023c),
	.w2(32'hbb200714),
	.w3(32'h3b186684),
	.w4(32'h3bd03eca),
	.w5(32'h3bece9dc),
	.w6(32'hbb80d7ad),
	.w7(32'hbb0d5e2b),
	.w8(32'hbb00e430),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d220e),
	.w1(32'h39d5ce68),
	.w2(32'hba749937),
	.w3(32'h3c023f03),
	.w4(32'hbc436abc),
	.w5(32'hbb90ea52),
	.w6(32'hb8d04855),
	.w7(32'hbb54682c),
	.w8(32'h3a2dfd5d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc1d62),
	.w1(32'hbc04173e),
	.w2(32'h3a804c55),
	.w3(32'hb9f270f4),
	.w4(32'hbb0796f5),
	.w5(32'hbb24e43a),
	.w6(32'hbb931465),
	.w7(32'h3af15a92),
	.w8(32'h3a8d1fec),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70e6ed),
	.w1(32'h3d41688f),
	.w2(32'hbb96ba70),
	.w3(32'hbb8e1867),
	.w4(32'hbbffd55a),
	.w5(32'h3b955abb),
	.w6(32'hbaa8d99b),
	.w7(32'hbbcb4b62),
	.w8(32'hbb71469e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23faa6),
	.w1(32'h3b432c03),
	.w2(32'hbb0f3778),
	.w3(32'hbba688ed),
	.w4(32'h3947060a),
	.w5(32'hbad9b2c0),
	.w6(32'hb999c677),
	.w7(32'hbbad1526),
	.w8(32'h3cb433ba),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e7d94),
	.w1(32'hbb021a31),
	.w2(32'hbb4c70ab),
	.w3(32'hbb98f504),
	.w4(32'hb65787a2),
	.w5(32'hbc32709b),
	.w6(32'hbabed9d1),
	.w7(32'h3c09f91d),
	.w8(32'h392fe73b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72e8b),
	.w1(32'h3a903127),
	.w2(32'hba862789),
	.w3(32'hbc8caffe),
	.w4(32'hbb937979),
	.w5(32'hbb4d4c51),
	.w6(32'h3bd16e4e),
	.w7(32'hbb98e500),
	.w8(32'hbbd95689),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47308b),
	.w1(32'hbb613fd1),
	.w2(32'hbb0181d5),
	.w3(32'hbb7c7f3b),
	.w4(32'hba366063),
	.w5(32'h3aa52e47),
	.w6(32'h3ac4883b),
	.w7(32'hba7ac8ff),
	.w8(32'h3b9edece),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b3465),
	.w1(32'h392abbde),
	.w2(32'hbb1c7b6a),
	.w3(32'hb8905171),
	.w4(32'hbae16a5c),
	.w5(32'h38939799),
	.w6(32'h3bfc7d5f),
	.w7(32'hbbe67cd5),
	.w8(32'hbb88c234),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d3c7b),
	.w1(32'h3b797d5d),
	.w2(32'h3bd3caf3),
	.w3(32'hbb8530d8),
	.w4(32'hba7d708c),
	.w5(32'hbb9e1e1d),
	.w6(32'hbb4012e2),
	.w7(32'h3cb1b9cc),
	.w8(32'hbb9fab91),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941f4a),
	.w1(32'hb9a7012a),
	.w2(32'h39a33369),
	.w3(32'hbc16b549),
	.w4(32'hbbbf56e9),
	.w5(32'hbb809a80),
	.w6(32'hbbb30799),
	.w7(32'h3a8ddf1d),
	.w8(32'h3ac5bacc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb3786),
	.w1(32'h3b8bc00f),
	.w2(32'h3d139e33),
	.w3(32'hb6e9e32b),
	.w4(32'h3b95b616),
	.w5(32'hbbd98846),
	.w6(32'h3a20976f),
	.w7(32'hba3c739c),
	.w8(32'hba99f159),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2f274),
	.w1(32'hb9a3e1c0),
	.w2(32'hbb8cec7e),
	.w3(32'hbb1f7ccc),
	.w4(32'h3c226a5c),
	.w5(32'h3b1eb45c),
	.w6(32'h3be363e8),
	.w7(32'hbba1670e),
	.w8(32'h3c470d0f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64b2941),
	.w1(32'hbc75918f),
	.w2(32'h3ba202b2),
	.w3(32'hbb84ca4f),
	.w4(32'h3a1c377c),
	.w5(32'h3b6bd91c),
	.w6(32'hbb05161a),
	.w7(32'hbbbf54e5),
	.w8(32'hba2b73b2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59b97a),
	.w1(32'h3a9cded6),
	.w2(32'hbadc9cff),
	.w3(32'hbbfce922),
	.w4(32'hbad142ac),
	.w5(32'h3a691f5e),
	.w6(32'h3bea8f0f),
	.w7(32'h3bde8c7c),
	.w8(32'h3c8b6b05),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43ef3d),
	.w1(32'hbba61de4),
	.w2(32'hbb82d325),
	.w3(32'h3af1a85b),
	.w4(32'h3a04a4b9),
	.w5(32'h3ac35f59),
	.w6(32'hbaad78ef),
	.w7(32'h3af24182),
	.w8(32'hbb87f025),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4394d5),
	.w1(32'h3b7ab65d),
	.w2(32'hbb9f0ec3),
	.w3(32'h3b09dc37),
	.w4(32'hbbbea1f4),
	.w5(32'h3c765c20),
	.w6(32'hbb449c79),
	.w7(32'hba1b06e7),
	.w8(32'hbb3cb694),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f613b),
	.w1(32'hba698efe),
	.w2(32'h39b5648e),
	.w3(32'h3af0dac7),
	.w4(32'h3b3f93fd),
	.w5(32'h3a74fa01),
	.w6(32'h3bbccd20),
	.w7(32'h3a7c8d64),
	.w8(32'hbac1ec4d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e1471),
	.w1(32'hbaa22282),
	.w2(32'h3a661971),
	.w3(32'hb9bd6e5a),
	.w4(32'hb94e02e8),
	.w5(32'hbaf45ad1),
	.w6(32'hbbfff61f),
	.w7(32'hb7bd4cc1),
	.w8(32'hb8a441d8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ba728),
	.w1(32'hbca9e58f),
	.w2(32'hbb95c665),
	.w3(32'h3a740326),
	.w4(32'h3a00ba7c),
	.w5(32'h3b833f11),
	.w6(32'hbc716593),
	.w7(32'hbac95768),
	.w8(32'h3c10a83a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a665048),
	.w1(32'hbb954acc),
	.w2(32'hbb09b7fd),
	.w3(32'h390d16f6),
	.w4(32'h3b42de52),
	.w5(32'hbb39e0bd),
	.w6(32'hba4ce70d),
	.w7(32'h3ab203ea),
	.w8(32'hbbdc346e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce894c),
	.w1(32'h3b54bf9e),
	.w2(32'hbadb7c1c),
	.w3(32'hba3c536a),
	.w4(32'hbbeac3de),
	.w5(32'hbc474054),
	.w6(32'h3bb6e04b),
	.w7(32'h3b8c1506),
	.w8(32'hb9a88c80),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32b517),
	.w1(32'hbafbbc17),
	.w2(32'hbbb70dce),
	.w3(32'h3a4c0668),
	.w4(32'hbb6240f6),
	.w5(32'hbbcfbfbe),
	.w6(32'hbbbda4d3),
	.w7(32'h39a37518),
	.w8(32'h39a05455),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256bfc),
	.w1(32'h3c12e1bc),
	.w2(32'h3b407353),
	.w3(32'hbb98ece5),
	.w4(32'hbaf8c6ad),
	.w5(32'hbb83550a),
	.w6(32'h3afb1663),
	.w7(32'hbba098ea),
	.w8(32'hbb9edf43),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b596),
	.w1(32'hbac1ad6b),
	.w2(32'hbb80e80a),
	.w3(32'hbc7d147b),
	.w4(32'hbafda62d),
	.w5(32'hba3d6477),
	.w6(32'h3a025eb1),
	.w7(32'hbb4f01ae),
	.w8(32'h3b0e3c5b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule