module layer_10_featuremap_208(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38481a9d),
	.w1(32'hbade737a),
	.w2(32'hbb3098d1),
	.w3(32'hb9137382),
	.w4(32'h38f2499c),
	.w5(32'hbae2c10d),
	.w6(32'hbb4ddee1),
	.w7(32'hba8f9e72),
	.w8(32'hba2c8ab2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf66d58),
	.w1(32'hbae8f8ea),
	.w2(32'hbb064387),
	.w3(32'hbafe97bd),
	.w4(32'hbac7e8b6),
	.w5(32'hbaf713db),
	.w6(32'hbaea77c6),
	.w7(32'hbaded5db),
	.w8(32'hbae52f51),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae87f90),
	.w1(32'hba562b33),
	.w2(32'hba6c2739),
	.w3(32'hbafbc290),
	.w4(32'hbaaa2dfe),
	.w5(32'hbaea166b),
	.w6(32'hba94a07b),
	.w7(32'hba9a4862),
	.w8(32'hba826e91),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e5719),
	.w1(32'hb9e342fe),
	.w2(32'hb9b7a368),
	.w3(32'hbacaf45f),
	.w4(32'hba86df2e),
	.w5(32'hba430c0a),
	.w6(32'hba1e5f2d),
	.w7(32'hba1bb67e),
	.w8(32'hb9867357),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eca5fb),
	.w1(32'h39ce912b),
	.w2(32'hb96b386f),
	.w3(32'hba8b0df7),
	.w4(32'h3a492024),
	.w5(32'h390db3b0),
	.w6(32'h3a54af0e),
	.w7(32'hba2f3f64),
	.w8(32'h3a740421),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa724b3),
	.w1(32'hb9f1f2b7),
	.w2(32'hb8dc8b67),
	.w3(32'h39a76fcf),
	.w4(32'hba040ad2),
	.w5(32'hb9ad3b4c),
	.w6(32'hba537c08),
	.w7(32'hba4f9e98),
	.w8(32'hba4ff28e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba103704),
	.w1(32'hbaefaf77),
	.w2(32'hbadffbf5),
	.w3(32'hba7ce706),
	.w4(32'hbab9b339),
	.w5(32'hbae1f9d2),
	.w6(32'hbac731bf),
	.w7(32'hbaec3d08),
	.w8(32'hbac5b450),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb924d),
	.w1(32'h391791a0),
	.w2(32'h39740375),
	.w3(32'hbace2ae8),
	.w4(32'h37ad414b),
	.w5(32'h39a186b7),
	.w6(32'hb8ef243d),
	.w7(32'hb894c9a3),
	.w8(32'h39842990),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397fe64d),
	.w1(32'hb97095bb),
	.w2(32'h38b47062),
	.w3(32'h391b801b),
	.w4(32'hba45f4f8),
	.w5(32'hba116308),
	.w6(32'hb9edb786),
	.w7(32'hb9de7665),
	.w8(32'hb9c57203),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0331e),
	.w1(32'hba5dd3cf),
	.w2(32'hba6e3425),
	.w3(32'hb9fae901),
	.w4(32'hba739223),
	.w5(32'hba8b527e),
	.w6(32'hba7ad742),
	.w7(32'hba88d288),
	.w8(32'hba6971e2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d35c0),
	.w1(32'h3a249f79),
	.w2(32'h3ae674b0),
	.w3(32'hba930f1f),
	.w4(32'hba85e9ec),
	.w5(32'hba4b0b01),
	.w6(32'hba6c856e),
	.w7(32'hba67c9d8),
	.w8(32'hb9129338),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0279c9),
	.w1(32'hb8ee5e92),
	.w2(32'h39a91aa4),
	.w3(32'hb8e91dc1),
	.w4(32'h3945d529),
	.w5(32'h39c4e7ed),
	.w6(32'h3adb95b9),
	.w7(32'h3b1e144f),
	.w8(32'h3ad49a5c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9850d51),
	.w1(32'h38b54cba),
	.w2(32'h39cd3c3a),
	.w3(32'hb985fd9d),
	.w4(32'hb94ae97b),
	.w5(32'h390156c6),
	.w6(32'h391f09f2),
	.w7(32'h392cafee),
	.w8(32'h394847a3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0580f),
	.w1(32'h3a8acc12),
	.w2(32'h3a810303),
	.w3(32'hb86c495c),
	.w4(32'h3a412364),
	.w5(32'h3a616716),
	.w6(32'h39d0b602),
	.w7(32'h3a33b9a7),
	.w8(32'h3acabe3f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4ce41),
	.w1(32'h39eaf936),
	.w2(32'h38e4f234),
	.w3(32'h3a86c652),
	.w4(32'h3af2f8c7),
	.w5(32'h3ad72d62),
	.w6(32'h3aca2433),
	.w7(32'h3b2f1134),
	.w8(32'h3b2195b7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80025ef),
	.w1(32'hb9ca4217),
	.w2(32'hb918aa5a),
	.w3(32'h384c13d8),
	.w4(32'hba1ac077),
	.w5(32'hba2bd599),
	.w6(32'hba39fb21),
	.w7(32'hba10dc0d),
	.w8(32'hba140b78),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f47d2),
	.w1(32'h3a02b3f2),
	.w2(32'hb9ccb200),
	.w3(32'hba3093eb),
	.w4(32'h39f1d400),
	.w5(32'hba6223ee),
	.w6(32'h3a006b58),
	.w7(32'hb8ac2be1),
	.w8(32'h38a9ed62),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5d60a),
	.w1(32'hba8f34c4),
	.w2(32'hba77b44b),
	.w3(32'hba25253b),
	.w4(32'hba8cb724),
	.w5(32'hbac78a1c),
	.w6(32'hba89edee),
	.w7(32'hba870897),
	.w8(32'hba83f635),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f21d8),
	.w1(32'hba65587a),
	.w2(32'hba7636c2),
	.w3(32'hbab5485e),
	.w4(32'hba319c24),
	.w5(32'hba888a72),
	.w6(32'hba550ba0),
	.w7(32'hba700e2a),
	.w8(32'hba558020),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855712),
	.w1(32'hb8faf441),
	.w2(32'h397297c2),
	.w3(32'hba782605),
	.w4(32'hb969dea1),
	.w5(32'hb9017069),
	.w6(32'hb98a6ea6),
	.w7(32'h37d35785),
	.w8(32'h38897985),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b99e16),
	.w1(32'hb93595d0),
	.w2(32'hb9089179),
	.w3(32'hb8f8ab1f),
	.w4(32'hb98ea35b),
	.w5(32'hb9bc5276),
	.w6(32'h38f50458),
	.w7(32'hb844bbfe),
	.w8(32'h371d006e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e8d11),
	.w1(32'hbb205890),
	.w2(32'hba2ad562),
	.w3(32'hb9a23061),
	.w4(32'hbac2d114),
	.w5(32'hba23ad26),
	.w6(32'hbaef2406),
	.w7(32'hb9d6c9a1),
	.w8(32'hba321358),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9806789),
	.w1(32'h39de6d78),
	.w2(32'h39b37feb),
	.w3(32'hbab96718),
	.w4(32'hb99bdc57),
	.w5(32'hba815e7e),
	.w6(32'h39ac792f),
	.w7(32'h388e43f9),
	.w8(32'hb93eb315),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb809902e),
	.w1(32'hb99ddb33),
	.w2(32'hb89a87e5),
	.w3(32'hba67056f),
	.w4(32'hb96f4d78),
	.w5(32'hb8d8254c),
	.w6(32'hb9efa673),
	.w7(32'hb961dea8),
	.w8(32'h375a985c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9bbaa),
	.w1(32'hba92ddeb),
	.w2(32'hbab3107b),
	.w3(32'hb9da5021),
	.w4(32'hb9832c87),
	.w5(32'hba5ca6e4),
	.w6(32'hbaadcf35),
	.w7(32'hbab052ec),
	.w8(32'hbaa94270),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cad99),
	.w1(32'h3a88c734),
	.w2(32'h3a2deb2c),
	.w3(32'hba0bc2c7),
	.w4(32'hba44ba81),
	.w5(32'hb9ee5052),
	.w6(32'h3a3fd49a),
	.w7(32'h3a73f9e5),
	.w8(32'h3a99f6cb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39add0c6),
	.w1(32'h382b0349),
	.w2(32'h39e98a21),
	.w3(32'hb98495b3),
	.w4(32'hb9115bfb),
	.w5(32'h39a16186),
	.w6(32'hb7c10970),
	.w7(32'h39a87d6e),
	.w8(32'h39b1cf6e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39956d69),
	.w1(32'hba6a1629),
	.w2(32'hba2a425d),
	.w3(32'h394dc580),
	.w4(32'hb9e5d9c5),
	.w5(32'hb9df5ffc),
	.w6(32'hba803309),
	.w7(32'hb9bf352e),
	.w8(32'hba56b083),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8775c7),
	.w1(32'hb9f28936),
	.w2(32'h39d509b3),
	.w3(32'hb9e1f85c),
	.w4(32'hba0c50a6),
	.w5(32'h3963d42c),
	.w6(32'hba9dfef4),
	.w7(32'hb9b4afcc),
	.w8(32'h39d7e107),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89a34b),
	.w1(32'h3a64fd53),
	.w2(32'hb97848d1),
	.w3(32'h3a14b79b),
	.w4(32'h3a882074),
	.w5(32'h38065327),
	.w6(32'h3a71f3cc),
	.w7(32'hb9088041),
	.w8(32'h3805e33b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f8af85),
	.w1(32'hb8b26d03),
	.w2(32'hb603240f),
	.w3(32'h39910881),
	.w4(32'hb8ceba42),
	.w5(32'hb9035f75),
	.w6(32'h37ff9ad4),
	.w7(32'hb78beb5f),
	.w8(32'h3706659d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3805f0e2),
	.w1(32'hb907fa12),
	.w2(32'h375d1f0f),
	.w3(32'hb77e8c6f),
	.w4(32'hb9a346f2),
	.w5(32'hb997be9a),
	.w6(32'hb904900e),
	.w7(32'hb94b7032),
	.w8(32'hb8714399),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97aaa2a),
	.w1(32'hb9ef7731),
	.w2(32'hba62054b),
	.w3(32'hba0e9e46),
	.w4(32'hba1f8a5b),
	.w5(32'hb9ed89b6),
	.w6(32'hb915a4ae),
	.w7(32'hba4e314b),
	.w8(32'hba853a66),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c887b),
	.w1(32'hbaa628c4),
	.w2(32'h39158adb),
	.w3(32'hba034707),
	.w4(32'hbab4d47c),
	.w5(32'h3a6f0257),
	.w6(32'hbb07df20),
	.w7(32'hb9513662),
	.w8(32'h3832ba7a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e29e8f),
	.w1(32'hbafba21e),
	.w2(32'hbaebe98f),
	.w3(32'hb9a269f8),
	.w4(32'hbb0389a8),
	.w5(32'hbb065eae),
	.w6(32'hbafc4b67),
	.w7(32'hbb0da11d),
	.w8(32'hbad2d3aa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6b16f),
	.w1(32'hb88cd822),
	.w2(32'h39994a7c),
	.w3(32'hbae7f4f5),
	.w4(32'hb86009ea),
	.w5(32'hb96dd9a4),
	.w6(32'h3907fc3e),
	.w7(32'h39c3a53a),
	.w8(32'h39f65008),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39228958),
	.w1(32'hbab18055),
	.w2(32'hbabe6dc0),
	.w3(32'hb916ee15),
	.w4(32'hba7b15ec),
	.w5(32'hbab79238),
	.w6(32'hba8c56ce),
	.w7(32'hbaa7de55),
	.w8(32'hba95d2ed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8169e),
	.w1(32'hbab516d6),
	.w2(32'hbabf8ba9),
	.w3(32'hbaba05c1),
	.w4(32'hba82e2f8),
	.w5(32'hbabd05a8),
	.w6(32'hbaa881d6),
	.w7(32'hba8be608),
	.w8(32'hba7a0dda),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbecee),
	.w1(32'hba0ead5d),
	.w2(32'hba0bc371),
	.w3(32'hbab99f0e),
	.w4(32'hb98108b5),
	.w5(32'hb9e9dd13),
	.w6(32'hba274192),
	.w7(32'hb9a8558f),
	.w8(32'hb9566ad8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8faa612),
	.w1(32'hba9bd407),
	.w2(32'hbab6f88d),
	.w3(32'hb9af728c),
	.w4(32'hba7ee4b4),
	.w5(32'hba9580ad),
	.w6(32'hbaa4983a),
	.w7(32'hbaa91116),
	.w8(32'hba8a55d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fae8a),
	.w1(32'h39e023ca),
	.w2(32'hb8dad5a5),
	.w3(32'hbaaea220),
	.w4(32'h3a5987e6),
	.w5(32'h39c4b83e),
	.w6(32'h39fe41f4),
	.w7(32'h38149436),
	.w8(32'h395d81be),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c33ed2),
	.w1(32'hba88276a),
	.w2(32'hbaa35658),
	.w3(32'h3a3cbbf9),
	.w4(32'hba9d1257),
	.w5(32'hbaad6dd7),
	.w6(32'hba701996),
	.w7(32'hba693744),
	.w8(32'hba6d203a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafe7e5),
	.w1(32'hb9905f6a),
	.w2(32'hb95050ff),
	.w3(32'hbad6678e),
	.w4(32'hba0f8d9b),
	.w5(32'hba0cb928),
	.w6(32'hb9c73e87),
	.w7(32'hb9c826f9),
	.w8(32'hb901b5b3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8661c12),
	.w1(32'hb9ddaa33),
	.w2(32'hb9fd0695),
	.w3(32'hba0ffc49),
	.w4(32'hb97fe265),
	.w5(32'hb9c26cea),
	.w6(32'hb9d9a84d),
	.w7(32'hb95bc7c5),
	.w8(32'hb94050d1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9d5d1),
	.w1(32'h396a7e0b),
	.w2(32'h38ba5800),
	.w3(32'hb9915ce0),
	.w4(32'h39c700e8),
	.w5(32'hb9bbca9e),
	.w6(32'h399e55fb),
	.w7(32'h3a2044a6),
	.w8(32'h3a67784a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a36192),
	.w1(32'hba61819e),
	.w2(32'hb8c2874a),
	.w3(32'hba2a3fac),
	.w4(32'hba71661f),
	.w5(32'hb9b5870e),
	.w6(32'hba067f48),
	.w7(32'hb9aacb32),
	.w8(32'hb983d01a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5d87d),
	.w1(32'hba6a17b9),
	.w2(32'hb92ccf89),
	.w3(32'hb9941bff),
	.w4(32'h3a3b08f5),
	.w5(32'h3a852b76),
	.w6(32'h3ae8ee59),
	.w7(32'h3ae5479a),
	.w8(32'h3a578b96),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eb194),
	.w1(32'h386d9ae4),
	.w2(32'h3959050f),
	.w3(32'hba04373f),
	.w4(32'hba6beb12),
	.w5(32'hba5ae11e),
	.w6(32'hba2e699a),
	.w7(32'hb9d347d0),
	.w8(32'h3a6095c5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7e46a),
	.w1(32'hb79506f9),
	.w2(32'h38b5c19f),
	.w3(32'h398180bc),
	.w4(32'hb93cdf2f),
	.w5(32'hb8e47b65),
	.w6(32'hb98a8591),
	.w7(32'hb8149020),
	.w8(32'h39836086),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b87d5),
	.w1(32'h393763da),
	.w2(32'h38c3e411),
	.w3(32'hb982167f),
	.w4(32'h388a909d),
	.w5(32'h38efa21d),
	.w6(32'hb92527f2),
	.w7(32'hb7a53669),
	.w8(32'h396a6b28),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1d09e),
	.w1(32'h390e9fbb),
	.w2(32'h39cb1215),
	.w3(32'h39b558e9),
	.w4(32'hb8ba1543),
	.w5(32'h37d79e22),
	.w6(32'h392a12c7),
	.w7(32'h3a07a9f2),
	.w8(32'h39cbfa09),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e43ff5),
	.w1(32'hb9d924b2),
	.w2(32'h37cf606f),
	.w3(32'h3a38c434),
	.w4(32'hbad01f12),
	.w5(32'hbaf63606),
	.w6(32'hba627b5d),
	.w7(32'hba46690c),
	.w8(32'hbaad8304),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bc562),
	.w1(32'hba0fe49b),
	.w2(32'hb9eb8c16),
	.w3(32'hba52869f),
	.w4(32'hb9073ee4),
	.w5(32'hba229698),
	.w6(32'hba493f57),
	.w7(32'hba557c63),
	.w8(32'hbaa935c9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80055d),
	.w1(32'h39d8c391),
	.w2(32'h36e87638),
	.w3(32'hba7c78dc),
	.w4(32'h3a6b2de7),
	.w5(32'h3955a179),
	.w6(32'h3a93bd58),
	.w7(32'hba8180e5),
	.w8(32'hb9b53fea),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f87f17),
	.w1(32'h37b416dd),
	.w2(32'hba351ae7),
	.w3(32'h388c3f71),
	.w4(32'h39ce5301),
	.w5(32'hb9c1df99),
	.w6(32'hb99a1ae5),
	.w7(32'hba0e83f3),
	.w8(32'hb935fc37),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98986ea),
	.w1(32'hb9c7d42e),
	.w2(32'hba1781e8),
	.w3(32'hba183437),
	.w4(32'h39d03dc1),
	.w5(32'h39f8068b),
	.w6(32'hb7bbb1c0),
	.w7(32'hba24c48b),
	.w8(32'hba0015a3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3774af0e),
	.w1(32'h3a141e2f),
	.w2(32'h3a643b04),
	.w3(32'h3a9dd217),
	.w4(32'h39db592f),
	.w5(32'h3a29e60e),
	.w6(32'h39f9380b),
	.w7(32'h3a643a8c),
	.w8(32'h3a79b0c1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4409),
	.w1(32'h39655c56),
	.w2(32'hbabdfb14),
	.w3(32'h3a1ffa25),
	.w4(32'h3855d9ad),
	.w5(32'hb95ada30),
	.w6(32'h3a96c406),
	.w7(32'hbaa3319f),
	.w8(32'h3ab7e278),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa12f8e),
	.w1(32'hbada3c87),
	.w2(32'hbb0280f2),
	.w3(32'h3aac476d),
	.w4(32'hba9d8393),
	.w5(32'hbae89d13),
	.w6(32'hbafa46c1),
	.w7(32'hbaf05074),
	.w8(32'hbad7cdf5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec9e4f),
	.w1(32'hb9dcf1d8),
	.w2(32'hb907e509),
	.w3(32'hbb043410),
	.w4(32'hb9dfe0ee),
	.w5(32'hb996d97c),
	.w6(32'hba3fca0f),
	.w7(32'hb9e3dc17),
	.w8(32'hb90cf41c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909365f),
	.w1(32'hbae93aee),
	.w2(32'hbaef6833),
	.w3(32'hb9a36d90),
	.w4(32'hbacd8d7a),
	.w5(32'hbaf24417),
	.w6(32'hbab57c85),
	.w7(32'hbab84a49),
	.w8(32'hbaac1fb8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3f723),
	.w1(32'hb9216a21),
	.w2(32'h38a48558),
	.w3(32'hbad7a7ee),
	.w4(32'hb974ed70),
	.w5(32'hb61814f9),
	.w6(32'hb9908c92),
	.w7(32'h390bc348),
	.w8(32'hb855178b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9278cd2),
	.w1(32'h389aedd6),
	.w2(32'hbae600ee),
	.w3(32'h378b238f),
	.w4(32'hbac919af),
	.w5(32'hbabbcd9c),
	.w6(32'hb9f90b81),
	.w7(32'hbaf25dc4),
	.w8(32'hba71c2d6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf81d18),
	.w1(32'hba1f4f26),
	.w2(32'hba1f7228),
	.w3(32'hbb1a955d),
	.w4(32'hb9ed58d1),
	.w5(32'hba1791d5),
	.w6(32'hb9b83bde),
	.w7(32'hb9b99f85),
	.w8(32'hb9b2b3a8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdd0de),
	.w1(32'hba805d8f),
	.w2(32'hba8f1743),
	.w3(32'hb9c3e61b),
	.w4(32'hba4acb7f),
	.w5(32'hba4f98e5),
	.w6(32'hba97aace),
	.w7(32'hba48b796),
	.w8(32'hba6709ed),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d91c),
	.w1(32'hb7d0cf17),
	.w2(32'hb9d7eb8a),
	.w3(32'hba9ad98b),
	.w4(32'hba4c76b7),
	.w5(32'hb93602b7),
	.w6(32'hb8aace1a),
	.w7(32'hba4dbd18),
	.w8(32'h393f57f5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeffa33),
	.w1(32'hb874e066),
	.w2(32'hba5bfd9d),
	.w3(32'h3a7312fb),
	.w4(32'h39d588c8),
	.w5(32'hb8df8131),
	.w6(32'h3a208371),
	.w7(32'hb871733b),
	.w8(32'hb9209a49),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65e81b),
	.w1(32'h3966ba72),
	.w2(32'h3a19da3d),
	.w3(32'hb885f836),
	.w4(32'hb9ce978f),
	.w5(32'hb9644746),
	.w6(32'h3a3c3783),
	.w7(32'h3a59b4c4),
	.w8(32'h3a8b12cb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a786374),
	.w1(32'hba0d504d),
	.w2(32'hb9900050),
	.w3(32'h38820350),
	.w4(32'hb99813ec),
	.w5(32'hb9ed11d1),
	.w6(32'hba023144),
	.w7(32'hb9bdbc07),
	.w8(32'hba0f1ca6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a684e),
	.w1(32'h3a2ee9e3),
	.w2(32'h39ae31b9),
	.w3(32'hba2ba35a),
	.w4(32'h3901def5),
	.w5(32'h39ffdc8a),
	.w6(32'h3a1e7ba6),
	.w7(32'h3a049b46),
	.w8(32'h3a8ce1ff),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4bd3),
	.w1(32'hbaa91509),
	.w2(32'hbabd4228),
	.w3(32'h3ae11cff),
	.w4(32'hbaa4a4dd),
	.w5(32'hbaddceba),
	.w6(32'hbaa640fe),
	.w7(32'hba99b925),
	.w8(32'hba8acbc4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9581ce),
	.w1(32'hb8c4cb83),
	.w2(32'h38e90fb2),
	.w3(32'hbac90a4c),
	.w4(32'hb732d1ea),
	.w5(32'h39306963),
	.w6(32'h3856eb72),
	.w7(32'h379eac90),
	.w8(32'h3951ffc1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b7a4e),
	.w1(32'hb9b2d481),
	.w2(32'hb8f9f763),
	.w3(32'h38f16b37),
	.w4(32'hb9a592ce),
	.w5(32'hb9936ee6),
	.w6(32'hba120897),
	.w7(32'hb9beac93),
	.w8(32'hb8f46974),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a51871),
	.w1(32'h36644cea),
	.w2(32'h3925a03f),
	.w3(32'hb97d2375),
	.w4(32'hb8e7b93a),
	.w5(32'hb9c8b152),
	.w6(32'hb8e4e012),
	.w7(32'hb8bdcdf1),
	.w8(32'hb7fec06e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398291c0),
	.w1(32'hbada6a5b),
	.w2(32'hbae06ed8),
	.w3(32'hb9b29d1a),
	.w4(32'hbab5a8ae),
	.w5(32'hbaed6c02),
	.w6(32'hbafab15d),
	.w7(32'hbaea4ab8),
	.w8(32'hbada7c84),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfbab9),
	.w1(32'hbac06ae9),
	.w2(32'hbabf3a22),
	.w3(32'hbad998e1),
	.w4(32'hbad1bce0),
	.w5(32'hbaae2d37),
	.w6(32'h3ab89f1b),
	.w7(32'h3ade2d81),
	.w8(32'h3910498c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbcf1a),
	.w1(32'h3a09a79c),
	.w2(32'h3a553d0e),
	.w3(32'hb9b45d91),
	.w4(32'h399c2c32),
	.w5(32'h3a3c5d83),
	.w6(32'h389e4267),
	.w7(32'h397b1887),
	.w8(32'h3a1aeecd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84a176),
	.w1(32'hba7b742a),
	.w2(32'hbab56f7d),
	.w3(32'h3a7e8f63),
	.w4(32'hbaa94f2f),
	.w5(32'hbabd11fa),
	.w6(32'hba680be2),
	.w7(32'hbac04302),
	.w8(32'hbaa79067),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5fb94),
	.w1(32'h3a8f48e3),
	.w2(32'h3901ffaa),
	.w3(32'hbac223aa),
	.w4(32'h39cdfba8),
	.w5(32'hba2b7218),
	.w6(32'h39d5813d),
	.w7(32'h37cadc0f),
	.w8(32'hb968697b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fe3b6),
	.w1(32'hb9ca038c),
	.w2(32'hb99149fd),
	.w3(32'hb88a24f0),
	.w4(32'hba0bd1a0),
	.w5(32'hb9f3566c),
	.w6(32'hb91555e9),
	.w7(32'hb9acf61a),
	.w8(32'hb8c8a5b2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb96c1),
	.w1(32'h38f101b4),
	.w2(32'h3a43b959),
	.w3(32'hb98f1a71),
	.w4(32'h38e55ed8),
	.w5(32'h39d9f602),
	.w6(32'h39d14660),
	.w7(32'h3a446b02),
	.w8(32'h3a5f1e8c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33c0bb),
	.w1(32'hba223e54),
	.w2(32'hba5e3722),
	.w3(32'h3a07c54c),
	.w4(32'hb9e71334),
	.w5(32'hba4cbb7c),
	.w6(32'hba38afcf),
	.w7(32'hba57cb2f),
	.w8(32'hba8545a4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75b6ed),
	.w1(32'h39b537cc),
	.w2(32'h39340ace),
	.w3(32'hba871a0c),
	.w4(32'h39f61b9d),
	.w5(32'h392fd001),
	.w6(32'h3816ad94),
	.w7(32'h391009d2),
	.w8(32'hb6c9e1c3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8def606),
	.w1(32'hbaf0ca2c),
	.w2(32'hbb06c535),
	.w3(32'hb8fcc22f),
	.w4(32'hba94f14a),
	.w5(32'hbacf780b),
	.w6(32'hbae3471d),
	.w7(32'hbae4bf56),
	.w8(32'hbacde56d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5cc22),
	.w1(32'hb73a0944),
	.w2(32'h3a983145),
	.w3(32'hbaf255c8),
	.w4(32'hbabd94b2),
	.w5(32'hba9096f9),
	.w6(32'hba68d2ab),
	.w7(32'hb998a297),
	.w8(32'h3a882c66),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8a92e),
	.w1(32'h39b070a9),
	.w2(32'hb8f282b6),
	.w3(32'h38e5cbc2),
	.w4(32'h39e16829),
	.w5(32'h3946213b),
	.w6(32'h3a1ae8c1),
	.w7(32'h39dc826a),
	.w8(32'h39f4f145),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f58388),
	.w1(32'hb987388f),
	.w2(32'h399c299a),
	.w3(32'h39e4ceec),
	.w4(32'hba6634f7),
	.w5(32'hb839f315),
	.w6(32'hb9c8396a),
	.w7(32'hb7df3ace),
	.w8(32'h39f34e12),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f837e3),
	.w1(32'hb9297072),
	.w2(32'hb8e53d90),
	.w3(32'h39c19024),
	.w4(32'hb981054c),
	.w5(32'hb98ae438),
	.w6(32'hb8bb9763),
	.w7(32'hb9421d94),
	.w8(32'hb9264bcb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9234dc3),
	.w1(32'hb9e42f97),
	.w2(32'hbaa413bd),
	.w3(32'hb9860b93),
	.w4(32'h390656c6),
	.w5(32'hba5195d0),
	.w6(32'hba0ec3fb),
	.w7(32'hba6d8b2a),
	.w8(32'hba18f686),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a6b69),
	.w1(32'hb8af6dcb),
	.w2(32'hb9b561fa),
	.w3(32'hba7696d7),
	.w4(32'hb987d7cd),
	.w5(32'hba189691),
	.w6(32'h38709207),
	.w7(32'hb99633b1),
	.w8(32'hb970c49d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca3425),
	.w1(32'hb8a10a8e),
	.w2(32'h38633423),
	.w3(32'hba09a31a),
	.w4(32'hb9395651),
	.w5(32'hb9a49985),
	.w6(32'hb89bb144),
	.w7(32'hb8c070f2),
	.w8(32'hb8b1e9c0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7080a),
	.w1(32'hba6374ea),
	.w2(32'hba5b16f7),
	.w3(32'hb9a6a89b),
	.w4(32'hba65ef46),
	.w5(32'hba73c29f),
	.w6(32'hb99df59b),
	.w7(32'hb9a7ddaa),
	.w8(32'hb9db1b2f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba257d4e),
	.w1(32'hbac89d5c),
	.w2(32'hbaed0252),
	.w3(32'hba51973f),
	.w4(32'hbaa268ef),
	.w5(32'hbae4c5a9),
	.w6(32'hbac3991c),
	.w7(32'hbabeff24),
	.w8(32'hbab4e179),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc9051),
	.w1(32'h39709682),
	.w2(32'h39d75cdc),
	.w3(32'hbaea9c3f),
	.w4(32'h3994fc94),
	.w5(32'h399fb9df),
	.w6(32'h3996f6ab),
	.w7(32'h39b31aaa),
	.w8(32'h39de9c52),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08559b),
	.w1(32'hba8aedbe),
	.w2(32'hba9ca192),
	.w3(32'h3a142622),
	.w4(32'hbac79a8d),
	.w5(32'hbacbf680),
	.w6(32'hbaac0900),
	.w7(32'hbacd2e0c),
	.w8(32'hba7ad12a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f80aa),
	.w1(32'hba6eb71a),
	.w2(32'hb9d57b00),
	.w3(32'hbac36304),
	.w4(32'hba29d3a8),
	.w5(32'h38327850),
	.w6(32'hb9fe0811),
	.w7(32'hba67baaf),
	.w8(32'hba96958a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d7fee),
	.w1(32'hba3262d7),
	.w2(32'hb97d79a6),
	.w3(32'hba066bea),
	.w4(32'hba8f0471),
	.w5(32'hbaa0e02a),
	.w6(32'hba067f1d),
	.w7(32'hb9e876c6),
	.w8(32'hb9fcf037),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13e842),
	.w1(32'hb9a1ec0d),
	.w2(32'hb99ead7f),
	.w3(32'hba786268),
	.w4(32'hba3e4f14),
	.w5(32'h37009a50),
	.w6(32'hba446212),
	.w7(32'hb820fe2e),
	.w8(32'hba051cad),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5dec),
	.w1(32'hbaa1c895),
	.w2(32'hbac16723),
	.w3(32'hb90c292e),
	.w4(32'hba849c41),
	.w5(32'hba915d5d),
	.w6(32'hbabc726a),
	.w7(32'hbab7423e),
	.w8(32'hbabdf99d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad701dd),
	.w1(32'hb8f57f32),
	.w2(32'hba379082),
	.w3(32'hbaec8706),
	.w4(32'hb98856ef),
	.w5(32'hba595b05),
	.w6(32'hba3e0314),
	.w7(32'hba6719ee),
	.w8(32'hba8a20ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50912a),
	.w1(32'h36a0acd7),
	.w2(32'hbafb57e5),
	.w3(32'hba51bbf1),
	.w4(32'hb9062426),
	.w5(32'h393bf087),
	.w6(32'h3908e6b0),
	.w7(32'hba997740),
	.w8(32'hb9a7cd24),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9517353),
	.w1(32'h3a0b9679),
	.w2(32'h3a950d7f),
	.w3(32'h387aaddc),
	.w4(32'hb918583d),
	.w5(32'h3ad68233),
	.w6(32'h3ad63088),
	.w7(32'h3a823f4e),
	.w8(32'h3ac7813a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6cd49),
	.w1(32'h3a76eb46),
	.w2(32'h3ab5cb0b),
	.w3(32'h3b386968),
	.w4(32'h3a11c00b),
	.w5(32'h3aa6c00e),
	.w6(32'h398029f8),
	.w7(32'h3a08d264),
	.w8(32'h3a8dbc19),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7512d),
	.w1(32'hb73a6967),
	.w2(32'h397c66f6),
	.w3(32'h3ac47a9f),
	.w4(32'h39944572),
	.w5(32'h39ab0b5d),
	.w6(32'hb8bada86),
	.w7(32'hb74173de),
	.w8(32'h395f43b3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d5fe0),
	.w1(32'h39cb34bc),
	.w2(32'h3a25d5a0),
	.w3(32'hb98808be),
	.w4(32'h395d0d7b),
	.w5(32'h3a0ae962),
	.w6(32'h382c1b6f),
	.w7(32'h3922bccc),
	.w8(32'h39b3d981),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b41fc),
	.w1(32'hb9a8b9d9),
	.w2(32'h38e30dc7),
	.w3(32'h3a1af739),
	.w4(32'hb9f06737),
	.w5(32'hb92b4bd1),
	.w6(32'hb9bebdcc),
	.w7(32'h3808831b),
	.w8(32'hb76cae22),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd73d7),
	.w1(32'hba805595),
	.w2(32'hba2d92e4),
	.w3(32'hb935d801),
	.w4(32'hbab3048d),
	.w5(32'hbadc754d),
	.w6(32'hba951673),
	.w7(32'hba9859a0),
	.w8(32'hbaa439bd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b4d7e),
	.w1(32'h391f50ac),
	.w2(32'hb6c7269e),
	.w3(32'hbae5fedc),
	.w4(32'h388a1154),
	.w5(32'hb92c9962),
	.w6(32'h38d9cfb2),
	.w7(32'hb8944413),
	.w8(32'hb86d15dd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a21848),
	.w1(32'h3a3b57d2),
	.w2(32'h3a60e12b),
	.w3(32'hb911adc2),
	.w4(32'h39f96778),
	.w5(32'h3a462daa),
	.w6(32'h389a9d47),
	.w7(32'h394586c9),
	.w8(32'h3a0c8f0d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a625e60),
	.w1(32'hb831117a),
	.w2(32'hb917b831),
	.w3(32'h3a55e348),
	.w4(32'hb8dd6280),
	.w5(32'hba7727d0),
	.w6(32'hb903114e),
	.w7(32'hb7ba8a8b),
	.w8(32'hb893437d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9012dda),
	.w1(32'hb93cbd9d),
	.w2(32'h3886fff7),
	.w3(32'hba16270e),
	.w4(32'hb9e4f985),
	.w5(32'hba29269d),
	.w6(32'hba411718),
	.w7(32'hb98e0adb),
	.w8(32'hb883a6c8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c54250),
	.w1(32'h39d1ba75),
	.w2(32'hbb227041),
	.w3(32'hb9d41506),
	.w4(32'hba23060d),
	.w5(32'hbb2b6552),
	.w6(32'hb7dc9d38),
	.w7(32'hbabbd5d9),
	.w8(32'hb9ea7d96),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd23ed),
	.w1(32'hb9eb723d),
	.w2(32'hb9847d11),
	.w3(32'hbb015b38),
	.w4(32'hb993c90e),
	.w5(32'hba144701),
	.w6(32'hba46a03e),
	.w7(32'hb9b4cba0),
	.w8(32'hb98e2fc7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1da3f),
	.w1(32'hba99f6f9),
	.w2(32'hba69c460),
	.w3(32'hba11570e),
	.w4(32'hbab0ecc6),
	.w5(32'hbace0d04),
	.w6(32'hba892dd2),
	.w7(32'hba461d91),
	.w8(32'hba3c2803),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa29c95),
	.w1(32'hb9dbe09d),
	.w2(32'hb987b3d2),
	.w3(32'hbacd6cd4),
	.w4(32'hba1e6e56),
	.w5(32'hba8c51b8),
	.w6(32'hb9cc96eb),
	.w7(32'hb8d9ea89),
	.w8(32'h39845412),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a76b8f),
	.w1(32'h3a1abebd),
	.w2(32'h3a6ed05c),
	.w3(32'hba22c97c),
	.w4(32'h39a570ae),
	.w5(32'h3a57d0cb),
	.w6(32'h38d381bc),
	.w7(32'h398f0de1),
	.w8(32'h3a3c07bb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a968dc8),
	.w1(32'hb846d946),
	.w2(32'h391c02a6),
	.w3(32'h3a8e5f94),
	.w4(32'hb8c4d4b6),
	.w5(32'h389b72fa),
	.w6(32'hb94eba20),
	.w7(32'hb8dac9cd),
	.w8(32'h38269c20),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d9fd3),
	.w1(32'h37c6ea20),
	.w2(32'h397e00be),
	.w3(32'h388ba189),
	.w4(32'hb908d2ec),
	.w5(32'h38c82869),
	.w6(32'hb9a71116),
	.w7(32'hb947b6fd),
	.w8(32'hb887400d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977d53b),
	.w1(32'hb99cfaa6),
	.w2(32'h38a70a9d),
	.w3(32'h38a9f53e),
	.w4(32'h39a5c27d),
	.w5(32'h399bab3c),
	.w6(32'hb9613445),
	.w7(32'h3a58909d),
	.w8(32'hb97b4c09),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9daff22),
	.w1(32'hbaab6319),
	.w2(32'hbadf82c0),
	.w3(32'hb9e7d18c),
	.w4(32'hba92fbfb),
	.w5(32'hbae78f1e),
	.w6(32'hba99cefc),
	.w7(32'hba95f2a9),
	.w8(32'hba1c1d66),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a05a9),
	.w1(32'h3a0cff45),
	.w2(32'h3a6f8d56),
	.w3(32'hba4c2ef3),
	.w4(32'h399c2593),
	.w5(32'h3a6ac61b),
	.w6(32'h3a0b8111),
	.w7(32'h39b7d805),
	.w8(32'h3a1c1291),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087069),
	.w1(32'hb84aef6d),
	.w2(32'h39d8e280),
	.w3(32'h39be5de3),
	.w4(32'h393154bd),
	.w5(32'h39b5c6d8),
	.w6(32'hb9a281fd),
	.w7(32'h3929b6d8),
	.w8(32'hb8b6c77a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f6b958),
	.w1(32'hb99a802d),
	.w2(32'hb8c6d492),
	.w3(32'h3982c08a),
	.w4(32'hb9a1d58f),
	.w5(32'hb961f87c),
	.w6(32'hba0e1a5f),
	.w7(32'hb9a6a36b),
	.w8(32'hb8e76ff2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bbf2e),
	.w1(32'hbac74bf0),
	.w2(32'hba57600a),
	.w3(32'hb982402f),
	.w4(32'h3a77ae99),
	.w5(32'h3ab8f463),
	.w6(32'hb7f0dbe3),
	.w7(32'h3abbe4ae),
	.w8(32'h3988d42b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf713),
	.w1(32'hba94e3bd),
	.w2(32'hba0b54f7),
	.w3(32'h39de9bd6),
	.w4(32'hba1c64e0),
	.w5(32'hba26fcc5),
	.w6(32'hbabfb660),
	.w7(32'hbab88b7c),
	.w8(32'hbad8cf48),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98e3b1),
	.w1(32'hb9957e58),
	.w2(32'h3912efa8),
	.w3(32'hbac7cfee),
	.w4(32'hb9a88574),
	.w5(32'hb84a7b21),
	.w6(32'hb9316194),
	.w7(32'hb8000934),
	.w8(32'hb8130f10),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fa5f74),
	.w1(32'hb9b6fbc1),
	.w2(32'hb9deb8b7),
	.w3(32'hb823f107),
	.w4(32'hb8f19327),
	.w5(32'hb96a1b57),
	.w6(32'hb8cc4c24),
	.w7(32'hb9a09667),
	.w8(32'hb90f4270),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9420e49),
	.w1(32'hb9c7f168),
	.w2(32'hb9d73c1c),
	.w3(32'hb939dcf7),
	.w4(32'hb95c2cd1),
	.w5(32'hb99bf3c3),
	.w6(32'hb9a471c0),
	.w7(32'hb9bc91b6),
	.w8(32'hb97c3132),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977b0d5),
	.w1(32'hb96287e7),
	.w2(32'h3a1c97a0),
	.w3(32'hb921e304),
	.w4(32'hb8216000),
	.w5(32'h388c1ff8),
	.w6(32'hb8355706),
	.w7(32'h39718b21),
	.w8(32'h391b348e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394473b2),
	.w1(32'h395c4bb4),
	.w2(32'h39c3672b),
	.w3(32'h39ee54bc),
	.w4(32'h392e34ea),
	.w5(32'h39a7e954),
	.w6(32'h390ac4c2),
	.w7(32'h39804c3e),
	.w8(32'h38c7e0c4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39328e58),
	.w1(32'h38ceaf8a),
	.w2(32'h391c38ec),
	.w3(32'h39a700f4),
	.w4(32'hb8d2be53),
	.w5(32'hb6a6bfba),
	.w6(32'h38ac77c1),
	.w7(32'h38ef59d9),
	.w8(32'hb85652ac),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e610ed),
	.w1(32'hb9a76f25),
	.w2(32'hba02964e),
	.w3(32'hb8e40f89),
	.w4(32'h3941b72f),
	.w5(32'hb8327231),
	.w6(32'hb85d74c6),
	.w7(32'hb63a3ff0),
	.w8(32'h38ada944),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9997657),
	.w1(32'hb8fce1ce),
	.w2(32'h394f19eb),
	.w3(32'hb9468db7),
	.w4(32'h3930ac62),
	.w5(32'h39a91bdb),
	.w6(32'hb99d59b1),
	.w7(32'h3951c70f),
	.w8(32'h39bb1cfb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac0ad5),
	.w1(32'hb9b50024),
	.w2(32'hb9c9bb9d),
	.w3(32'hb8c5cd69),
	.w4(32'h36ac2f10),
	.w5(32'hb974883f),
	.w6(32'hb9bea5b0),
	.w7(32'hb9f67638),
	.w8(32'hb9a8d443),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8d48f),
	.w1(32'h386e3543),
	.w2(32'h393c9863),
	.w3(32'hb982791b),
	.w4(32'h382a6dfd),
	.w5(32'h39833d5a),
	.w6(32'h38bc49eb),
	.w7(32'h396a862f),
	.w8(32'h3739a798),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d4d0f6),
	.w1(32'hb9860360),
	.w2(32'hb9e25c33),
	.w3(32'h39228dac),
	.w4(32'hb7b01cc1),
	.w5(32'hb95e6c75),
	.w6(32'hb934b75c),
	.w7(32'hb99e7a14),
	.w8(32'hb927b84d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98875eb),
	.w1(32'hb9caf5e3),
	.w2(32'hb9df96cd),
	.w3(32'hb9010d4e),
	.w4(32'hb99cef8d),
	.w5(32'hb9f41fec),
	.w6(32'hb9a04996),
	.w7(32'hb9ccc23c),
	.w8(32'hb999ed45),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99173d2),
	.w1(32'h3a5f7f26),
	.w2(32'h3a2d0099),
	.w3(32'hb97c7b3c),
	.w4(32'h3a6d1fd6),
	.w5(32'h3a285bd2),
	.w6(32'h3a511f80),
	.w7(32'h3a1181a8),
	.w8(32'h39d80eaa),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c72b23),
	.w1(32'hba0ae760),
	.w2(32'hb9a9444e),
	.w3(32'h3a17d79a),
	.w4(32'hb909649f),
	.w5(32'h371db3e6),
	.w6(32'hba027809),
	.w7(32'hb95d0993),
	.w8(32'hb8d4bbfe),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9178d3b),
	.w1(32'hb99d8e7f),
	.w2(32'hba19e469),
	.w3(32'h38992687),
	.w4(32'hb9456b95),
	.w5(32'hba0bb825),
	.w6(32'hb983d770),
	.w7(32'hb990db78),
	.w8(32'hb92db195),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b9f0f),
	.w1(32'hb9ff2b6e),
	.w2(32'hb9a87441),
	.w3(32'hba1d819d),
	.w4(32'hb98d30a0),
	.w5(32'hb9598cbc),
	.w6(32'hb993f29b),
	.w7(32'hb99d29ca),
	.w8(32'hb9795d45),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9368f1c),
	.w1(32'hb99d2669),
	.w2(32'hba0f9f13),
	.w3(32'hb97a1a3d),
	.w4(32'hb7b2ef15),
	.w5(32'hb9889946),
	.w6(32'hb9117772),
	.w7(32'hb9e26ec6),
	.w8(32'hb953d5ec),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1fd16),
	.w1(32'hb8ba5ff2),
	.w2(32'hb87b0b65),
	.w3(32'hb8914485),
	.w4(32'h39f9238b),
	.w5(32'h3935736b),
	.w6(32'hb998be73),
	.w7(32'h39aec472),
	.w8(32'h3a0db046),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b55c3),
	.w1(32'hb9883bb2),
	.w2(32'hb9b4ffa2),
	.w3(32'hb964aaed),
	.w4(32'hb92d4a34),
	.w5(32'hb98cfd57),
	.w6(32'hb9847a44),
	.w7(32'hb998588c),
	.w8(32'hb932a84c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966e63f),
	.w1(32'h394bc95f),
	.w2(32'h38c9133a),
	.w3(32'hb8ea2dc6),
	.w4(32'h37865770),
	.w5(32'h38919ad8),
	.w6(32'h3842c276),
	.w7(32'h386b707e),
	.w8(32'h383abc77),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783e4d1),
	.w1(32'h39aaeeca),
	.w2(32'h39e04799),
	.w3(32'hb8e67472),
	.w4(32'h39a6f506),
	.w5(32'h39cfff76),
	.w6(32'h39bdf8bf),
	.w7(32'h39e0ffba),
	.w8(32'h39a66441),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1d011),
	.w1(32'h370062b0),
	.w2(32'h392630be),
	.w3(32'h398bf803),
	.w4(32'h37c6808a),
	.w5(32'h375d1fa3),
	.w6(32'hb8776cb0),
	.w7(32'h375d8fae),
	.w8(32'hb916319d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b69895),
	.w1(32'hb9c56860),
	.w2(32'hb9bc7b83),
	.w3(32'hb7e82aeb),
	.w4(32'hb99d3e7e),
	.w5(32'hb9c4dcc6),
	.w6(32'hb9c8d139),
	.w7(32'hb9ce8da2),
	.w8(32'hb989a8c0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a30ee3),
	.w1(32'hb9c85f79),
	.w2(32'hba52b23c),
	.w3(32'hb98de06e),
	.w4(32'hb9845604),
	.w5(32'hba0af5ec),
	.w6(32'hb929c412),
	.w7(32'hba19d656),
	.w8(32'hb980b830),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e00a79),
	.w1(32'hba8618de),
	.w2(32'hba5687ac),
	.w3(32'hb9b50c48),
	.w4(32'hba4926e0),
	.w5(32'hba154da0),
	.w6(32'hb99a37c4),
	.w7(32'hb9671882),
	.w8(32'hb9b6f7ed),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2f59),
	.w1(32'hb72e8c5c),
	.w2(32'hb938e12d),
	.w3(32'hba2c4479),
	.w4(32'hb9112769),
	.w5(32'hb99932ac),
	.w6(32'h3935965e),
	.w7(32'hb7daf40a),
	.w8(32'h3911bc8f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398edd68),
	.w1(32'hb9bab6b5),
	.w2(32'hb9faf49c),
	.w3(32'hb87c6f4b),
	.w4(32'hb8e7ea07),
	.w5(32'hb984564b),
	.w6(32'hb96236a6),
	.w7(32'hb9a96e19),
	.w8(32'hb9629a5f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995941e),
	.w1(32'hb8437139),
	.w2(32'hb992b97f),
	.w3(32'hb90b82d5),
	.w4(32'h399cd2ab),
	.w5(32'h391278fb),
	.w6(32'hb9797bab),
	.w7(32'hb94c4646),
	.w8(32'hb899cbd6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9392394),
	.w1(32'h39810668),
	.w2(32'h39972117),
	.w3(32'h391c792e),
	.w4(32'hb8269d4e),
	.w5(32'hb79681f8),
	.w6(32'hb6246cef),
	.w7(32'h394660a5),
	.w8(32'h37ec7609),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39550f8d),
	.w1(32'hb961f1eb),
	.w2(32'hb974df5c),
	.w3(32'h398c02dc),
	.w4(32'hb93733c0),
	.w5(32'hb9a7e270),
	.w6(32'hb9691d8c),
	.w7(32'hb962032c),
	.w8(32'hb7dc9a1d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9657343),
	.w1(32'hb8edcdf0),
	.w2(32'h3900f09d),
	.w3(32'hb933dbc5),
	.w4(32'h385d689f),
	.w5(32'h378e13b5),
	.w6(32'hb98a3075),
	.w7(32'hb95c005d),
	.w8(32'hb92c82c6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2ee1d),
	.w1(32'h39093a31),
	.w2(32'hba0af989),
	.w3(32'h37da7b82),
	.w4(32'hb785f546),
	.w5(32'hb9c47e51),
	.w6(32'h391d561f),
	.w7(32'hb9e25d3e),
	.w8(32'hb94bfe76),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ab784),
	.w1(32'h39a5d37b),
	.w2(32'hb946e692),
	.w3(32'hb8d5fd66),
	.w4(32'h39a9e0f5),
	.w5(32'hb8ade086),
	.w6(32'h39852bc9),
	.w7(32'hb97f574c),
	.w8(32'hb9c6100e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940c40d),
	.w1(32'hb999a117),
	.w2(32'hb9e11840),
	.w3(32'hb8721c1e),
	.w4(32'hb93996e4),
	.w5(32'hb98e6553),
	.w6(32'hb96356b9),
	.w7(32'hb9c65cfa),
	.w8(32'hb920da75),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d25e8),
	.w1(32'hb9c3dc70),
	.w2(32'hb9bdd827),
	.w3(32'hb9129381),
	.w4(32'hb96d0f37),
	.w5(32'hb992a1a9),
	.w6(32'hb9a8b37c),
	.w7(32'hb9dc1118),
	.w8(32'hb9856b2d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977071d),
	.w1(32'hb9e283e3),
	.w2(32'hb9981620),
	.w3(32'hb95004af),
	.w4(32'hba0df802),
	.w5(32'hba248316),
	.w6(32'hb9b4a07c),
	.w7(32'hba1effab),
	.w8(32'hb9c901de),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0885c9),
	.w1(32'h39254f3c),
	.w2(32'h3991e202),
	.w3(32'hb9acc466),
	.w4(32'h3991d7c4),
	.w5(32'h3954cf31),
	.w6(32'h39676cbe),
	.w7(32'hb939ba7d),
	.w8(32'hba22f6f5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba156ba7),
	.w1(32'h39d6a5dc),
	.w2(32'h39ecc688),
	.w3(32'hb9ba15fe),
	.w4(32'h3a09da98),
	.w5(32'h39e3f08a),
	.w6(32'h39a40bdf),
	.w7(32'h399cde27),
	.w8(32'h396599da),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966f5bd),
	.w1(32'hb9b28c77),
	.w2(32'hb9bd8882),
	.w3(32'h39ee347b),
	.w4(32'hb94c9ff9),
	.w5(32'hb9a65b4d),
	.w6(32'hb97d140b),
	.w7(32'hb9c2fda0),
	.w8(32'hb9394b3a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0895e),
	.w1(32'hb8f4adc4),
	.w2(32'hb7abaf9a),
	.w3(32'hb9aedcad),
	.w4(32'h392c4a56),
	.w5(32'h39005169),
	.w6(32'hb94ff815),
	.w7(32'h38d972ab),
	.w8(32'h38d0b224),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eeb86d),
	.w1(32'h39d7d489),
	.w2(32'h39ed7dd3),
	.w3(32'h38963d66),
	.w4(32'h39aba369),
	.w5(32'h39f315f4),
	.w6(32'h39a2e463),
	.w7(32'h39d2c93e),
	.w8(32'h3908756d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f19b5),
	.w1(32'hb9b6f52f),
	.w2(32'hb9e1032f),
	.w3(32'h3984ec8b),
	.w4(32'hb958c998),
	.w5(32'hb9ae5d09),
	.w6(32'hb97793cc),
	.w7(32'hb9baf48c),
	.w8(32'hb977c9dc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c282ed),
	.w1(32'h38b45a48),
	.w2(32'h399947e6),
	.w3(32'hb97dbc88),
	.w4(32'h38e43db8),
	.w5(32'h396333f8),
	.w6(32'hb76f1e37),
	.w7(32'h39703347),
	.w8(32'h38aac4a5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3826b69f),
	.w1(32'h3957fe7a),
	.w2(32'hb939f425),
	.w3(32'h38242bcf),
	.w4(32'h38d842d9),
	.w5(32'hb960ca96),
	.w6(32'h39981a11),
	.w7(32'hb990da3c),
	.w8(32'hba0126dd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c94c37),
	.w1(32'hb9562060),
	.w2(32'hb952ced6),
	.w3(32'hb943581f),
	.w4(32'h391663fc),
	.w5(32'h390cbeb5),
	.w6(32'hb99f8fc4),
	.w7(32'hb8263a37),
	.w8(32'hb89a538e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d1229),
	.w1(32'hb9bd8094),
	.w2(32'hb98d648f),
	.w3(32'hb90d7876),
	.w4(32'hb9ac9a71),
	.w5(32'hb9bd08bf),
	.w6(32'hb9984824),
	.w7(32'hb9d1f3d6),
	.w8(32'hb9bb3f77),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb13cf),
	.w1(32'h3ab05e12),
	.w2(32'h3a7c1693),
	.w3(32'hb9932d90),
	.w4(32'h3ac01cae),
	.w5(32'h3a9c9e29),
	.w6(32'h3acc68f4),
	.w7(32'h3aa76199),
	.w8(32'h3a843478),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e2d23),
	.w1(32'h384e78ad),
	.w2(32'h39126767),
	.w3(32'h3a82e4f8),
	.w4(32'h37a88415),
	.w5(32'h390523ca),
	.w6(32'h39a84971),
	.w7(32'h391a897a),
	.w8(32'h389f4b4e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997777c),
	.w1(32'hb9ae3c01),
	.w2(32'hb95fa356),
	.w3(32'hb894680a),
	.w4(32'hb9187147),
	.w5(32'hb91bf2a2),
	.w6(32'hb906d6b1),
	.w7(32'h3892cc41),
	.w8(32'h390a8fa2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a340d8),
	.w1(32'h38d155d9),
	.w2(32'hb9c63b64),
	.w3(32'hb964f440),
	.w4(32'h39bada88),
	.w5(32'h36ed2737),
	.w6(32'h3908f730),
	.w7(32'h39daca82),
	.w8(32'h39a45c43),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a4e201),
	.w1(32'h393421e0),
	.w2(32'hb9c26370),
	.w3(32'hb9911d37),
	.w4(32'h38e9b262),
	.w5(32'hb9780403),
	.w6(32'h3987b2fe),
	.w7(32'hb9a4109a),
	.w8(32'hb9b0d58d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2f221),
	.w1(32'hba02dd9f),
	.w2(32'hb9b93a61),
	.w3(32'hb9b83678),
	.w4(32'hb9c8d8a6),
	.w5(32'hb9c621c7),
	.w6(32'hb9f5e28c),
	.w7(32'hba0a7c88),
	.w8(32'hb9d4b01b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c56edd),
	.w1(32'hb9a5ce02),
	.w2(32'hb9db23eb),
	.w3(32'hb9a91fa8),
	.w4(32'hb8f12efc),
	.w5(32'hb931bc52),
	.w6(32'hb9329dd2),
	.w7(32'hb980a130),
	.w8(32'hb823120f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917641a),
	.w1(32'h39a604aa),
	.w2(32'h38e76f27),
	.w3(32'h35fe3ff3),
	.w4(32'h394fc3ca),
	.w5(32'h39297b50),
	.w6(32'h3971c5fd),
	.w7(32'h39b20ded),
	.w8(32'h39eda6a7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fe31e),
	.w1(32'h398751bb),
	.w2(32'h390f2e02),
	.w3(32'h39a97902),
	.w4(32'h39141234),
	.w5(32'hb8ebe259),
	.w6(32'h39b391e1),
	.w7(32'h39e39078),
	.w8(32'h39824dac),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ab024),
	.w1(32'h3928e1ae),
	.w2(32'h36b0a179),
	.w3(32'h39d9ee74),
	.w4(32'h39d18062),
	.w5(32'h3931b2f3),
	.w6(32'hb4b9deb3),
	.w7(32'hb907f44f),
	.w8(32'h391536c3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c3410),
	.w1(32'hba150a8e),
	.w2(32'hb99a0126),
	.w3(32'h39a112e6),
	.w4(32'hb9cfca06),
	.w5(32'hb8310d6f),
	.w6(32'hba03f6b2),
	.w7(32'hb98cd079),
	.w8(32'hb9296fcb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d028c2),
	.w1(32'h39c3871e),
	.w2(32'h39e9ebe5),
	.w3(32'hb941a19f),
	.w4(32'h39c6ee93),
	.w5(32'h39db61b5),
	.w6(32'h3910eddb),
	.w7(32'h394431e0),
	.w8(32'h374a3fa5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e20b93),
	.w1(32'h393d2375),
	.w2(32'hb9d9dbee),
	.w3(32'h393744ed),
	.w4(32'h39ac66d8),
	.w5(32'hb8a806bb),
	.w6(32'h39c9d57c),
	.w7(32'hb9c6768b),
	.w8(32'hb89234b7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37be3e0b),
	.w1(32'h3a0bcd76),
	.w2(32'h3a4eb88c),
	.w3(32'h398269b1),
	.w4(32'h39b28de1),
	.w5(32'h3a334bea),
	.w6(32'h39913996),
	.w7(32'h3a0b68ec),
	.w8(32'h39b7b0eb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997a649),
	.w1(32'hba0eac5c),
	.w2(32'hb7c0ec4a),
	.w3(32'h39ae3d25),
	.w4(32'hb96dbc82),
	.w5(32'hb86fcb42),
	.w6(32'hba37be62),
	.w7(32'hb8d4669c),
	.w8(32'h383d80b5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984409f),
	.w1(32'h37e9c0b3),
	.w2(32'h3946c3d0),
	.w3(32'h3800b9c5),
	.w4(32'h38d72327),
	.w5(32'h3946bf67),
	.w6(32'hb70df95e),
	.w7(32'h38f0caed),
	.w8(32'hb8c6584c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852f1eb),
	.w1(32'hb9c725fa),
	.w2(32'hba00968c),
	.w3(32'h3963df37),
	.w4(32'hb95b6212),
	.w5(32'hb9edb7c0),
	.w6(32'hb9883a18),
	.w7(32'hb9fed877),
	.w8(32'hb9d7f678),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99533bc),
	.w1(32'h393179d4),
	.w2(32'h3987bf09),
	.w3(32'hb9564421),
	.w4(32'h37eaf3f2),
	.w5(32'h3916e8b1),
	.w6(32'h37c89673),
	.w7(32'h398061bf),
	.w8(32'hb8cdaa4d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377112c1),
	.w1(32'hba0c410f),
	.w2(32'hb9f1f941),
	.w3(32'h39356482),
	.w4(32'hb99bf4d2),
	.w5(32'hb994f16f),
	.w6(32'hb9305e86),
	.w7(32'hb937c17a),
	.w8(32'hb7a43f8d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a8183),
	.w1(32'hb9ab5fad),
	.w2(32'h3a04beea),
	.w3(32'hb93e1032),
	.w4(32'hba0ccc39),
	.w5(32'hb9a6ee0e),
	.w6(32'hb9310237),
	.w7(32'hb8b2113c),
	.w8(32'hb985c9db),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963983b),
	.w1(32'h3a52da8b),
	.w2(32'h3a154f73),
	.w3(32'hb9b33825),
	.w4(32'h3a5e3d8e),
	.w5(32'h3a2a9193),
	.w6(32'h3a759e90),
	.w7(32'h3a3cc1d1),
	.w8(32'h3a052d1d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd2b00),
	.w1(32'hb916ecbe),
	.w2(32'hb4f39894),
	.w3(32'h3a2424e5),
	.w4(32'hb85eb191),
	.w5(32'h36c0ddc2),
	.w6(32'hb8c5bab8),
	.w7(32'hb8f12950),
	.w8(32'hb80e1dd7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c58df7),
	.w1(32'hb9a7dbb7),
	.w2(32'hb9140a1f),
	.w3(32'hb74561c7),
	.w4(32'hb9509beb),
	.w5(32'hb900ff17),
	.w6(32'hb935d92f),
	.w7(32'hb8a3d269),
	.w8(32'hb9823d73),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee3cd3),
	.w1(32'h392ff99f),
	.w2(32'h38802b53),
	.w3(32'hb92ebb6f),
	.w4(32'h3911de57),
	.w5(32'hb886f1fe),
	.w6(32'h387d8341),
	.w7(32'hb889708c),
	.w8(32'hb9a40c48),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913d2d9),
	.w1(32'h3994cd69),
	.w2(32'hb9f0126a),
	.w3(32'hb92dcc22),
	.w4(32'h398c799d),
	.w5(32'hb98ddc40),
	.w6(32'h39f23840),
	.w7(32'hb98a2153),
	.w8(32'hb9b33134),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b31871),
	.w1(32'hb9b23baa),
	.w2(32'hba0a6ed0),
	.w3(32'hb9d10470),
	.w4(32'hb952ce32),
	.w5(32'hb9b7d5df),
	.w6(32'hb9a63fdb),
	.w7(32'hb9d3ffa9),
	.w8(32'hb979dd48),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cea5d2),
	.w1(32'hb9624690),
	.w2(32'hb8ce3f25),
	.w3(32'hb94254c9),
	.w4(32'h385d4f2f),
	.w5(32'h38908939),
	.w6(32'hb9562711),
	.w7(32'h394f60fa),
	.w8(32'h3a0a9c8e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05432a),
	.w1(32'h39554674),
	.w2(32'h39d3238e),
	.w3(32'h3a01c162),
	.w4(32'h396c61ea),
	.w5(32'h39b94f12),
	.w6(32'h3971aac6),
	.w7(32'h39aa7007),
	.w8(32'h395c815e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395fcd53),
	.w1(32'hb9bc2abb),
	.w2(32'hb9cb26ff),
	.w3(32'h39444094),
	.w4(32'hb98a918c),
	.w5(32'hb9753b83),
	.w6(32'hb99ab7d6),
	.w7(32'hb9b5bcb1),
	.w8(32'hb93d8559),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9759039),
	.w1(32'hb9ab618b),
	.w2(32'hb9d9fd4c),
	.w3(32'hb956ca27),
	.w4(32'hb954f9b2),
	.w5(32'hb9a46cba),
	.w6(32'hb955512b),
	.w7(32'hb9ba4042),
	.w8(32'hb97a8d33),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a11f45),
	.w1(32'hb9f03de2),
	.w2(32'hba0f7a81),
	.w3(32'hb9576b40),
	.w4(32'hb9b1eba8),
	.w5(32'hb9e87822),
	.w6(32'hb9d9375c),
	.w7(32'hba18ec8d),
	.w8(32'hb9be2422),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2ccc8),
	.w1(32'h37e92db4),
	.w2(32'h3797ca59),
	.w3(32'hb9a05ab7),
	.w4(32'h394b8980),
	.w5(32'h39427171),
	.w6(32'hb8892656),
	.w7(32'h37dee87a),
	.w8(32'hb7ebe1aa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f4926),
	.w1(32'h371af25c),
	.w2(32'hba814b38),
	.w3(32'h392ffa1c),
	.w4(32'hb9127295),
	.w5(32'hb9e0017e),
	.w6(32'hb7d572f7),
	.w7(32'h38d830d2),
	.w8(32'hb8f422fd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77e753),
	.w1(32'hb99a5dc0),
	.w2(32'hba26f240),
	.w3(32'hb938e8c1),
	.w4(32'h385c8cff),
	.w5(32'hb981ff43),
	.w6(32'hb79f0b7e),
	.w7(32'hb997fb19),
	.w8(32'h368fb802),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9852dfb),
	.w1(32'hb8853386),
	.w2(32'h398a82b4),
	.w3(32'hb830f02e),
	.w4(32'hb8e2e77a),
	.w5(32'h37fb0181),
	.w6(32'hb7ede13a),
	.w7(32'h38b462dd),
	.w8(32'hb902f047),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5222759),
	.w1(32'h3923ede3),
	.w2(32'h399a831c),
	.w3(32'h38b5709a),
	.w4(32'hb8cb9912),
	.w5(32'hb7615c95),
	.w6(32'hb84e9247),
	.w7(32'h392f4365),
	.w8(32'hb92d764e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7a6d7),
	.w1(32'hb9baf999),
	.w2(32'hba1bca52),
	.w3(32'hb952da38),
	.w4(32'hb98fcc87),
	.w5(32'hb9dd2ff2),
	.w6(32'hb99a218d),
	.w7(32'hba14919a),
	.w8(32'hb975dfaa),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968d3e2),
	.w1(32'h39ecffdc),
	.w2(32'hb96b96d3),
	.w3(32'hb91e2107),
	.w4(32'h3a14d441),
	.w5(32'hb79654da),
	.w6(32'h3a19a302),
	.w7(32'hb91d9c61),
	.w8(32'hb8f1ba6d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969b16d),
	.w1(32'h389d78be),
	.w2(32'h38e5d23f),
	.w3(32'hb92041b7),
	.w4(32'h3954eee2),
	.w5(32'h39b109b5),
	.w6(32'hb8c2b988),
	.w7(32'hb8714073),
	.w8(32'hb8cd32ce),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373dcbd7),
	.w1(32'h38a8693b),
	.w2(32'hb895c5fe),
	.w3(32'h3967db67),
	.w4(32'h3918f162),
	.w5(32'h36a92ec5),
	.w6(32'h38040d3e),
	.w7(32'hb8dcc3a6),
	.w8(32'hb6e4807b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8400a32),
	.w1(32'h38c2d536),
	.w2(32'h399f7f83),
	.w3(32'h391a2165),
	.w4(32'h3912f2ae),
	.w5(32'h395a4b7f),
	.w6(32'h386c2388),
	.w7(32'h390aa461),
	.w8(32'hb8448eb3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9554325),
	.w1(32'h38f02459),
	.w2(32'hb9b3cc19),
	.w3(32'h3886c1f9),
	.w4(32'h39904ae3),
	.w5(32'hb969f620),
	.w6(32'hb90a5350),
	.w7(32'hba11382c),
	.w8(32'hb97ec7bb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7857358),
	.w1(32'h39d5df19),
	.w2(32'h39fe5c4d),
	.w3(32'hb930ed3c),
	.w4(32'h39a6d88e),
	.w5(32'h39eb0478),
	.w6(32'h39a932e3),
	.w7(32'h39dd6a6b),
	.w8(32'h398e19c8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b591e6),
	.w1(32'h39e93d1f),
	.w2(32'h3a190d44),
	.w3(32'h39df3e43),
	.w4(32'h3a10794e),
	.w5(32'h39f50fd6),
	.w6(32'h39db7d48),
	.w7(32'h39c8f5af),
	.w8(32'h39996b3c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c10197),
	.w1(32'hb988dc8b),
	.w2(32'hb9eb243d),
	.w3(32'h39e2c606),
	.w4(32'hb9309753),
	.w5(32'hb991235f),
	.w6(32'hb9214d72),
	.w7(32'hb9beb824),
	.w8(32'hb9127f22),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cd32e),
	.w1(32'h39858343),
	.w2(32'h39773dbc),
	.w3(32'hb8e6c987),
	.w4(32'h39aab40e),
	.w5(32'h39a8d2ed),
	.w6(32'h35089aec),
	.w7(32'h37088910),
	.w8(32'hb892e625),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a18dd),
	.w1(32'hb9befc1e),
	.w2(32'hb9e15efe),
	.w3(32'h38803f8b),
	.w4(32'hb94250e2),
	.w5(32'hb9a0be05),
	.w6(32'hb90cc835),
	.w7(32'hb99327c7),
	.w8(32'hb89c5e90),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941d96f),
	.w1(32'hb993f2a6),
	.w2(32'hb9f7f30b),
	.w3(32'hb8c6109a),
	.w4(32'hb919e930),
	.w5(32'hb98fb5f4),
	.w6(32'hb9688cd6),
	.w7(32'hb9df3ff2),
	.w8(32'hb990d063),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d55f5),
	.w1(32'h3a3cda8c),
	.w2(32'h3a26a7df),
	.w3(32'hb927a8d8),
	.w4(32'h3a2c383e),
	.w5(32'h3a18f4c7),
	.w6(32'h3a351b80),
	.w7(32'h3a288077),
	.w8(32'h39ddc671),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b29eb5),
	.w1(32'h375dec52),
	.w2(32'hb7d84867),
	.w3(32'h39b07d6f),
	.w4(32'h38858fe0),
	.w5(32'h38353a2c),
	.w6(32'hb844d1b4),
	.w7(32'hb8fcba73),
	.w8(32'hb86729ee),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ef9dc),
	.w1(32'h399df67d),
	.w2(32'hb9e0dae3),
	.w3(32'h38ed19ca),
	.w4(32'h39a2f567),
	.w5(32'hb996317c),
	.w6(32'h39f87eed),
	.w7(32'hb9a4d8a8),
	.w8(32'hb918ff4a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9312cf4),
	.w1(32'h36e7340f),
	.w2(32'h39310a9f),
	.w3(32'hb89b43b6),
	.w4(32'hb89f2027),
	.w5(32'hb7f1d6e1),
	.w6(32'hb8960ec4),
	.w7(32'h381e6b90),
	.w8(32'hb8444916),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3848a91d),
	.w1(32'hba1715b0),
	.w2(32'hba108525),
	.w3(32'h37b5109e),
	.w4(32'hb9aa47b4),
	.w5(32'hb8ec9790),
	.w6(32'hb9c0697e),
	.w7(32'hba0c087c),
	.w8(32'hb9f6ff5b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cd4c3),
	.w1(32'h39e8aaed),
	.w2(32'h39ef87cb),
	.w3(32'hb42f270e),
	.w4(32'h3966c5f6),
	.w5(32'h3940f58f),
	.w6(32'h39e8917b),
	.w7(32'h3a0b68f5),
	.w8(32'h39abf09f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d16f69),
	.w1(32'hb927008c),
	.w2(32'h37e859f9),
	.w3(32'h37c27e12),
	.w4(32'hb9b441de),
	.w5(32'hb9ee629f),
	.w6(32'h37fea17f),
	.w7(32'h385fe588),
	.w8(32'hb97a434c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad9757),
	.w1(32'hb92c9ef0),
	.w2(32'h392da52e),
	.w3(32'hb97bccfb),
	.w4(32'hb83b5126),
	.w5(32'h391961a6),
	.w6(32'hb9906e72),
	.w7(32'hb71ef66e),
	.w8(32'hb90265a7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853c226),
	.w1(32'h391f6c19),
	.w2(32'hb8f4c9b1),
	.w3(32'h3809e676),
	.w4(32'h39bd5994),
	.w5(32'h3836cbf4),
	.w6(32'h38352368),
	.w7(32'hb97cf52f),
	.w8(32'hb8d32e64),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d4b70c),
	.w1(32'hba0a134c),
	.w2(32'h3a0b03f2),
	.w3(32'h39428acf),
	.w4(32'hb9aedc5c),
	.w5(32'h39d2de6f),
	.w6(32'hba3eb4b4),
	.w7(32'h397ee321),
	.w8(32'hb7d65ba0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39955ad6),
	.w1(32'hba6e7115),
	.w2(32'hba7e797e),
	.w3(32'h38b7688b),
	.w4(32'hba0940ac),
	.w5(32'hba02a271),
	.w6(32'hba4546ab),
	.w7(32'hb98f8de8),
	.w8(32'hb653e876),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18dc20),
	.w1(32'hb9e86f01),
	.w2(32'hba6b353f),
	.w3(32'h38a14780),
	.w4(32'h37eb9908),
	.w5(32'hb9cf04ba),
	.w6(32'hb8400394),
	.w7(32'hba089769),
	.w8(32'hb90123c4),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cec4e9),
	.w1(32'hb9ed7402),
	.w2(32'hb9c71053),
	.w3(32'hb8b6503e),
	.w4(32'hb9984323),
	.w5(32'hb9a665fe),
	.w6(32'hb9ea13cb),
	.w7(32'hb9cbead4),
	.w8(32'hb958e556),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98212fc),
	.w1(32'hb95d80e9),
	.w2(32'hb9f52e32),
	.w3(32'hb989dd5d),
	.w4(32'h36b60de4),
	.w5(32'hb967fffb),
	.w6(32'hb7ff395f),
	.w7(32'hb98df0ac),
	.w8(32'hb8527e98),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969651a),
	.w1(32'hb9cf5940),
	.w2(32'hb9da1a1c),
	.w3(32'hb8852721),
	.w4(32'hb9b0dec4),
	.w5(32'hb9e233a8),
	.w6(32'hb9bfa690),
	.w7(32'hb9dc4f06),
	.w8(32'hb9995956),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf5068),
	.w1(32'h38784746),
	.w2(32'h3950c8eb),
	.w3(32'hb9bf2bf8),
	.w4(32'hb8b750e7),
	.w5(32'h38caaa4e),
	.w6(32'hb8d1d491),
	.w7(32'hb7a409a2),
	.w8(32'hb946a107),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e9ba7b),
	.w1(32'hb9995bd4),
	.w2(32'hba26c399),
	.w3(32'hb8d6033a),
	.w4(32'hb95967b0),
	.w5(32'hb9c4d041),
	.w6(32'hb960adbe),
	.w7(32'hba0ec510),
	.w8(32'hb9a76627),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3015b),
	.w1(32'hb95a6799),
	.w2(32'hb9f4684a),
	.w3(32'hb9791446),
	.w4(32'h37963dc6),
	.w5(32'hb9591dff),
	.w6(32'hb7b77a5b),
	.w7(32'hb98ba732),
	.w8(32'hb812d828),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952776e),
	.w1(32'h38cfb83f),
	.w2(32'h390e8181),
	.w3(32'hb83e4484),
	.w4(32'hb882977d),
	.w5(32'h3655f99e),
	.w6(32'hb75fc8aa),
	.w7(32'hb8ec3d66),
	.w8(32'hb9785bc2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f4cc2),
	.w1(32'hb99fe8a7),
	.w2(32'hb9dfacda),
	.w3(32'hb89199b8),
	.w4(32'hb9327b58),
	.w5(32'hb9ddb042),
	.w6(32'hb98cc5a0),
	.w7(32'hb9b574db),
	.w8(32'hb998a870),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be6ece),
	.w1(32'hba4d9d08),
	.w2(32'hb87c74ae),
	.w3(32'hb929ef16),
	.w4(32'hba593950),
	.w5(32'hba2e76b3),
	.w6(32'hb9d18fa2),
	.w7(32'hb9facfbc),
	.w8(32'hba004a2b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13f9ac),
	.w1(32'hb9340551),
	.w2(32'hb991afaf),
	.w3(32'hba07775f),
	.w4(32'hb7c096b7),
	.w5(32'hb9136d59),
	.w6(32'hb98f804d),
	.w7(32'hb9887a03),
	.w8(32'hb92b3679),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984c1d8),
	.w1(32'h38045c9d),
	.w2(32'h38f941ce),
	.w3(32'hb897c69a),
	.w4(32'h3918c735),
	.w5(32'h387bfa38),
	.w6(32'hb89888bc),
	.w7(32'h38c5695e),
	.w8(32'h38b7bcf5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37842984),
	.w1(32'hba06e23f),
	.w2(32'hb9aa6548),
	.w3(32'hb8900186),
	.w4(32'hba0b2794),
	.w5(32'hb9fc7c16),
	.w6(32'hb9b017de),
	.w7(32'hb9a4d4fd),
	.w8(32'hb93f6e67),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f7526),
	.w1(32'hb99c1907),
	.w2(32'hba31c0f4),
	.w3(32'hb95e6c7a),
	.w4(32'h37aaf6af),
	.w5(32'hb9a23b9b),
	.w6(32'hb7de4d8c),
	.w7(32'hb9c91885),
	.w8(32'hb8721871),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b2376),
	.w1(32'hb9a7bd60),
	.w2(32'hba0111f3),
	.w3(32'hb853d104),
	.w4(32'hb910f60c),
	.w5(32'hb98ffd3b),
	.w6(32'hb947555e),
	.w7(32'hb9c2e17d),
	.w8(32'hb94faad6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a082b4),
	.w1(32'hb9bd49a0),
	.w2(32'hba1240c3),
	.w3(32'hb972eb59),
	.w4(32'hb908063b),
	.w5(32'hb99ce10c),
	.w6(32'hb97d7f07),
	.w7(32'hb9dca5aa),
	.w8(32'hb9693b4d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982e4cd),
	.w1(32'hba57c161),
	.w2(32'hba091847),
	.w3(32'hb93053bb),
	.w4(32'hba391a60),
	.w5(32'hb9c6f8fb),
	.w6(32'hb9ae8a6c),
	.w7(32'hb9edded7),
	.w8(32'hba15c444),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba733c8f),
	.w1(32'hb90a4673),
	.w2(32'hb5de4204),
	.w3(32'hba2b32a7),
	.w4(32'hb922b9f6),
	.w5(32'hb88776e4),
	.w6(32'hb8bc9e57),
	.w7(32'h37cb40c7),
	.w8(32'hb992fdb2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bc7a1),
	.w1(32'hb9de92c3),
	.w2(32'hb9cebf91),
	.w3(32'hb9170a4b),
	.w4(32'hb98b6374),
	.w5(32'hb9e3007c),
	.w6(32'hba1a2579),
	.w7(32'hba14937c),
	.w8(32'hb982108f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9044c5a),
	.w1(32'hb9a3d971),
	.w2(32'hb9b4776a),
	.w3(32'hb9980e55),
	.w4(32'hb916a026),
	.w5(32'hb9b14394),
	.w6(32'hb9edd363),
	.w7(32'hb9fdb8e8),
	.w8(32'hb9922ce2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92dbbcd),
	.w1(32'hb9ce6313),
	.w2(32'hb9fcc1e9),
	.w3(32'hb915f7bd),
	.w4(32'hb947be26),
	.w5(32'hb993fd68),
	.w6(32'hb94fb8f4),
	.w7(32'hb9b3d58f),
	.w8(32'hb955fb70),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a05a46),
	.w1(32'hba526794),
	.w2(32'hba71e1db),
	.w3(32'hb91f1711),
	.w4(32'hba3bdc48),
	.w5(32'hba123e90),
	.w6(32'hb9d45484),
	.w7(32'hba05b3be),
	.w8(32'hba173d8c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a875f),
	.w1(32'h36a037ee),
	.w2(32'hb9740372),
	.w3(32'hb9c72aa3),
	.w4(32'h39b05666),
	.w5(32'h392ffe09),
	.w6(32'hb90ee977),
	.w7(32'hb9e46230),
	.w8(32'hb884e161),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4809b),
	.w1(32'hb99c1990),
	.w2(32'hba1a07a1),
	.w3(32'h39998ef4),
	.w4(32'hb8f58a71),
	.w5(32'hb9bc4b73),
	.w6(32'hb9427c71),
	.w7(32'hb9f812aa),
	.w8(32'hb912ffb4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978a024),
	.w1(32'h396bf4c4),
	.w2(32'h391e1c64),
	.w3(32'hb9401b97),
	.w4(32'h393d6c12),
	.w5(32'h38f3b9e9),
	.w6(32'h39b86757),
	.w7(32'h3920eeff),
	.w8(32'h3885af4b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b922ce),
	.w1(32'h399dcd0b),
	.w2(32'h39c72ad3),
	.w3(32'h39189cea),
	.w4(32'h3977a71b),
	.w5(32'h39717dc3),
	.w6(32'h398c3b12),
	.w7(32'h39a1c8b9),
	.w8(32'h394af5ee),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule