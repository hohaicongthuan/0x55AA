module layer_10_featuremap_232(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012022),
	.w1(32'hbd024675),
	.w2(32'hbbbeea45),
	.w3(32'hbb6fba4d),
	.w4(32'hba6c2643),
	.w5(32'h3b9a16a8),
	.w6(32'h3babc5ab),
	.w7(32'h3adc73b7),
	.w8(32'hbc06f974),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a61fb),
	.w1(32'hbc273f70),
	.w2(32'hbc0f78d8),
	.w3(32'hbcab45c7),
	.w4(32'h3bf37b73),
	.w5(32'hbc169abe),
	.w6(32'hbb72bd0d),
	.w7(32'hbc741f0b),
	.w8(32'h3c0d16b2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82134e),
	.w1(32'hbb260ad6),
	.w2(32'h3cc38aa6),
	.w3(32'hbb858c48),
	.w4(32'h3cba319f),
	.w5(32'h3b9955f6),
	.w6(32'h3b3a93e3),
	.w7(32'hbc8f5c03),
	.w8(32'hbb79a893),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc613b94),
	.w1(32'h3a6157ee),
	.w2(32'hb9e9cb94),
	.w3(32'h3c1e638e),
	.w4(32'h3ab44f86),
	.w5(32'hbbd78878),
	.w6(32'hbb91967a),
	.w7(32'hbc0d45b3),
	.w8(32'h3d137a62),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b24d4),
	.w1(32'hb9187ab8),
	.w2(32'hbbeb0524),
	.w3(32'h3b270792),
	.w4(32'hbbb37eaa),
	.w5(32'hbabdb239),
	.w6(32'hbc499c65),
	.w7(32'h3aae70f1),
	.w8(32'hbbf8bb02),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d0ee5),
	.w1(32'hbc9e207d),
	.w2(32'hbb855489),
	.w3(32'hbc02e725),
	.w4(32'h3b2497b1),
	.w5(32'h3d94569d),
	.w6(32'h3c8ab5ef),
	.w7(32'h3c83c1a2),
	.w8(32'hbcb8ecf4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023cf2),
	.w1(32'hbd7e8bdb),
	.w2(32'hbc6c8080),
	.w3(32'hb79d7214),
	.w4(32'h3c77cbd7),
	.w5(32'hba13379a),
	.w6(32'hbb247045),
	.w7(32'hbccb485a),
	.w8(32'h3bb54a2c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad76d1),
	.w1(32'hbc29b092),
	.w2(32'h3aa6c9e6),
	.w3(32'hba938e4d),
	.w4(32'hba1f6e6c),
	.w5(32'h3bdb7a77),
	.w6(32'h3c889e2d),
	.w7(32'hba60b9e9),
	.w8(32'hb8fe5e21),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ecd38),
	.w1(32'hbcc282b6),
	.w2(32'hbc7b9839),
	.w3(32'hbbea6430),
	.w4(32'hbd52db9d),
	.w5(32'h3b02c523),
	.w6(32'hbbdbe3d7),
	.w7(32'hbb8b64eb),
	.w8(32'hbac9aede),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f258b),
	.w1(32'h397851ed),
	.w2(32'hbc00b03c),
	.w3(32'h3c81d73f),
	.w4(32'h3b7ea613),
	.w5(32'hbc8bb818),
	.w6(32'h3c194fd0),
	.w7(32'h3c31a520),
	.w8(32'h3c81faf9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8aa98),
	.w1(32'hbb8791e8),
	.w2(32'hbb6c1404),
	.w3(32'h3c6bbf42),
	.w4(32'hbba500f0),
	.w5(32'hbb994870),
	.w6(32'h3cf6292b),
	.w7(32'h3c096d3c),
	.w8(32'hbc1f1a82),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf978e),
	.w1(32'h3b96f891),
	.w2(32'h3c25de97),
	.w3(32'h3c092f5b),
	.w4(32'h3ba19083),
	.w5(32'hba057006),
	.w6(32'hba913e08),
	.w7(32'h37c94b95),
	.w8(32'h3c7cd2da),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb2bf),
	.w1(32'h3bd62fd7),
	.w2(32'h3ad597d4),
	.w3(32'hbb5d57d2),
	.w4(32'hbb8c520f),
	.w5(32'h3cc51e56),
	.w6(32'h3c12cd6b),
	.w7(32'h3c34330c),
	.w8(32'h3bdf0369),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bdfd6),
	.w1(32'hbb75e4fd),
	.w2(32'h3b038ef3),
	.w3(32'hbb52d12c),
	.w4(32'h3c181cce),
	.w5(32'h3ba533dc),
	.w6(32'hbbc52143),
	.w7(32'h3bbf4adf),
	.w8(32'hb992746d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00daac),
	.w1(32'hbb2eeb6f),
	.w2(32'hbcc595b4),
	.w3(32'hbc0acbd3),
	.w4(32'hbafb15ca),
	.w5(32'hbc601483),
	.w6(32'hbb8f4371),
	.w7(32'h3cbf6d69),
	.w8(32'h3c1254b7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba91f8f),
	.w1(32'h3c8345dd),
	.w2(32'h3c84429a),
	.w3(32'h3c97b86b),
	.w4(32'h3b8ae581),
	.w5(32'h3b0b1394),
	.w6(32'hbbfeab38),
	.w7(32'hbb65d473),
	.w8(32'hba97145b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae791),
	.w1(32'h3cabc9a1),
	.w2(32'h3ad63e29),
	.w3(32'hbb3c7e50),
	.w4(32'h35e2553f),
	.w5(32'hbc753725),
	.w6(32'hbc29d79e),
	.w7(32'hbbe1a333),
	.w8(32'h3c28fe15),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceaf46a),
	.w1(32'hbc0b4786),
	.w2(32'h3c28243a),
	.w3(32'h3a2c79c6),
	.w4(32'h3c864124),
	.w5(32'h3b43b751),
	.w6(32'h3c195072),
	.w7(32'h3ba32d7a),
	.w8(32'hbc3e52c7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b34c),
	.w1(32'hba9304d3),
	.w2(32'hbc3c7a56),
	.w3(32'h3c8631c4),
	.w4(32'hbacbc8f6),
	.w5(32'h3abd8293),
	.w6(32'h3c86adfc),
	.w7(32'h3bb37b2a),
	.w8(32'hbc0bb035),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a2d4a),
	.w1(32'hbcadaddb),
	.w2(32'hbb9f6b2c),
	.w3(32'hbc1907fe),
	.w4(32'h3c0ea6f0),
	.w5(32'hbb8e433b),
	.w6(32'h3c700354),
	.w7(32'hbc573f1e),
	.w8(32'hb9a75b44),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39810c28),
	.w1(32'h3ba64089),
	.w2(32'hbb94c5eb),
	.w3(32'hbc4e8d26),
	.w4(32'h3ab12154),
	.w5(32'hbc0079a5),
	.w6(32'h3b669fa3),
	.w7(32'hbb1166d0),
	.w8(32'h3b76bfb4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5def96),
	.w1(32'h3c4f5d23),
	.w2(32'h3b7a9bba),
	.w3(32'hba9af351),
	.w4(32'h3a826fe8),
	.w5(32'h3bb9230f),
	.w6(32'hbc381686),
	.w7(32'hb9ee18c4),
	.w8(32'hbb0698b4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc42e),
	.w1(32'hb9c26be4),
	.w2(32'hbc05f7ae),
	.w3(32'h3cb7ddc3),
	.w4(32'h3c16456d),
	.w5(32'h3bbf1b8b),
	.w6(32'h385ebb0c),
	.w7(32'h3c6c0b99),
	.w8(32'h3ba7fca6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc177d04),
	.w1(32'h3c549c6b),
	.w2(32'hbc59a512),
	.w3(32'h3bebd366),
	.w4(32'hbc7b3880),
	.w5(32'h3c1bc06f),
	.w6(32'hbc0cf63b),
	.w7(32'hbc26b26a),
	.w8(32'h3c5a5982),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86e1d3),
	.w1(32'h3a5ff00f),
	.w2(32'hbb305e2b),
	.w3(32'h3cc0095d),
	.w4(32'h3c4d09a7),
	.w5(32'h3c0b279b),
	.w6(32'h3c1e4b44),
	.w7(32'hbb49038a),
	.w8(32'h3bb904a5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a6704),
	.w1(32'hba9d26ee),
	.w2(32'hbc3d52c4),
	.w3(32'hba949aad),
	.w4(32'hbdee7601),
	.w5(32'h3c6a9162),
	.w6(32'hbb1d584a),
	.w7(32'h3a1b3637),
	.w8(32'hbcdb6ca6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf4be05),
	.w1(32'hbc2e0e59),
	.w2(32'hba083af4),
	.w3(32'hbc761228),
	.w4(32'h3b6c4360),
	.w5(32'hbb58bdca),
	.w6(32'h392ae73d),
	.w7(32'hbca08863),
	.w8(32'hbbd54db3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98758e),
	.w1(32'hbbedef1a),
	.w2(32'h3c591653),
	.w3(32'h3c490e5e),
	.w4(32'hbc805b01),
	.w5(32'hbd0d331e),
	.w6(32'hbc1e5f74),
	.w7(32'h3bf8557f),
	.w8(32'hba10ad68),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb462e53),
	.w1(32'h3b9bc800),
	.w2(32'h3cf1c674),
	.w3(32'h3b95a35e),
	.w4(32'hbbd89b55),
	.w5(32'h3c1af2c1),
	.w6(32'hbb8a841f),
	.w7(32'hba641938),
	.w8(32'h3b0cf9df),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eeb449),
	.w1(32'h3ba5034a),
	.w2(32'h3c1136b3),
	.w3(32'hbbb3b052),
	.w4(32'h3bec0c09),
	.w5(32'h3a541832),
	.w6(32'h3ce31cd7),
	.w7(32'hbb04ecd4),
	.w8(32'h3b0b4200),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821606),
	.w1(32'h3c15afb7),
	.w2(32'hbb768a15),
	.w3(32'hba6bb7a1),
	.w4(32'h3c004cb0),
	.w5(32'h3b50a26e),
	.w6(32'hbb332aa4),
	.w7(32'h3aa373ce),
	.w8(32'h3b34f507),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3810bc),
	.w1(32'h3b3afd06),
	.w2(32'hbb14e37b),
	.w3(32'hbcbc4820),
	.w4(32'hbc26fdbe),
	.w5(32'h3c9b4721),
	.w6(32'h3c257b59),
	.w7(32'hbc7d4df0),
	.w8(32'h3c0f1ada),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69bd75),
	.w1(32'hbbf25a7e),
	.w2(32'hbc50fe05),
	.w3(32'h3b3a74ca),
	.w4(32'hbc1b5d88),
	.w5(32'h3bc67f61),
	.w6(32'h3b5d3914),
	.w7(32'hbbcbbc2f),
	.w8(32'hbba2d69d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa53bb6),
	.w1(32'hbcceabcd),
	.w2(32'h3c88d40e),
	.w3(32'hbbe2ee23),
	.w4(32'h3bac5e70),
	.w5(32'h3c7ba56a),
	.w6(32'h3b22ca93),
	.w7(32'hbc8f6f1a),
	.w8(32'h3b65279c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf72a97),
	.w1(32'h3a3aae50),
	.w2(32'h3b70a82f),
	.w3(32'hba1a783b),
	.w4(32'hbaa3d264),
	.w5(32'h3ad529bf),
	.w6(32'h3c87b94b),
	.w7(32'hbd0779ad),
	.w8(32'h3d171060),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc304194),
	.w1(32'h3caf93c9),
	.w2(32'hbc81cf81),
	.w3(32'hb95d8b8b),
	.w4(32'h386fb94c),
	.w5(32'hb9f41176),
	.w6(32'h393a66b5),
	.w7(32'hbb5a24a6),
	.w8(32'h3b07a271),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6662d2),
	.w1(32'hbbbd3516),
	.w2(32'h3ba05cc4),
	.w3(32'h3c097a91),
	.w4(32'hba43a12d),
	.w5(32'hbc0acfd7),
	.w6(32'hba3bcff6),
	.w7(32'h3c12c733),
	.w8(32'h3a92e3e9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff99ab),
	.w1(32'h3a63ae24),
	.w2(32'h3d279526),
	.w3(32'h3a561e25),
	.w4(32'h3a49dfbf),
	.w5(32'hb90b039e),
	.w6(32'h3b0d6bc3),
	.w7(32'h3c3c0c84),
	.w8(32'hbb3cba99),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe727d9),
	.w1(32'h3cb345bb),
	.w2(32'h3c8fd0d0),
	.w3(32'h3c325ecb),
	.w4(32'hbaa0982d),
	.w5(32'h3ba2e649),
	.w6(32'hbbfee5dc),
	.w7(32'hbb8e4f84),
	.w8(32'h39edb65c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5657e5),
	.w1(32'hbc55b441),
	.w2(32'h3b2483c3),
	.w3(32'hb982058b),
	.w4(32'h3c01e910),
	.w5(32'h3ba0ab98),
	.w6(32'hbb9f95d0),
	.w7(32'h3bb3cd68),
	.w8(32'h3c47002e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53890d3),
	.w1(32'h3c819a27),
	.w2(32'hbb8ede67),
	.w3(32'hbbbaa6a2),
	.w4(32'hbb05dcdf),
	.w5(32'hbc3f8665),
	.w6(32'hba9d7816),
	.w7(32'h3ae74901),
	.w8(32'h38f86b84),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2a98e),
	.w1(32'h3a23d405),
	.w2(32'h3ba9ed80),
	.w3(32'hb9c865e5),
	.w4(32'h3c822d57),
	.w5(32'hbb2f12ee),
	.w6(32'h3c99f118),
	.w7(32'hbc6e72ba),
	.w8(32'hbc124216),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1a3ef),
	.w1(32'h3ae960a5),
	.w2(32'hbc2fbc3a),
	.w3(32'hbc86beb3),
	.w4(32'hbba18863),
	.w5(32'h3bd0a7aa),
	.w6(32'h3b880a80),
	.w7(32'hbc4811f5),
	.w8(32'h3c01bcbd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c8b34),
	.w1(32'h3af03ff1),
	.w2(32'h39d8b106),
	.w3(32'h3b0484d5),
	.w4(32'hbbf5765b),
	.w5(32'h3a295d55),
	.w6(32'h37a9a758),
	.w7(32'h3c396bbf),
	.w8(32'h3b8c707b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2de65),
	.w1(32'h3cedae8e),
	.w2(32'hbc0f8240),
	.w3(32'h3b0cfbbb),
	.w4(32'h3b96102a),
	.w5(32'h3c6c66e2),
	.w6(32'hbb0285f5),
	.w7(32'h3bc64b46),
	.w8(32'hb63f3731),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3349),
	.w1(32'hbc11fe51),
	.w2(32'h3d07d659),
	.w3(32'hbb3926e7),
	.w4(32'hbc04d814),
	.w5(32'hbaf158a8),
	.w6(32'hbb8e49cb),
	.w7(32'hbb88c5ee),
	.w8(32'h3c01dc5b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a6eb6),
	.w1(32'hb99de273),
	.w2(32'hbb9b9231),
	.w3(32'hbc0160b4),
	.w4(32'hbc041476),
	.w5(32'h3b6b799c),
	.w6(32'hb9130963),
	.w7(32'h3c9a0861),
	.w8(32'hbb1faa16),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf308),
	.w1(32'h3b0965a7),
	.w2(32'hbb4d6263),
	.w3(32'hbc88c62a),
	.w4(32'h3b990de5),
	.w5(32'hbb6a01bf),
	.w6(32'hbccc2e7f),
	.w7(32'hbaf39dc5),
	.w8(32'h3c8fa5fa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaca16),
	.w1(32'hbabb0bda),
	.w2(32'h3bec5bb8),
	.w3(32'hbb8f3b29),
	.w4(32'hbbe8dbc7),
	.w5(32'hbbe215f7),
	.w6(32'hbbb7d68d),
	.w7(32'hbc8a8aca),
	.w8(32'hbaa8f642),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb3e75),
	.w1(32'h3abcc593),
	.w2(32'h3be9b9da),
	.w3(32'h3c4df083),
	.w4(32'h3c26547d),
	.w5(32'hbbbd41ca),
	.w6(32'hbbe6e20e),
	.w7(32'h3aa3e310),
	.w8(32'h3ba718b9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9432313),
	.w1(32'h39e872f9),
	.w2(32'h3b0fd1d0),
	.w3(32'hb9e37904),
	.w4(32'h3a8bca33),
	.w5(32'h39ab7bd7),
	.w6(32'hb8e5cd93),
	.w7(32'hbba82916),
	.w8(32'hbb83e670),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14090c),
	.w1(32'h3b82d5aa),
	.w2(32'h3b3ecbef),
	.w3(32'hbc880c5d),
	.w4(32'h3c4951bc),
	.w5(32'h3c86c58b),
	.w6(32'h3b438848),
	.w7(32'h3b07052d),
	.w8(32'hbba15e53),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf3934),
	.w1(32'h3b5e373d),
	.w2(32'hbb2a03d4),
	.w3(32'hbc1adfe5),
	.w4(32'hbbc9c3ae),
	.w5(32'hbb36e552),
	.w6(32'hbbf388d1),
	.w7(32'h3bc23335),
	.w8(32'hbb78b3b3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bcabb),
	.w1(32'h3cc18675),
	.w2(32'hbbaa639c),
	.w3(32'hbb9d2767),
	.w4(32'h3a43901d),
	.w5(32'hbab4c981),
	.w6(32'h3c853919),
	.w7(32'h3c012b55),
	.w8(32'hbc6efc13),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca626),
	.w1(32'h3b2cee2b),
	.w2(32'h3aaf19d0),
	.w3(32'h3cb7e47f),
	.w4(32'h38b99055),
	.w5(32'h3ba955f4),
	.w6(32'h3c1956c2),
	.w7(32'hbacde3ec),
	.w8(32'h3be52900),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1515d5),
	.w1(32'h3b91389c),
	.w2(32'h3b134f42),
	.w3(32'h3c10b037),
	.w4(32'hbc8e0ee4),
	.w5(32'hbbfd1682),
	.w6(32'h3aff1cdb),
	.w7(32'h3ba6d34d),
	.w8(32'h3c0006b5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44116d),
	.w1(32'h39d5036b),
	.w2(32'h3aeda555),
	.w3(32'hbb379dbe),
	.w4(32'hbc6de4d8),
	.w5(32'h3bfd38d4),
	.w6(32'hbb0f883b),
	.w7(32'h3b982661),
	.w8(32'hbc1fd938),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf399fd),
	.w1(32'h39402729),
	.w2(32'hbcf81069),
	.w3(32'h3b65bfdf),
	.w4(32'h3bafb18c),
	.w5(32'h3b225967),
	.w6(32'h39fc02c7),
	.w7(32'h3b514176),
	.w8(32'hbba1b82a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8429f0),
	.w1(32'h3c96c188),
	.w2(32'hbc02ea71),
	.w3(32'hb99e71e7),
	.w4(32'hbc59f655),
	.w5(32'hbc84dc6b),
	.w6(32'hbc0db4df),
	.w7(32'hbb8211c8),
	.w8(32'hbb392fe1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b011670),
	.w1(32'h3c67c09f),
	.w2(32'hbae065d7),
	.w3(32'hbb29551a),
	.w4(32'h3ad357c3),
	.w5(32'h3c062480),
	.w6(32'hbaf917e6),
	.w7(32'hbbb987cf),
	.w8(32'h3ca6775a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324967),
	.w1(32'hba604336),
	.w2(32'h3ccde923),
	.w3(32'h3c23c1ef),
	.w4(32'hbbf96a63),
	.w5(32'h3c3c78d4),
	.w6(32'hbc086743),
	.w7(32'hbc0359da),
	.w8(32'hbc7a08cc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39198),
	.w1(32'hbbd6d31c),
	.w2(32'hba7572af),
	.w3(32'h3ade406f),
	.w4(32'h3c312f34),
	.w5(32'hbc722b5a),
	.w6(32'hb9ebbd19),
	.w7(32'h3b433cf1),
	.w8(32'h3b6b3c61),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f990f),
	.w1(32'h3adc9d63),
	.w2(32'hbcce6e95),
	.w3(32'hbbb8bd3f),
	.w4(32'h3c8385fd),
	.w5(32'hbc00e344),
	.w6(32'hbc3952fb),
	.w7(32'hbae8a77f),
	.w8(32'hbb8425e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95cfb15),
	.w1(32'hbc82e518),
	.w2(32'h3b89c1d3),
	.w3(32'h3c778cdb),
	.w4(32'h3c0f2b3e),
	.w5(32'hbc1303be),
	.w6(32'h3b927d32),
	.w7(32'h3a36435a),
	.w8(32'h3c4b97b3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f9aa1),
	.w1(32'hbb8999d8),
	.w2(32'hbc472591),
	.w3(32'hbc3d5dc1),
	.w4(32'hbc8c7d2c),
	.w5(32'hbc38e548),
	.w6(32'h3c851346),
	.w7(32'hbb8c9499),
	.w8(32'hbc22f90d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c509776),
	.w1(32'hba2f22f4),
	.w2(32'h3c1bcf27),
	.w3(32'hbc20b186),
	.w4(32'h3bf5d914),
	.w5(32'hba92b618),
	.w6(32'h3c4bb17a),
	.w7(32'hbc749d14),
	.w8(32'hbc7bddac),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ae61d),
	.w1(32'hbc0e3529),
	.w2(32'hbb18a493),
	.w3(32'hbc1d4151),
	.w4(32'h3b9485f8),
	.w5(32'h3ce60b1c),
	.w6(32'h39b47060),
	.w7(32'hbc559e84),
	.w8(32'h3bb51d96),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8d11e),
	.w1(32'hbc450da3),
	.w2(32'hbb9fd1f9),
	.w3(32'h3ad35864),
	.w4(32'hbb172ca4),
	.w5(32'h3c3378a7),
	.w6(32'hba7ead66),
	.w7(32'h3bae803c),
	.w8(32'hbbb0471b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5f6d2),
	.w1(32'h3bc41c6f),
	.w2(32'hb9e608ce),
	.w3(32'h3b96d040),
	.w4(32'h38843a1e),
	.w5(32'hbd139409),
	.w6(32'hbbab99e1),
	.w7(32'hbb8d7ac9),
	.w8(32'hbb24e171),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7df3),
	.w1(32'hba9a4848),
	.w2(32'h3bfe8240),
	.w3(32'hbc53fb79),
	.w4(32'hbbbb4f8d),
	.w5(32'h3b677596),
	.w6(32'h3acd1df6),
	.w7(32'hbbd67a8c),
	.w8(32'h39a6b7cd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4cb35),
	.w1(32'hbc0a147c),
	.w2(32'hbbe6cf0a),
	.w3(32'hbc1af0fd),
	.w4(32'hbab214b4),
	.w5(32'h3b605368),
	.w6(32'h3c0139d9),
	.w7(32'hbcd127a7),
	.w8(32'hbccbd52f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005b27),
	.w1(32'hbbaa7285),
	.w2(32'h3b90f1da),
	.w3(32'h3d7589d7),
	.w4(32'h3c586e90),
	.w5(32'h3b9e8256),
	.w6(32'hbc6620cc),
	.w7(32'h3c88bdc5),
	.w8(32'hbbd7485c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52c2b7),
	.w1(32'h3b15039b),
	.w2(32'h3aa04265),
	.w3(32'hbb044c29),
	.w4(32'hbb8c3910),
	.w5(32'hba9edca4),
	.w6(32'h3b84de0d),
	.w7(32'h3bd25587),
	.w8(32'hb9c5eebe),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bdd08),
	.w1(32'h37742e1e),
	.w2(32'hbc8256cb),
	.w3(32'h3b8d142c),
	.w4(32'h3c374598),
	.w5(32'hbc4d0dcd),
	.w6(32'h3c5a02f3),
	.w7(32'hbb1e96a0),
	.w8(32'h3bacb87d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3c127),
	.w1(32'h3b9fc85d),
	.w2(32'h3adfd834),
	.w3(32'hbc2e966e),
	.w4(32'hb9fd2b54),
	.w5(32'h3b48220c),
	.w6(32'hbaec2db3),
	.w7(32'hbcaa2470),
	.w8(32'h3c442752),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e86db),
	.w1(32'hbc4191e8),
	.w2(32'hbbf48cdc),
	.w3(32'h3c1d6aab),
	.w4(32'h3b93d9d4),
	.w5(32'hbc59b29c),
	.w6(32'hbb96b306),
	.w7(32'hbc46a13c),
	.w8(32'hbbbb76b9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51f928),
	.w1(32'h3b521828),
	.w2(32'hbb95bf93),
	.w3(32'h3c7bba7c),
	.w4(32'h3b0c8c21),
	.w5(32'h3a29c5bf),
	.w6(32'h3bd28aa8),
	.w7(32'hbbab3ed6),
	.w8(32'h3b19bd82),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e110),
	.w1(32'h3cae5f5b),
	.w2(32'hbaa58614),
	.w3(32'hbbb4dc48),
	.w4(32'hbba49434),
	.w5(32'hbbbdd7a4),
	.w6(32'h39bf1c26),
	.w7(32'hbcbb34d6),
	.w8(32'h3c07b70e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87fee16),
	.w1(32'h3c6f9568),
	.w2(32'h3aeb8696),
	.w3(32'hbc9d5b45),
	.w4(32'hba0d7762),
	.w5(32'h3c94502a),
	.w6(32'h3af2f2d3),
	.w7(32'h3ad96fba),
	.w8(32'h3ca54738),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9f150),
	.w1(32'hba216881),
	.w2(32'h39c5d400),
	.w3(32'h3b73951f),
	.w4(32'h3b2f1ebd),
	.w5(32'hbb289f4d),
	.w6(32'h3a435d7e),
	.w7(32'hbc13a408),
	.w8(32'hbc193518),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba24e96),
	.w1(32'h3b9c050b),
	.w2(32'hbb2b3603),
	.w3(32'hbae7c70f),
	.w4(32'hbc3c42a8),
	.w5(32'h3b9a628a),
	.w6(32'hbb117244),
	.w7(32'hbc5b50bd),
	.w8(32'h3bc86e8b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9efa4),
	.w1(32'h398fa649),
	.w2(32'hba03a5c3),
	.w3(32'h3b39a4ac),
	.w4(32'hbbfddd6b),
	.w5(32'hbcab25b9),
	.w6(32'h3887c9fe),
	.w7(32'hbaf978f7),
	.w8(32'hbbaebdc4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20d1ed),
	.w1(32'h3c8cca91),
	.w2(32'hbbff61ba),
	.w3(32'hbb04cd73),
	.w4(32'h3b9e7038),
	.w5(32'hba7ee394),
	.w6(32'h3c619fc5),
	.w7(32'hbb00ff21),
	.w8(32'h3cc570a9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c7a9f),
	.w1(32'hb7c8de7b),
	.w2(32'h39395282),
	.w3(32'h3bb69cd2),
	.w4(32'hbb3dd555),
	.w5(32'hbbe080f4),
	.w6(32'hbc50fe9b),
	.w7(32'hbaf57bfd),
	.w8(32'hb9a2984f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f37b),
	.w1(32'hbaf45718),
	.w2(32'h3b8d8041),
	.w3(32'hba44d56d),
	.w4(32'hbc2410f7),
	.w5(32'hbb10bd25),
	.w6(32'hbba40c1b),
	.w7(32'h3c3094bb),
	.w8(32'hbbbd0343),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b9028),
	.w1(32'h3aa58e3f),
	.w2(32'hbc24d66d),
	.w3(32'h3c1cba98),
	.w4(32'hb9f07095),
	.w5(32'h3be0039e),
	.w6(32'h3c4ecfff),
	.w7(32'hbc159879),
	.w8(32'h3a1b013f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a91c),
	.w1(32'hbc69f225),
	.w2(32'hbc1c394a),
	.w3(32'h3c505807),
	.w4(32'h3bc13158),
	.w5(32'h3c58d90c),
	.w6(32'h398c7a3a),
	.w7(32'hbbee6992),
	.w8(32'hbc41a83f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88c005),
	.w1(32'hbafadd1b),
	.w2(32'h3b547375),
	.w3(32'h3af46a33),
	.w4(32'hbb10eb96),
	.w5(32'hba946b1c),
	.w6(32'h3c060f4d),
	.w7(32'hba8ed1aa),
	.w8(32'h3af6ab82),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65fb81),
	.w1(32'hba6ba1a5),
	.w2(32'h3bf638f4),
	.w3(32'hbbce9aa8),
	.w4(32'hbacd33cd),
	.w5(32'h3bd694f4),
	.w6(32'h3beacb20),
	.w7(32'h3a8060b2),
	.w8(32'h3bc05bb7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba277fb0),
	.w1(32'hbbaa7eea),
	.w2(32'h3be35e85),
	.w3(32'h3ab9c853),
	.w4(32'hbb0ec2a0),
	.w5(32'h3a76b360),
	.w6(32'hbc4a8a74),
	.w7(32'h3b9f195c),
	.w8(32'hbb1a5aca),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c646aaa),
	.w1(32'h3ba0e321),
	.w2(32'hbc2821af),
	.w3(32'h3a5f4f21),
	.w4(32'hb94f9c40),
	.w5(32'hbb33dad6),
	.w6(32'h3b9cd7b1),
	.w7(32'hbaf279cc),
	.w8(32'hbbc4cf03),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8192e),
	.w1(32'hbb215343),
	.w2(32'h3c862c63),
	.w3(32'hb9d7e0af),
	.w4(32'h3c98a2e2),
	.w5(32'hb8ba83db),
	.w6(32'h3c06bc8a),
	.w7(32'hbb086a78),
	.w8(32'hb983b2f5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18696e),
	.w1(32'hbc0437cb),
	.w2(32'h3c02eb37),
	.w3(32'h3bddc6b5),
	.w4(32'hbb381f70),
	.w5(32'hbc01df27),
	.w6(32'h3b870adc),
	.w7(32'hbbc0dad2),
	.w8(32'hba556956),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00b5b6),
	.w1(32'h3b9b39df),
	.w2(32'h3c1ab876),
	.w3(32'h3b842347),
	.w4(32'hb9055ba5),
	.w5(32'hbc30fe3d),
	.w6(32'h3b6150e3),
	.w7(32'hbc18bbea),
	.w8(32'h3bd608ed),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e25f),
	.w1(32'h3ae8ff45),
	.w2(32'hb8929656),
	.w3(32'hbafa793c),
	.w4(32'h3b071ff1),
	.w5(32'hba9cd0d0),
	.w6(32'h39109de7),
	.w7(32'hbbeaa041),
	.w8(32'h3a9af658),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a8654),
	.w1(32'h3bb459e9),
	.w2(32'hbba69503),
	.w3(32'h3b455d72),
	.w4(32'h3d231b89),
	.w5(32'hbc31b55c),
	.w6(32'h3abd776c),
	.w7(32'hbb07bb24),
	.w8(32'hbab048e8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bf8ee),
	.w1(32'hbb9740f2),
	.w2(32'h3b230c64),
	.w3(32'hbb51a61f),
	.w4(32'h3c062634),
	.w5(32'hbc2ac383),
	.w6(32'h3a75da41),
	.w7(32'hbad02a66),
	.w8(32'h350058c8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f4d7c),
	.w1(32'hbc867cbe),
	.w2(32'h3a3f48fc),
	.w3(32'hba3d3777),
	.w4(32'h3a93a6f9),
	.w5(32'h3b85f016),
	.w6(32'hbc830d74),
	.w7(32'h3b858e92),
	.w8(32'h3ae3f9cf),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c206632),
	.w1(32'hbb69a31f),
	.w2(32'h39c1de9b),
	.w3(32'hbaa7b884),
	.w4(32'h3b762755),
	.w5(32'hbc24851e),
	.w6(32'h3baab7c3),
	.w7(32'hba65f234),
	.w8(32'hbbb68194),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f613),
	.w1(32'hbc2c8a5b),
	.w2(32'hbc036d82),
	.w3(32'h3b0c8bda),
	.w4(32'hbaf21d2b),
	.w5(32'h3b594570),
	.w6(32'h3ad16c0a),
	.w7(32'h3bb0d9c5),
	.w8(32'h3c8a219a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cddbc),
	.w1(32'h3b837427),
	.w2(32'h3b3e7c66),
	.w3(32'h3b0324dc),
	.w4(32'h3c46e47e),
	.w5(32'h3a9cdb82),
	.w6(32'h38face36),
	.w7(32'h3a5b7982),
	.w8(32'hbbc4d847),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3af03d),
	.w1(32'h3c55f6dc),
	.w2(32'h3bae5199),
	.w3(32'h3998915a),
	.w4(32'h3c3bdd41),
	.w5(32'hb7549573),
	.w6(32'hbb5ef8e5),
	.w7(32'hbae58ba5),
	.w8(32'h3b5f9606),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8167e35),
	.w1(32'hbbd15bdf),
	.w2(32'hbc526323),
	.w3(32'hbbbf1776),
	.w4(32'hbbac1b55),
	.w5(32'h3b67bfad),
	.w6(32'h3bbea02c),
	.w7(32'h3b9d4b86),
	.w8(32'hba98d533),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc13992),
	.w1(32'hbb0f25cc),
	.w2(32'hbc15e22f),
	.w3(32'h39b2b084),
	.w4(32'h3ac319d0),
	.w5(32'h3b829c94),
	.w6(32'h3b9ea91a),
	.w7(32'h3c163c35),
	.w8(32'hbc8c8f70),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c175f04),
	.w1(32'hbc3d36bd),
	.w2(32'h3c011535),
	.w3(32'hbb176189),
	.w4(32'h3b183100),
	.w5(32'hbb779960),
	.w6(32'hbb7d808d),
	.w7(32'h3c06b257),
	.w8(32'h3c77be1a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ff96),
	.w1(32'h3b974fd3),
	.w2(32'h3ac846ff),
	.w3(32'hb8bf4078),
	.w4(32'hbc5571bf),
	.w5(32'h3b625a1d),
	.w6(32'hbbf7d102),
	.w7(32'hb9b983cb),
	.w8(32'hbb0c233d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8859c2),
	.w1(32'hbc3b5f78),
	.w2(32'h3ba0ce39),
	.w3(32'hbc155e2b),
	.w4(32'h3b174dd2),
	.w5(32'h3b5cae47),
	.w6(32'h3abcbf48),
	.w7(32'hbba595c6),
	.w8(32'h3921d4b6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e1f1),
	.w1(32'h3bfea707),
	.w2(32'hb8253ef6),
	.w3(32'hbb391277),
	.w4(32'hba781c48),
	.w5(32'h3bc56366),
	.w6(32'hbba44a91),
	.w7(32'h3b0f4ee7),
	.w8(32'h3a2182b9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba88409),
	.w1(32'hbb98a200),
	.w2(32'hbabcc073),
	.w3(32'hbb4cf4bc),
	.w4(32'h3beeebca),
	.w5(32'h3c0fa4f5),
	.w6(32'hbbc37d33),
	.w7(32'h3bf5561a),
	.w8(32'hbba35547),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc842f00),
	.w1(32'h3bb07780),
	.w2(32'hbb87a8c2),
	.w3(32'h3c10da91),
	.w4(32'h3b484128),
	.w5(32'hbb1e9f44),
	.w6(32'hba0ec7f9),
	.w7(32'hbc2c8015),
	.w8(32'h3b2f8e80),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93d25b),
	.w1(32'hbc4cb51c),
	.w2(32'hbc0dfd67),
	.w3(32'hba3ae04f),
	.w4(32'hbbb7d7e7),
	.w5(32'hbc93c32f),
	.w6(32'hbc914568),
	.w7(32'hbb0c989d),
	.w8(32'h3a4d87f4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f5f74),
	.w1(32'hba702f63),
	.w2(32'h3af8bc5d),
	.w3(32'h3b31e30d),
	.w4(32'hbb94dbc4),
	.w5(32'hbc226b80),
	.w6(32'h3b17476e),
	.w7(32'h3bed6703),
	.w8(32'h3c337658),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31a976),
	.w1(32'h3c4d2396),
	.w2(32'h3bdf9aa1),
	.w3(32'hbb5e165a),
	.w4(32'hbb825eb6),
	.w5(32'hbb8cb7ba),
	.w6(32'hbb593fe7),
	.w7(32'h3ac526ea),
	.w8(32'hbbab9a5d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2abf),
	.w1(32'h3bd6df02),
	.w2(32'hbaf9d98f),
	.w3(32'h3a32be01),
	.w4(32'h3a1a45f2),
	.w5(32'h3b319f7c),
	.w6(32'h39a864d7),
	.w7(32'hbb9cc39f),
	.w8(32'h3a57d799),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32c6f9),
	.w1(32'h3bdf3558),
	.w2(32'hbbcfcdf5),
	.w3(32'hbb3dbb6c),
	.w4(32'hbb83046a),
	.w5(32'h3b0be4c5),
	.w6(32'h3c3c0110),
	.w7(32'hbb1bf5fd),
	.w8(32'hbbf27a22),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f7cf7),
	.w1(32'h3b9c41af),
	.w2(32'hbc279013),
	.w3(32'hbab361fc),
	.w4(32'hbba81ebb),
	.w5(32'h3c3a97e5),
	.w6(32'h3bd5abb3),
	.w7(32'h3be31511),
	.w8(32'hbb33ac92),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b740b57),
	.w1(32'hb9a362a0),
	.w2(32'h3b77279c),
	.w3(32'h3c2a908d),
	.w4(32'h3b8a25cc),
	.w5(32'hbaaf236e),
	.w6(32'h3ac3eeff),
	.w7(32'h3c1129ef),
	.w8(32'h3b9d1f0b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81f99),
	.w1(32'hbad445ca),
	.w2(32'h39814c99),
	.w3(32'hbb97f02a),
	.w4(32'h3a174123),
	.w5(32'hbc2b9fb8),
	.w6(32'hbc27883a),
	.w7(32'h3d010757),
	.w8(32'h3bb7e1ad),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a2125),
	.w1(32'hbaa05966),
	.w2(32'h3c2fba79),
	.w3(32'h3c5e7466),
	.w4(32'h3bdd9531),
	.w5(32'hbb7101b6),
	.w6(32'hb9b17c2c),
	.w7(32'hb8900a40),
	.w8(32'hbb1e2bdd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3f520),
	.w1(32'hb9c69e20),
	.w2(32'hbc0bdc7e),
	.w3(32'hbb3f5439),
	.w4(32'hba294f6f),
	.w5(32'hba91c947),
	.w6(32'h3b310d7c),
	.w7(32'h3cda6887),
	.w8(32'hbbad51d9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03bb4),
	.w1(32'hbc0bea99),
	.w2(32'hbb8cd2ab),
	.w3(32'hbc9ffdfa),
	.w4(32'hba9481fe),
	.w5(32'hba9a7294),
	.w6(32'h3c0f26e3),
	.w7(32'hbc26fed3),
	.w8(32'h3b9f8f8e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb083d44),
	.w1(32'h3bb7cc24),
	.w2(32'hba73cc6d),
	.w3(32'hbb6c4b86),
	.w4(32'hbb0a8140),
	.w5(32'hbc42e985),
	.w6(32'hbb97cdfb),
	.w7(32'hba3e051d),
	.w8(32'hbbd4d316),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393becff),
	.w1(32'hbb9064de),
	.w2(32'hba5d748c),
	.w3(32'h38509620),
	.w4(32'h39f5f110),
	.w5(32'h3b45bf5e),
	.w6(32'hbc871ffb),
	.w7(32'h3b0f1d78),
	.w8(32'h3b1b1aff),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe982c0),
	.w1(32'hbc0b109c),
	.w2(32'h3b6273b9),
	.w3(32'h390c04f0),
	.w4(32'h3c8340cf),
	.w5(32'hbc0b1f49),
	.w6(32'hbb3d5e03),
	.w7(32'h3bf8cc9e),
	.w8(32'h3a7fb8d0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d2405),
	.w1(32'hbc0fd621),
	.w2(32'hbc8cb262),
	.w3(32'hbc0875bb),
	.w4(32'h3b369dac),
	.w5(32'h3b5ecfa1),
	.w6(32'h3b367049),
	.w7(32'h3a9d2929),
	.w8(32'h3b00caf4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3edd0f),
	.w1(32'hb2f6f205),
	.w2(32'hbbb52907),
	.w3(32'hba323966),
	.w4(32'hbb7b933b),
	.w5(32'hbc61222d),
	.w6(32'h3b989f96),
	.w7(32'hba56f931),
	.w8(32'h3b5f3ee7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6a331),
	.w1(32'hb8615953),
	.w2(32'hbbd5bcdc),
	.w3(32'hba3c0ac5),
	.w4(32'hbc05159e),
	.w5(32'h3bbc525b),
	.w6(32'hbae0ba11),
	.w7(32'h3c71b185),
	.w8(32'hbb89eccb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8281aa),
	.w1(32'h3b7bb332),
	.w2(32'h3c2ad6c4),
	.w3(32'h3bfc8870),
	.w4(32'h3c3bdc30),
	.w5(32'hbb0e079a),
	.w6(32'hbc1f0380),
	.w7(32'h3c99feaf),
	.w8(32'hbbb25856),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b166),
	.w1(32'hba8ef205),
	.w2(32'h3b49128d),
	.w3(32'h3bb70c3a),
	.w4(32'hbbc7dd7e),
	.w5(32'hbc803a0a),
	.w6(32'hbb1575a2),
	.w7(32'hbb24fa01),
	.w8(32'h3b3b5c13),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc308573),
	.w1(32'hbb9a5afa),
	.w2(32'hbaa56e06),
	.w3(32'hbb487cf6),
	.w4(32'hbaebd929),
	.w5(32'hbc4fc96f),
	.w6(32'h3b7099c3),
	.w7(32'h3b18012a),
	.w8(32'hbbaa15b6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf7a54),
	.w1(32'h3b4f7371),
	.w2(32'hbb26bde2),
	.w3(32'h3c0c400c),
	.w4(32'hbc249580),
	.w5(32'h3c8713c1),
	.w6(32'h373c9151),
	.w7(32'h3b1b14f8),
	.w8(32'h3b3ba37f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc220c8a),
	.w1(32'hbbbd9219),
	.w2(32'hbbcbd8ea),
	.w3(32'h3c069633),
	.w4(32'h3afe199f),
	.w5(32'hb85499ae),
	.w6(32'h3aa4303c),
	.w7(32'h38e54b2c),
	.w8(32'h3c584ce6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff670b),
	.w1(32'h3c971b2b),
	.w2(32'h3be209bd),
	.w3(32'h3ad3837b),
	.w4(32'hb9f10efb),
	.w5(32'hbaba9c98),
	.w6(32'h3b2338d5),
	.w7(32'hbc3b1009),
	.w8(32'hb9de74ce),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8c59),
	.w1(32'hbbd3b2d7),
	.w2(32'h3c7c5d5f),
	.w3(32'h3bd447bc),
	.w4(32'h3a0c04c4),
	.w5(32'h3ac9ed7b),
	.w6(32'h391606a3),
	.w7(32'h3b995da5),
	.w8(32'hbafc574f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07aa6),
	.w1(32'h3af0c408),
	.w2(32'h3bfea8d4),
	.w3(32'hbbd0b28f),
	.w4(32'hbbb760b7),
	.w5(32'hbc7433f4),
	.w6(32'hba9bf0a6),
	.w7(32'h3bd8535d),
	.w8(32'hb95e94d4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0ecc),
	.w1(32'hb8ee90bf),
	.w2(32'hbbf21fd8),
	.w3(32'h3c5c2d8f),
	.w4(32'hba7901fe),
	.w5(32'h3b08aead),
	.w6(32'hba840c54),
	.w7(32'hb998feb1),
	.w8(32'h3a04ea8d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad06692),
	.w1(32'hbbd5d9dd),
	.w2(32'h3c614a51),
	.w3(32'hb9663c92),
	.w4(32'h3a81d1ec),
	.w5(32'hbafebd0a),
	.w6(32'hbae81944),
	.w7(32'h3bd4fdbe),
	.w8(32'hbc36d03b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d428),
	.w1(32'hba8b6848),
	.w2(32'hbafe8c94),
	.w3(32'hba0df4f7),
	.w4(32'h3b73ec86),
	.w5(32'hbbdebf4d),
	.w6(32'hbbe963c5),
	.w7(32'hbb048c65),
	.w8(32'h3b7fdb02),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba29bf4),
	.w1(32'hbba58d9b),
	.w2(32'hbc0af3a2),
	.w3(32'h3d0f807b),
	.w4(32'h3c1ea61f),
	.w5(32'h3b331c86),
	.w6(32'hbc2902eb),
	.w7(32'hb9dafd98),
	.w8(32'h3acd4d55),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9687b9e),
	.w1(32'hbb4c0d50),
	.w2(32'h3c15f75d),
	.w3(32'h39b62163),
	.w4(32'hbbfecee3),
	.w5(32'hbbb04d19),
	.w6(32'hbbf0ac14),
	.w7(32'h3c28fbd6),
	.w8(32'hbb8134c9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda5427),
	.w1(32'hba416ae1),
	.w2(32'h3a8274ad),
	.w3(32'hbb987bdb),
	.w4(32'hba816297),
	.w5(32'hbba8d01f),
	.w6(32'hbbad290b),
	.w7(32'hbaa1cbc8),
	.w8(32'h3ae811de),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8a38e),
	.w1(32'h38af120a),
	.w2(32'h3cab30dd),
	.w3(32'h3b74b810),
	.w4(32'hbc906943),
	.w5(32'hbb1d6a3c),
	.w6(32'h3c57aaa0),
	.w7(32'hbbd8f796),
	.w8(32'h3b099144),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8698b4),
	.w1(32'hb9e899e9),
	.w2(32'hbc0e7f71),
	.w3(32'h3b882b63),
	.w4(32'hba0dd1a5),
	.w5(32'hbbbdd3c8),
	.w6(32'hba4a575e),
	.w7(32'hbac5a3bb),
	.w8(32'h3b1dc993),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab664b),
	.w1(32'hbc189be5),
	.w2(32'hbb0bafd5),
	.w3(32'h3a874db6),
	.w4(32'hba33dbb8),
	.w5(32'hb94e183c),
	.w6(32'hbb16d1fd),
	.w7(32'hbb6b86f5),
	.w8(32'h3a84eac1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103a46),
	.w1(32'hbb1ac116),
	.w2(32'h3b04446c),
	.w3(32'h3bc09e71),
	.w4(32'h3c13315e),
	.w5(32'h3c0f7ba3),
	.w6(32'hbc86f290),
	.w7(32'hbba9603d),
	.w8(32'hbc39fec8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fa9b6),
	.w1(32'hbc205f00),
	.w2(32'h3bc91265),
	.w3(32'hbbf2bd4a),
	.w4(32'hbc0d5963),
	.w5(32'h3ab0c41e),
	.w6(32'h3b12e908),
	.w7(32'hbbe0b306),
	.w8(32'hbaec753b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50afa9),
	.w1(32'h3b7b6dca),
	.w2(32'hb984c9c2),
	.w3(32'h3a158301),
	.w4(32'hbc5200ff),
	.w5(32'h39dfbf47),
	.w6(32'h3cb3a735),
	.w7(32'h3aa08063),
	.w8(32'hbbb387e4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e43c),
	.w1(32'hbb8be804),
	.w2(32'h3a671351),
	.w3(32'h3bf04398),
	.w4(32'h3c0d8f4e),
	.w5(32'hbbdf0255),
	.w6(32'hbc18bb13),
	.w7(32'hbbad565f),
	.w8(32'h3b7d0495),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e1fdb),
	.w1(32'h3b8d1a83),
	.w2(32'h3bb504dd),
	.w3(32'hbb943bf5),
	.w4(32'h3bebcfa5),
	.w5(32'h3b59a8fe),
	.w6(32'hba62f520),
	.w7(32'hbc907cbd),
	.w8(32'h3bcf0aa6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59db0d),
	.w1(32'h3be92191),
	.w2(32'h3b69c125),
	.w3(32'hbb7a7a24),
	.w4(32'h3a9322ab),
	.w5(32'hbbd85575),
	.w6(32'h3c07308c),
	.w7(32'hbb66e596),
	.w8(32'h3b82fe7c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3bb19),
	.w1(32'hbb98555c),
	.w2(32'hbc6e2ab8),
	.w3(32'h3b034a5e),
	.w4(32'hbbd56551),
	.w5(32'hbafa8673),
	.w6(32'hbb764fff),
	.w7(32'h3b5ff407),
	.w8(32'hbc0501c1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dece3),
	.w1(32'hbbdfe9f8),
	.w2(32'h3c465ae8),
	.w3(32'hba1f4fb5),
	.w4(32'hbc005a35),
	.w5(32'hbb70385d),
	.w6(32'h3b2f6bd1),
	.w7(32'h38b0d674),
	.w8(32'hbbe357f8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc723d9),
	.w1(32'hbb0bb43a),
	.w2(32'h3b9a4503),
	.w3(32'h3c465b93),
	.w4(32'hbb8af5c1),
	.w5(32'hbba46e4c),
	.w6(32'hbbb482a2),
	.w7(32'h3bfeaeb4),
	.w8(32'hbaa38c75),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a5655),
	.w1(32'h3a0ff0b0),
	.w2(32'h39f9224f),
	.w3(32'hbb864f8f),
	.w4(32'h3b42534e),
	.w5(32'hb7551e5a),
	.w6(32'hbaa94ada),
	.w7(32'hbb6be0ab),
	.w8(32'hbbfac164),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba865e35),
	.w1(32'hbbfd7517),
	.w2(32'hbad17ada),
	.w3(32'h3bfb9750),
	.w4(32'h3bbd6239),
	.w5(32'hbc03f06d),
	.w6(32'hbc6580be),
	.w7(32'h3ae67a1d),
	.w8(32'hbb494bed),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2f51f),
	.w1(32'hbba127e6),
	.w2(32'h3adf8eaf),
	.w3(32'h3b9ebe84),
	.w4(32'hbb839add),
	.w5(32'h3b083c7b),
	.w6(32'h3ad2dce3),
	.w7(32'h3c357ea4),
	.w8(32'hb98bfb8b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba08fd),
	.w1(32'hbc0a3aa6),
	.w2(32'hbb223648),
	.w3(32'h3ce113e8),
	.w4(32'h39ad79f5),
	.w5(32'h3b1e8647),
	.w6(32'hbc66ecfb),
	.w7(32'hbc329a66),
	.w8(32'hbb9ffbe3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6241c),
	.w1(32'hbb32df52),
	.w2(32'hbaf16af6),
	.w3(32'h3b2b5dc7),
	.w4(32'h3ac4c97f),
	.w5(32'hbbcea851),
	.w6(32'h3aeea0e0),
	.w7(32'hbb23e752),
	.w8(32'h3b90429a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61fcc4),
	.w1(32'hbb7b063b),
	.w2(32'h37c01a5e),
	.w3(32'hbab80726),
	.w4(32'hbb3d057f),
	.w5(32'h3b29484f),
	.w6(32'hbbed0ab9),
	.w7(32'hbb255fbd),
	.w8(32'hbbcb2d1b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaa9b2),
	.w1(32'h3af30439),
	.w2(32'h3acd5699),
	.w3(32'hbba3140e),
	.w4(32'h3c23353f),
	.w5(32'hbb972058),
	.w6(32'h3c8d4f68),
	.w7(32'hba8f0c27),
	.w8(32'hbbe249df),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b14282),
	.w1(32'hbc43829a),
	.w2(32'h3b8b485a),
	.w3(32'hbbf7dbf6),
	.w4(32'hbc29c238),
	.w5(32'hbc3bae51),
	.w6(32'hbb2495c9),
	.w7(32'hba6c7a6f),
	.w8(32'hbba4ccb7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda0838),
	.w1(32'h3b58cb1d),
	.w2(32'h3b97658e),
	.w3(32'hba0f5762),
	.w4(32'h3d20ef5c),
	.w5(32'h3bd693de),
	.w6(32'hbae3ad4e),
	.w7(32'h3c49d979),
	.w8(32'hbc25c506),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc266010),
	.w1(32'hbbd2d0eb),
	.w2(32'hb90b97ac),
	.w3(32'hbc0f90db),
	.w4(32'h3adb8e6d),
	.w5(32'h3a863c5d),
	.w6(32'hbbca16f3),
	.w7(32'hbb87c153),
	.w8(32'hbbc661f2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8840d7),
	.w1(32'hba286988),
	.w2(32'h3b3eb9f6),
	.w3(32'h3be89f66),
	.w4(32'h3b8b33dc),
	.w5(32'hb898fce3),
	.w6(32'hbad4fbd1),
	.w7(32'h3be5cdd5),
	.w8(32'h3ac3f98b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7358e),
	.w1(32'h3aa59289),
	.w2(32'hbb1e6b65),
	.w3(32'hbc43932f),
	.w4(32'hb9982233),
	.w5(32'hbc333a39),
	.w6(32'hbc63000c),
	.w7(32'h3a0d316a),
	.w8(32'hbb8f41a6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d07c8),
	.w1(32'hbb804868),
	.w2(32'hbbf84a01),
	.w3(32'h3c87b8bc),
	.w4(32'h3b0e5502),
	.w5(32'hbc20d258),
	.w6(32'h3ac86bce),
	.w7(32'h3b5662a9),
	.w8(32'hb9f9a386),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bbacc),
	.w1(32'h3af1c711),
	.w2(32'hbc70e103),
	.w3(32'hbbcbc939),
	.w4(32'h3c5c8b22),
	.w5(32'hbbaba7d7),
	.w6(32'hbbab2e21),
	.w7(32'h3c2131f2),
	.w8(32'hbaaebf9a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b937b),
	.w1(32'h3c8b153e),
	.w2(32'h3b93790a),
	.w3(32'h3ab3044b),
	.w4(32'h3b493f39),
	.w5(32'h3b837472),
	.w6(32'hbc188928),
	.w7(32'h3b783d36),
	.w8(32'hbb488a32),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c889b0d),
	.w1(32'hbc04e642),
	.w2(32'hba69cb41),
	.w3(32'hbbdd2de4),
	.w4(32'h3c471206),
	.w5(32'hbbc698fd),
	.w6(32'hbb55f34e),
	.w7(32'hbb1b7f70),
	.w8(32'h3b416a5d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb165),
	.w1(32'hbaaa6ee4),
	.w2(32'h3b6da325),
	.w3(32'hbc291853),
	.w4(32'h3b20e747),
	.w5(32'h3bf635f5),
	.w6(32'hbc209dba),
	.w7(32'hbb36adef),
	.w8(32'h3b2bbfc8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a848772),
	.w1(32'h3ad99d8c),
	.w2(32'hbbb5405c),
	.w3(32'h3aefc1d3),
	.w4(32'hbc918314),
	.w5(32'hbaea934e),
	.w6(32'h3bf97ec7),
	.w7(32'hbc3cffb1),
	.w8(32'h3c6f4856),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc3890),
	.w1(32'hbc1f36ee),
	.w2(32'h3bd628df),
	.w3(32'hbbb85d06),
	.w4(32'hbcd869d1),
	.w5(32'h3b51f63a),
	.w6(32'hbbcc4f43),
	.w7(32'hbbc49a7d),
	.w8(32'hbc290138),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf82d63),
	.w1(32'hbb22c09e),
	.w2(32'hbc36b31f),
	.w3(32'hbbd0136e),
	.w4(32'h3995423e),
	.w5(32'hb9a8e16d),
	.w6(32'hbb0bd35b),
	.w7(32'hbb672fe4),
	.w8(32'hbb83b962),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0fe52),
	.w1(32'h3cec1c7d),
	.w2(32'h3b63a8e2),
	.w3(32'hbc0cbb7c),
	.w4(32'h3c06514b),
	.w5(32'h3a25df72),
	.w6(32'h3bf7578b),
	.w7(32'h3abfd409),
	.w8(32'hba580570),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ddaa3),
	.w1(32'hb9d861c3),
	.w2(32'h3b650037),
	.w3(32'hbbf2337c),
	.w4(32'hbb4ab0d8),
	.w5(32'hbc05da5e),
	.w6(32'hbc82fcb1),
	.w7(32'h3bdf33dc),
	.w8(32'h3bc7985a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275d05),
	.w1(32'h3c0e1430),
	.w2(32'hbb22f176),
	.w3(32'h3b074a02),
	.w4(32'hb6ba8af1),
	.w5(32'h3cc19aba),
	.w6(32'h3b1574ff),
	.w7(32'hbb93663a),
	.w8(32'hbc02f07e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93be8a),
	.w1(32'hbb894d38),
	.w2(32'h3a296baa),
	.w3(32'h3a9bd0da),
	.w4(32'hbc819a2e),
	.w5(32'h3c349624),
	.w6(32'h3bf76d32),
	.w7(32'hbbb2377a),
	.w8(32'hbc58ca10),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c9f8d),
	.w1(32'hbc192629),
	.w2(32'hbac0a165),
	.w3(32'hbb6a1455),
	.w4(32'h3bd347e3),
	.w5(32'hbc0afef1),
	.w6(32'hbc68cee0),
	.w7(32'h3b62deff),
	.w8(32'hbcaee939),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aec4f),
	.w1(32'h3bab357f),
	.w2(32'hbb0d51cd),
	.w3(32'h3b9045e9),
	.w4(32'hba86a746),
	.w5(32'h3af6b1bf),
	.w6(32'h3c07c2f0),
	.w7(32'h3a051606),
	.w8(32'hbb972956),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ab4ea),
	.w1(32'hb9c93e13),
	.w2(32'h3a834d3e),
	.w3(32'hbc0744b1),
	.w4(32'h3bf076cd),
	.w5(32'h3ae96551),
	.w6(32'h3b8afff4),
	.w7(32'h3acdda2e),
	.w8(32'hbba0fd59),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e2170),
	.w1(32'hbc1618ed),
	.w2(32'h3c8f1959),
	.w3(32'hbc460b9a),
	.w4(32'h3b993e0a),
	.w5(32'hbc59da3d),
	.w6(32'hbb0f8dab),
	.w7(32'hbb51e7fd),
	.w8(32'h3c573f17),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4f47),
	.w1(32'hbb27f4b9),
	.w2(32'h3a8e496b),
	.w3(32'h3c1d8eb4),
	.w4(32'h3b35a0fb),
	.w5(32'h3abfd070),
	.w6(32'h39068ed0),
	.w7(32'h3bf0fc4f),
	.w8(32'hbaafcab5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc37c68),
	.w1(32'h3b6296e8),
	.w2(32'h3cb31586),
	.w3(32'hbbba9ced),
	.w4(32'h3a960774),
	.w5(32'hb96c6f8e),
	.w6(32'h35754691),
	.w7(32'h3b076659),
	.w8(32'hbc9ddb41),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855a7c),
	.w1(32'h3c80a104),
	.w2(32'h3ad19179),
	.w3(32'hbb0de759),
	.w4(32'hbc8134b1),
	.w5(32'hbb193fdc),
	.w6(32'hbc23fdd3),
	.w7(32'hba985a6c),
	.w8(32'hbc1b46f1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01dd00),
	.w1(32'h3cfc14ad),
	.w2(32'h3b8fd7ff),
	.w3(32'h3c07d4f9),
	.w4(32'hbaba37ea),
	.w5(32'hbc17037f),
	.w6(32'h3af8f2ac),
	.w7(32'h3b6ba63a),
	.w8(32'h3d1e5fbd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ac2e9),
	.w1(32'h3ad9d951),
	.w2(32'hbc5ba773),
	.w3(32'hbbe1d822),
	.w4(32'h3cc6f5d7),
	.w5(32'hbbc5831a),
	.w6(32'h3bb40d7b),
	.w7(32'hbb301937),
	.w8(32'hba15f670),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bfba7),
	.w1(32'hbc23bf03),
	.w2(32'h3b2329b0),
	.w3(32'hbaa0d677),
	.w4(32'hbbaaf349),
	.w5(32'hbb8f227f),
	.w6(32'h3c8d91ff),
	.w7(32'hbb9657e6),
	.w8(32'h3b85dbf7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf049c),
	.w1(32'hbad6033b),
	.w2(32'h39a1a959),
	.w3(32'h3856e251),
	.w4(32'hbb97bddf),
	.w5(32'h3b2d302d),
	.w6(32'hbb75a10a),
	.w7(32'hbbc5a5d1),
	.w8(32'h3b7713a8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ad232),
	.w1(32'h3ab5b3dd),
	.w2(32'h3adc2d21),
	.w3(32'hbb0903b0),
	.w4(32'hb99376b7),
	.w5(32'h3aaa63bf),
	.w6(32'h36713671),
	.w7(32'h3b296586),
	.w8(32'h3b2201f2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0b5a5),
	.w1(32'hbb850cd4),
	.w2(32'h3b158223),
	.w3(32'hbb2f9b0b),
	.w4(32'hbb9b5a0e),
	.w5(32'h3c473765),
	.w6(32'hbaf2bf1f),
	.w7(32'hbc227b14),
	.w8(32'h3bcb0ee4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb764331),
	.w1(32'hbb842d7f),
	.w2(32'h3b6d6c6a),
	.w3(32'h3c2f0997),
	.w4(32'hba083bb8),
	.w5(32'h3b92dc0d),
	.w6(32'hbb34ac88),
	.w7(32'hbc341ca2),
	.w8(32'h3b4db8eb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b825ca),
	.w1(32'h3bac4bac),
	.w2(32'h3bd23375),
	.w3(32'hbb1d2bc4),
	.w4(32'h3d0809c4),
	.w5(32'hb9b45ba2),
	.w6(32'h3a05337b),
	.w7(32'hbc003a8c),
	.w8(32'hbc98002f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f268f),
	.w1(32'h3aee67d4),
	.w2(32'hbb8d9f53),
	.w3(32'hb947de09),
	.w4(32'hb89dbfd1),
	.w5(32'hbba757cb),
	.w6(32'hb990b886),
	.w7(32'hbb9b7f48),
	.w8(32'hba88a072),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a629fd3),
	.w1(32'h3bbc02bb),
	.w2(32'h3b685e12),
	.w3(32'h3a925c9a),
	.w4(32'hbb39203a),
	.w5(32'h3b4e6903),
	.w6(32'h3c0a8a5e),
	.w7(32'hbb7b361b),
	.w8(32'hbbf588e5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba30d0e),
	.w1(32'h3ca32a38),
	.w2(32'h3a9c87b5),
	.w3(32'hbbfc27dc),
	.w4(32'h3b90ff61),
	.w5(32'hbbeb6c2d),
	.w6(32'h3baf6b6f),
	.w7(32'h3c212287),
	.w8(32'h3a69f8af),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76cb7c),
	.w1(32'hbb39bda1),
	.w2(32'hbbb72e8e),
	.w3(32'h3b161f15),
	.w4(32'hbb9b4434),
	.w5(32'hbc5f1f5f),
	.w6(32'hbc497d18),
	.w7(32'h3a03fc76),
	.w8(32'hbb36bb4f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b488ca5),
	.w1(32'h3b8709e9),
	.w2(32'hbabd61de),
	.w3(32'hbbeca12b),
	.w4(32'hbc2bbdf9),
	.w5(32'h3ba2d87f),
	.w6(32'h3a326866),
	.w7(32'h3c34deca),
	.w8(32'hbb72ff64),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2149b),
	.w1(32'h3c184aa0),
	.w2(32'hba934d4b),
	.w3(32'h3b9afe9c),
	.w4(32'hbb1d388b),
	.w5(32'h3ac54580),
	.w6(32'hbb9e271f),
	.w7(32'h3bba485d),
	.w8(32'h3b9aa095),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4b084),
	.w1(32'hbc15d1cf),
	.w2(32'h3b8a2d89),
	.w3(32'hbb2d6aff),
	.w4(32'h3c51d90d),
	.w5(32'h3bdd4e1f),
	.w6(32'hbb48e574),
	.w7(32'h3bb2ead6),
	.w8(32'h3a16bfa9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7f58e),
	.w1(32'hbb618fac),
	.w2(32'h3ba10e7c),
	.w3(32'hba5fba3f),
	.w4(32'hbc886390),
	.w5(32'h3bd88346),
	.w6(32'h3bf5509e),
	.w7(32'hbabfad76),
	.w8(32'hb9eac703),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e2cef),
	.w1(32'hbb5659ec),
	.w2(32'h3c01ddc0),
	.w3(32'h38d7d165),
	.w4(32'h3c721638),
	.w5(32'h3b12efb1),
	.w6(32'hbc28874d),
	.w7(32'hbb64dfe9),
	.w8(32'hba91348d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f783c),
	.w1(32'h3c02c718),
	.w2(32'h3b09f473),
	.w3(32'h3b56a983),
	.w4(32'hbb8c80b1),
	.w5(32'hbc348a3e),
	.w6(32'h3b1552da),
	.w7(32'h3ae953ea),
	.w8(32'hbc3034ff),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ecf8a),
	.w1(32'hbc0c6fb8),
	.w2(32'hbbce480c),
	.w3(32'hbbc9813b),
	.w4(32'hbbf9dda9),
	.w5(32'hbaceccf0),
	.w6(32'hba13b039),
	.w7(32'hbac58cdb),
	.w8(32'hbb103f4e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ccb77),
	.w1(32'hbbcafa62),
	.w2(32'hba5e7a4e),
	.w3(32'h3c4a6c0e),
	.w4(32'h3a3226b4),
	.w5(32'hbb8df7a3),
	.w6(32'h3c3e67f9),
	.w7(32'hbc1af0b4),
	.w8(32'h3969a55e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb535a0),
	.w1(32'hbb0f54bb),
	.w2(32'h3c330c90),
	.w3(32'h3aaa57dc),
	.w4(32'hbb987123),
	.w5(32'h3b969b11),
	.w6(32'hbb80f6ed),
	.w7(32'hbab2d558),
	.w8(32'h3c91846a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9337cf),
	.w1(32'h3bd42eef),
	.w2(32'hba419407),
	.w3(32'h3a677c5b),
	.w4(32'hbcfdc862),
	.w5(32'h3c0e6f1b),
	.w6(32'h3c9c58cc),
	.w7(32'hbc696052),
	.w8(32'hbb29283a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0a38c),
	.w1(32'hba9e47fa),
	.w2(32'hbb206465),
	.w3(32'h3c48d2ab),
	.w4(32'h3c23c5bb),
	.w5(32'h3bca482d),
	.w6(32'hbb1ce806),
	.w7(32'h3b6207a5),
	.w8(32'hbac8d21c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c028237),
	.w1(32'hba80ef8e),
	.w2(32'hba45bf89),
	.w3(32'hbb76a480),
	.w4(32'hbbc13a04),
	.w5(32'h3c36bd5e),
	.w6(32'h3c17d9d8),
	.w7(32'hbc828b74),
	.w8(32'h39bf920d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01a58a),
	.w1(32'h3ba0b022),
	.w2(32'hbaa26270),
	.w3(32'h3c6d920a),
	.w4(32'h38f3a28f),
	.w5(32'hbc413030),
	.w6(32'h3a907fa5),
	.w7(32'h3c03c123),
	.w8(32'h3c0b57c9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0daca1),
	.w1(32'hbbf84c22),
	.w2(32'h3c5485ba),
	.w3(32'hbbf03e2c),
	.w4(32'hba8f0276),
	.w5(32'h376c1bce),
	.w6(32'h3b8a0bb0),
	.w7(32'h3c1da38f),
	.w8(32'hbab0cf8d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00a2b3),
	.w1(32'hb8b3c326),
	.w2(32'h34bb9a8f),
	.w3(32'h3a574026),
	.w4(32'h3c137791),
	.w5(32'hbc283908),
	.w6(32'hbc1acb85),
	.w7(32'h3a0431a1),
	.w8(32'hbb95c6bc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e2894),
	.w1(32'h3c498a07),
	.w2(32'h3aa94115),
	.w3(32'hbb564e86),
	.w4(32'hba9a9fc2),
	.w5(32'h3b94e550),
	.w6(32'hbb438a70),
	.w7(32'hbbc64caf),
	.w8(32'hbb6e75a2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f33c),
	.w1(32'h3b6b70d2),
	.w2(32'h3b48b120),
	.w3(32'h3a9e1e8d),
	.w4(32'hba2c64ba),
	.w5(32'h3ca13c26),
	.w6(32'hba9d5eb3),
	.w7(32'hbaf0f855),
	.w8(32'h3baaaed4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6a34a),
	.w1(32'h3a5a3dbd),
	.w2(32'h3c62951b),
	.w3(32'h3bd98eec),
	.w4(32'hbb48ebe8),
	.w5(32'hbc2951b5),
	.w6(32'hbc512d94),
	.w7(32'hbba013a3),
	.w8(32'hbabb30ca),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9922102),
	.w1(32'h3c7ff5cb),
	.w2(32'h3c345056),
	.w3(32'hbc07ef1c),
	.w4(32'h3b8f4068),
	.w5(32'hba1bb651),
	.w6(32'hbb0114c2),
	.w7(32'hbae2d744),
	.w8(32'h3b03bf0f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c202559),
	.w1(32'h3c2572cd),
	.w2(32'hbc6d822d),
	.w3(32'hbade6657),
	.w4(32'h3abe4164),
	.w5(32'h3ba4e82b),
	.w6(32'hbb9c8e8a),
	.w7(32'h369e0156),
	.w8(32'hbb1833af),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6b45e),
	.w1(32'hbcf4e79a),
	.w2(32'h39156526),
	.w3(32'h39d08f7c),
	.w4(32'h3c18ed54),
	.w5(32'hbc4c7cfc),
	.w6(32'hbb3e9472),
	.w7(32'h3b08ffc8),
	.w8(32'hba2a3440),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ce60d),
	.w1(32'h3c960ee9),
	.w2(32'h3b974ac5),
	.w3(32'h3b2f6877),
	.w4(32'hbbc8e671),
	.w5(32'hbc1d7328),
	.w6(32'hbb24cce5),
	.w7(32'h3c6f8d01),
	.w8(32'hbc0d8335),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa9782),
	.w1(32'hbb29c4bf),
	.w2(32'h3b1d2dcb),
	.w3(32'h3a616542),
	.w4(32'h381b056e),
	.w5(32'h3b0baa1e),
	.w6(32'hbb439eb4),
	.w7(32'h3b7f38a4),
	.w8(32'hbb922aee),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf94012),
	.w1(32'hbb3d665e),
	.w2(32'h3b3a4739),
	.w3(32'hbc1aa1d8),
	.w4(32'hba6462db),
	.w5(32'h3ae0f6eb),
	.w6(32'h3bac5b95),
	.w7(32'hbb753a78),
	.w8(32'hb9f51e38),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fe8ca),
	.w1(32'h3a5249d5),
	.w2(32'hb9018502),
	.w3(32'h3a14dcc0),
	.w4(32'h3c0ac7a3),
	.w5(32'h3bcf43da),
	.w6(32'hbad13072),
	.w7(32'h3a4b4c52),
	.w8(32'h3a0aba73),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f669),
	.w1(32'hb857e190),
	.w2(32'h3b8ee816),
	.w3(32'hbaed1d90),
	.w4(32'h388247dd),
	.w5(32'h3be3882b),
	.w6(32'hbb575a57),
	.w7(32'h3b5c945d),
	.w8(32'hbc5a277f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50dc1f),
	.w1(32'hbb5291a4),
	.w2(32'h3ba9e72e),
	.w3(32'h3b70a884),
	.w4(32'hbcba4fa0),
	.w5(32'h3bf06e01),
	.w6(32'h3c133458),
	.w7(32'h3b249adb),
	.w8(32'hbada877d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800edc),
	.w1(32'h3c397d44),
	.w2(32'h3c3c8129),
	.w3(32'hbb96218a),
	.w4(32'h3c3478d5),
	.w5(32'hbc0201d1),
	.w6(32'hba09629e),
	.w7(32'h3bf64a0d),
	.w8(32'hbb675640),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8af78),
	.w1(32'h3bd82549),
	.w2(32'h3c43938a),
	.w3(32'hbc4d1370),
	.w4(32'h3d0742bf),
	.w5(32'hbbd4b512),
	.w6(32'hbbe41055),
	.w7(32'hbb68bc81),
	.w8(32'h3c221d62),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdef52e),
	.w1(32'h3911c273),
	.w2(32'hbb29f6c6),
	.w3(32'h3c2365bb),
	.w4(32'h3b1379e7),
	.w5(32'hbc0d5f33),
	.w6(32'hbac90a37),
	.w7(32'h3c2327c8),
	.w8(32'hb93fe9de),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7438a9),
	.w1(32'hbc1ffc42),
	.w2(32'hbb5cd932),
	.w3(32'hbc2b6b1c),
	.w4(32'hbbf7fab2),
	.w5(32'hbb612b17),
	.w6(32'hbbe22322),
	.w7(32'h3bb3a2e9),
	.w8(32'h3b6ce765),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b70c5),
	.w1(32'hbac1f52f),
	.w2(32'h3ab4fb9f),
	.w3(32'h3a8cdcea),
	.w4(32'hbb58c203),
	.w5(32'h3bd086a6),
	.w6(32'hbbef76b0),
	.w7(32'hbba63c8f),
	.w8(32'h3c3b03d6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a057f),
	.w1(32'hbd9da7b0),
	.w2(32'h3c142764),
	.w3(32'h3b88a90b),
	.w4(32'h3b1f8f5d),
	.w5(32'h3a9cb0b1),
	.w6(32'hbc118874),
	.w7(32'hbbd2c2ff),
	.w8(32'hbbd5f5df),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc660579),
	.w1(32'h3b6e48d7),
	.w2(32'hbb889b4d),
	.w3(32'hbb57a99d),
	.w4(32'hbbd8d4e6),
	.w5(32'h3baa5276),
	.w6(32'hbad3e730),
	.w7(32'hbc185e48),
	.w8(32'hbc578598),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3914a),
	.w1(32'h3be7d09a),
	.w2(32'h3b89f52b),
	.w3(32'hbbab91ef),
	.w4(32'h3b221034),
	.w5(32'h3c500d83),
	.w6(32'h3c170624),
	.w7(32'h3c19ad10),
	.w8(32'h3c23b6c6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcb100),
	.w1(32'h3c53779d),
	.w2(32'h3ba77014),
	.w3(32'h3b809050),
	.w4(32'hbb91a0e9),
	.w5(32'hbc1d1427),
	.w6(32'h3b01cd4b),
	.w7(32'h3b47f1e9),
	.w8(32'h3afb41b2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4897bb),
	.w1(32'hbb70d07c),
	.w2(32'hbc0d2d4d),
	.w3(32'hbc299af7),
	.w4(32'h3bd05cfe),
	.w5(32'h3bb1c2b1),
	.w6(32'h3c0dcd02),
	.w7(32'h3c0dc026),
	.w8(32'hbbaa6119),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbed81),
	.w1(32'hbd2db260),
	.w2(32'hbbda3878),
	.w3(32'hbb93389f),
	.w4(32'h3c0d0c35),
	.w5(32'hbc9ccb76),
	.w6(32'h3bdaa176),
	.w7(32'hba078a0b),
	.w8(32'h3b6c5a90),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62952a),
	.w1(32'h3a57186b),
	.w2(32'hbbf37b5a),
	.w3(32'h3bffb3da),
	.w4(32'h3ae61381),
	.w5(32'h3c29c862),
	.w6(32'hbc28ad6c),
	.w7(32'h3b587484),
	.w8(32'hbc3b5630),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bb734),
	.w1(32'hba57471b),
	.w2(32'hbc0fe9eb),
	.w3(32'h3bb4cf5b),
	.w4(32'h3c8f7192),
	.w5(32'hbb091068),
	.w6(32'h3ca3a93f),
	.w7(32'h3be50e0d),
	.w8(32'h3b0de6ff),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d5a2),
	.w1(32'hba233d4a),
	.w2(32'hb9f6f92f),
	.w3(32'hbc13bac5),
	.w4(32'h3aac828f),
	.w5(32'hbbc9e037),
	.w6(32'h3c6b9d1f),
	.w7(32'hbb9d6a04),
	.w8(32'h3a0aba41),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf6d25),
	.w1(32'hba80080b),
	.w2(32'hbc855575),
	.w3(32'hbb6c5286),
	.w4(32'hbc5b99eb),
	.w5(32'h3b7b138d),
	.w6(32'h3d076ce7),
	.w7(32'h3c1f7e73),
	.w8(32'h3b5f1793),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69c033),
	.w1(32'hbb0df7d2),
	.w2(32'hbc314ab8),
	.w3(32'h3b833ef5),
	.w4(32'h3c43b024),
	.w5(32'hbbc51a6b),
	.w6(32'hbae9484c),
	.w7(32'hbaaaaaf9),
	.w8(32'hbbaa5dd7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972731),
	.w1(32'hbb518e2e),
	.w2(32'hbb9fa249),
	.w3(32'h36c7161b),
	.w4(32'h3c859d2f),
	.w5(32'hbce656e9),
	.w6(32'hbaa1f222),
	.w7(32'h3ce46aea),
	.w8(32'h3b40bbfd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03daa1),
	.w1(32'h3b8eba85),
	.w2(32'h3a78c53d),
	.w3(32'h3b06fb3a),
	.w4(32'hba03d593),
	.w5(32'h3a8fcf50),
	.w6(32'h3c41d259),
	.w7(32'h3bf4fe39),
	.w8(32'h3bd7fbda),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831c47),
	.w1(32'hbb96088a),
	.w2(32'hba076b46),
	.w3(32'h394b3835),
	.w4(32'hbbbf912a),
	.w5(32'h3cd91e97),
	.w6(32'h3b30969b),
	.w7(32'h3c3d911e),
	.w8(32'hbc113206),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba41c03),
	.w1(32'h3ae22df6),
	.w2(32'hbb97db43),
	.w3(32'hbbe0fd89),
	.w4(32'hbafa1ce6),
	.w5(32'hbbe05d07),
	.w6(32'hbba6b593),
	.w7(32'h39962ee7),
	.w8(32'hbc10509f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931e9f),
	.w1(32'hbac0fa7d),
	.w2(32'hbc154455),
	.w3(32'hbace36d2),
	.w4(32'h3b9422b3),
	.w5(32'hbc744d3f),
	.w6(32'hbb12d711),
	.w7(32'hbc1f110d),
	.w8(32'h3aa53f06),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350a3cc0),
	.w1(32'h3b11f598),
	.w2(32'h3b34d888),
	.w3(32'hbb80d529),
	.w4(32'h3b74f930),
	.w5(32'h3c0839d1),
	.w6(32'hbc4e1cae),
	.w7(32'hbc41717e),
	.w8(32'hbba9201f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96eb06),
	.w1(32'hbaa5b4f9),
	.w2(32'hbc950379),
	.w3(32'h3b9bd95d),
	.w4(32'hb9f7e4af),
	.w5(32'hbbed2e77),
	.w6(32'h3c137d83),
	.w7(32'hbc19c801),
	.w8(32'hbb72ef50),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aa3d9),
	.w1(32'h3c2a56c8),
	.w2(32'h3c706fd2),
	.w3(32'hbb155e15),
	.w4(32'hbc2e60f2),
	.w5(32'h3bb178d5),
	.w6(32'hbbd43b4d),
	.w7(32'hbb025f13),
	.w8(32'hbb4d124d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc2094),
	.w1(32'hba5e81a5),
	.w2(32'h3c3b8254),
	.w3(32'h3b2e614d),
	.w4(32'hbb3a26f4),
	.w5(32'h3c9752b7),
	.w6(32'hbc916346),
	.w7(32'hbbb69bc8),
	.w8(32'h3ae6a543),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a1d94),
	.w1(32'h3d3eb590),
	.w2(32'h3a576cc6),
	.w3(32'h3af621dc),
	.w4(32'hbbe8f5a1),
	.w5(32'h3c279ea7),
	.w6(32'hbb843a07),
	.w7(32'h3bff9b5b),
	.w8(32'hbaded20d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37dd2a),
	.w1(32'h3adf3af8),
	.w2(32'h399b3a8a),
	.w3(32'hb9d69223),
	.w4(32'hbcabee15),
	.w5(32'hbb9026de),
	.w6(32'hbad4d9c1),
	.w7(32'hbc812ed5),
	.w8(32'h3ace3cf0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0cb0),
	.w1(32'hbbbff7d4),
	.w2(32'h3b17aece),
	.w3(32'h3bf3eea4),
	.w4(32'hbb97844f),
	.w5(32'h3b3d79f4),
	.w6(32'hba1d2766),
	.w7(32'hbab89d86),
	.w8(32'hbbe3e0ee),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78cc4d),
	.w1(32'h3bc197aa),
	.w2(32'hbc3c0e1b),
	.w3(32'h3c11c743),
	.w4(32'hbbcf6bcd),
	.w5(32'h3c4ea43b),
	.w6(32'h3bfd93cd),
	.w7(32'hba203275),
	.w8(32'h3a889ae1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd8de1),
	.w1(32'hbc14a18c),
	.w2(32'h3bd6a80f),
	.w3(32'hbc190c86),
	.w4(32'h3ac024ff),
	.w5(32'hbc1f6790),
	.w6(32'hbc2896ff),
	.w7(32'h3b85ed57),
	.w8(32'h3c1de707),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd21e29),
	.w1(32'hbbd53255),
	.w2(32'h3b53d1c9),
	.w3(32'hbc605fdd),
	.w4(32'hba5a1d23),
	.w5(32'hbc4721e3),
	.w6(32'hbcb8c08e),
	.w7(32'h3b277894),
	.w8(32'h3b8d0a09),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97186a),
	.w1(32'h3abf57d6),
	.w2(32'h3a2ebc69),
	.w3(32'hbc6509f9),
	.w4(32'hbb89d321),
	.w5(32'h3b75a343),
	.w6(32'hbbcf0683),
	.w7(32'hbc271319),
	.w8(32'h3b99589b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92169d),
	.w1(32'hbc16e295),
	.w2(32'hb6fae548),
	.w3(32'hba1d6e6e),
	.w4(32'hba329fc7),
	.w5(32'h3b06d34b),
	.w6(32'h3b850d13),
	.w7(32'h3a050eb0),
	.w8(32'hbbb20ad4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule