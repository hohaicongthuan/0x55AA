module layer_8_featuremap_242(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8efe84),
	.w1(32'hbc13c10b),
	.w2(32'hbccad646),
	.w3(32'h3c3f3102),
	.w4(32'hbbc98b72),
	.w5(32'hbc7a850e),
	.w6(32'hbbddfe04),
	.w7(32'hbc22fa67),
	.w8(32'hbb9d258e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c9169),
	.w1(32'hbbd4388a),
	.w2(32'hbbe3212c),
	.w3(32'hbc8f1e20),
	.w4(32'hbbde42ea),
	.w5(32'hbba00b12),
	.w6(32'hbbd66d2c),
	.w7(32'hbbb9c9b5),
	.w8(32'hbb7efdf4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88282),
	.w1(32'hbc60ebf1),
	.w2(32'hbc889821),
	.w3(32'hbb383daa),
	.w4(32'hbbb32256),
	.w5(32'hbc1b4c76),
	.w6(32'h3b9cbc2c),
	.w7(32'h3b561c57),
	.w8(32'h3bd9d6b2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66290d),
	.w1(32'hbc2c307c),
	.w2(32'hbc50b0c4),
	.w3(32'hbba50ae0),
	.w4(32'hbbe835ee),
	.w5(32'hbc4ba785),
	.w6(32'h3b3e4d73),
	.w7(32'h3beb49c7),
	.w8(32'h3b65d393),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab21d97),
	.w1(32'hbb32de49),
	.w2(32'hbbbbf909),
	.w3(32'hbc3ae988),
	.w4(32'hbb75f9f9),
	.w5(32'hbb400581),
	.w6(32'hba4d83f8),
	.w7(32'h389f8504),
	.w8(32'h39a29ae9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5267a),
	.w1(32'h3ab72850),
	.w2(32'hbc339ed8),
	.w3(32'hba34c816),
	.w4(32'hbb8c31b0),
	.w5(32'hbc0ba036),
	.w6(32'h3b81cf36),
	.w7(32'h39c2cd81),
	.w8(32'hbbc430b0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20dbff),
	.w1(32'hbb5fbb53),
	.w2(32'hbbe99e30),
	.w3(32'h3ac2aba9),
	.w4(32'hbb9a682b),
	.w5(32'hbbdbfd29),
	.w6(32'hbb5d76b7),
	.w7(32'hbb51ba0e),
	.w8(32'hbb5f19f5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33bc16),
	.w1(32'hbab75562),
	.w2(32'hbc19d28b),
	.w3(32'hbb9e7369),
	.w4(32'hbc452ebf),
	.w5(32'hbc6d3f6c),
	.w6(32'h3c380e63),
	.w7(32'h3c0719d9),
	.w8(32'hbb01cd2e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ac8a),
	.w1(32'h3b8e2798),
	.w2(32'hba0450f1),
	.w3(32'hbca295c7),
	.w4(32'h3acfbf4c),
	.w5(32'hba284f98),
	.w6(32'h3bda852b),
	.w7(32'h3b84f828),
	.w8(32'h3bfa0a55),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7c32),
	.w1(32'hbc396e2a),
	.w2(32'hbc5fa2f6),
	.w3(32'h3ab23142),
	.w4(32'h3b8d3d9b),
	.w5(32'hba3e6e69),
	.w6(32'hbc8b432c),
	.w7(32'hbbf2f0ae),
	.w8(32'hbb876256),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075c2e),
	.w1(32'hbc32f0ca),
	.w2(32'hbc2863e3),
	.w3(32'hbbbf3a54),
	.w4(32'hbbdcf441),
	.w5(32'hbc6cf4ea),
	.w6(32'hbbf87093),
	.w7(32'hbbc822eb),
	.w8(32'hbb6ad5b6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c2ce9),
	.w1(32'hbb0d6b2b),
	.w2(32'hbc0efb7a),
	.w3(32'hbc246aa5),
	.w4(32'hbb921e32),
	.w5(32'hbc07b761),
	.w6(32'hbb37b2a7),
	.w7(32'hbb8f8abf),
	.w8(32'hbbb3e238),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93fc5e),
	.w1(32'hbb84530e),
	.w2(32'hbbf8ab98),
	.w3(32'hbb4abf8a),
	.w4(32'hbbb725cd),
	.w5(32'hbb3b024f),
	.w6(32'h39282a9b),
	.w7(32'hbaf21ff9),
	.w8(32'hbbc0a30a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f20bf),
	.w1(32'hbb3fa356),
	.w2(32'hbc28425f),
	.w3(32'hbb8c33c5),
	.w4(32'h3b63cbd6),
	.w5(32'hb9b679e6),
	.w6(32'hbb370090),
	.w7(32'hbbd94488),
	.w8(32'h3bf3de67),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa51b6e),
	.w1(32'h3b000701),
	.w2(32'h3c1bcb1d),
	.w3(32'hb95dff36),
	.w4(32'h3acc0b6a),
	.w5(32'h3bbb1bdd),
	.w6(32'hbb899797),
	.w7(32'hba3720ef),
	.w8(32'hbb02e50a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf5bf1),
	.w1(32'hbb81c6aa),
	.w2(32'hbc8d3dec),
	.w3(32'h39720441),
	.w4(32'hbbf0c33f),
	.w5(32'hbc1c18b4),
	.w6(32'hbc201687),
	.w7(32'hbc7a6936),
	.w8(32'hbbb1d922),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc123799),
	.w1(32'hbc02e919),
	.w2(32'hbc52d465),
	.w3(32'hba926677),
	.w4(32'h3bb354a9),
	.w5(32'hbaa3a1e6),
	.w6(32'hbab59d88),
	.w7(32'hbbf7d4b4),
	.w8(32'hbb5cdc01),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b3d03),
	.w1(32'h3a4f8628),
	.w2(32'hba3de71f),
	.w3(32'hbb847ca0),
	.w4(32'hba25c7a2),
	.w5(32'h3aedeaa6),
	.w6(32'hbb987ae3),
	.w7(32'hbbbb6bb6),
	.w8(32'h3b00c7e9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f8618),
	.w1(32'hbac0eeea),
	.w2(32'hbb9299bb),
	.w3(32'h3b4f9de6),
	.w4(32'hbbd7298a),
	.w5(32'hbbcb76c9),
	.w6(32'hbc500c97),
	.w7(32'hbbcf5d35),
	.w8(32'h3b6386dc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f5c15),
	.w1(32'hbbd02317),
	.w2(32'hbc1f6456),
	.w3(32'hbb1b477a),
	.w4(32'hbb6651a6),
	.w5(32'hbc22a138),
	.w6(32'hbb553dcd),
	.w7(32'hbbd68720),
	.w8(32'hbb834455),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb8dd6),
	.w1(32'hbbf704f9),
	.w2(32'hbc6c4a3b),
	.w3(32'hbbf83415),
	.w4(32'h3af2c509),
	.w5(32'hbc5fe095),
	.w6(32'hbc38e72b),
	.w7(32'hbc89f0c6),
	.w8(32'hbc4e1dbb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b1fc),
	.w1(32'h3b9a9c61),
	.w2(32'hba0f01fe),
	.w3(32'hbbbcd351),
	.w4(32'h3b8c712e),
	.w5(32'h3b8ac00a),
	.w6(32'h3bbc0064),
	.w7(32'hbacb0d82),
	.w8(32'h3afac532),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa11d6b),
	.w1(32'hbb8bb087),
	.w2(32'hbc7dcb35),
	.w3(32'h39b5480a),
	.w4(32'hbc21a7cc),
	.w5(32'hbc2efb36),
	.w6(32'hbb156709),
	.w7(32'hbbc2bbf0),
	.w8(32'hbc0f44fa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd6bed),
	.w1(32'h3c507e44),
	.w2(32'h3c014880),
	.w3(32'h3b502f65),
	.w4(32'h3b93ba88),
	.w5(32'h3b930b72),
	.w6(32'h3b3a7661),
	.w7(32'hba48e13b),
	.w8(32'h3b3b1306),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0906),
	.w1(32'hbba80e94),
	.w2(32'hbbd1894a),
	.w3(32'h3baab785),
	.w4(32'hbb332d99),
	.w5(32'h3a46c4aa),
	.w6(32'hbb80fbb8),
	.w7(32'hbb12e241),
	.w8(32'hbae66948),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb382328),
	.w1(32'hbc6626d7),
	.w2(32'hbcdb1abe),
	.w3(32'h3bb4c3bb),
	.w4(32'hbc504c86),
	.w5(32'hbc1a81bb),
	.w6(32'hbc95cd6e),
	.w7(32'hbce559b6),
	.w8(32'hbc92666b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc0ca6),
	.w1(32'hbc432099),
	.w2(32'hbca70b2f),
	.w3(32'hbc8044e5),
	.w4(32'hbc434bd2),
	.w5(32'hbc90afca),
	.w6(32'h3b2b62d3),
	.w7(32'h3ab7c535),
	.w8(32'h3ab59179),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca154b3),
	.w1(32'hbbd71dcc),
	.w2(32'hbbf562a3),
	.w3(32'hbbd344f5),
	.w4(32'h3bb362a7),
	.w5(32'hbba338c3),
	.w6(32'hbbaf35fe),
	.w7(32'h3bc8af75),
	.w8(32'h3b4df222),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed80dc),
	.w1(32'hb9e15628),
	.w2(32'hbbcec28a),
	.w3(32'hbbbeed04),
	.w4(32'h3a70ca4b),
	.w5(32'hbb599181),
	.w6(32'h3b0b9fa3),
	.w7(32'hba47e028),
	.w8(32'h3ad77019),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e7fa),
	.w1(32'h3bbc617d),
	.w2(32'h3be0117f),
	.w3(32'hb98158f7),
	.w4(32'hb9e8e690),
	.w5(32'h3b0461d8),
	.w6(32'h3b013591),
	.w7(32'h3af934f1),
	.w8(32'h3c7f2f3e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb22b97),
	.w1(32'hbbef8f1b),
	.w2(32'hbc03172b),
	.w3(32'h3c82ccdf),
	.w4(32'hbb34c43e),
	.w5(32'hbaa54b46),
	.w6(32'hbb921c06),
	.w7(32'hbb32e515),
	.w8(32'hbac431b0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b77df),
	.w1(32'h3c1d2201),
	.w2(32'h3c2c5806),
	.w3(32'h3ad4be22),
	.w4(32'h3b66d322),
	.w5(32'h3bd3d3c0),
	.w6(32'h3b3bfebf),
	.w7(32'h3c040988),
	.w8(32'h3b0a4570),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3b8d),
	.w1(32'hbb9ef6d6),
	.w2(32'hbc81184e),
	.w3(32'h3aeee218),
	.w4(32'hbb63f91c),
	.w5(32'hbbe4ef0f),
	.w6(32'hbc8b5056),
	.w7(32'hbc93a580),
	.w8(32'hbb2fcd0d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a49b9),
	.w1(32'h3bbbb871),
	.w2(32'h3c2ce715),
	.w3(32'hbbc71620),
	.w4(32'h3b0d2792),
	.w5(32'h3ba36f3d),
	.w6(32'hbb0d3e69),
	.w7(32'h3bed2c51),
	.w8(32'h3ba63e59),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5db6c2),
	.w1(32'h3b2a2e24),
	.w2(32'h39c27a5f),
	.w3(32'h3bf04285),
	.w4(32'hbb68a01c),
	.w5(32'hba702ff6),
	.w6(32'hb8abe531),
	.w7(32'hbb0aef9d),
	.w8(32'h3b02eca8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b361863),
	.w1(32'h39ea027b),
	.w2(32'h3c05fb64),
	.w3(32'h3bb72b42),
	.w4(32'h3b241750),
	.w5(32'h3be3ca26),
	.w6(32'h3c76bd3b),
	.w7(32'h3bf5d40a),
	.w8(32'h3c067d1f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa90ab),
	.w1(32'hbab17ea1),
	.w2(32'h3b49722d),
	.w3(32'h3c0dea15),
	.w4(32'hbb4f1670),
	.w5(32'hbaac9446),
	.w6(32'h39d4151b),
	.w7(32'h3ba54e3d),
	.w8(32'h3bf352c7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3e488),
	.w1(32'h3c0b45d0),
	.w2(32'h3cc1b007),
	.w3(32'h3b02b1cd),
	.w4(32'h3b81c3f2),
	.w5(32'h3c9d5df4),
	.w6(32'hbaea0c73),
	.w7(32'h3c0ae402),
	.w8(32'h3bb3e476),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9da65c),
	.w1(32'h3bb25cc9),
	.w2(32'h3c5b4ed7),
	.w3(32'h3c33b270),
	.w4(32'h3bdb663f),
	.w5(32'h3c70946f),
	.w6(32'h3b13043e),
	.w7(32'h3c366d46),
	.w8(32'h3c6ac790),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f477f),
	.w1(32'h3c3eda8a),
	.w2(32'h3c485e35),
	.w3(32'h3c036145),
	.w4(32'h3b900093),
	.w5(32'h3bb0e44d),
	.w6(32'h3b835017),
	.w7(32'h3b987d7d),
	.w8(32'h3bb0983a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02af34),
	.w1(32'hbb20f671),
	.w2(32'hba52a23a),
	.w3(32'h3bbb3abd),
	.w4(32'hbb261af9),
	.w5(32'hbb1e3953),
	.w6(32'hbb3db603),
	.w7(32'hbaed5ec5),
	.w8(32'hbb0eb4a2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad164b0),
	.w1(32'hbbfb6b3b),
	.w2(32'hba93cdda),
	.w3(32'hbb0fb445),
	.w4(32'hbbb84694),
	.w5(32'hbb075e85),
	.w6(32'hbc1c0c8f),
	.w7(32'h3b831a95),
	.w8(32'h3aa601fd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4748),
	.w1(32'hbb107fc9),
	.w2(32'hbb5d346c),
	.w3(32'hbb44ba37),
	.w4(32'hbb00b931),
	.w5(32'hbb1c6013),
	.w6(32'hbb575f71),
	.w7(32'hba0df26d),
	.w8(32'h3c25498a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3e2de),
	.w1(32'h3b8e6436),
	.w2(32'h3c580453),
	.w3(32'h3b3e17ec),
	.w4(32'h3ba4efe9),
	.w5(32'h3c7a9b05),
	.w6(32'h3aca68ea),
	.w7(32'h3c3a8b07),
	.w8(32'h3b80da56),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be516b2),
	.w1(32'hbab2de54),
	.w2(32'hbc61b4be),
	.w3(32'h3c28e16b),
	.w4(32'hba202e24),
	.w5(32'hbc809b9c),
	.w6(32'h3b959e80),
	.w7(32'hbbbd3cc0),
	.w8(32'h3b032b6f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e0cf),
	.w1(32'hbb07afae),
	.w2(32'hbbef7a43),
	.w3(32'hbc12613b),
	.w4(32'hbadf84c2),
	.w5(32'hbbc46b36),
	.w6(32'hb89461ee),
	.w7(32'hbba8cd0c),
	.w8(32'hbb1ab6da),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4cab),
	.w1(32'hbbcd50dc),
	.w2(32'hbc38918b),
	.w3(32'hbb94ef13),
	.w4(32'hb9f55388),
	.w5(32'hbbad3afc),
	.w6(32'hbb82f02c),
	.w7(32'hbb23f932),
	.w8(32'hbb0190ff),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfafce7),
	.w1(32'h3bf23388),
	.w2(32'h3c179561),
	.w3(32'hbbab570d),
	.w4(32'h3adba428),
	.w5(32'hba711494),
	.w6(32'h3c02a9ea),
	.w7(32'h3c024898),
	.w8(32'h3c010e7a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7890bf),
	.w1(32'h3bc644d4),
	.w2(32'hba2f8e52),
	.w3(32'h3bd76516),
	.w4(32'h3b2a73af),
	.w5(32'hbaf10d4f),
	.w6(32'h3c174c4a),
	.w7(32'h3ba49b4d),
	.w8(32'h3b52fcd1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1248fe),
	.w1(32'h3c0e09d1),
	.w2(32'h3a28ee3c),
	.w3(32'h3b894cad),
	.w4(32'h3a832579),
	.w5(32'hbb4b14a6),
	.w6(32'h3b9de806),
	.w7(32'h3ae2cec3),
	.w8(32'h3bd1b377),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af61e1e),
	.w1(32'hbb4ee438),
	.w2(32'h3b533976),
	.w3(32'h3ab223bf),
	.w4(32'hba83bad5),
	.w5(32'h3b9caa86),
	.w6(32'hbb43fb17),
	.w7(32'h3b08e555),
	.w8(32'hbb323178),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32e7e4),
	.w1(32'h3bfe2deb),
	.w2(32'h3b6230ee),
	.w3(32'h3a0ea74d),
	.w4(32'h3b2edb90),
	.w5(32'h3b509278),
	.w6(32'h3c06879b),
	.w7(32'h3ba24982),
	.w8(32'h3a299c6e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2347a5),
	.w1(32'hbbaa187f),
	.w2(32'h3c19b797),
	.w3(32'h3a444152),
	.w4(32'hbbced502),
	.w5(32'h3c21dd15),
	.w6(32'hbc28eed8),
	.w7(32'hbae54778),
	.w8(32'hbb6cffe5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0271a6),
	.w1(32'hbb80960b),
	.w2(32'hbc2fe46b),
	.w3(32'h3bbc8a2b),
	.w4(32'hbc27def2),
	.w5(32'hbc2afa14),
	.w6(32'hbb20cd72),
	.w7(32'hbc15503d),
	.w8(32'hbc3828e3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324f17),
	.w1(32'hbad8c7aa),
	.w2(32'hbbc8d933),
	.w3(32'hbc7b2c26),
	.w4(32'h3b76983d),
	.w5(32'hbb9c33e0),
	.w6(32'hbc2e7285),
	.w7(32'hbc85ee88),
	.w8(32'h3b0a7249),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2306a4),
	.w1(32'h3baf71e4),
	.w2(32'h3c1c1d96),
	.w3(32'hbb8f6885),
	.w4(32'h3b1b7e28),
	.w5(32'h3c342ce1),
	.w6(32'h3bb48bbf),
	.w7(32'h3b8c460c),
	.w8(32'h3b19d28c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cdc8c),
	.w1(32'hbb728571),
	.w2(32'hbba26ec1),
	.w3(32'h3b8fd26c),
	.w4(32'hbba74cf8),
	.w5(32'hbb8666aa),
	.w6(32'hba868e5e),
	.w7(32'hbbd36825),
	.w8(32'hbb8a6170),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c81ae),
	.w1(32'hb9b350fb),
	.w2(32'h3a6d1aec),
	.w3(32'hbb2244d9),
	.w4(32'hbafe6307),
	.w5(32'hba5f333c),
	.w6(32'hbb054390),
	.w7(32'hb9965fa0),
	.w8(32'h3b7ea7f0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8349e6),
	.w1(32'h3b21d1d3),
	.w2(32'h3b15b4b3),
	.w3(32'hb81769bf),
	.w4(32'h39c73367),
	.w5(32'h3b9698be),
	.w6(32'hb9927a8f),
	.w7(32'h3a6608ee),
	.w8(32'h3a7024b7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48046d),
	.w1(32'h3b2e04b0),
	.w2(32'h3aa2ab78),
	.w3(32'h3b2b4055),
	.w4(32'h3bb15451),
	.w5(32'h3b4dd6f9),
	.w6(32'h3a778fa5),
	.w7(32'h39ae0c94),
	.w8(32'hba488b48),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6fb93),
	.w1(32'hbc146345),
	.w2(32'hbc07918b),
	.w3(32'h3b9d2be6),
	.w4(32'hbb8c962c),
	.w5(32'hbbf1e2c4),
	.w6(32'hbbc1a77a),
	.w7(32'h3b6b3c37),
	.w8(32'h3b91eda9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258bbb),
	.w1(32'h3b2aae46),
	.w2(32'h3be8d79f),
	.w3(32'hbb1f3e25),
	.w4(32'hbb9dc850),
	.w5(32'hba492a42),
	.w6(32'h3accb0c9),
	.w7(32'h3c07caea),
	.w8(32'h3c1e952c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cd34f),
	.w1(32'h3b9815af),
	.w2(32'h3cb16b81),
	.w3(32'h3b0519a1),
	.w4(32'hbb0b03c9),
	.w5(32'h3c31f341),
	.w6(32'h3983bb81),
	.w7(32'h3c76a9eb),
	.w8(32'h3c3d5ed8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c971983),
	.w1(32'hbb8bf577),
	.w2(32'hbba1c710),
	.w3(32'h3c21a255),
	.w4(32'hbac946bc),
	.w5(32'hbb28abb6),
	.w6(32'hbb426d3a),
	.w7(32'hbb87a0e1),
	.w8(32'hbb13d8d4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63ea89),
	.w1(32'hb92f4fc6),
	.w2(32'h3c1b3b5e),
	.w3(32'hbad922f9),
	.w4(32'hbaae4995),
	.w5(32'h3bda2ddb),
	.w6(32'hbbc92a42),
	.w7(32'hb91790be),
	.w8(32'hbb873fa3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f6434),
	.w1(32'h3c208372),
	.w2(32'h3c2f2c5e),
	.w3(32'h39bfd148),
	.w4(32'h3c320652),
	.w5(32'h3bff11b3),
	.w6(32'h3c1b4c2e),
	.w7(32'h3c21047b),
	.w8(32'h3bda2cef),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c226186),
	.w1(32'hbcd7e43f),
	.w2(32'hbd26d57c),
	.w3(32'h3bfc7a8d),
	.w4(32'hbc2cc763),
	.w5(32'hbcb2408d),
	.w6(32'hbc95436c),
	.w7(32'hbc9a6699),
	.w8(32'hbcb8627a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce906a9),
	.w1(32'hbc3b6751),
	.w2(32'hbcc65bf5),
	.w3(32'hbbae89d4),
	.w4(32'hbc088402),
	.w5(32'hbc5b84c4),
	.w6(32'hbbbd8d0c),
	.w7(32'hbc67fc0a),
	.w8(32'hbc3be1b3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc802efa),
	.w1(32'h3b679903),
	.w2(32'h3ad7b658),
	.w3(32'hbc14cbfe),
	.w4(32'hbb862d0e),
	.w5(32'h3bc788dc),
	.w6(32'h39f305a0),
	.w7(32'h3b36b8fe),
	.w8(32'h3bea54b5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba96e6f),
	.w1(32'hbbceabea),
	.w2(32'hbc896487),
	.w3(32'h3bc0abb0),
	.w4(32'hbc4140ca),
	.w5(32'hbc60d644),
	.w6(32'h3b6a12df),
	.w7(32'hbc0370fc),
	.w8(32'hbc1d14db),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2669b2),
	.w1(32'h3b9d0151),
	.w2(32'h3be87d66),
	.w3(32'hbafeb7bc),
	.w4(32'h3b9c84f2),
	.w5(32'h3bc8128f),
	.w6(32'h3a203afa),
	.w7(32'h3ab31f0a),
	.w8(32'h3ac2a4a7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2536ec),
	.w1(32'h3bb3b599),
	.w2(32'h3c009b18),
	.w3(32'hba89ccf7),
	.w4(32'h3c245fda),
	.w5(32'h3b1a634c),
	.w6(32'h3c0eef1f),
	.w7(32'h3c409970),
	.w8(32'h3c253ee7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2177b4),
	.w1(32'h3bbbad2e),
	.w2(32'h3bdca415),
	.w3(32'h3b618a9f),
	.w4(32'h3b0ee204),
	.w5(32'h3b954ec1),
	.w6(32'h3c8e267c),
	.w7(32'h3c65ed8f),
	.w8(32'h3c923929),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe3206),
	.w1(32'h3abeb188),
	.w2(32'hbb4e37a4),
	.w3(32'h3c2bb14c),
	.w4(32'h3b821fe7),
	.w5(32'hbb4009ae),
	.w6(32'h3b29e11b),
	.w7(32'hbb1e425d),
	.w8(32'h3b436b39),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad00eaa),
	.w1(32'hba8be6ee),
	.w2(32'h39f952ce),
	.w3(32'h3b02acc9),
	.w4(32'hbb98cc21),
	.w5(32'h3af03555),
	.w6(32'h3b31b92b),
	.w7(32'hb9bc39a9),
	.w8(32'hbb0edf4d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2286c2),
	.w1(32'h3bf31dc2),
	.w2(32'h3b0780a1),
	.w3(32'h3c162634),
	.w4(32'h3be00f5e),
	.w5(32'h3b5d4b60),
	.w6(32'h3854f286),
	.w7(32'hbac1e3b6),
	.w8(32'hbbd930db),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81898d),
	.w1(32'h3a6b94b3),
	.w2(32'h39ad00c6),
	.w3(32'h399f18dc),
	.w4(32'hbac82f4d),
	.w5(32'hbac5eff1),
	.w6(32'h3bbe0308),
	.w7(32'hb90802a8),
	.w8(32'h3b66ba79),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d100c),
	.w1(32'hbb1cc719),
	.w2(32'h3b56e157),
	.w3(32'h3ba1c9d0),
	.w4(32'hba5943d5),
	.w5(32'h3b004487),
	.w6(32'hba3082e2),
	.w7(32'h3b58a792),
	.w8(32'h3bca9f39),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0229b),
	.w1(32'hbad5b8e6),
	.w2(32'hbbdd0585),
	.w3(32'h3ba9085c),
	.w4(32'h3b57a462),
	.w5(32'hbba4eab5),
	.w6(32'hbbc24e97),
	.w7(32'hbba9c220),
	.w8(32'h3adf3335),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f3122),
	.w1(32'h3b3d76d5),
	.w2(32'hbab1461a),
	.w3(32'hbc22829b),
	.w4(32'h3bfbdeb3),
	.w5(32'h3c156a26),
	.w6(32'hb9693ec3),
	.w7(32'h3b60e780),
	.w8(32'h39d1a5b4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b826e11),
	.w1(32'hbc17cc40),
	.w2(32'hbc6c5b53),
	.w3(32'h3ba1c5d7),
	.w4(32'hbb12a454),
	.w5(32'hbb95eb3e),
	.w6(32'hbbbfdf0e),
	.w7(32'hbc057404),
	.w8(32'h3a9a0355),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca1831),
	.w1(32'h3c0f71a3),
	.w2(32'h3c232e2a),
	.w3(32'hbb4b7e50),
	.w4(32'h3bd24297),
	.w5(32'h3b6a6449),
	.w6(32'hbab66c24),
	.w7(32'h3bcd8d5d),
	.w8(32'h3bea64e8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd07d77),
	.w1(32'hbb5773a6),
	.w2(32'hbc34e00c),
	.w3(32'h3bce05f2),
	.w4(32'hbb3e6267),
	.w5(32'hbc0092d5),
	.w6(32'hbb133af0),
	.w7(32'hbc4e5dd9),
	.w8(32'hbc03d4f1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc233b6),
	.w1(32'hb9f2ab51),
	.w2(32'hbc999383),
	.w3(32'hbbe6b465),
	.w4(32'hbc344207),
	.w5(32'hbc5c5e0f),
	.w6(32'h3a91f788),
	.w7(32'hbc148312),
	.w8(32'hbc05a720),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6621e),
	.w1(32'hbc865f7d),
	.w2(32'hbc87de15),
	.w3(32'hbb17b1ec),
	.w4(32'h3af64bc9),
	.w5(32'hbc119c81),
	.w6(32'hbc65014d),
	.w7(32'hbc59b9ee),
	.w8(32'h3b04ffbf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc276fcc),
	.w1(32'hbb7f95cc),
	.w2(32'hbc588380),
	.w3(32'hbc197222),
	.w4(32'hbb982475),
	.w5(32'hbc35d0ee),
	.w6(32'h3b3eeab4),
	.w7(32'h3b1b7bf5),
	.w8(32'hbc04b3ba),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e2b0d),
	.w1(32'h3b2a03ef),
	.w2(32'h39ccff0b),
	.w3(32'h397fa7a6),
	.w4(32'h3bf3676b),
	.w5(32'h3bddf7c5),
	.w6(32'hb988efbe),
	.w7(32'hbae7d79c),
	.w8(32'hb7ab78e0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1486a),
	.w1(32'hbb33e389),
	.w2(32'hbbec7054),
	.w3(32'h3b8480eb),
	.w4(32'hbbc39cfb),
	.w5(32'hbbc53c67),
	.w6(32'h39e5e41b),
	.w7(32'hba92a0fd),
	.w8(32'hba615e20),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00afef),
	.w1(32'hbab8301c),
	.w2(32'hbb5a1bb9),
	.w3(32'hbbf2b5d6),
	.w4(32'h38102eb7),
	.w5(32'hbb175c54),
	.w6(32'h3b0f386d),
	.w7(32'hbb0ae138),
	.w8(32'hbae9c326),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba412405),
	.w1(32'hbc8037cc),
	.w2(32'hbc99341a),
	.w3(32'hba46cace),
	.w4(32'hbb86b522),
	.w5(32'hbb5b3812),
	.w6(32'h3b0285bd),
	.w7(32'hbc266df1),
	.w8(32'hbc220c76),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83d7bc),
	.w1(32'h3c0be864),
	.w2(32'h3b636eda),
	.w3(32'h3ba01343),
	.w4(32'h3c10a991),
	.w5(32'h3b98da8e),
	.w6(32'h3c2f16d5),
	.w7(32'h3c290d2e),
	.w8(32'h3bfb1d58),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c406d6d),
	.w1(32'h3c6ccce7),
	.w2(32'h3c6b9237),
	.w3(32'h3bf59508),
	.w4(32'h3bb2080c),
	.w5(32'h3c5ca033),
	.w6(32'h3c13a8c1),
	.w7(32'h3c19f11c),
	.w8(32'h3b62afb6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c0686),
	.w1(32'h3a62f7ff),
	.w2(32'hbb15a546),
	.w3(32'h3c597faa),
	.w4(32'h3aefa7f6),
	.w5(32'hba9e969e),
	.w6(32'h3adf0e39),
	.w7(32'h3913d554),
	.w8(32'h3a0d3284),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bbe8b),
	.w1(32'hbb08a27d),
	.w2(32'hbb9c3cce),
	.w3(32'h370c1b0a),
	.w4(32'hba67923a),
	.w5(32'hbadf34f2),
	.w6(32'hba847d91),
	.w7(32'hba9e5fd3),
	.w8(32'hbabc6512),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b043d),
	.w1(32'h3bdd563c),
	.w2(32'hbc37b5d3),
	.w3(32'hba669cdd),
	.w4(32'hbbecb006),
	.w5(32'hbc425955),
	.w6(32'h3b9b1192),
	.w7(32'hbc67fa4d),
	.w8(32'hbaaee35d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a26b5),
	.w1(32'h39d62e84),
	.w2(32'h3bb7a50c),
	.w3(32'h3a298552),
	.w4(32'h3b24276d),
	.w5(32'h3bc65ff5),
	.w6(32'h3aefbc1b),
	.w7(32'h3b68c1d9),
	.w8(32'h3be48974),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce5038),
	.w1(32'hbc467287),
	.w2(32'hbbf3e8d3),
	.w3(32'h3bb60690),
	.w4(32'hbc4ae765),
	.w5(32'h3aa86403),
	.w6(32'h3a85d419),
	.w7(32'hbc2d0fa5),
	.w8(32'hbbf316fc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3582b7),
	.w1(32'h3c02fda8),
	.w2(32'h3c4b43ca),
	.w3(32'h3c054ba6),
	.w4(32'h3be031e0),
	.w5(32'h3c002e73),
	.w6(32'h3bace384),
	.w7(32'h3c395b44),
	.w8(32'h3be582d0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6d36f),
	.w1(32'h3c5f7d88),
	.w2(32'h3c718baf),
	.w3(32'h3bffa18e),
	.w4(32'h3c5cb29c),
	.w5(32'h3c8df9ec),
	.w6(32'h3c46e8da),
	.w7(32'h3c53feca),
	.w8(32'h3bae1691),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095f40),
	.w1(32'hbb7dc93c),
	.w2(32'hbc28f469),
	.w3(32'h3c7208c4),
	.w4(32'h3c1246c7),
	.w5(32'hbbaea73c),
	.w6(32'hbc04b94e),
	.w7(32'hbb334bbc),
	.w8(32'hba5d4149),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8eead),
	.w1(32'hbc542556),
	.w2(32'hbc8a3ac9),
	.w3(32'hbc3774fe),
	.w4(32'h3b05bb0c),
	.w5(32'hbc23ee77),
	.w6(32'hbc723793),
	.w7(32'hbc26a309),
	.w8(32'hbc7fd2a4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3edb37),
	.w1(32'hbc15a446),
	.w2(32'hbc39556f),
	.w3(32'hbc7dec84),
	.w4(32'hbc74583b),
	.w5(32'hbc68b20d),
	.w6(32'hbc29e0d6),
	.w7(32'hbc5ae459),
	.w8(32'hbc11a810),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dd99d),
	.w1(32'h3c874d69),
	.w2(32'h3c4375ed),
	.w3(32'hbc842b1f),
	.w4(32'h3c05837c),
	.w5(32'h3c239fd7),
	.w6(32'h3bee7d13),
	.w7(32'h3ba0e740),
	.w8(32'h3c4f428d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11bf3c),
	.w1(32'hbc73b496),
	.w2(32'hbc089cca),
	.w3(32'h3be2b760),
	.w4(32'hbbb67e29),
	.w5(32'h3a558b61),
	.w6(32'hbc0c109b),
	.w7(32'hbc4308fc),
	.w8(32'hbc217428),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74502e),
	.w1(32'hbb5d66e9),
	.w2(32'hbbff4eae),
	.w3(32'hbbb33bd4),
	.w4(32'h39b665ab),
	.w5(32'hbb7e2265),
	.w6(32'hbb853932),
	.w7(32'hbb00b67f),
	.w8(32'hbbdb8e08),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68129b),
	.w1(32'hbbbf7559),
	.w2(32'h39baf0fe),
	.w3(32'hbafba559),
	.w4(32'hbb62d264),
	.w5(32'h38a5c022),
	.w6(32'hbbf2c6ea),
	.w7(32'hbc093da1),
	.w8(32'hbc26ea90),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e30674),
	.w1(32'hbbe1c6b3),
	.w2(32'hbbad0de9),
	.w3(32'hbb0f831e),
	.w4(32'hbb4fd8b2),
	.w5(32'hbadace11),
	.w6(32'hbb8c0e80),
	.w7(32'hbbf1cb30),
	.w8(32'hbbd1d8a2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915f850),
	.w1(32'hbbaf87cb),
	.w2(32'hbb665320),
	.w3(32'h3b5c124e),
	.w4(32'hbab065b0),
	.w5(32'hbb8faa88),
	.w6(32'hbbc88207),
	.w7(32'hba690e09),
	.w8(32'h3c02cf6b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d5f77),
	.w1(32'hb9f36d64),
	.w2(32'h3c15e611),
	.w3(32'hbbf4ba7a),
	.w4(32'hbb97799f),
	.w5(32'hbb1a251b),
	.w6(32'hbc052526),
	.w7(32'h3b7f9a96),
	.w8(32'h3a12c983),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62a703),
	.w1(32'h3b1a14a7),
	.w2(32'h3c0cfd59),
	.w3(32'hbbb8553c),
	.w4(32'h3a9b4a39),
	.w5(32'h3c13c40a),
	.w6(32'h3a6c23ac),
	.w7(32'h3bd69976),
	.w8(32'h3b7b8d41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedb39a),
	.w1(32'h3b6cdc5f),
	.w2(32'h3ba70f3e),
	.w3(32'h3bddf28d),
	.w4(32'h3c21da6a),
	.w5(32'h3bf895b0),
	.w6(32'hb8eaa117),
	.w7(32'h3bfa0437),
	.w8(32'h3c2e07cc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced0de),
	.w1(32'hbbe4e36b),
	.w2(32'hbbf0f4c9),
	.w3(32'h3b89e1f7),
	.w4(32'hbba3b984),
	.w5(32'hbc0abb96),
	.w6(32'hbb5e9398),
	.w7(32'hbbbd706a),
	.w8(32'hbbd8fd1a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f709),
	.w1(32'hbb228a5e),
	.w2(32'h3b238d1f),
	.w3(32'hbc0b54e1),
	.w4(32'hbbbbd911),
	.w5(32'hbb2481ba),
	.w6(32'hbc085392),
	.w7(32'hbb51a330),
	.w8(32'hbb210932),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2254),
	.w1(32'hbc16749d),
	.w2(32'hbc78fe1e),
	.w3(32'hbc18baa0),
	.w4(32'hb9e51fe1),
	.w5(32'hbb29d553),
	.w6(32'hbc005886),
	.w7(32'hbc5ad7dc),
	.w8(32'hbc2c23e2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb4b6),
	.w1(32'h3ad07a08),
	.w2(32'h3b1f5213),
	.w3(32'h3abc205c),
	.w4(32'h3b1df211),
	.w5(32'hba9c8063),
	.w6(32'h3a4bdbe4),
	.w7(32'h3b5e080e),
	.w8(32'h3b9b71dc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982adcc),
	.w1(32'h3b702592),
	.w2(32'h3c4c493f),
	.w3(32'hbbb36de0),
	.w4(32'h3b03fe90),
	.w5(32'h3c3a7d48),
	.w6(32'h3853d351),
	.w7(32'h3bdef0fa),
	.w8(32'h3b841756),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c134c7d),
	.w1(32'h3b8e2c8e),
	.w2(32'h3becfdbe),
	.w3(32'h3bf31c8e),
	.w4(32'hbb545d3a),
	.w5(32'hb9a65bc0),
	.w6(32'hbb639cbf),
	.w7(32'h3b019263),
	.w8(32'h3b98344e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc06a65),
	.w1(32'hbb0480f5),
	.w2(32'h3a4b9421),
	.w3(32'hbacab3bc),
	.w4(32'hbbab4df7),
	.w5(32'hbb4480d7),
	.w6(32'hbbd6006d),
	.w7(32'hba67cea6),
	.w8(32'hbbdf6e1f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe72215),
	.w1(32'h3b09aeb2),
	.w2(32'hbbf18537),
	.w3(32'hbb4926d5),
	.w4(32'hba8466e9),
	.w5(32'hbb664e50),
	.w6(32'hbb38fcbd),
	.w7(32'hbbd035bd),
	.w8(32'hbbc39424),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb39e8f),
	.w1(32'h3ad5fdd3),
	.w2(32'h3b9c5e53),
	.w3(32'hbbd4a5fe),
	.w4(32'h3b1b42a5),
	.w5(32'h3bc74df3),
	.w6(32'h3b3d108c),
	.w7(32'h3b7c63aa),
	.w8(32'h3b83ddb8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf42912),
	.w1(32'h3c140d0f),
	.w2(32'h3be13556),
	.w3(32'h3c285c43),
	.w4(32'h3b81a17b),
	.w5(32'h3c0edc3f),
	.w6(32'h3bd66903),
	.w7(32'h3b995642),
	.w8(32'h3b9cb221),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b915eb7),
	.w1(32'h3b7ce61c),
	.w2(32'h3a85f10b),
	.w3(32'h3c0a216d),
	.w4(32'h3c066cc0),
	.w5(32'h3b84fdd7),
	.w6(32'h3bccc3ca),
	.w7(32'h3bdf3ab2),
	.w8(32'h3a4a1ce5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38153db3),
	.w1(32'hb9b0a3c8),
	.w2(32'hbb7f3b28),
	.w3(32'h3b247d68),
	.w4(32'hba3bfa54),
	.w5(32'hbb2468eb),
	.w6(32'h3a746ff9),
	.w7(32'h3a33729b),
	.w8(32'h3a7b8bd2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea788),
	.w1(32'h3a85d6cb),
	.w2(32'hbabc5061),
	.w3(32'hbafe5d39),
	.w4(32'hba2a5408),
	.w5(32'hbb267197),
	.w6(32'hba9b7f88),
	.w7(32'h3814d37d),
	.w8(32'hbb9bfe4a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00e777),
	.w1(32'h3ac7294e),
	.w2(32'hbc1ad581),
	.w3(32'h3b973783),
	.w4(32'h3c063704),
	.w5(32'h3b84e06a),
	.w6(32'hbc3b53ef),
	.w7(32'hbc4442d0),
	.w8(32'h3ae98c41),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39353462),
	.w1(32'h3b8b5fa1),
	.w2(32'h3b97f215),
	.w3(32'hbb11bfa2),
	.w4(32'h3ab85cef),
	.w5(32'hba234dd2),
	.w6(32'h3be4ae51),
	.w7(32'h3bf8e0c7),
	.w8(32'h3ae0973f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c125ffd),
	.w1(32'hbace1d02),
	.w2(32'hbb6563dd),
	.w3(32'h3bc8a51d),
	.w4(32'h372bf03e),
	.w5(32'hbae575db),
	.w6(32'h3961819a),
	.w7(32'hbac40b6d),
	.w8(32'h3a7e3f0f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac57779),
	.w1(32'h3c2acf31),
	.w2(32'hbb359cb5),
	.w3(32'h3a055052),
	.w4(32'h3bb06431),
	.w5(32'hbbafbfa9),
	.w6(32'h3c90e8cf),
	.w7(32'h3b9d5f61),
	.w8(32'hba026325),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule