module layer_8_featuremap_143(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cfdcf),
	.w1(32'hbb3d7a3c),
	.w2(32'h3bad569f),
	.w3(32'hbbc659af),
	.w4(32'h3c76bd6a),
	.w5(32'hbc35c44a),
	.w6(32'hbbc33141),
	.w7(32'h3ca2ae2b),
	.w8(32'hbc8f0487),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd72d8d),
	.w1(32'h3c8e0188),
	.w2(32'hbc432a24),
	.w3(32'h3c49e58b),
	.w4(32'hbc2ce3fa),
	.w5(32'hbc55b51c),
	.w6(32'h3ccbf96a),
	.w7(32'hbafd1f0c),
	.w8(32'h3cdf42cd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd464b),
	.w1(32'hbca5f83e),
	.w2(32'h3baf7e56),
	.w3(32'hbc6c8e42),
	.w4(32'h3c017eb3),
	.w5(32'h3c398a2f),
	.w6(32'hb957b93f),
	.w7(32'h3c113e19),
	.w8(32'hbbe71a27),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeb650),
	.w1(32'hbb553d8a),
	.w2(32'h3c29edf4),
	.w3(32'hbc0bf48f),
	.w4(32'h3b184ea3),
	.w5(32'h3b1d25ca),
	.w6(32'hbd091044),
	.w7(32'hbc10ebc6),
	.w8(32'hbcb13f58),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66ea47),
	.w1(32'h3c529d04),
	.w2(32'h394199e1),
	.w3(32'h3cef3d86),
	.w4(32'h3b3b62e8),
	.w5(32'h3c1b5e78),
	.w6(32'h3cbcf24e),
	.w7(32'hbb26fdcf),
	.w8(32'hbb38dd79),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148b5a),
	.w1(32'h3b80a77c),
	.w2(32'hbcaa2b69),
	.w3(32'h3a0cb933),
	.w4(32'h3b0d2adb),
	.w5(32'h3bcf6573),
	.w6(32'hbc60a2e1),
	.w7(32'hbc704be5),
	.w8(32'h3d72ad6c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9371cc),
	.w1(32'hbc01eb71),
	.w2(32'h3c5a592c),
	.w3(32'hbcb50c37),
	.w4(32'h3c47d258),
	.w5(32'h3a533a27),
	.w6(32'h3bd1dfa3),
	.w7(32'h3bd7ea6b),
	.w8(32'hba903e6a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82585a),
	.w1(32'h3c631e19),
	.w2(32'h3ada0f54),
	.w3(32'h3c922539),
	.w4(32'h3cb15be6),
	.w5(32'h3be51794),
	.w6(32'h3bcba9dc),
	.w7(32'h3a971158),
	.w8(32'h3ccc82e6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16f530),
	.w1(32'h3c42c21c),
	.w2(32'h3a8e1f1b),
	.w3(32'hbc2ecd4c),
	.w4(32'hbc140665),
	.w5(32'hbb89db38),
	.w6(32'h3b51ac68),
	.w7(32'h3b503406),
	.w8(32'hbc3dc126),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e34141),
	.w1(32'h3c4cbfca),
	.w2(32'h3c2eff85),
	.w3(32'h3b924ecb),
	.w4(32'hbbfbc362),
	.w5(32'h3b90003f),
	.w6(32'h3c23e07f),
	.w7(32'h3c0d8e56),
	.w8(32'h3cfee2d3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf3f4b),
	.w1(32'hbc574f84),
	.w2(32'h3bb61235),
	.w3(32'hbb81ddb2),
	.w4(32'h3b9d31b4),
	.w5(32'h3b4f0c6c),
	.w6(32'hbcf00c04),
	.w7(32'h3b6992b5),
	.w8(32'hbc7f1500),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f029a),
	.w1(32'h3a9e539c),
	.w2(32'h3c1cf6bd),
	.w3(32'h3bb879f2),
	.w4(32'hbacb44a6),
	.w5(32'h3cc9ca0f),
	.w6(32'h3c7f5729),
	.w7(32'hbc4dbc85),
	.w8(32'h3cfaa797),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00b62e),
	.w1(32'h3ca534b9),
	.w2(32'hba126ba3),
	.w3(32'h3a99d8e5),
	.w4(32'h3b796605),
	.w5(32'h3bfef3a6),
	.w6(32'h3cd22f13),
	.w7(32'h3adeedc9),
	.w8(32'h3b4510c6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b940215),
	.w1(32'h3bd1a616),
	.w2(32'hbb1490d7),
	.w3(32'h3b21f98d),
	.w4(32'hb9601d8a),
	.w5(32'h3b2179a7),
	.w6(32'h3baedcd1),
	.w7(32'hbb753d04),
	.w8(32'h3b6af68e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a342e),
	.w1(32'h3bd4aa14),
	.w2(32'hbb6f7755),
	.w3(32'h3b4da785),
	.w4(32'hbaf3ec94),
	.w5(32'h3b6adbed),
	.w6(32'h3b3d8193),
	.w7(32'hbbb6062f),
	.w8(32'h3b08b880),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77d809),
	.w1(32'h3bc8c186),
	.w2(32'hbbb7258a),
	.w3(32'h3ba168f4),
	.w4(32'h3b2f5a90),
	.w5(32'h3b16ec94),
	.w6(32'h3b7647a5),
	.w7(32'hba3059af),
	.w8(32'hbb55f434),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd49fd),
	.w1(32'hbbb0e1b7),
	.w2(32'hbb99ba84),
	.w3(32'h3c8db414),
	.w4(32'hbc31763b),
	.w5(32'h3af50948),
	.w6(32'h3b8f3447),
	.w7(32'hbabec84c),
	.w8(32'h3bffd277),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7797f),
	.w1(32'hbc242483),
	.w2(32'hbc6bdc59),
	.w3(32'hbce7750a),
	.w4(32'hbb1f6e0b),
	.w5(32'hba7c77ad),
	.w6(32'hbc172e93),
	.w7(32'hbc3dc7b4),
	.w8(32'h3c243a6d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11d7c6),
	.w1(32'h3c3ce580),
	.w2(32'hbc4ee509),
	.w3(32'hbbb0b79d),
	.w4(32'hbc269427),
	.w5(32'h3b82a8df),
	.w6(32'h3aa7bb3c),
	.w7(32'hbc8ec50d),
	.w8(32'h3b0d28d6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8f2c),
	.w1(32'hbbc9f901),
	.w2(32'h3c8fca67),
	.w3(32'hbaca030d),
	.w4(32'h3bdcc5e4),
	.w5(32'hbc5f8b1a),
	.w6(32'hbc0fa634),
	.w7(32'h3c211270),
	.w8(32'hbcd76fbd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47cb2f),
	.w1(32'h3bc792c3),
	.w2(32'hbb49f53c),
	.w3(32'hba9cf4f9),
	.w4(32'hbc4ad317),
	.w5(32'h3cec0541),
	.w6(32'h3bfcb950),
	.w7(32'hbc94182a),
	.w8(32'h3bf9114c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40a6d0),
	.w1(32'h3bfa9f7f),
	.w2(32'h3bc0b560),
	.w3(32'hbc5a4419),
	.w4(32'h3bcc4590),
	.w5(32'hbbc558d8),
	.w6(32'hbbd293d7),
	.w7(32'h3a699156),
	.w8(32'hbc06b3f5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec1290),
	.w1(32'hbc517f58),
	.w2(32'h3a43a039),
	.w3(32'hbbd8ffb0),
	.w4(32'hbb2e6697),
	.w5(32'hbbe3305e),
	.w6(32'hbc7be126),
	.w7(32'hbb7b6918),
	.w8(32'hbc113e15),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57d0f8),
	.w1(32'h3a66be7a),
	.w2(32'h3c0aefc5),
	.w3(32'h3c025084),
	.w4(32'h3c57063e),
	.w5(32'hbc949e97),
	.w6(32'h3c56510a),
	.w7(32'h3c59fc73),
	.w8(32'hbbcfb148),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d15b8),
	.w1(32'h3b774b50),
	.w2(32'hb98e78ac),
	.w3(32'h3b6fc7d4),
	.w4(32'h3ab433f4),
	.w5(32'h3be70169),
	.w6(32'h3be205d2),
	.w7(32'hbb7027bc),
	.w8(32'h3bef6d87),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43208),
	.w1(32'h3ba3049c),
	.w2(32'h3c51c0dd),
	.w3(32'h3b5cef8f),
	.w4(32'h3c1b6059),
	.w5(32'hbc344570),
	.w6(32'h3b3ec8a3),
	.w7(32'h3ac96cd7),
	.w8(32'hbc06bd94),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b2a3e),
	.w1(32'h3ba6e8cd),
	.w2(32'hbb8e9be3),
	.w3(32'h3b53bb14),
	.w4(32'h3b394278),
	.w5(32'h3b67b9e6),
	.w6(32'h3bd1d711),
	.w7(32'h3b673d0e),
	.w8(32'hbb307db1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e677b),
	.w1(32'h3bc05626),
	.w2(32'h3aae4983),
	.w3(32'hbb462884),
	.w4(32'h3c552939),
	.w5(32'hbc6d1eae),
	.w6(32'hbb2953cd),
	.w7(32'h3a85a6fe),
	.w8(32'hbcd0180e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae307e8),
	.w1(32'hbac400dd),
	.w2(32'hbc21a9e7),
	.w3(32'h3b33d07b),
	.w4(32'hbba06fcd),
	.w5(32'hbb3d35c7),
	.w6(32'hbb6969dd),
	.w7(32'hbbeaf8f4),
	.w8(32'hbbb419aa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81eeec),
	.w1(32'h3bb34bb8),
	.w2(32'hbc979459),
	.w3(32'h3c7af26a),
	.w4(32'hbb978407),
	.w5(32'h3ce24437),
	.w6(32'h3c1056e4),
	.w7(32'hbc53e099),
	.w8(32'h3d80b1e0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d16d152),
	.w1(32'hbc21a70e),
	.w2(32'h3bfdcd17),
	.w3(32'hbd05587b),
	.w4(32'h3c14c699),
	.w5(32'h3c4acde0),
	.w6(32'hbce08ebb),
	.w7(32'h3bcf4706),
	.w8(32'h3c3461fa),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c443bad),
	.w1(32'h3c4c8ed5),
	.w2(32'hbc254948),
	.w3(32'h3c58b013),
	.w4(32'h3ae87b3e),
	.w5(32'hbc0ea910),
	.w6(32'h3c44393c),
	.w7(32'hb846d926),
	.w8(32'hbcb39dec),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b01f8),
	.w1(32'hb9905cd1),
	.w2(32'hbc56cbf7),
	.w3(32'hbb94fff8),
	.w4(32'hbb17441c),
	.w5(32'h3c6198f3),
	.w6(32'hbbb339a6),
	.w7(32'hbc796bc2),
	.w8(32'hbbe1b83f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2117e),
	.w1(32'h3c586d4d),
	.w2(32'hbbeaa4df),
	.w3(32'hbc6151b8),
	.w4(32'h3a0d9c01),
	.w5(32'h3cd5f684),
	.w6(32'h3c714041),
	.w7(32'h3b34d6a4),
	.w8(32'h3d8b688b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda9c16),
	.w1(32'hbae9380e),
	.w2(32'hbb65c67a),
	.w3(32'hbc37b425),
	.w4(32'hbbb8f1bd),
	.w5(32'hbb45969f),
	.w6(32'h3c01b576),
	.w7(32'hbbb3363b),
	.w8(32'hbb8f3ffb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1ef2),
	.w1(32'hb9fb4cdf),
	.w2(32'hbc4e752f),
	.w3(32'hbbebd58b),
	.w4(32'hbc4559af),
	.w5(32'h3ce36a20),
	.w6(32'hbb951920),
	.w7(32'hbc90ceed),
	.w8(32'h3ce7a662),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d0bd4),
	.w1(32'hbc2f0127),
	.w2(32'hbb3b0237),
	.w3(32'hbc105f1f),
	.w4(32'hbc15e9c8),
	.w5(32'hbbd96993),
	.w6(32'hbb2df338),
	.w7(32'hbbb95cef),
	.w8(32'hbc1fd604),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68c34f),
	.w1(32'h3b4af923),
	.w2(32'hbc0d553d),
	.w3(32'hbb4c68ac),
	.w4(32'hbc35b9ee),
	.w5(32'hbbf37ad2),
	.w6(32'h3ae3d310),
	.w7(32'h38878504),
	.w8(32'h3c8dc60f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04a371),
	.w1(32'hbbb2ac71),
	.w2(32'hbc6b6a5c),
	.w3(32'h3bd5aec2),
	.w4(32'hbc72479c),
	.w5(32'h373f5766),
	.w6(32'h3bbb7085),
	.w7(32'hbc5e96ff),
	.w8(32'hbc1f82df),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63fcab),
	.w1(32'h3bffce1c),
	.w2(32'hba8f4792),
	.w3(32'h3c3a09ed),
	.w4(32'hba4642db),
	.w5(32'h3ae7cfab),
	.w6(32'h3c07c3c0),
	.w7(32'h3b67c8b6),
	.w8(32'hbba32ba2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe274a0),
	.w1(32'h3b2c256f),
	.w2(32'h3bc99865),
	.w3(32'h3bbf8f95),
	.w4(32'h3b45f80c),
	.w5(32'hbbc16c64),
	.w6(32'h3a50d946),
	.w7(32'h3b7f481e),
	.w8(32'hbc32f12a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3997),
	.w1(32'hbc06a2ef),
	.w2(32'hbc02022f),
	.w3(32'hb9aa8832),
	.w4(32'hbbf1fcd2),
	.w5(32'h3a040351),
	.w6(32'hbc820fc6),
	.w7(32'hbc10d61a),
	.w8(32'hbc6dee19),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f992e),
	.w1(32'h3c16d2a4),
	.w2(32'hbbce37f2),
	.w3(32'hbb9a8c62),
	.w4(32'hbc74db20),
	.w5(32'h3b9573b0),
	.w6(32'h3b68fcdc),
	.w7(32'hbba89448),
	.w8(32'h3c5abc42),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70c03d),
	.w1(32'h3c1b85a5),
	.w2(32'hbabf49c7),
	.w3(32'h3a6df091),
	.w4(32'h3b32596b),
	.w5(32'h3bf80e01),
	.w6(32'hbad65e6f),
	.w7(32'h3a4f1585),
	.w8(32'h3bbf6ced),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19065f),
	.w1(32'h3c07b819),
	.w2(32'hbb40e7f4),
	.w3(32'h3a944862),
	.w4(32'h3a0ea4cc),
	.w5(32'h3c8f4dbf),
	.w6(32'h3bd9d358),
	.w7(32'hbbd06f23),
	.w8(32'hbbce330e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ebd50),
	.w1(32'hbc1c13de),
	.w2(32'h3c5ce43b),
	.w3(32'hbb4526ab),
	.w4(32'h3be04130),
	.w5(32'hbd079b0a),
	.w6(32'hbc16a8d4),
	.w7(32'h3c4fa4d7),
	.w8(32'hbcb313e4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd2ee),
	.w1(32'hbb8eb308),
	.w2(32'h3b19cc0b),
	.w3(32'h3bbe765c),
	.w4(32'h3c08ac14),
	.w5(32'hba46af72),
	.w6(32'h3b83c6c9),
	.w7(32'h3b7f2eb2),
	.w8(32'hbc66f098),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ec46f),
	.w1(32'h3c5ff302),
	.w2(32'hbc3a0b37),
	.w3(32'hbc225e11),
	.w4(32'h3b5d2840),
	.w5(32'h3c65592f),
	.w6(32'hbb982cce),
	.w7(32'hbb49085c),
	.w8(32'h3c5f44bc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2e337),
	.w1(32'hbc9496d5),
	.w2(32'hbbcbd0d7),
	.w3(32'hbc5cff54),
	.w4(32'hbbba8c6d),
	.w5(32'h3b381b76),
	.w6(32'hbca384ab),
	.w7(32'hbc56469e),
	.w8(32'hbc270b80),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8caa9b),
	.w1(32'h3c763338),
	.w2(32'hbc8b2372),
	.w3(32'h3b5a1352),
	.w4(32'hbc9cedbc),
	.w5(32'hbc7591d8),
	.w6(32'h3c765533),
	.w7(32'hbc733ac7),
	.w8(32'hbc8ee7d3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc864a89),
	.w1(32'hbc882137),
	.w2(32'hbc8050e6),
	.w3(32'hbc625ff1),
	.w4(32'hb96d84d1),
	.w5(32'hbce9191f),
	.w6(32'hbc87b22e),
	.w7(32'hbc013c90),
	.w8(32'h3c051875),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3a589),
	.w1(32'hbc526c4e),
	.w2(32'h3c841cbb),
	.w3(32'h3c5d3e0e),
	.w4(32'h3c35f8fb),
	.w5(32'h382ad3ef),
	.w6(32'h3c18370e),
	.w7(32'h3cc77663),
	.w8(32'hbc15cea5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3741dc),
	.w1(32'hbc0eaef1),
	.w2(32'hb9e18ad4),
	.w3(32'hbc0c19c4),
	.w4(32'h3bf4b1b2),
	.w5(32'hbb39eb83),
	.w6(32'hbbd2388c),
	.w7(32'h3c052737),
	.w8(32'hbb1cdae2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d70d26),
	.w1(32'hbc0711b6),
	.w2(32'hbab2b28a),
	.w3(32'hbc832b0b),
	.w4(32'h3b24a914),
	.w5(32'h3bc507d4),
	.w6(32'hbc90a152),
	.w7(32'hba39e16a),
	.w8(32'h3b832c58),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0166e4),
	.w1(32'h3b7306be),
	.w2(32'hba24b5d6),
	.w3(32'h3af3ecee),
	.w4(32'hbc5384e3),
	.w5(32'h3c36c02f),
	.w6(32'h3b57967b),
	.w7(32'h3b840f66),
	.w8(32'h3c599834),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4de1ad),
	.w1(32'hbba8bb09),
	.w2(32'hbb7a1360),
	.w3(32'hbc0f4322),
	.w4(32'hbc222792),
	.w5(32'hbc8ee7d2),
	.w6(32'hbba17886),
	.w7(32'hbb7a94b9),
	.w8(32'hbc803d45),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2487d5),
	.w1(32'hbcbe84f4),
	.w2(32'h398736b2),
	.w3(32'hbbd01ac5),
	.w4(32'hbbe0e84f),
	.w5(32'h3ac3a952),
	.w6(32'hbc632cfe),
	.w7(32'hbb2d8cbf),
	.w8(32'h3bd25645),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae78b2),
	.w1(32'h3c29c19c),
	.w2(32'h3c03aa1c),
	.w3(32'h3c124d4a),
	.w4(32'h3c0474d1),
	.w5(32'hbcd1927b),
	.w6(32'h3c0f52cc),
	.w7(32'h3aa0631c),
	.w8(32'hbc2ba6bb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37b020),
	.w1(32'hbb229660),
	.w2(32'hbaaa68a1),
	.w3(32'h3c30316b),
	.w4(32'h3b2c7f35),
	.w5(32'h3bf609a6),
	.w6(32'h3b00395e),
	.w7(32'h39231fd9),
	.w8(32'h3bd647b4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b52cb),
	.w1(32'h3bc3fcd3),
	.w2(32'h3cc22277),
	.w3(32'h3aa8a0ce),
	.w4(32'h3c714af7),
	.w5(32'hbd3b5711),
	.w6(32'h3bb70467),
	.w7(32'h3cb37cd7),
	.w8(32'hbd9df750),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd68aae9),
	.w1(32'h3c8ec63b),
	.w2(32'hbc779d8e),
	.w3(32'h3d18cdd5),
	.w4(32'hbbe78f97),
	.w5(32'h3bee4899),
	.w6(32'h3d09a057),
	.w7(32'hbbaffbf4),
	.w8(32'h3d527611),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d584c3c),
	.w1(32'hbcc56561),
	.w2(32'hbc427e27),
	.w3(32'h393ee547),
	.w4(32'hbbe318ee),
	.w5(32'h3b9d5d81),
	.w6(32'hbc926833),
	.w7(32'hbc21a8fe),
	.w8(32'h3aa24951),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca719),
	.w1(32'hbb076cb1),
	.w2(32'h3c4ede81),
	.w3(32'h3b8a81be),
	.w4(32'h3c06f601),
	.w5(32'hbc169bd1),
	.w6(32'h3b1135ce),
	.w7(32'h3c6d739c),
	.w8(32'hbba5bd76),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be21af2),
	.w1(32'hbc20a417),
	.w2(32'h395b8aad),
	.w3(32'hbc0d6520),
	.w4(32'h3a981090),
	.w5(32'hbbbf8b74),
	.w6(32'hbc869a74),
	.w7(32'h3b91a132),
	.w8(32'hbc5a0f34),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da74d3),
	.w1(32'h3c12dfdd),
	.w2(32'h3b88db7f),
	.w3(32'h3c41bdcd),
	.w4(32'h3bc2afb5),
	.w5(32'hbb0b477d),
	.w6(32'h3c45cd2c),
	.w7(32'h3b9e4475),
	.w8(32'h3a933bbb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade5f50),
	.w1(32'h3be3dd3a),
	.w2(32'hbc1149a6),
	.w3(32'h3ba7d85b),
	.w4(32'hbbb5e118),
	.w5(32'hba3840f0),
	.w6(32'h3b83fb3a),
	.w7(32'hbbfb1481),
	.w8(32'h3cb541c3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9805bc),
	.w1(32'hbc605a4e),
	.w2(32'h3bf188b2),
	.w3(32'hbbc59cce),
	.w4(32'h3abfbfd8),
	.w5(32'h38ec256c),
	.w6(32'h3a79e43c),
	.w7(32'h3c168dfd),
	.w8(32'hbafa1076),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee2ab),
	.w1(32'hbb49ae84),
	.w2(32'h3b39313f),
	.w3(32'h3b93262b),
	.w4(32'h3b1ef21f),
	.w5(32'h3b9e2334),
	.w6(32'hbbac611b),
	.w7(32'h3bf6fe3c),
	.w8(32'hbc01ce75),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad45a46),
	.w1(32'hbb8b83a3),
	.w2(32'hba8de3c3),
	.w3(32'hbc9bafdd),
	.w4(32'hbb8df528),
	.w5(32'hbb5206bf),
	.w6(32'hbca0f9de),
	.w7(32'hbb1b744e),
	.w8(32'hbca04e22),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5d3b9),
	.w1(32'hbbc37ecf),
	.w2(32'h3cc7c6cd),
	.w3(32'h3b94f938),
	.w4(32'hbc1bb19e),
	.w5(32'hbb4d510d),
	.w6(32'h3a7e6526),
	.w7(32'hbb82bf6e),
	.w8(32'hbc6f798f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20e7be),
	.w1(32'hbc63e176),
	.w2(32'h3abca645),
	.w3(32'hbb40525b),
	.w4(32'h3a106706),
	.w5(32'h3aebc394),
	.w6(32'hbbefa3ff),
	.w7(32'h3a926c9c),
	.w8(32'hbbf93989),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0d030),
	.w1(32'h3c3b1742),
	.w2(32'hbc4010cd),
	.w3(32'h3c0cc9e3),
	.w4(32'h3bc8d25d),
	.w5(32'h3bd48508),
	.w6(32'h3bc276c7),
	.w7(32'hbc1566a4),
	.w8(32'hbb32cda6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100c30),
	.w1(32'h3a0b3826),
	.w2(32'h3c06e65b),
	.w3(32'h3c37d732),
	.w4(32'h3c1d6e0a),
	.w5(32'hbbf6ae26),
	.w6(32'h3c657972),
	.w7(32'h3c2fcb81),
	.w8(32'hbc50dfdc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02a83),
	.w1(32'h3ae70d9d),
	.w2(32'hbb07b9a1),
	.w3(32'h38f9ba5d),
	.w4(32'h3bfb9d60),
	.w5(32'hbbf6e9c6),
	.w6(32'h3af0dd98),
	.w7(32'h3b060f58),
	.w8(32'hbc0f58c6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8e230),
	.w1(32'h3cd27473),
	.w2(32'h3afbaf49),
	.w3(32'h3b6ca7a0),
	.w4(32'hbaa5f330),
	.w5(32'hbc95417a),
	.w6(32'h3ca2828f),
	.w7(32'h3aa8a5ad),
	.w8(32'hbccce3fc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ce799),
	.w1(32'hbc57aefc),
	.w2(32'h3aaa4e7d),
	.w3(32'hbc825cbc),
	.w4(32'hbc69bd24),
	.w5(32'h3b06bdb3),
	.w6(32'hbc839b6e),
	.w7(32'hbc5d43a5),
	.w8(32'hbb8877ba),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8df903),
	.w1(32'hbca117d6),
	.w2(32'h39ee7b89),
	.w3(32'hbc7abea6),
	.w4(32'h3b3a04c0),
	.w5(32'h3c14ff60),
	.w6(32'hbcb3cdf8),
	.w7(32'hbb41f275),
	.w8(32'hbbb70183),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00f344),
	.w1(32'hb97eb164),
	.w2(32'h39b79dc3),
	.w3(32'h3c91f6e4),
	.w4(32'hbb41b31a),
	.w5(32'h39c9a46e),
	.w6(32'h3a294450),
	.w7(32'hbb64f6dd),
	.w8(32'hbc186705),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5b37e),
	.w1(32'h3b15dac0),
	.w2(32'h3ba7e47c),
	.w3(32'h3b05baee),
	.w4(32'h3b548e3c),
	.w5(32'hbb74543b),
	.w6(32'h3a114157),
	.w7(32'h3b5d2bf3),
	.w8(32'hbbba5371),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512a25),
	.w1(32'h3b4669be),
	.w2(32'hbb68012e),
	.w3(32'hba5df853),
	.w4(32'hbc1af188),
	.w5(32'hbc11bf33),
	.w6(32'hba761a4f),
	.w7(32'hbc3f0020),
	.w8(32'hbc5f39e9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9faaaa1),
	.w1(32'hba2cb9d0),
	.w2(32'h3b21be4b),
	.w3(32'hba01cc29),
	.w4(32'hbbeb6f55),
	.w5(32'hbb0ffe5f),
	.w6(32'hbc1271c8),
	.w7(32'hbc505d56),
	.w8(32'hbb8200a3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897a9c),
	.w1(32'h3c2f740b),
	.w2(32'h3adc86ae),
	.w3(32'h3c8118f0),
	.w4(32'h3c074f60),
	.w5(32'hbb2326d9),
	.w6(32'h3c5c2230),
	.w7(32'h3c0157e6),
	.w8(32'h3b404d41),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea6fd2),
	.w1(32'hbc0328f3),
	.w2(32'h3c012287),
	.w3(32'hb912d260),
	.w4(32'hbbf7ea17),
	.w5(32'hbbe16be7),
	.w6(32'h3b1af3b6),
	.w7(32'hbb2091b0),
	.w8(32'hbac5924f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa944ee),
	.w1(32'h3b2c4748),
	.w2(32'hbc2764b4),
	.w3(32'h3c9bb339),
	.w4(32'hbc80193a),
	.w5(32'hbb49b48d),
	.w6(32'h3cb0fec9),
	.w7(32'h3bc9376e),
	.w8(32'h3c2eb7ba),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1999a),
	.w1(32'hbc43e1d7),
	.w2(32'h3b45c338),
	.w3(32'h3ca04abb),
	.w4(32'h3a773a34),
	.w5(32'hbb88ef4c),
	.w6(32'hbb560ec5),
	.w7(32'hbb974430),
	.w8(32'h3c31bdbd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c974c86),
	.w1(32'h3c98eb2f),
	.w2(32'hbbf789d5),
	.w3(32'hbcf5e2ae),
	.w4(32'h3a1befc6),
	.w5(32'h3c4bb3f6),
	.w6(32'hbc0d6934),
	.w7(32'hbc3efdfc),
	.w8(32'h3b61245e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e658c),
	.w1(32'h3bbd2062),
	.w2(32'hbca8b355),
	.w3(32'h3ba70688),
	.w4(32'hbbd8daa2),
	.w5(32'hbb3a81a7),
	.w6(32'h3d02891e),
	.w7(32'hbbfec1aa),
	.w8(32'h3c85ad64),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6d9ec),
	.w1(32'hbac5fc2f),
	.w2(32'hbc6df76a),
	.w3(32'h3b0153b0),
	.w4(32'hbb70f920),
	.w5(32'h3c4cfbf8),
	.w6(32'hbbd2e2b5),
	.w7(32'hbc1d8e35),
	.w8(32'h3c3d66a0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d38d7),
	.w1(32'h3b819994),
	.w2(32'hbb576cd9),
	.w3(32'h3c620dba),
	.w4(32'hbb9eb422),
	.w5(32'hbba7eea8),
	.w6(32'h3c212a6c),
	.w7(32'hbba51520),
	.w8(32'hbb4897ec),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c47d),
	.w1(32'h3c64e248),
	.w2(32'hbb1f27b2),
	.w3(32'h3b93067c),
	.w4(32'hbc4ec79a),
	.w5(32'hbc9088e4),
	.w6(32'h3af810ff),
	.w7(32'hbbcd6de5),
	.w8(32'h3ae03f06),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b3472),
	.w1(32'h3a13595b),
	.w2(32'h3b617a6b),
	.w3(32'h3c000e5d),
	.w4(32'hbc28677c),
	.w5(32'h3bcf119e),
	.w6(32'hb92c164e),
	.w7(32'hb9c2a6d5),
	.w8(32'hbc4fcb16),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e3282),
	.w1(32'hbcb9c758),
	.w2(32'hbcaca4c0),
	.w3(32'hbbe5a58a),
	.w4(32'hbccd2cc5),
	.w5(32'h3bda9dde),
	.w6(32'hbccec1e7),
	.w7(32'hbcfa9ab7),
	.w8(32'hbb86c14c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc6aac),
	.w1(32'h3c58bdfe),
	.w2(32'hbc379f77),
	.w3(32'h3d0bf8f6),
	.w4(32'h3c226886),
	.w5(32'h3c5ca033),
	.w6(32'h3cec4b9b),
	.w7(32'h3c73e7f5),
	.w8(32'h3c045004),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391219),
	.w1(32'hbc0716e9),
	.w2(32'h3bd002db),
	.w3(32'hbc70f78c),
	.w4(32'hbc008ec9),
	.w5(32'hbbe2c1d1),
	.w6(32'h3ad1a120),
	.w7(32'hbb5817e8),
	.w8(32'h3cdde11a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5787cc),
	.w1(32'h3c206e78),
	.w2(32'h3c2779a9),
	.w3(32'hbc9517fa),
	.w4(32'h3b4380e9),
	.w5(32'h3aa1a2c0),
	.w6(32'hbab0e980),
	.w7(32'h3bc739fc),
	.w8(32'h3b7e7561),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e792),
	.w1(32'h3bb686d6),
	.w2(32'hbc0597ab),
	.w3(32'hbb17a7aa),
	.w4(32'hbbd67a0a),
	.w5(32'hbb69d23b),
	.w6(32'h396037e7),
	.w7(32'hbc524c57),
	.w8(32'hbcf73cd8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc219445),
	.w1(32'h3ad476af),
	.w2(32'h3c1dfac5),
	.w3(32'h3d1af517),
	.w4(32'h3c0cf93a),
	.w5(32'hbc036875),
	.w6(32'h3ba64e94),
	.w7(32'h3c64d82d),
	.w8(32'hbbd16fea),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb258ac5),
	.w1(32'hbc04dd92),
	.w2(32'h3c0db699),
	.w3(32'hbcb58a92),
	.w4(32'h3c25ddd1),
	.w5(32'h3b4f04fb),
	.w6(32'hbcc34ae5),
	.w7(32'h3c0562e3),
	.w8(32'h3c45faa7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c666790),
	.w1(32'hbab8435c),
	.w2(32'h3c3e1bc3),
	.w3(32'hba41daf7),
	.w4(32'h3c459f97),
	.w5(32'h3a9f9888),
	.w6(32'hbcfa8ad2),
	.w7(32'h3c7f70d4),
	.w8(32'h3c7d80f5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60bbc8),
	.w1(32'h3b7a325d),
	.w2(32'h3bf8ec63),
	.w3(32'hbc679366),
	.w4(32'h3c27d46f),
	.w5(32'h3c3a5c61),
	.w6(32'hbba18d48),
	.w7(32'h3cf23458),
	.w8(32'h3d5705b1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdea287),
	.w1(32'hbcc0baef),
	.w2(32'hbba3db7d),
	.w3(32'h3908c855),
	.w4(32'hbb9c8bdb),
	.w5(32'h3c0ad4f1),
	.w6(32'h3bbde0f3),
	.w7(32'h3960e3de),
	.w8(32'hbb08999c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb239),
	.w1(32'h3b10ee61),
	.w2(32'hbbfd8b81),
	.w3(32'h3bce951a),
	.w4(32'hbb2f117d),
	.w5(32'h3c3164f2),
	.w6(32'h3c097ebb),
	.w7(32'hbb2283b6),
	.w8(32'hbbacb677),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb34f56),
	.w1(32'hbb8bb3ce),
	.w2(32'hbc91d51f),
	.w3(32'h3b8abff7),
	.w4(32'hbba26fae),
	.w5(32'hb9e95028),
	.w6(32'hbb31630e),
	.w7(32'hbb7a166d),
	.w8(32'hbc3af216),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7ebd0),
	.w1(32'hbcaa856e),
	.w2(32'hbb74ec50),
	.w3(32'h3d4acda4),
	.w4(32'hba85504a),
	.w5(32'hbb2e0914),
	.w6(32'h3aaa7a71),
	.w7(32'hbb640761),
	.w8(32'h3ace85d5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6511f0),
	.w1(32'hbb6021e9),
	.w2(32'hbc840805),
	.w3(32'hbab1d604),
	.w4(32'hbca454af),
	.w5(32'hbc423533),
	.w6(32'hbc6ddc25),
	.w7(32'hbcc274da),
	.w8(32'hbce5b5df),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a0dc2),
	.w1(32'h3bf06008),
	.w2(32'h3bb5edd0),
	.w3(32'h3b11df84),
	.w4(32'h3c4779f5),
	.w5(32'hba1bb936),
	.w6(32'hbad4d232),
	.w7(32'h3c23070a),
	.w8(32'h3c7e0cc6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96b4eb),
	.w1(32'hba8a4139),
	.w2(32'hbbdfaf8b),
	.w3(32'hbc6188f0),
	.w4(32'hbb862277),
	.w5(32'hbb919326),
	.w6(32'h3bde8b72),
	.w7(32'h3ad51c2a),
	.w8(32'h3c00e472),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a159d),
	.w1(32'hbc038630),
	.w2(32'h3a00b663),
	.w3(32'hbbac074d),
	.w4(32'h3a14c95a),
	.w5(32'h3c4e2c1b),
	.w6(32'hbb415b40),
	.w7(32'hbbd71700),
	.w8(32'hbb91ea75),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d9a32),
	.w1(32'hbb2778f4),
	.w2(32'hbc2d7cc4),
	.w3(32'h3c9be022),
	.w4(32'hbb7dd109),
	.w5(32'hbb828ad4),
	.w6(32'h3b201f9e),
	.w7(32'hbc243b34),
	.w8(32'hbc6312ea),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3951e6),
	.w1(32'hbc2061ef),
	.w2(32'h3acade98),
	.w3(32'hbc2af014),
	.w4(32'h3c16506d),
	.w5(32'hbb1bcd90),
	.w6(32'h3bbdeb27),
	.w7(32'h3c3ee2b6),
	.w8(32'hbc7b289b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f731),
	.w1(32'hbc638c97),
	.w2(32'hbba1e7f6),
	.w3(32'h3c306787),
	.w4(32'hbbbeab45),
	.w5(32'hbc5e4034),
	.w6(32'h3c182bfd),
	.w7(32'hbb9dbdc2),
	.w8(32'hbc845e6a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb977),
	.w1(32'hbc8d3dbb),
	.w2(32'hbc33ac9d),
	.w3(32'h3c0cd99d),
	.w4(32'hbcaa459b),
	.w5(32'hbc37d5bb),
	.w6(32'hb90efce0),
	.w7(32'hbb7118ed),
	.w8(32'hbc86a415),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce181f1),
	.w1(32'hbc80487d),
	.w2(32'hbc118cff),
	.w3(32'hbc041957),
	.w4(32'hba6f96d3),
	.w5(32'hbb2c0a91),
	.w6(32'h3c02b730),
	.w7(32'hbc9f3fd4),
	.w8(32'hbcf34f61),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc919555),
	.w1(32'hbb026d42),
	.w2(32'hbd30be25),
	.w3(32'h3cbf407e),
	.w4(32'hbcbec252),
	.w5(32'h3c31d148),
	.w6(32'h3d174bab),
	.w7(32'hbd2f3c29),
	.w8(32'hbd14317e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd32ecde),
	.w1(32'hbc81f852),
	.w2(32'hba8753b1),
	.w3(32'h3d5e7b2d),
	.w4(32'hbc0957cf),
	.w5(32'hbab46f8a),
	.w6(32'h3d20c024),
	.w7(32'h3c1bdf91),
	.w8(32'h3c2774c6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d3d05),
	.w1(32'hbb7f8a87),
	.w2(32'h3c2fde5d),
	.w3(32'h3c14c05d),
	.w4(32'h3b893cbe),
	.w5(32'hbcbd5da8),
	.w6(32'h3a219a0a),
	.w7(32'hbb65fc97),
	.w8(32'hbca18d5c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c743324),
	.w1(32'h3ca23481),
	.w2(32'hbc609831),
	.w3(32'hbd16dee3),
	.w4(32'hbc26aa10),
	.w5(32'hbc1a1da2),
	.w6(32'hbcd72741),
	.w7(32'hbc9ef963),
	.w8(32'hbc85468b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20efd1),
	.w1(32'h3b9cf121),
	.w2(32'h3acb0395),
	.w3(32'h3bb4a665),
	.w4(32'hbaef8f54),
	.w5(32'h3c04e113),
	.w6(32'h3b8207ac),
	.w7(32'hbbd2a574),
	.w8(32'hbb1a121d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867620e),
	.w1(32'hbb2b9ce3),
	.w2(32'hbc4e689e),
	.w3(32'h3c09c50b),
	.w4(32'hbca2e576),
	.w5(32'hbc0f52f9),
	.w6(32'h3acf7bd2),
	.w7(32'hbc3f151e),
	.w8(32'hbb397b38),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba4904),
	.w1(32'hbb6b6a5b),
	.w2(32'hbc1a38e1),
	.w3(32'h3c354f72),
	.w4(32'hbc01fa21),
	.w5(32'h3c81693d),
	.w6(32'hbb75933f),
	.w7(32'hbc6f02bd),
	.w8(32'hbceeba62),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec1547),
	.w1(32'hbc28b1c1),
	.w2(32'h3c428a48),
	.w3(32'h3d0cb9ad),
	.w4(32'h3c8eab31),
	.w5(32'h3bd378d0),
	.w6(32'h3d0244d0),
	.w7(32'h3c5e8622),
	.w8(32'h3a8b9d8c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb6384),
	.w1(32'h3b2b304a),
	.w2(32'hbad567fe),
	.w3(32'h38dfff2e),
	.w4(32'hbc7a7973),
	.w5(32'h3b0debb1),
	.w6(32'hbaaa5e4e),
	.w7(32'h3b0311a4),
	.w8(32'h3d865088),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1932b),
	.w1(32'hba76fc86),
	.w2(32'h3a9662ed),
	.w3(32'hbba82cf3),
	.w4(32'hb9ce784c),
	.w5(32'h3c36b9f9),
	.w6(32'h3c6ab029),
	.w7(32'hbbd5dad5),
	.w8(32'hbb41071c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd0605),
	.w1(32'hbb1e124a),
	.w2(32'hbb6c6897),
	.w3(32'h3c66e75a),
	.w4(32'h3b11565f),
	.w5(32'hbb2d8d15),
	.w6(32'h3b0685c6),
	.w7(32'h3b08f774),
	.w8(32'hbcbd16c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38675f),
	.w1(32'hbc401032),
	.w2(32'hbc35016d),
	.w3(32'h3c1a2684),
	.w4(32'hbc541f9c),
	.w5(32'h3c97e5c2),
	.w6(32'h3aa9c696),
	.w7(32'h3c100d3c),
	.w8(32'h3d14b3c0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36bcda),
	.w1(32'h3b8b2035),
	.w2(32'h39e9183e),
	.w3(32'h3b454d88),
	.w4(32'h3bb6a732),
	.w5(32'h3ac83819),
	.w6(32'h3c8ac7c6),
	.w7(32'h3c1dfa34),
	.w8(32'h3b783941),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334617),
	.w1(32'h3be5dff6),
	.w2(32'h3a8bd17f),
	.w3(32'h3c0a4c77),
	.w4(32'hbbe3c14e),
	.w5(32'h3cbaf3b8),
	.w6(32'h3bc22f16),
	.w7(32'hbaa124b3),
	.w8(32'hbc98fb42),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd140b5),
	.w1(32'hba928d86),
	.w2(32'h3b051748),
	.w3(32'hbb4f20df),
	.w4(32'h3bb3cb9d),
	.w5(32'h3b1ed9f4),
	.w6(32'h3bbc235c),
	.w7(32'h3983ca8d),
	.w8(32'hbc341ee7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule