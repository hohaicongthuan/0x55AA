module layer_10_featuremap_41(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075b40),
	.w1(32'h391082d0),
	.w2(32'h3b995240),
	.w3(32'hbbffea02),
	.w4(32'h3a9113ee),
	.w5(32'h3aa69647),
	.w6(32'hbbf36b57),
	.w7(32'hba55a979),
	.w8(32'h3a1fff12),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd62b13),
	.w1(32'hbb3ca693),
	.w2(32'hbba94f14),
	.w3(32'h3b8bd6f0),
	.w4(32'h3a09c9e3),
	.w5(32'hbbaa72e4),
	.w6(32'h3c143d24),
	.w7(32'hb955308f),
	.w8(32'hba95da2f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b841),
	.w1(32'hbb669f3c),
	.w2(32'h3b353105),
	.w3(32'hb89a6cc2),
	.w4(32'hbb875caa),
	.w5(32'hbb00fd87),
	.w6(32'hbc0ef360),
	.w7(32'hbbb7cbb1),
	.w8(32'hbaaf2cb5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5542dc),
	.w1(32'h3ab9129a),
	.w2(32'h3c1f2b37),
	.w3(32'h3b1bfdfa),
	.w4(32'hbadc6d58),
	.w5(32'h3b243293),
	.w6(32'h3b13ffc5),
	.w7(32'h3b2c8db7),
	.w8(32'h3a7057cb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c1dc),
	.w1(32'h3b097b3f),
	.w2(32'h3b331fb3),
	.w3(32'h3b93dee4),
	.w4(32'h3b2a4bc7),
	.w5(32'h3bba6d94),
	.w6(32'h3b0874f4),
	.w7(32'hbba8f78a),
	.w8(32'h3b8316b7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30abfd),
	.w1(32'h3ac51258),
	.w2(32'hbc410de0),
	.w3(32'hba2a9c32),
	.w4(32'hba767122),
	.w5(32'h39e5979d),
	.w6(32'hbaee18a0),
	.w7(32'hba496f9d),
	.w8(32'hbc3a5059),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c063fce),
	.w1(32'h3ab51847),
	.w2(32'h3aa230d0),
	.w3(32'h3cca4c44),
	.w4(32'h3c2b5de7),
	.w5(32'h3bc7885b),
	.w6(32'h3c145838),
	.w7(32'hbaf36153),
	.w8(32'h3b01bf97),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71a538),
	.w1(32'hbad9d2df),
	.w2(32'h3a7e8f1d),
	.w3(32'hbc01e034),
	.w4(32'h39b6ccff),
	.w5(32'h3b32061e),
	.w6(32'h3c359808),
	.w7(32'h3b19b66a),
	.w8(32'hba74379b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5df283),
	.w1(32'h3bb51647),
	.w2(32'h3a8f38b1),
	.w3(32'h3c3fe048),
	.w4(32'h3c113127),
	.w5(32'hbbbcf819),
	.w6(32'h3c41d203),
	.w7(32'h3bc3dc06),
	.w8(32'hba814868),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa140a1),
	.w1(32'h39d2f541),
	.w2(32'hbcdda2a0),
	.w3(32'hbb9e6aab),
	.w4(32'hbaefce76),
	.w5(32'hbd214599),
	.w6(32'hb96133da),
	.w7(32'hba61e7bb),
	.w8(32'hbcc44a61),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06a4d7),
	.w1(32'hbc9c4f38),
	.w2(32'hba369d66),
	.w3(32'hbd6bcb90),
	.w4(32'hbd28ce49),
	.w5(32'h39fa160b),
	.w6(32'hbd2695ca),
	.w7(32'hbcd6507f),
	.w8(32'hbb950a91),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba74bdd),
	.w1(32'h3c44296c),
	.w2(32'hbcd60d0b),
	.w3(32'h3af61ec7),
	.w4(32'h3bfc4a61),
	.w5(32'hbcca4dd8),
	.w6(32'h389e8846),
	.w7(32'h3c1fe2c8),
	.w8(32'hbcc04371),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd3ab0),
	.w1(32'hbcc9d054),
	.w2(32'hbc6a92fe),
	.w3(32'hbc9b83c6),
	.w4(32'hbc9fa76a),
	.w5(32'hbc82c351),
	.w6(32'hbc72a68a),
	.w7(32'hbc8a6ff0),
	.w8(32'hbc3a86cf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeed082),
	.w1(32'hbc1c0df0),
	.w2(32'hbb44e329),
	.w3(32'hbc2f7b51),
	.w4(32'hbc3d4b6d),
	.w5(32'hbba84e1b),
	.w6(32'hbbc786cc),
	.w7(32'hbc349810),
	.w8(32'hbb331e79),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b880ee6),
	.w1(32'h3b89dcfb),
	.w2(32'hbb351f05),
	.w3(32'hb8ceb124),
	.w4(32'hbaadf221),
	.w5(32'h3baaa54a),
	.w6(32'hbb383360),
	.w7(32'h3a4bb504),
	.w8(32'h3b4d1ead),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb090e),
	.w1(32'hbc4cde07),
	.w2(32'hbce3ad08),
	.w3(32'h3bcfc25d),
	.w4(32'hbb9af443),
	.w5(32'hbd02c1ae),
	.w6(32'h3b2beca8),
	.w7(32'hbb56d0e9),
	.w8(32'hbc9640bb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1a47c),
	.w1(32'hbc4f8105),
	.w2(32'h39a8f710),
	.w3(32'hbd2c56e0),
	.w4(32'hbcfc71e1),
	.w5(32'hbb4b256a),
	.w6(32'hbcf1ce43),
	.w7(32'hbca0b346),
	.w8(32'h3b3b03c8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a512c5c),
	.w1(32'h3b68fe84),
	.w2(32'hbc7f0d8a),
	.w3(32'hbbd4ce23),
	.w4(32'hb9684d8a),
	.w5(32'hbc75fa63),
	.w6(32'h3c21ce25),
	.w7(32'h3c4fa0d7),
	.w8(32'hbb7f0e68),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ccf1),
	.w1(32'hbbdc7ee1),
	.w2(32'hbc62308f),
	.w3(32'hbbc43776),
	.w4(32'hbc060f2b),
	.w5(32'hbc31f7ea),
	.w6(32'hbb295c1e),
	.w7(32'hbab2dc9c),
	.w8(32'hbb07d45d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d0583),
	.w1(32'h3c0bdfb0),
	.w2(32'h3b9b9ce1),
	.w3(32'h3b501807),
	.w4(32'h3a02881c),
	.w5(32'h3b8141fe),
	.w6(32'hbb30e627),
	.w7(32'hbb069513),
	.w8(32'h3b9f5bd8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acecfab),
	.w1(32'hbaa398e2),
	.w2(32'hbb21805c),
	.w3(32'hb93303cc),
	.w4(32'hb99f55f4),
	.w5(32'hbb8bf12f),
	.w6(32'h3b456833),
	.w7(32'h3a8ac652),
	.w8(32'hbb9331f7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387cea20),
	.w1(32'h3b821676),
	.w2(32'hbba8f5e5),
	.w3(32'hbaca50d8),
	.w4(32'h3ab4977d),
	.w5(32'hbbe7c194),
	.w6(32'h3af81301),
	.w7(32'h3aa084d4),
	.w8(32'hbbb5c1fd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ed607),
	.w1(32'h3b6e08fa),
	.w2(32'h3b8ba3ae),
	.w3(32'hbbf98a2f),
	.w4(32'hbb9d632b),
	.w5(32'h3b050772),
	.w6(32'h3a229ba1),
	.w7(32'h3c3a70e2),
	.w8(32'h3c8fab1a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c2e3),
	.w1(32'h3c19b5c6),
	.w2(32'hbbaf924e),
	.w3(32'hbc17faf6),
	.w4(32'h3ac76af2),
	.w5(32'hbbcac7df),
	.w6(32'h3b78eb40),
	.w7(32'h3c5aae36),
	.w8(32'h3a852713),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1dec6),
	.w1(32'hbbc01614),
	.w2(32'h3b0fa70d),
	.w3(32'hbc60c705),
	.w4(32'hbbec034f),
	.w5(32'h3b0a4774),
	.w6(32'hbc40d694),
	.w7(32'hbbf8be93),
	.w8(32'h3b6c8af8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c236de0),
	.w1(32'h3c66ad2e),
	.w2(32'h3b8b7877),
	.w3(32'h3c14e7d0),
	.w4(32'h3bc544ae),
	.w5(32'h3ba00460),
	.w6(32'h3c002870),
	.w7(32'h3beebfd9),
	.w8(32'h3bae04b5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099899),
	.w1(32'hbb914b1f),
	.w2(32'h3a9e7c30),
	.w3(32'h39d8d70a),
	.w4(32'hbbcd6c59),
	.w5(32'hb9436b52),
	.w6(32'hbad0a41f),
	.w7(32'hbb02295b),
	.w8(32'hb73b2d16),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5939d6),
	.w1(32'h3b283c6f),
	.w2(32'h3c8083bf),
	.w3(32'hbc47e065),
	.w4(32'hb9f7e51a),
	.w5(32'h3ce6f39c),
	.w6(32'hbc7537f7),
	.w7(32'hbba86aaa),
	.w8(32'h3ca277ce),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc585fd2),
	.w1(32'h3b55b0bc),
	.w2(32'h3c2e7791),
	.w3(32'hbc02d264),
	.w4(32'h3c00ea9b),
	.w5(32'h3b815c07),
	.w6(32'hbc21ae65),
	.w7(32'hbbeac702),
	.w8(32'hbbd8df95),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc20732),
	.w1(32'h3bd03363),
	.w2(32'hbb997fbf),
	.w3(32'hbbc64eb3),
	.w4(32'hbbe2a01c),
	.w5(32'hbbd08b3f),
	.w6(32'hbbb6ddd5),
	.w7(32'hbc73e278),
	.w8(32'hbc44ee3a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025b75),
	.w1(32'hbb98e33b),
	.w2(32'h3b6d9c23),
	.w3(32'h3a6b3fdb),
	.w4(32'hbb41a35d),
	.w5(32'hbb0120df),
	.w6(32'hba1385aa),
	.w7(32'hbb483a84),
	.w8(32'hbc01ab11),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a3b83),
	.w1(32'h3bd1b221),
	.w2(32'h3aa2fe70),
	.w3(32'hbc145092),
	.w4(32'h3bee28d9),
	.w5(32'hbc1553e8),
	.w6(32'hbc03588c),
	.w7(32'h3c3ff3f5),
	.w8(32'hbbd2c4b3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba300522),
	.w1(32'hbb76c7d2),
	.w2(32'hbbae1371),
	.w3(32'hbb5d945e),
	.w4(32'hbb315948),
	.w5(32'hbaf46cfc),
	.w6(32'hbbf359b0),
	.w7(32'h3b5a1bf5),
	.w8(32'hba971b7b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6002a7),
	.w1(32'hbb784b6a),
	.w2(32'hbbccee5f),
	.w3(32'hbaef869a),
	.w4(32'hba64a8d0),
	.w5(32'hbc3ece7f),
	.w6(32'hbb4ced1c),
	.w7(32'hbb897252),
	.w8(32'hbc6a3803),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14c86f),
	.w1(32'h3bb6cdce),
	.w2(32'hba8789aa),
	.w3(32'h3c3dd0dc),
	.w4(32'h3c58fe8a),
	.w5(32'hba9b5e23),
	.w6(32'h3c92e4cf),
	.w7(32'h3c282c53),
	.w8(32'h3b11826d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967f37),
	.w1(32'h3b09d481),
	.w2(32'hbbbd21b4),
	.w3(32'hbbd10dba),
	.w4(32'h39c9cdd2),
	.w5(32'hbc94e7da),
	.w6(32'hba1cece2),
	.w7(32'h3b9cd2ab),
	.w8(32'hbc84751d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b4357),
	.w1(32'h3be9d681),
	.w2(32'hbc03f9c4),
	.w3(32'hbc0a293b),
	.w4(32'hbbe28139),
	.w5(32'hbba45fd5),
	.w6(32'hbc48ec82),
	.w7(32'hbbfdf1a9),
	.w8(32'hbb070aa6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e1075),
	.w1(32'h3bbbbc3a),
	.w2(32'h3c1b0c51),
	.w3(32'hbc6d5bf0),
	.w4(32'h3c72b232),
	.w5(32'h3c54195a),
	.w6(32'hbc6c4f92),
	.w7(32'h3c009009),
	.w8(32'h3bc45127),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee6f83),
	.w1(32'h3c12aa64),
	.w2(32'h3cc307f7),
	.w3(32'hbb90bac5),
	.w4(32'h3c3c5bde),
	.w5(32'h3cb4ba0c),
	.w6(32'hbc583b8f),
	.w7(32'hbb44c98c),
	.w8(32'h3ba8a632),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a60c8),
	.w1(32'hbb6eb54c),
	.w2(32'hbc0555ab),
	.w3(32'hba0d284c),
	.w4(32'hbc6ac12a),
	.w5(32'hbabfad9a),
	.w6(32'h3bb334e3),
	.w7(32'hbc738ceb),
	.w8(32'h3b54c0ea),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb209a),
	.w1(32'hbb5b7e21),
	.w2(32'hbb3a05fe),
	.w3(32'h3c555b2f),
	.w4(32'hb98792c4),
	.w5(32'hbc347a8e),
	.w6(32'h3c968cae),
	.w7(32'h3b9c270e),
	.w8(32'h3a8700d9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94579f),
	.w1(32'hbb5233eb),
	.w2(32'h3c03fea1),
	.w3(32'h39b18420),
	.w4(32'hbba4cf47),
	.w5(32'hbb43ff60),
	.w6(32'h386f7bca),
	.w7(32'h3ae17125),
	.w8(32'hb94bcb88),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19648d),
	.w1(32'h3b26bb9c),
	.w2(32'hba2e1144),
	.w3(32'hbc0c218d),
	.w4(32'h3b2534ed),
	.w5(32'h3aa6b0e2),
	.w6(32'hbb896259),
	.w7(32'h3b9a79c9),
	.w8(32'h3b4a7d06),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc253f5),
	.w1(32'hbc0db601),
	.w2(32'hbb0aa6e6),
	.w3(32'hbc396c5b),
	.w4(32'hba787670),
	.w5(32'h3bf4a37d),
	.w6(32'hbc08f210),
	.w7(32'h3ad09390),
	.w8(32'h3c19205c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc002f23),
	.w1(32'h3ba04d07),
	.w2(32'h3bf55ef3),
	.w3(32'hbbd06d73),
	.w4(32'hbb9a9ebf),
	.w5(32'h3c32fc06),
	.w6(32'h3b9de698),
	.w7(32'hbbeb7232),
	.w8(32'h3c6255f5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18b4ec),
	.w1(32'h3b958227),
	.w2(32'hbc46a9a9),
	.w3(32'hbc7c1de2),
	.w4(32'h3c7a2b9e),
	.w5(32'hbc48b4f0),
	.w6(32'hbae11154),
	.w7(32'h3ca00116),
	.w8(32'hbc4d1bbf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c288006),
	.w1(32'hbbdf32e0),
	.w2(32'hbd15f7c1),
	.w3(32'hba36c6ba),
	.w4(32'hbc7ec99f),
	.w5(32'hbd008202),
	.w6(32'hbbe14ab8),
	.w7(32'hbc2bbd16),
	.w8(32'hbcb8b416),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0908ce),
	.w1(32'hbc1f0c46),
	.w2(32'hbc4b0dd8),
	.w3(32'h3cce5f46),
	.w4(32'h3b2e5dd3),
	.w5(32'hbc1f5725),
	.w6(32'h3c1d32c7),
	.w7(32'h3b78f911),
	.w8(32'hbb80fa02),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab4668),
	.w1(32'hba5cf089),
	.w2(32'h3ae9d790),
	.w3(32'hbbf987f7),
	.w4(32'h3ad4a93d),
	.w5(32'h3c34859e),
	.w6(32'hbbaeff76),
	.w7(32'h39c18ffd),
	.w8(32'h3c026413),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdc4a6),
	.w1(32'h3b8af187),
	.w2(32'h3b0243f5),
	.w3(32'h3c0c6312),
	.w4(32'h3c44f49f),
	.w5(32'h3ba0ff23),
	.w6(32'h3b1c7c9e),
	.w7(32'h3c0ef4e6),
	.w8(32'hba8c48af),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fb834),
	.w1(32'h3b2cf50c),
	.w2(32'hbbc78d96),
	.w3(32'h3be3b69f),
	.w4(32'hbb337ca5),
	.w5(32'hbb0f018e),
	.w6(32'h3c33e770),
	.w7(32'h3b85f16c),
	.w8(32'h3b333bca),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37454c),
	.w1(32'hbc66c8f5),
	.w2(32'hbc0b3c64),
	.w3(32'hbbc617d0),
	.w4(32'hbc1bb022),
	.w5(32'h3b1fea29),
	.w6(32'h396096d5),
	.w7(32'hbb67b7f7),
	.w8(32'h3c16b216),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f7454),
	.w1(32'hbbcc7b61),
	.w2(32'hbb445377),
	.w3(32'hbc8608b0),
	.w4(32'hbba1ca13),
	.w5(32'hbc176078),
	.w6(32'hbbc9e5e2),
	.w7(32'hbc152086),
	.w8(32'hbbbeea95),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1a7be),
	.w1(32'h3a36c379),
	.w2(32'h3b883613),
	.w3(32'hba9150bc),
	.w4(32'h3afc849c),
	.w5(32'h3b370483),
	.w6(32'h3bd4fbe0),
	.w7(32'h3c591ca9),
	.w8(32'h3bd866b5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff3bbe),
	.w1(32'hbb9e9337),
	.w2(32'h3c8ffe5f),
	.w3(32'h3b4ca665),
	.w4(32'hbb80667c),
	.w5(32'h3c354e95),
	.w6(32'h3be281df),
	.w7(32'h3b413b6f),
	.w8(32'h3c11a068),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c9ed8),
	.w1(32'h3c383ab8),
	.w2(32'hba6eecad),
	.w3(32'h3c23da19),
	.w4(32'h3c809db9),
	.w5(32'hba04253b),
	.w6(32'h3ba37425),
	.w7(32'h3caa9f45),
	.w8(32'hbb40c502),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca20763),
	.w1(32'h3b4f931d),
	.w2(32'h3ad626ab),
	.w3(32'hbc7fc0fb),
	.w4(32'h3b88c927),
	.w5(32'h3c042d1d),
	.w6(32'hbc1283ce),
	.w7(32'hbb6a76f6),
	.w8(32'h3bf5046f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e59fb),
	.w1(32'hba1a47d1),
	.w2(32'h3b868c0b),
	.w3(32'h3b2d1be3),
	.w4(32'hbb0b915b),
	.w5(32'h3afdc64b),
	.w6(32'h39db39d9),
	.w7(32'hb9866f25),
	.w8(32'h3b7e4a43),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06687f),
	.w1(32'hbb9ec48a),
	.w2(32'hb8ec88dd),
	.w3(32'hbbc73083),
	.w4(32'hbb38d50f),
	.w5(32'h3b8184d9),
	.w6(32'h3a587bd5),
	.w7(32'h3b40d126),
	.w8(32'h3c062d75),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95f5b1),
	.w1(32'h3b2397ff),
	.w2(32'hb9e3916b),
	.w3(32'h3aa41670),
	.w4(32'h3b3df31f),
	.w5(32'h3abbffbd),
	.w6(32'hba578a76),
	.w7(32'h3c2b4476),
	.w8(32'hbb1606c4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002882),
	.w1(32'hbbbbcc42),
	.w2(32'h3c632a8f),
	.w3(32'h3c5059f8),
	.w4(32'hbb14c9b1),
	.w5(32'h3c57a1c4),
	.w6(32'h3c27aa3f),
	.w7(32'h3aa61941),
	.w8(32'h3c223e7d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1c050),
	.w1(32'h3a441af7),
	.w2(32'hbad68506),
	.w3(32'h3cc98be4),
	.w4(32'h3c170287),
	.w5(32'hb936181d),
	.w6(32'h3c871713),
	.w7(32'h3b5c10d6),
	.w8(32'hbac4f7ed),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8852d67),
	.w1(32'hba7ea317),
	.w2(32'h3b29bece),
	.w3(32'hbaaaefd3),
	.w4(32'h3b84b29b),
	.w5(32'h39fb03e7),
	.w6(32'hbb16dcc3),
	.w7(32'h3bf830d7),
	.w8(32'hbb484931),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea48a5),
	.w1(32'h3ab3fa0e),
	.w2(32'h399c65e7),
	.w3(32'hbc19be20),
	.w4(32'h3bd156b5),
	.w5(32'hbc209aa5),
	.w6(32'hbc1ef600),
	.w7(32'h3b0ee7cd),
	.w8(32'hbafcffa8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc029aa1),
	.w1(32'h3b9419ce),
	.w2(32'h3b832110),
	.w3(32'hbc5519a5),
	.w4(32'h3c1b03c8),
	.w5(32'h3b6f4af2),
	.w6(32'hbc99835b),
	.w7(32'h3a51eb81),
	.w8(32'h3bdddea8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3a190),
	.w1(32'h3bb478d4),
	.w2(32'h3b08a49d),
	.w3(32'hbac71157),
	.w4(32'h3b13734b),
	.w5(32'h3bc3c2f8),
	.w6(32'hbab73582),
	.w7(32'h3a925eb6),
	.w8(32'h3c05104d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea165),
	.w1(32'hbbb6c3cc),
	.w2(32'hbd0022c6),
	.w3(32'h3b51df64),
	.w4(32'h3b2a8763),
	.w5(32'hbc83852a),
	.w6(32'hbac5f954),
	.w7(32'h39f49083),
	.w8(32'hbb9563df),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98b2c6),
	.w1(32'hbcb5b71a),
	.w2(32'h3acdf9d5),
	.w3(32'hbb15c34b),
	.w4(32'hbcce29a2),
	.w5(32'h3b5d3049),
	.w6(32'h3ca49758),
	.w7(32'hbc418fe6),
	.w8(32'h3c903f97),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75561e),
	.w1(32'h3c0aef97),
	.w2(32'hbb56c3e8),
	.w3(32'hbc7b2869),
	.w4(32'h3c399d80),
	.w5(32'h3b171967),
	.w6(32'hbb67db9c),
	.w7(32'h3c9ac3c5),
	.w8(32'h3c56be24),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd4f9a),
	.w1(32'h3ba89357),
	.w2(32'hbbbec6b3),
	.w3(32'hbbe177b8),
	.w4(32'h3ba20b7b),
	.w5(32'hbbc0e64c),
	.w6(32'hbad091b3),
	.w7(32'h3c2b3b30),
	.w8(32'hbbb09005),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e9d3e),
	.w1(32'hbc0f7ba8),
	.w2(32'h3b7304a4),
	.w3(32'h3b76332a),
	.w4(32'hbc06b02a),
	.w5(32'h3b8dc4d1),
	.w6(32'h3984325a),
	.w7(32'hbb9cc695),
	.w8(32'hba7a5c41),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f6f1),
	.w1(32'hbafdac0f),
	.w2(32'h3abad2f6),
	.w3(32'hbbeaa36d),
	.w4(32'hbc2a4649),
	.w5(32'h3b656bf6),
	.w6(32'h3b119cf4),
	.w7(32'hbc500354),
	.w8(32'hbc04137b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d22e267),
	.w1(32'hbc6f50b4),
	.w2(32'h3c476b14),
	.w3(32'h3d60d8be),
	.w4(32'hbb86fa5d),
	.w5(32'h3c435a11),
	.w6(32'h3d2a58e1),
	.w7(32'hbb9e5354),
	.w8(32'h3c5dd001),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d787e),
	.w1(32'h3c8d8fbd),
	.w2(32'h3aa42aa8),
	.w3(32'hbd54f250),
	.w4(32'h3ca5926d),
	.w5(32'h3ab1dd06),
	.w6(32'hbd18be6d),
	.w7(32'h3bab8d6e),
	.w8(32'h3ba92f1a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecdc27),
	.w1(32'hba8d34ba),
	.w2(32'h3acda3bf),
	.w3(32'hbc3e1659),
	.w4(32'hb938a3f6),
	.w5(32'h3b458966),
	.w6(32'hbc004eb2),
	.w7(32'hb9f1455f),
	.w8(32'h3af94ca4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf26a6),
	.w1(32'h3afcc64e),
	.w2(32'h3b6906e2),
	.w3(32'hbb1e08f4),
	.w4(32'h3b638277),
	.w5(32'h3bcf4518),
	.w6(32'hb9cd625e),
	.w7(32'h3aab4bea),
	.w8(32'h3bf6b9e0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25d54e),
	.w1(32'h3b3ed836),
	.w2(32'hbba8dff0),
	.w3(32'hbc42aabe),
	.w4(32'h3b910525),
	.w5(32'hb9625ddc),
	.w6(32'hbbe434e9),
	.w7(32'hb9bddec2),
	.w8(32'h3bf15422),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5665b),
	.w1(32'h3c2f058f),
	.w2(32'hbcbf41c6),
	.w3(32'hbc399c40),
	.w4(32'h3c3fcf44),
	.w5(32'hbc86fb98),
	.w6(32'hbc56f655),
	.w7(32'h3b3d85c0),
	.w8(32'hbc4867d7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42a71c),
	.w1(32'hbc08c954),
	.w2(32'hbb11b1ad),
	.w3(32'hbc99b6dd),
	.w4(32'hbc5c31f5),
	.w5(32'hb9a91e9f),
	.w6(32'hbc5b9041),
	.w7(32'hbc06084e),
	.w8(32'hba17414e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c031bf3),
	.w1(32'h39308484),
	.w2(32'hbc3a9f18),
	.w3(32'h3c4389c6),
	.w4(32'hbab2e3cb),
	.w5(32'hbc4740a9),
	.w6(32'h3c2267b5),
	.w7(32'hbb413d37),
	.w8(32'hbc2deadc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4fb98),
	.w1(32'h39212efe),
	.w2(32'h3a79ce63),
	.w3(32'h3aa79d8c),
	.w4(32'h3ac09aa7),
	.w5(32'h3b0c8a9c),
	.w6(32'hbb75cc7a),
	.w7(32'h3ada638e),
	.w8(32'h3a09fb23),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf86c),
	.w1(32'hbb3b6f10),
	.w2(32'hbcb3ae2a),
	.w3(32'hb9fa0eef),
	.w4(32'hbb69c31a),
	.w5(32'hbcf4cee7),
	.w6(32'hb8b29ad2),
	.w7(32'hbb02b9ba),
	.w8(32'hbcb9a9dd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfcb4f),
	.w1(32'hbc87e339),
	.w2(32'h3b950e54),
	.w3(32'h3d008bba),
	.w4(32'hbc7ad489),
	.w5(32'h3c562d12),
	.w6(32'h3cd281a7),
	.w7(32'hbc2a9523),
	.w8(32'h3c484b7c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d9cf5),
	.w1(32'h3c6b7667),
	.w2(32'hbbc87f4f),
	.w3(32'hbb92b9c8),
	.w4(32'h3cb4807f),
	.w5(32'hbc289069),
	.w6(32'hbc2eaf63),
	.w7(32'h3bacdc8e),
	.w8(32'hbc688407),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e887e),
	.w1(32'hbc2c29cf),
	.w2(32'h3c51d8fc),
	.w3(32'h3cdb2ece),
	.w4(32'hbbe07a5d),
	.w5(32'h3c45143d),
	.w6(32'h3c4b681c),
	.w7(32'hbbb7f8e9),
	.w8(32'h3c02ecec),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16811c),
	.w1(32'h3bc7aff8),
	.w2(32'h3a62b963),
	.w3(32'hbbcaceeb),
	.w4(32'h3c52a912),
	.w5(32'hb9ed5f55),
	.w6(32'hba515b04),
	.w7(32'h3bfc6212),
	.w8(32'h3abbafc3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8861d0),
	.w1(32'h3c19d663),
	.w2(32'h3b981fad),
	.w3(32'hbb5c4d08),
	.w4(32'h3c066a31),
	.w5(32'h3b310bfe),
	.w6(32'hbbe4e84f),
	.w7(32'h3bc77bb4),
	.w8(32'h3bca87c4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d58323),
	.w1(32'h39906fdb),
	.w2(32'hbc18eed8),
	.w3(32'hbaddb133),
	.w4(32'hbb0b8215),
	.w5(32'hbc4efecf),
	.w6(32'hb9fb45a6),
	.w7(32'h3800e0a3),
	.w8(32'h392d1f37),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ded9a),
	.w1(32'hbc1bb8af),
	.w2(32'h3ac2d097),
	.w3(32'hbca200ef),
	.w4(32'hbc47a0ea),
	.w5(32'hbbc7e46d),
	.w6(32'hbc344d12),
	.w7(32'hbc06e256),
	.w8(32'hbc1fe64a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53efe3),
	.w1(32'hbc048424),
	.w2(32'h3c088496),
	.w3(32'h3a702dfe),
	.w4(32'hbc754768),
	.w5(32'h3bdee89a),
	.w6(32'h3b371a33),
	.w7(32'h3b8316ee),
	.w8(32'h3c2ade57),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91d48b),
	.w1(32'h3bc199cf),
	.w2(32'h3c165f61),
	.w3(32'hbc0b6fcb),
	.w4(32'h3c14ab20),
	.w5(32'h3c571866),
	.w6(32'hbc1899cb),
	.w7(32'h3bc13f82),
	.w8(32'h3c095e90),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f414),
	.w1(32'h3ae1d8b0),
	.w2(32'hbb95c6f0),
	.w3(32'h3c031a86),
	.w4(32'h3c2881e6),
	.w5(32'h3b511299),
	.w6(32'h3c4b8520),
	.w7(32'h3c0ade0f),
	.w8(32'h3c5c8d56),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea1e1d),
	.w1(32'h3a021397),
	.w2(32'h3aa44428),
	.w3(32'h3b4b049b),
	.w4(32'h3b9ee410),
	.w5(32'h3b94f4b5),
	.w6(32'h3c27536a),
	.w7(32'h3c5e782b),
	.w8(32'h3bc5e7f0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a3ec9),
	.w1(32'hbc4a7f78),
	.w2(32'h3ac24d3b),
	.w3(32'h3b8a5469),
	.w4(32'hbb3e3920),
	.w5(32'h3c28bd12),
	.w6(32'h3b9796e4),
	.w7(32'h3a8618bb),
	.w8(32'h3c9a264e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26ee5a),
	.w1(32'h3c01d33f),
	.w2(32'hbc12ca53),
	.w3(32'hbafe6508),
	.w4(32'h3bfb778f),
	.w5(32'hbaf0b890),
	.w6(32'hbb2d3763),
	.w7(32'h3b8d8726),
	.w8(32'h3c252cd0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99246),
	.w1(32'hbc3dba99),
	.w2(32'h3c061f43),
	.w3(32'hbbfefa37),
	.w4(32'hbc6c524d),
	.w5(32'hbb893716),
	.w6(32'hbc6516a7),
	.w7(32'hbc847129),
	.w8(32'hbc0e02da),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a627),
	.w1(32'hbc49cff6),
	.w2(32'hba570d4c),
	.w3(32'hbc3571ad),
	.w4(32'hbc081945),
	.w5(32'hbcb2650f),
	.w6(32'hbb4ee35d),
	.w7(32'hbc05a9c0),
	.w8(32'hbc80f6b0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156c8d),
	.w1(32'hbc3ca068),
	.w2(32'hbc0c8f7f),
	.w3(32'hbc9d8001),
	.w4(32'hbc51225f),
	.w5(32'hbbe94008),
	.w6(32'hbc73c237),
	.w7(32'h3ba544d9),
	.w8(32'hbc003560),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9915601),
	.w1(32'h3c3255ef),
	.w2(32'hbb2eaa73),
	.w3(32'hbc1fbd8b),
	.w4(32'h3c9f56af),
	.w5(32'h3bf2a90a),
	.w6(32'hbb944c6e),
	.w7(32'h3cb570d1),
	.w8(32'h3c57163f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f34eb),
	.w1(32'h3bb8c925),
	.w2(32'hbbb43735),
	.w3(32'hbc2de074),
	.w4(32'h3ac00402),
	.w5(32'hbb99c69a),
	.w6(32'h38c6fbd0),
	.w7(32'h3c708935),
	.w8(32'hbb8971c7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16eccc),
	.w1(32'h3cd622f8),
	.w2(32'h3c607890),
	.w3(32'hbc3aa203),
	.w4(32'h3d0efbb6),
	.w5(32'h3c82f3b6),
	.w6(32'hbc9e2b13),
	.w7(32'h3cc8a422),
	.w8(32'h3c723758),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8ff3),
	.w1(32'h3b1ff664),
	.w2(32'hbb25103e),
	.w3(32'hbba60d47),
	.w4(32'h3c40b3e0),
	.w5(32'hbc0ee7b8),
	.w6(32'hbb77059d),
	.w7(32'h3c134eec),
	.w8(32'hbb0b80a3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f14d9),
	.w1(32'h3c84b14c),
	.w2(32'hbb065211),
	.w3(32'hbc715317),
	.w4(32'h3c7ecda1),
	.w5(32'hb901160d),
	.w6(32'hbc530cc9),
	.w7(32'h3ca4fe66),
	.w8(32'hbbe737a9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab22dc),
	.w1(32'h3bc7955d),
	.w2(32'h3c16ae53),
	.w3(32'h3b6f542f),
	.w4(32'h3c3e8442),
	.w5(32'h3b992ed6),
	.w6(32'hbaa625fa),
	.w7(32'h3c6f13db),
	.w8(32'hbc3fedb5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4047a3),
	.w1(32'hbcdded1c),
	.w2(32'h3ad306b3),
	.w3(32'h3b970d3c),
	.w4(32'hbcb0189a),
	.w5(32'hbbbbe851),
	.w6(32'h3bd8907b),
	.w7(32'hbc711a40),
	.w8(32'h3a208973),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f14ef),
	.w1(32'h3b02d369),
	.w2(32'h3be85be2),
	.w3(32'h3a6ccceb),
	.w4(32'h3a511c2f),
	.w5(32'h3b25cecc),
	.w6(32'h3bc8fc36),
	.w7(32'h3b6bd3af),
	.w8(32'hbaf2e37b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade3eca),
	.w1(32'hbadf141c),
	.w2(32'hbc34ce5e),
	.w3(32'hb9cb187d),
	.w4(32'hbb687610),
	.w5(32'hbc1f7dd1),
	.w6(32'hbb084f5e),
	.w7(32'hbbb1419a),
	.w8(32'hbae50b2a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc363a1),
	.w1(32'h3bfcaa72),
	.w2(32'h3c565a93),
	.w3(32'h3bd518b4),
	.w4(32'h3bbfa27a),
	.w5(32'hba9fe9f1),
	.w6(32'hba7bd62f),
	.w7(32'h3ade0195),
	.w8(32'hbc30a5fc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab74f2),
	.w1(32'hbba929c0),
	.w2(32'h3b443aa9),
	.w3(32'h3cc34fef),
	.w4(32'hbc9c2eca),
	.w5(32'h3c323e76),
	.w6(32'h3cb92ddd),
	.w7(32'hbc584c3d),
	.w8(32'h3c7cdf26),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ac095),
	.w1(32'h3c7b08b1),
	.w2(32'h3c5a3f30),
	.w3(32'h3bd84582),
	.w4(32'h3cd6935f),
	.w5(32'hbabaf4b7),
	.w6(32'h3bf5d5e8),
	.w7(32'h3ca70af9),
	.w8(32'h3b8e2b22),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba766a3),
	.w1(32'h38382f90),
	.w2(32'h3b2c179c),
	.w3(32'hbb53c156),
	.w4(32'h3bb69e61),
	.w5(32'h3b71da10),
	.w6(32'h3b586a09),
	.w7(32'h3b25d4ea),
	.w8(32'hbae551f3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed42e),
	.w1(32'hbc17ad8b),
	.w2(32'hbaeedaa0),
	.w3(32'h3cdbe643),
	.w4(32'hbb434d70),
	.w5(32'h39a68660),
	.w6(32'h3c9e69c6),
	.w7(32'hbc172541),
	.w8(32'h3b3274a3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88008cb),
	.w1(32'h3b1664d4),
	.w2(32'hbb8993b6),
	.w3(32'h3b6d9e18),
	.w4(32'h3b84be3b),
	.w5(32'hbc1b5416),
	.w6(32'h3c424a75),
	.w7(32'h3c9af6cd),
	.w8(32'h39f00201),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0ad95),
	.w1(32'hbc1723f1),
	.w2(32'h3a82b21d),
	.w3(32'hbb58820a),
	.w4(32'hbb3ed99b),
	.w5(32'h399152b3),
	.w6(32'h38c4f310),
	.w7(32'h3bb4f6e7),
	.w8(32'h3aa501af),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23db2e),
	.w1(32'h3c2cca47),
	.w2(32'hbb9b9ff0),
	.w3(32'hbc9bda45),
	.w4(32'h3b2f870f),
	.w5(32'h3b28f3a8),
	.w6(32'hbc9b514c),
	.w7(32'hba16cbfb),
	.w8(32'h3babe993),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b411e95),
	.w1(32'h3bfd1e3c),
	.w2(32'h3b5aa82e),
	.w3(32'h3ae92b64),
	.w4(32'h3b6e54aa),
	.w5(32'h3a24b6c1),
	.w6(32'hba6090c1),
	.w7(32'hba563ae8),
	.w8(32'hb7609528),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34ec90),
	.w1(32'hbad9b847),
	.w2(32'hbb12f6e0),
	.w3(32'h3aacd398),
	.w4(32'hbbbdd95a),
	.w5(32'hbb412c32),
	.w6(32'h3a2c844c),
	.w7(32'hbab806b5),
	.w8(32'h393a638f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02dba6),
	.w1(32'h3b775722),
	.w2(32'hbc040801),
	.w3(32'hbaf3225e),
	.w4(32'hb9947c59),
	.w5(32'hbc2376f2),
	.w6(32'h3b23f0f9),
	.w7(32'h3b321dbb),
	.w8(32'hbb9b50ed),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014341),
	.w1(32'hbc04d596),
	.w2(32'hbba46f4b),
	.w3(32'hbc0d14a3),
	.w4(32'h3b05b6a2),
	.w5(32'hbad099cb),
	.w6(32'hbc445ae0),
	.w7(32'h3933b389),
	.w8(32'h3bb0f46f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e2cf),
	.w1(32'h3b85a1fb),
	.w2(32'h3ba19329),
	.w3(32'hbc459e12),
	.w4(32'h3c56b81f),
	.w5(32'h3bef0452),
	.w6(32'hbc2de3b3),
	.w7(32'h3c66a098),
	.w8(32'h3bfd52d0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f350a4),
	.w1(32'h3a9f63a0),
	.w2(32'hbac358da),
	.w3(32'hbaf4fdeb),
	.w4(32'h3a50fe27),
	.w5(32'hbb5f8fdd),
	.w6(32'hb8c9f223),
	.w7(32'h3bfe7e75),
	.w8(32'hbb5b47d3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061bad),
	.w1(32'h3ac5c7e4),
	.w2(32'hbbdf1297),
	.w3(32'hbbe4ff19),
	.w4(32'h3906cb38),
	.w5(32'hbb8ef599),
	.w6(32'hbb2872a9),
	.w7(32'h3ad6b9a0),
	.w8(32'hbb809b55),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3466b8),
	.w1(32'hbafdeb45),
	.w2(32'hbbb7131c),
	.w3(32'h3b64019d),
	.w4(32'hbbbf5ecc),
	.w5(32'hbc045103),
	.w6(32'hbafd5184),
	.w7(32'hbbc3cf08),
	.w8(32'hbc8f1c44),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaa251),
	.w1(32'hbc3783a4),
	.w2(32'h3bd87f9f),
	.w3(32'hbc859682),
	.w4(32'hbcb04da0),
	.w5(32'h3c0cb839),
	.w6(32'hbc90e81d),
	.w7(32'hbcb2901d),
	.w8(32'h3afa15ca),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf44c06),
	.w1(32'h3b9e42b1),
	.w2(32'h3bd7d6f8),
	.w3(32'h39e1626b),
	.w4(32'h3b1d94e1),
	.w5(32'hbae336b6),
	.w6(32'hbb77ccbf),
	.w7(32'hbb07e076),
	.w8(32'hbbaec46d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa28530),
	.w1(32'hbcae32f3),
	.w2(32'hbc21fc15),
	.w3(32'h3bde1eb2),
	.w4(32'hbcd14bc7),
	.w5(32'hbc55fd4a),
	.w6(32'hbbd35fae),
	.w7(32'hbc45e28e),
	.w8(32'hbca5043a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadbf25),
	.w1(32'hbc5f57d9),
	.w2(32'hbbb4a687),
	.w3(32'h3d0b2cf1),
	.w4(32'hbcabb25c),
	.w5(32'hbb6dd791),
	.w6(32'h3d17efcc),
	.w7(32'hbc57cab6),
	.w8(32'hbc081d7e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c215716),
	.w1(32'hbca01992),
	.w2(32'h3bff4b0a),
	.w3(32'h3c7d5187),
	.w4(32'hbcdd36c9),
	.w5(32'h3b1a7534),
	.w6(32'h3cfefe7f),
	.w7(32'hbbe95cc8),
	.w8(32'h3aae4d22),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d717),
	.w1(32'hbb0b568f),
	.w2(32'hbc719cc4),
	.w3(32'h3bc73494),
	.w4(32'hbc71317d),
	.w5(32'hbc274532),
	.w6(32'h3c470bff),
	.w7(32'hbc77e695),
	.w8(32'h3a55e36f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a1992),
	.w1(32'hbc4f9b1e),
	.w2(32'h3bccd19b),
	.w3(32'h3bde7240),
	.w4(32'hbbdeaae5),
	.w5(32'h3c441606),
	.w6(32'hbc0b3c6c),
	.w7(32'hbad0289f),
	.w8(32'h3c3d38f4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8befed),
	.w1(32'h3c6a89ae),
	.w2(32'h3ba7da6d),
	.w3(32'hbd0290e4),
	.w4(32'h3d03021b),
	.w5(32'h3c3f6d8e),
	.w6(32'hbc766f67),
	.w7(32'h3cb481ee),
	.w8(32'h3bc48d38),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2797ba),
	.w1(32'h3b7bfd40),
	.w2(32'hbc384cb0),
	.w3(32'h3b583607),
	.w4(32'h3c5e61b0),
	.w5(32'hbc6c2bca),
	.w6(32'h3abc9a4b),
	.w7(32'h3c120c2e),
	.w8(32'hbb0934e0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9c4e),
	.w1(32'hbb9c4e30),
	.w2(32'hbbaeb029),
	.w3(32'hbc53745b),
	.w4(32'h3927d1a9),
	.w5(32'hbc1c7441),
	.w6(32'hbc5d87f6),
	.w7(32'hbbd2cbb1),
	.w8(32'hbb9c0f36),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16bc10),
	.w1(32'h3c4a1352),
	.w2(32'hbb9ebac3),
	.w3(32'hbb589d95),
	.w4(32'h3c0f73b2),
	.w5(32'hb9acffa9),
	.w6(32'hbb834c24),
	.w7(32'h3c05d809),
	.w8(32'h3a2014d5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5d9c5),
	.w1(32'hbaad4a8d),
	.w2(32'hbbe0a2de),
	.w3(32'hbbd4ee4c),
	.w4(32'hbb0068a0),
	.w5(32'h3a039569),
	.w6(32'hbbc0cc2a),
	.w7(32'hb7e502ca),
	.w8(32'h3ab08ca8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b47a8),
	.w1(32'h3b82b012),
	.w2(32'h3c46b92e),
	.w3(32'hbb2cb77c),
	.w4(32'h3c034eb5),
	.w5(32'h3c00d1e9),
	.w6(32'hbc04ca60),
	.w7(32'h3b69adf6),
	.w8(32'h3baa8ebf),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac0171),
	.w1(32'h3c6037c5),
	.w2(32'h3b1f5074),
	.w3(32'hbbe4ffea),
	.w4(32'hb9ee603e),
	.w5(32'h3baa9204),
	.w6(32'hbb9bddec),
	.w7(32'h3c005e88),
	.w8(32'h3bd69c07),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af235ff),
	.w1(32'hbb409114),
	.w2(32'hba2012c4),
	.w3(32'h386e94bf),
	.w4(32'hbb8b5a8f),
	.w5(32'h3a0415b3),
	.w6(32'hbaa13041),
	.w7(32'hbac66103),
	.w8(32'h3b516a91),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f7672),
	.w1(32'h3aa7ada6),
	.w2(32'h3bb15457),
	.w3(32'h3bf8a47f),
	.w4(32'h3a0cc207),
	.w5(32'hbbc83ac0),
	.w6(32'h3c1b77d4),
	.w7(32'h3b820e97),
	.w8(32'hbb4c7a86),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcc07b),
	.w1(32'hba858e29),
	.w2(32'hbbd68d01),
	.w3(32'hbbce3477),
	.w4(32'h3b735450),
	.w5(32'hba63c680),
	.w6(32'hbc011398),
	.w7(32'h3bd0975c),
	.w8(32'h3a8d1124),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb5ebc),
	.w1(32'hbb527e32),
	.w2(32'hba2c2d7f),
	.w3(32'hba25b932),
	.w4(32'hbba8ab92),
	.w5(32'hb8b8eb07),
	.w6(32'hbad86703),
	.w7(32'hbb822d81),
	.w8(32'h3a086aef),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3004ce),
	.w1(32'h3c5d515c),
	.w2(32'h3b91913c),
	.w3(32'hbba3fa09),
	.w4(32'h39b984d5),
	.w5(32'h3a7d7736),
	.w6(32'hbc4b67c4),
	.w7(32'hbbd921e6),
	.w8(32'h3b1e9149),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe854b),
	.w1(32'h3c3d3a3c),
	.w2(32'hbb029152),
	.w3(32'hbb16f3c5),
	.w4(32'h3c94050c),
	.w5(32'hbb49d98a),
	.w6(32'hbb81a04f),
	.w7(32'h3bedd078),
	.w8(32'h3b992f88),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a808b28),
	.w1(32'h3a9d3569),
	.w2(32'hb9f8aa08),
	.w3(32'hbaf29cbc),
	.w4(32'hb99873bc),
	.w5(32'h3ae65bd0),
	.w6(32'h39a44133),
	.w7(32'h3a0a74c2),
	.w8(32'h3a59254d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58ee1c),
	.w1(32'hbb38d55e),
	.w2(32'h3a8bf22d),
	.w3(32'h3c0f8ebb),
	.w4(32'hbb3b11a9),
	.w5(32'h3a6368a8),
	.w6(32'h3bdb3f40),
	.w7(32'hbb1c6992),
	.w8(32'hba5ecfdf),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cb0e8),
	.w1(32'h3ba85831),
	.w2(32'h3b51b49d),
	.w3(32'hbabe7437),
	.w4(32'h3c1e410e),
	.w5(32'h3b696749),
	.w6(32'hbb94d75b),
	.w7(32'h3c36a7c4),
	.w8(32'hbba4ce68),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3642b),
	.w1(32'h3ad7546f),
	.w2(32'hbb98d5f0),
	.w3(32'h3a24b94f),
	.w4(32'hba8bb780),
	.w5(32'hbc056fca),
	.w6(32'hbb0b7095),
	.w7(32'hbb10edec),
	.w8(32'hba5f785c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6aa993),
	.w1(32'hbc281c3e),
	.w2(32'hbc12bdc8),
	.w3(32'h3c911f02),
	.w4(32'h3ba00e4b),
	.w5(32'hbc2b9050),
	.w6(32'h3c85389f),
	.w7(32'h3c1653e0),
	.w8(32'hbbed0427),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43ee8),
	.w1(32'h39e7e0a2),
	.w2(32'h39824aa4),
	.w3(32'h3b05c52f),
	.w4(32'h3ba57bed),
	.w5(32'hbbc6bd78),
	.w6(32'hbb503219),
	.w7(32'h3ba6a6e7),
	.w8(32'hbbdf34c9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef78c1),
	.w1(32'hbc5a6c86),
	.w2(32'hbbab3563),
	.w3(32'h3bfd5246),
	.w4(32'hbc234808),
	.w5(32'hbb9ec825),
	.w6(32'hbb95cbd7),
	.w7(32'h3b665170),
	.w8(32'hbb5b745b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6848),
	.w1(32'hbc681012),
	.w2(32'hbc02944c),
	.w3(32'h3c7c6f1f),
	.w4(32'hbca667e8),
	.w5(32'hbbef3671),
	.w6(32'h3c3cc746),
	.w7(32'hbc0af455),
	.w8(32'hbbdae816),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5693),
	.w1(32'hbc306ac5),
	.w2(32'hbc479175),
	.w3(32'hbbe8c032),
	.w4(32'hbc2bc0a9),
	.w5(32'hbbd75bfa),
	.w6(32'hbb5819d6),
	.w7(32'hbb934631),
	.w8(32'hbc1cfc9b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8134ca),
	.w1(32'h3aceb6da),
	.w2(32'hbc36750c),
	.w3(32'hbc3fcb51),
	.w4(32'h3aa0cf88),
	.w5(32'hbbca0c93),
	.w6(32'hbc4f1001),
	.w7(32'hbc07fc7d),
	.w8(32'hbb8c39d5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5127ad),
	.w1(32'hbb55d083),
	.w2(32'h3bc69389),
	.w3(32'hbce6e86a),
	.w4(32'hbb07df7e),
	.w5(32'h3c48bec8),
	.w6(32'hbc8a32c4),
	.w7(32'hbbb23934),
	.w8(32'h3c8e3dd8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d9d87),
	.w1(32'h3c500175),
	.w2(32'h3aab8662),
	.w3(32'h3b1814d4),
	.w4(32'h3c3fcf72),
	.w5(32'h3b8b23f2),
	.w6(32'h3b86d1fe),
	.w7(32'h3bafdac4),
	.w8(32'h3b3d8ea8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac7400),
	.w1(32'h3b46b74e),
	.w2(32'hbc1fa122),
	.w3(32'h3bd15223),
	.w4(32'h3bd20637),
	.w5(32'hbca164f8),
	.w6(32'h3b1fdd50),
	.w7(32'h3b9103c1),
	.w8(32'hbc8b9465),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace13ee),
	.w1(32'h3be9fbcf),
	.w2(32'h3c21d570),
	.w3(32'h3b8dabeb),
	.w4(32'h3cc19077),
	.w5(32'h3c278df2),
	.w6(32'hbb781e47),
	.w7(32'h3ccb34b9),
	.w8(32'h3c57ee32),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a47f7),
	.w1(32'h3ab01a72),
	.w2(32'h3b394166),
	.w3(32'hbbc9be22),
	.w4(32'hbb936064),
	.w5(32'h3b1f228d),
	.w6(32'hbaa783d1),
	.w7(32'hbb9c3576),
	.w8(32'h3bb4039b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb210c88),
	.w1(32'hba85ebe2),
	.w2(32'hbba08547),
	.w3(32'hbbc41df0),
	.w4(32'hbbac42d0),
	.w5(32'hba25ae8e),
	.w6(32'hba9adeae),
	.w7(32'hbb008d70),
	.w8(32'hb7e47c6c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beab910),
	.w1(32'h3a068f9b),
	.w2(32'h3a075638),
	.w3(32'h3b1966c5),
	.w4(32'h3bb24c4b),
	.w5(32'h3b8aa65d),
	.w6(32'hbb32964d),
	.w7(32'hbb47de62),
	.w8(32'hbc6c1261),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb744b4c),
	.w1(32'hbc876c51),
	.w2(32'hbbb494c7),
	.w3(32'h3b8c58be),
	.w4(32'hbc06bc31),
	.w5(32'hbb638c31),
	.w6(32'hbb8236ca),
	.w7(32'hbbf60552),
	.w8(32'hbb921feb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaef569),
	.w1(32'hbb818b52),
	.w2(32'hbc465fd7),
	.w3(32'h3b19c9cc),
	.w4(32'hbb9885af),
	.w5(32'hbc1f43df),
	.w6(32'h3b1a0a67),
	.w7(32'hb9f08452),
	.w8(32'hbbee8ed1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b5135),
	.w1(32'h3a83c678),
	.w2(32'hbaccecae),
	.w3(32'hbc5f6973),
	.w4(32'h3a74d487),
	.w5(32'hbb435318),
	.w6(32'hbcb88fd5),
	.w7(32'hbb1f45a0),
	.w8(32'hbbacd5db),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf22803),
	.w1(32'hbb910f14),
	.w2(32'h3b280f71),
	.w3(32'h3b62aa16),
	.w4(32'hba28c39a),
	.w5(32'hb988c818),
	.w6(32'h3a2572fb),
	.w7(32'hb97202df),
	.w8(32'hbc18f70a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4beb93),
	.w1(32'hbc51a165),
	.w2(32'hbc17959a),
	.w3(32'hbc05bf9a),
	.w4(32'hbc609ad6),
	.w5(32'hbc8a90ef),
	.w6(32'hba9b118b),
	.w7(32'hbb14d50d),
	.w8(32'hbca4cdf5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39debb58),
	.w1(32'hbc4b2500),
	.w2(32'h3c59a851),
	.w3(32'h3bedcd1e),
	.w4(32'hbc279d4c),
	.w5(32'h3bb89bff),
	.w6(32'h3bf34bfc),
	.w7(32'hbac1c322),
	.w8(32'h39a65bf1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf52f9),
	.w1(32'hbbde8e24),
	.w2(32'hbc435b36),
	.w3(32'hbba5cca4),
	.w4(32'hbccc6ba3),
	.w5(32'hbbdcb205),
	.w6(32'hbb6b46b4),
	.w7(32'hbc89dfad),
	.w8(32'h3c296db2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2458d),
	.w1(32'hbb161fe1),
	.w2(32'h3ae4fed5),
	.w3(32'hbd199b38),
	.w4(32'hbb394ec2),
	.w5(32'h3a4475bd),
	.w6(32'hbcc4d55c),
	.w7(32'hbc233715),
	.w8(32'h3a4f1994),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42c46f),
	.w1(32'h3c8095e3),
	.w2(32'h3c0f8bf6),
	.w3(32'h3b0a49c8),
	.w4(32'h3c51fee2),
	.w5(32'h3c3b50f7),
	.w6(32'h3b983ff7),
	.w7(32'h3c80fb01),
	.w8(32'h3c4ca5c0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e954c),
	.w1(32'h3b60d046),
	.w2(32'hbc45755c),
	.w3(32'h3ca6264a),
	.w4(32'h3a49d0c3),
	.w5(32'hbc0313df),
	.w6(32'h3c176ad8),
	.w7(32'hbb589726),
	.w8(32'hbb8a8bb6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec6df9),
	.w1(32'h3b786032),
	.w2(32'hbc48e904),
	.w3(32'hbb3f75f8),
	.w4(32'hbc4fb359),
	.w5(32'hbc66ed76),
	.w6(32'hbc3cd8f3),
	.w7(32'hbbdf80e7),
	.w8(32'hbc8dbb20),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28edb0),
	.w1(32'hbb79e803),
	.w2(32'hb6f81381),
	.w3(32'h3c3855f4),
	.w4(32'h3b512af1),
	.w5(32'h377730f6),
	.w6(32'h3bc9ee2d),
	.w7(32'h3b906f5c),
	.w8(32'hba71f301),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e142c),
	.w1(32'hbbd81a09),
	.w2(32'hbc4736d6),
	.w3(32'hbb4ded17),
	.w4(32'hbbc707c2),
	.w5(32'hbb5410dd),
	.w6(32'h3af839f1),
	.w7(32'h3adaf20c),
	.w8(32'h3ad01ea5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8a2fa),
	.w1(32'h39784fe3),
	.w2(32'hbbceb74a),
	.w3(32'hba804ac4),
	.w4(32'h3a157f35),
	.w5(32'hba469adb),
	.w6(32'h3b2216d9),
	.w7(32'hba75a51a),
	.w8(32'h3b25e255),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe9690),
	.w1(32'hbc472904),
	.w2(32'h3c1a5f87),
	.w3(32'hbc08935c),
	.w4(32'h3bd69576),
	.w5(32'h3cb5c2a7),
	.w6(32'hbc11bcb0),
	.w7(32'h3b06a6b0),
	.w8(32'h3cabde11),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbb493),
	.w1(32'hbc87f4f9),
	.w2(32'hbc1e524c),
	.w3(32'h3c8f881a),
	.w4(32'hbc57c84d),
	.w5(32'hbc31fa21),
	.w6(32'h3c65b65b),
	.w7(32'hbc0b62e0),
	.w8(32'hbc3e9410),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b589403),
	.w1(32'hbbd59fb1),
	.w2(32'hbc13b53f),
	.w3(32'h3bfa453f),
	.w4(32'h3b39f95b),
	.w5(32'h3a0c3d9e),
	.w6(32'h3b9a1497),
	.w7(32'h3b15dc5a),
	.w8(32'h3ad9e559),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb693c),
	.w1(32'h3bace5eb),
	.w2(32'hbb587b82),
	.w3(32'h3b7566ef),
	.w4(32'hb96e8efd),
	.w5(32'hbc1c1650),
	.w6(32'hbb04aa52),
	.w7(32'hbbd408e3),
	.w8(32'hbbcf1f56),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39168d83),
	.w1(32'hbb3f9c1e),
	.w2(32'h3b87c78a),
	.w3(32'hbbab635c),
	.w4(32'hbc0dd0f0),
	.w5(32'h3c181cd4),
	.w6(32'hbc319b32),
	.w7(32'hb9da2aa8),
	.w8(32'h3c58f0a1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d80a1),
	.w1(32'hbcad9c61),
	.w2(32'h3ba202cf),
	.w3(32'hbb302b9d),
	.w4(32'hbc9abd23),
	.w5(32'hbb6a16fc),
	.w6(32'hb97a66af),
	.w7(32'hbcbcbab0),
	.w8(32'hbb88721c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e7a9),
	.w1(32'hba3d7e4c),
	.w2(32'hbc483ba7),
	.w3(32'hbaf9e024),
	.w4(32'h3b69e4b8),
	.w5(32'hbc1d309b),
	.w6(32'hb9f012f3),
	.w7(32'h3a232280),
	.w8(32'hbbc59107),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73d665),
	.w1(32'hbc22bf28),
	.w2(32'hb9d5d003),
	.w3(32'h3b53442c),
	.w4(32'h3ba76da5),
	.w5(32'hbc295a81),
	.w6(32'h3a83df0c),
	.w7(32'h3c0e87cf),
	.w8(32'hbc5407f9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397675d6),
	.w1(32'h3c446ffa),
	.w2(32'hbb83d15f),
	.w3(32'hbae10d3f),
	.w4(32'h3c80b275),
	.w5(32'hbc4164c0),
	.w6(32'h3b9fe2aa),
	.w7(32'h3c3fd680),
	.w8(32'hbbc64eb1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb372f8b),
	.w1(32'hbb9643b5),
	.w2(32'hbbdef6eb),
	.w3(32'hbc5b350b),
	.w4(32'hbbc06cb3),
	.w5(32'hbbe4bf5e),
	.w6(32'hbbad760e),
	.w7(32'hbacd7cf8),
	.w8(32'hbc100303),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bd77d),
	.w1(32'hbc9495a2),
	.w2(32'hbcb49e54),
	.w3(32'h3ce2e5f3),
	.w4(32'hbbc181e1),
	.w5(32'hbd0009a6),
	.w6(32'h3caa6319),
	.w7(32'h3bc9288d),
	.w8(32'hbcb8e347),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6bb0d),
	.w1(32'h3d14cd39),
	.w2(32'hbb5bdf9a),
	.w3(32'hbc7904c5),
	.w4(32'h3d2c668d),
	.w5(32'hbbdd4db7),
	.w6(32'hbc67010f),
	.w7(32'h3d1fa025),
	.w8(32'h3a80e4dc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f874),
	.w1(32'hbbade36e),
	.w2(32'h3c00a26f),
	.w3(32'h3b8a34af),
	.w4(32'hbb51ab0e),
	.w5(32'h3bb9381c),
	.w6(32'h3c601805),
	.w7(32'h3c3df3c7),
	.w8(32'hb8a31fe8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe97c9f),
	.w1(32'hbbaf73fa),
	.w2(32'hbcd2397d),
	.w3(32'hbc2b9786),
	.w4(32'hbc956b8f),
	.w5(32'hbcc5052e),
	.w6(32'h3b1aa652),
	.w7(32'hbc039a3d),
	.w8(32'h3b020a42),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc381a54),
	.w1(32'h3c364aa1),
	.w2(32'h3bbca195),
	.w3(32'hbd07ada9),
	.w4(32'hba2f22b8),
	.w5(32'h3b624582),
	.w6(32'hbccc821e),
	.w7(32'h3a2f323b),
	.w8(32'h3bd97098),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c350f58),
	.w1(32'hbb2d3312),
	.w2(32'h3b79d4dc),
	.w3(32'h3cbb4628),
	.w4(32'h3c26459e),
	.w5(32'h3b78af9c),
	.w6(32'h3cb4685f),
	.w7(32'h3b827804),
	.w8(32'h3b349177),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc829e5),
	.w1(32'h3c1d10ac),
	.w2(32'hbae0a9ba),
	.w3(32'hbabe666a),
	.w4(32'h3b9ac315),
	.w5(32'h3a147aac),
	.w6(32'h3be5c917),
	.w7(32'h3b0d7111),
	.w8(32'h3a87d29b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a5ce1),
	.w1(32'h3c2340fc),
	.w2(32'hbbd69ce8),
	.w3(32'h3c595554),
	.w4(32'h3c592228),
	.w5(32'h3b4b644b),
	.w6(32'h39c60489),
	.w7(32'h3c2704bc),
	.w8(32'hbb74152a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83dab2),
	.w1(32'hbbcb8fdd),
	.w2(32'hbc59d28b),
	.w3(32'hbb448069),
	.w4(32'hbae84a4f),
	.w5(32'hbca3f1eb),
	.w6(32'hbbcbcf9d),
	.w7(32'hbb0fa48e),
	.w8(32'hbcb1c038),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c076a27),
	.w1(32'h3cb143a7),
	.w2(32'hbbc926d3),
	.w3(32'h3b68bb44),
	.w4(32'h3cb1591b),
	.w5(32'hbbe7b7f5),
	.w6(32'hb9cf8819),
	.w7(32'h3c67a6f2),
	.w8(32'hbc336537),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50149d),
	.w1(32'hbbe6792c),
	.w2(32'h396db190),
	.w3(32'h3c82246e),
	.w4(32'h3ac1503b),
	.w5(32'hbb02d260),
	.w6(32'h3c4f5f7d),
	.w7(32'h3bae4af6),
	.w8(32'hbbad8848),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd68e8f),
	.w1(32'hbc8c924d),
	.w2(32'hbbf9032d),
	.w3(32'hbc593570),
	.w4(32'hbc983c39),
	.w5(32'hbc077730),
	.w6(32'hbc751b16),
	.w7(32'hbc7ea718),
	.w8(32'hbbff36c9),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f722),
	.w1(32'hb9bc9f4a),
	.w2(32'h3b533107),
	.w3(32'hbb342d37),
	.w4(32'h3b10cdc2),
	.w5(32'h3b557e33),
	.w6(32'hbb05bdc4),
	.w7(32'h3ab6d27f),
	.w8(32'h3b774174),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a9191),
	.w1(32'hbbdeaf96),
	.w2(32'h3ca4adeb),
	.w3(32'hbb860be6),
	.w4(32'hbbe38e21),
	.w5(32'h3d16f8ad),
	.w6(32'h3ac2681a),
	.w7(32'hbb128a1b),
	.w8(32'h3d147245),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fb3b4),
	.w1(32'hbce5f78d),
	.w2(32'hbc3f4c80),
	.w3(32'hbb1d8891),
	.w4(32'hbd35e1ed),
	.w5(32'hbcdb3d24),
	.w6(32'h3c80c055),
	.w7(32'hbcec1763),
	.w8(32'hbcbbcf35),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dcd31),
	.w1(32'h3ca27d0b),
	.w2(32'hbc0fb836),
	.w3(32'hbb900a14),
	.w4(32'h3cb8884f),
	.w5(32'hbbe914fd),
	.w6(32'hbba1252a),
	.w7(32'h3c3348e1),
	.w8(32'hbc0f13ec),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3aafe),
	.w1(32'hbc4ce3ec),
	.w2(32'hbc3173da),
	.w3(32'hbb95a4d7),
	.w4(32'hbc714502),
	.w5(32'hbca33381),
	.w6(32'hbb8771f5),
	.w7(32'hbc9f0615),
	.w8(32'hbc84da85),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a696ba3),
	.w1(32'hbc07b81c),
	.w2(32'h3b0820fd),
	.w3(32'h3adb438d),
	.w4(32'hbbcbafe3),
	.w5(32'h3a0856e0),
	.w6(32'hbadd5b49),
	.w7(32'h39ab517b),
	.w8(32'h3b94f569),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72801f),
	.w1(32'hbb81d089),
	.w2(32'hbc32cf95),
	.w3(32'hb9fa9f56),
	.w4(32'hbb3c4ad5),
	.w5(32'hbc291d4a),
	.w6(32'h3b4d1230),
	.w7(32'h3b3279cf),
	.w8(32'hbc0661de),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc283dda),
	.w1(32'hba3f31cb),
	.w2(32'h3bcd190c),
	.w3(32'h3a391360),
	.w4(32'h3b9db70d),
	.w5(32'h3b9ffa14),
	.w6(32'h3b0f6706),
	.w7(32'h3c2bb91f),
	.w8(32'h3bae98ad),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa86c9e),
	.w1(32'h3bfbe924),
	.w2(32'hbb0102ec),
	.w3(32'h3a360eee),
	.w4(32'h3c1462ba),
	.w5(32'hbbdc4516),
	.w6(32'hbb4feb04),
	.w7(32'hbb25c364),
	.w8(32'hbb76e1a2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5256d),
	.w1(32'h3b84a2f8),
	.w2(32'hbbd84b9a),
	.w3(32'hbad03b88),
	.w4(32'hbb489f37),
	.w5(32'hbc27a56d),
	.w6(32'hbb4ec9c1),
	.w7(32'h3bcb9757),
	.w8(32'hbc132f28),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132824),
	.w1(32'hba7e6e73),
	.w2(32'h39806929),
	.w3(32'h3bd67202),
	.w4(32'h3c34a422),
	.w5(32'h3b39070d),
	.w6(32'hbbc35da7),
	.w7(32'h3c4eb408),
	.w8(32'h3b8b83ba),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb000bf3),
	.w1(32'h39842bb8),
	.w2(32'h3b4dd775),
	.w3(32'hba16dd47),
	.w4(32'hba3134d2),
	.w5(32'h3c527ce2),
	.w6(32'hb994283c),
	.w7(32'h3a46ace9),
	.w8(32'h3c84b0cc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91bf51),
	.w1(32'hbd074f35),
	.w2(32'hbbfc56e1),
	.w3(32'hbc197084),
	.w4(32'hbd2237a8),
	.w5(32'hbbdb6c57),
	.w6(32'h3b1ba37e),
	.w7(32'hbcc71f3d),
	.w8(32'hbb8d76c7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb339d7e),
	.w1(32'hbb684b73),
	.w2(32'h3b3498cb),
	.w3(32'hbab6fa20),
	.w4(32'hbb7c149e),
	.w5(32'hb98fbc84),
	.w6(32'h3b02388b),
	.w7(32'hbaff11a9),
	.w8(32'hbb22927d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbe58a),
	.w1(32'hbbc6dcab),
	.w2(32'hbbd465e1),
	.w3(32'h39aceece),
	.w4(32'hbc047682),
	.w5(32'hbb45ffaa),
	.w6(32'h3b7589c4),
	.w7(32'hbc3bc559),
	.w8(32'hbc19077a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb927c0c),
	.w1(32'h3adf389e),
	.w2(32'hbbb41f27),
	.w3(32'h3c3f6d4d),
	.w4(32'hbc1e3a90),
	.w5(32'hbc2839e0),
	.w6(32'h3c93b9e8),
	.w7(32'hba57db5f),
	.w8(32'hb4903800),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44abe1),
	.w1(32'hbc598736),
	.w2(32'h3c09a49a),
	.w3(32'hba9d2724),
	.w4(32'hbb220722),
	.w5(32'hbb9570ce),
	.w6(32'h3bd72192),
	.w7(32'h3b222eac),
	.w8(32'hbc48eb10),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabb1f4),
	.w1(32'h3c3ad6d1),
	.w2(32'hbcdc12d8),
	.w3(32'h3cfd7674),
	.w4(32'h3c908546),
	.w5(32'hbd17afb0),
	.w6(32'h3c58ca4e),
	.w7(32'h3c6f4cc5),
	.w8(32'hbd0a716a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1e9c1),
	.w1(32'h3c9889ee),
	.w2(32'hbba2ce3c),
	.w3(32'h3acf4f31),
	.w4(32'h3c97f9ae),
	.w5(32'hbaa71327),
	.w6(32'h39bcad00),
	.w7(32'h3ca1fd29),
	.w8(32'h3ab0802c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac0c9d),
	.w1(32'hbbd31129),
	.w2(32'h3aa24aa7),
	.w3(32'hbb01fbe3),
	.w4(32'hbb673786),
	.w5(32'hbbaf1a4b),
	.w6(32'h3a4ecfcc),
	.w7(32'hbb1502f5),
	.w8(32'hbc2740a5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9123b8),
	.w1(32'h3b3d2cf0),
	.w2(32'hbbe15a3a),
	.w3(32'hbc0d935d),
	.w4(32'hbc0ad730),
	.w5(32'hbb590127),
	.w6(32'h3aa32252),
	.w7(32'hba509d15),
	.w8(32'hbb5729d4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9a688),
	.w1(32'h3c339e87),
	.w2(32'hbc275b75),
	.w3(32'hbbb546c0),
	.w4(32'hbb27e5b4),
	.w5(32'hbced6de9),
	.w6(32'h3c6c4a85),
	.w7(32'h3c6ff38b),
	.w8(32'hbc9f229e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ddb26),
	.w1(32'hbb8ca9dc),
	.w2(32'hbc6da731),
	.w3(32'hbc2cfa38),
	.w4(32'hba83112f),
	.w5(32'hbc968740),
	.w6(32'hbbcdee4f),
	.w7(32'h3c09b2fc),
	.w8(32'hbb534880),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74a387),
	.w1(32'h3c366c74),
	.w2(32'h3b5fa076),
	.w3(32'hbd059ec3),
	.w4(32'hbb7a39be),
	.w5(32'h3bd0614f),
	.w6(32'hbcab0f3e),
	.w7(32'hb9361067),
	.w8(32'h3c09767f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbad010),
	.w1(32'h3baa96eb),
	.w2(32'h3bd78588),
	.w3(32'h3bd4db1c),
	.w4(32'h3bfa8278),
	.w5(32'h3be0c9c2),
	.w6(32'h3bd31d56),
	.w7(32'h3c0a3c15),
	.w8(32'h3c0d52f6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0776b3),
	.w1(32'hbb2d77ef),
	.w2(32'hbbae247a),
	.w3(32'hbc271bcd),
	.w4(32'hbb2f195f),
	.w5(32'hbc0fe412),
	.w6(32'hbbd6ac25),
	.w7(32'hbb1f498a),
	.w8(32'h3ab2256f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980f8cd),
	.w1(32'h3b870e15),
	.w2(32'h3c0be353),
	.w3(32'hbb2e466b),
	.w4(32'hba7924fa),
	.w5(32'h3ba4e625),
	.w6(32'hbc004274),
	.w7(32'hbafeea9b),
	.w8(32'h3b9331d3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be904c8),
	.w1(32'h3b029f3d),
	.w2(32'hbc09634f),
	.w3(32'hbb350473),
	.w4(32'h3aa36b49),
	.w5(32'h3a7d7a8c),
	.w6(32'hbba67367),
	.w7(32'hba991300),
	.w8(32'hbb8fb8cd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab82f),
	.w1(32'hbc8ae652),
	.w2(32'hbbc95d16),
	.w3(32'h3c1f80f2),
	.w4(32'hbb78f829),
	.w5(32'hbbb72d38),
	.w6(32'h3bbde705),
	.w7(32'hba9ecd3e),
	.w8(32'hbb908dcc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49a6b0),
	.w1(32'hbb71be67),
	.w2(32'hbaecdd82),
	.w3(32'hbbd42b5d),
	.w4(32'hbc48e0ea),
	.w5(32'hbba9dab3),
	.w6(32'hbb8d5c1f),
	.w7(32'hbc580288),
	.w8(32'hbaa90d75),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcf6b9),
	.w1(32'hba7bd651),
	.w2(32'h3c948701),
	.w3(32'h3bfadf62),
	.w4(32'h3b07c332),
	.w5(32'h3cc7204e),
	.w6(32'h3be8161a),
	.w7(32'hb89e1bf5),
	.w8(32'h3c8f3255),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90122c),
	.w1(32'hbca0c37f),
	.w2(32'hbbc25478),
	.w3(32'h3c4c0bd6),
	.w4(32'hbcd467a7),
	.w5(32'hbba27084),
	.w6(32'h3cc1d0d4),
	.w7(32'hbc441ec7),
	.w8(32'hbc08d2e0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f5bba),
	.w1(32'hbbd631e2),
	.w2(32'h3a2a7daf),
	.w3(32'hbad4f92f),
	.w4(32'hbb7a7752),
	.w5(32'hbb83e7c3),
	.w6(32'hba6d4be0),
	.w7(32'hb9df9a58),
	.w8(32'hbc48db1f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22c07),
	.w1(32'hbba0390a),
	.w2(32'hbab9c1ba),
	.w3(32'hbaf49f18),
	.w4(32'hba153546),
	.w5(32'hbbc6df61),
	.w6(32'hbbf8effe),
	.w7(32'h3b401913),
	.w8(32'hbc0e912c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea3cd6),
	.w1(32'h3a9c9152),
	.w2(32'h3bbf9f84),
	.w3(32'h3bc18e5c),
	.w4(32'hbb08ca6c),
	.w5(32'h3c12d2d1),
	.w6(32'h3c3679b7),
	.w7(32'h3bac845a),
	.w8(32'h3c8af60b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d71a),
	.w1(32'hbc0b8fac),
	.w2(32'h3c485c44),
	.w3(32'h3a1fff37),
	.w4(32'hbc35e1ef),
	.w5(32'h3c0a8868),
	.w6(32'h3c819709),
	.w7(32'hbc3d40b2),
	.w8(32'h3c4202ae),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb14d72),
	.w1(32'hbb8a1c54),
	.w2(32'hbbf07734),
	.w3(32'h3c006f5b),
	.w4(32'hba3d555c),
	.w5(32'hbc96f068),
	.w6(32'h3c2b050e),
	.w7(32'hbba6787d),
	.w8(32'hbc41f333),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3bc70),
	.w1(32'h3be547d2),
	.w2(32'hbc583fe3),
	.w3(32'hb94bcf51),
	.w4(32'h3c4c0691),
	.w5(32'hbc852e6c),
	.w6(32'hbb719ef8),
	.w7(32'h3c83a3eb),
	.w8(32'hbc458f2f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bac87),
	.w1(32'h39fb0b7a),
	.w2(32'h3c06be38),
	.w3(32'h3bcb9c51),
	.w4(32'h3c1e5f51),
	.w5(32'h3cc1a6df),
	.w6(32'h3bea2f55),
	.w7(32'h3c35d7c1),
	.w8(32'h3c7f199e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd44b7b),
	.w1(32'hbcd9892a),
	.w2(32'hbabf4c84),
	.w3(32'h3c5ae80a),
	.w4(32'hbcdad226),
	.w5(32'h3bf31523),
	.w6(32'h3c63bb2e),
	.w7(32'hbba5b85d),
	.w8(32'hbc07a2e0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc295533),
	.w1(32'hbc435006),
	.w2(32'hbb60ffa3),
	.w3(32'hbb8f9899),
	.w4(32'hbc65e5be),
	.w5(32'h3b0c9680),
	.w6(32'hbb1258a6),
	.w7(32'hbc23b4e2),
	.w8(32'hbb86b70e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda267e),
	.w1(32'hb9de38f0),
	.w2(32'hbb90fa16),
	.w3(32'h3c606ac6),
	.w4(32'h3bdc33a4),
	.w5(32'hbb552d74),
	.w6(32'h3b96eb04),
	.w7(32'h3ae5a6e1),
	.w8(32'hbb85a88f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de96c),
	.w1(32'h3c3e62f9),
	.w2(32'h3bddd895),
	.w3(32'h3888dd1f),
	.w4(32'hbb8a14f5),
	.w5(32'h3c565a58),
	.w6(32'hbba7a6cb),
	.w7(32'hbb9ebabd),
	.w8(32'h3c27ff3b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf04e3e),
	.w1(32'hbcbd7042),
	.w2(32'hbbf58058),
	.w3(32'h3c3d3007),
	.w4(32'hbcb56bf3),
	.w5(32'h3adf96c1),
	.w6(32'h39331d05),
	.w7(32'hbc8e9036),
	.w8(32'hba113895),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22b971),
	.w1(32'hbc2bb6fc),
	.w2(32'hbc44bd47),
	.w3(32'h3c658607),
	.w4(32'hbb2f56b3),
	.w5(32'hbab7fcfc),
	.w6(32'h3c211d40),
	.w7(32'hbb8e206c),
	.w8(32'h3b715f9b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d04bc),
	.w1(32'hbc214124),
	.w2(32'hbc277e6a),
	.w3(32'h3aae9af7),
	.w4(32'hbc484c55),
	.w5(32'h3b8d345f),
	.w6(32'h3b97035a),
	.w7(32'hbbe16283),
	.w8(32'hbb91b137),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07abb3),
	.w1(32'hbb1e71f6),
	.w2(32'h3c825772),
	.w3(32'h3c21a139),
	.w4(32'h3b5604d9),
	.w5(32'h3ca4d576),
	.w6(32'h3c04b408),
	.w7(32'hb9c31449),
	.w8(32'h3c8adef6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380b6c),
	.w1(32'hbc60e5bb),
	.w2(32'hbc7a44da),
	.w3(32'hbb2bb74b),
	.w4(32'hbca2e7a7),
	.w5(32'hbc6da9e1),
	.w6(32'hbaa2f3a1),
	.w7(32'hbc4a86f5),
	.w8(32'hbc550c8f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55473f),
	.w1(32'h3c21eb12),
	.w2(32'h3b3cabaf),
	.w3(32'h3b9fb489),
	.w4(32'h3ce2f8b5),
	.w5(32'h3bbbba9b),
	.w6(32'hbc3c58cd),
	.w7(32'h3c331ffc),
	.w8(32'h3a9c1862),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa691d3),
	.w1(32'hbb82a876),
	.w2(32'hbaa009bd),
	.w3(32'h3a2ca56a),
	.w4(32'hbc2f6ca8),
	.w5(32'h3bb65bad),
	.w6(32'hbb879a0f),
	.w7(32'hbc09c138),
	.w8(32'h3a41e41f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d4a9),
	.w1(32'hbc56efc0),
	.w2(32'hbc61f1da),
	.w3(32'hbbf630c9),
	.w4(32'hbc0fc3a2),
	.w5(32'hbb14d4bc),
	.w6(32'hbb93a0df),
	.w7(32'hbb72c89e),
	.w8(32'hbac1fef5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97e7ab),
	.w1(32'hbb87e852),
	.w2(32'h3c061d64),
	.w3(32'hbb85df72),
	.w4(32'hbab5ab68),
	.w5(32'h39751171),
	.w6(32'hbb367f52),
	.w7(32'hbb197c6e),
	.w8(32'h3ad029b4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accc7bf),
	.w1(32'h3b981d45),
	.w2(32'h3b7500a7),
	.w3(32'h3b02f9ca),
	.w4(32'hbb01b4e4),
	.w5(32'h3b8d40fe),
	.w6(32'hbb3d300b),
	.w7(32'hbb91df68),
	.w8(32'h3b8bd930),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab46858),
	.w1(32'hbb6dee57),
	.w2(32'hbafbc582),
	.w3(32'hbb29ce13),
	.w4(32'hbb8e0e88),
	.w5(32'hba04bfd8),
	.w6(32'hbb1e0dbe),
	.w7(32'hbb66c250),
	.w8(32'h3b1563d6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6230f6),
	.w1(32'h3a137c98),
	.w2(32'hbcbaf4a1),
	.w3(32'hbb9451ac),
	.w4(32'hba467776),
	.w5(32'hbd2173a5),
	.w6(32'hbb7b6549),
	.w7(32'h39c32c87),
	.w8(32'hbce244bc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56726e),
	.w1(32'hbb99f5c1),
	.w2(32'hbc250a2b),
	.w3(32'hbc8ff317),
	.w4(32'h3c49fd84),
	.w5(32'hbc6b5561),
	.w6(32'hbca951db),
	.w7(32'h3c2e36fd),
	.w8(32'hbc6b8692),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8207d9),
	.w1(32'h3c2ea63e),
	.w2(32'hb9ff09c4),
	.w3(32'h3a3cdaa0),
	.w4(32'h3c4eadb6),
	.w5(32'hbc0376bc),
	.w6(32'hbb3b1ca2),
	.w7(32'h3c6e73da),
	.w8(32'hbbac8b00),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc142cc8),
	.w1(32'hbc4d9250),
	.w2(32'hbce66b05),
	.w3(32'hbc43ba39),
	.w4(32'hbbae1fef),
	.w5(32'hbc93da20),
	.w6(32'hbc5b22c0),
	.w7(32'h3b77230e),
	.w8(32'hbc02e62e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17c2a1),
	.w1(32'hbc38fc92),
	.w2(32'hbc2f3959),
	.w3(32'h3b9e5641),
	.w4(32'hbc80aa73),
	.w5(32'hbc0a1791),
	.w6(32'hbb323e14),
	.w7(32'hbc3481d1),
	.w8(32'hbc28bbce),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabef00c),
	.w1(32'hbbc4dd79),
	.w2(32'hba34c0b7),
	.w3(32'h39bc91c5),
	.w4(32'hbbf9c4fb),
	.w5(32'h3b8ceffb),
	.w6(32'h3a1f2f9f),
	.w7(32'hbaf36c8a),
	.w8(32'h3b4365a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule