module layer_10_featuremap_477(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023298),
	.w1(32'h3a3e683f),
	.w2(32'hba12a3bb),
	.w3(32'h3b7d9bd0),
	.w4(32'hba3ebf45),
	.w5(32'h374ffe89),
	.w6(32'hbaaf094a),
	.w7(32'hba018e97),
	.w8(32'h3acc9a40),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eaf8e),
	.w1(32'hb9230d65),
	.w2(32'hbbaf9179),
	.w3(32'hba90363c),
	.w4(32'hbb55b28b),
	.w5(32'hbb8632a9),
	.w6(32'h3abfcbeb),
	.w7(32'hbb845689),
	.w8(32'hba3c219f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad23c01),
	.w1(32'hba4fa140),
	.w2(32'hbabcf5fe),
	.w3(32'h3b1e2326),
	.w4(32'hb9885732),
	.w5(32'hbb8c7540),
	.w6(32'h3b2cf234),
	.w7(32'hbad0689b),
	.w8(32'hba09ffab),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3c33f),
	.w1(32'hb97cca32),
	.w2(32'hb9833db9),
	.w3(32'h3b815b44),
	.w4(32'hbb5f93c2),
	.w5(32'h3aea8185),
	.w6(32'h3b95ae83),
	.w7(32'hba3f742b),
	.w8(32'hb8c2e27c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9633d6a),
	.w1(32'h3b9f783e),
	.w2(32'h3b19e3e3),
	.w3(32'h3b948a71),
	.w4(32'h3a027d79),
	.w5(32'h3ba371f5),
	.w6(32'hba04eaff),
	.w7(32'hbb22c31e),
	.w8(32'h3a966059),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb1eaf),
	.w1(32'hbb0436dd),
	.w2(32'hbb11ce9d),
	.w3(32'hb90390d1),
	.w4(32'h3a1598cc),
	.w5(32'h3a12dfe1),
	.w6(32'h3b1853d4),
	.w7(32'hbaebc365),
	.w8(32'hbb6554f7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9ee6f),
	.w1(32'h3a7b1e37),
	.w2(32'h3c0e9d7e),
	.w3(32'h3b0ad16e),
	.w4(32'h3c033159),
	.w5(32'h3c48b05c),
	.w6(32'h3b788c4b),
	.w7(32'h3c25bb92),
	.w8(32'h3c5a10f0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178fb0),
	.w1(32'hbc591bad),
	.w2(32'hbbd001fc),
	.w3(32'h3b94bff3),
	.w4(32'h3b5427ae),
	.w5(32'hbc0768cb),
	.w6(32'hba1b7eeb),
	.w7(32'hbade221f),
	.w8(32'hbbba0a94),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5537be),
	.w1(32'hbb7dd3e5),
	.w2(32'hb9ff5e63),
	.w3(32'h3ac52a44),
	.w4(32'hbb594a8e),
	.w5(32'h3acf6181),
	.w6(32'h3ab30293),
	.w7(32'hbb8bc744),
	.w8(32'hbbccedd5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a2eb),
	.w1(32'h3b86a472),
	.w2(32'h3bc20a72),
	.w3(32'hbbb4fb31),
	.w4(32'h3a846ff9),
	.w5(32'h3acc1503),
	.w6(32'hbbc53c58),
	.w7(32'h3b879d74),
	.w8(32'h3be91ce2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a397a99),
	.w1(32'h3ab77f12),
	.w2(32'h3b0201f8),
	.w3(32'hbb451a33),
	.w4(32'h3ac92c5c),
	.w5(32'h3c1ef5e0),
	.w6(32'h3a327f3b),
	.w7(32'h3b698d26),
	.w8(32'h3ba20d7f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885a73),
	.w1(32'h3b5d53c1),
	.w2(32'h3c8156f5),
	.w3(32'h3b69c2a8),
	.w4(32'h3a180213),
	.w5(32'h3c733a36),
	.w6(32'h3c00db36),
	.w7(32'h3ba70b71),
	.w8(32'h3c3467bf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c43ad),
	.w1(32'hb982e0cd),
	.w2(32'h3bca43b6),
	.w3(32'h3914d6f3),
	.w4(32'h3b0d5e52),
	.w5(32'h3bb24af1),
	.w6(32'hbb8da863),
	.w7(32'h3b28219f),
	.w8(32'h3adf8508),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89a471),
	.w1(32'h3c24dfe8),
	.w2(32'h3af0f03d),
	.w3(32'h3b227a15),
	.w4(32'h3b9eb6b6),
	.w5(32'h3aa6618d),
	.w6(32'hba682cac),
	.w7(32'h3abcdc16),
	.w8(32'h3bfcf93a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadae456),
	.w1(32'hbb0c640f),
	.w2(32'hbbe48567),
	.w3(32'hbaf163a1),
	.w4(32'hbbaa8f35),
	.w5(32'hba2f00ab),
	.w6(32'h3aba5f33),
	.w7(32'hbbaeab81),
	.w8(32'hbb8c585c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab218b2),
	.w1(32'hbb1cb9e2),
	.w2(32'hbbc061cc),
	.w3(32'hbbfa1e5b),
	.w4(32'hbbd87f43),
	.w5(32'hbb47c01f),
	.w6(32'hbb51a877),
	.w7(32'hbbd4ebe2),
	.w8(32'hbbe7be9c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b502ab7),
	.w1(32'h3a95d1f7),
	.w2(32'hb9d9b3d3),
	.w3(32'hba7e3601),
	.w4(32'hbb2ac53f),
	.w5(32'hbb1d4d8a),
	.w6(32'hb9c8f046),
	.w7(32'h3add5e41),
	.w8(32'h3b02d46a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b040),
	.w1(32'h3bcdc732),
	.w2(32'h3c539ea4),
	.w3(32'hbae37e43),
	.w4(32'h3ba7f798),
	.w5(32'h3ba5d104),
	.w6(32'h3ba8f5ec),
	.w7(32'h3c3b2899),
	.w8(32'h3a0c9b64),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dd776),
	.w1(32'h3b0eebbc),
	.w2(32'h3c3ebbc8),
	.w3(32'hbb53ebf3),
	.w4(32'h3b09250e),
	.w5(32'h3c831328),
	.w6(32'h395db098),
	.w7(32'h3b86317d),
	.w8(32'h3b349216),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d66bb4),
	.w1(32'hbb12fdfe),
	.w2(32'hba4731af),
	.w3(32'hbae3b367),
	.w4(32'hbb2600eb),
	.w5(32'h3a88a18e),
	.w6(32'hbaa2d6f2),
	.w7(32'h39c5dcc0),
	.w8(32'hbb510b26),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1047c9),
	.w1(32'hb97eaf4f),
	.w2(32'h3b09ce9f),
	.w3(32'h38934e75),
	.w4(32'h39db72bc),
	.w5(32'h38a88b36),
	.w6(32'hbb5a72e7),
	.w7(32'hb9fb62b4),
	.w8(32'h39d58a64),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec8dda),
	.w1(32'hbb0b4a2c),
	.w2(32'h3a709107),
	.w3(32'h3b0e1583),
	.w4(32'hba955a80),
	.w5(32'hb9f16872),
	.w6(32'h3b2ad2f2),
	.w7(32'hba883462),
	.w8(32'hbaea6dd6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc398429),
	.w1(32'hb9c37707),
	.w2(32'h3c643944),
	.w3(32'hbc084bf4),
	.w4(32'hbbbd08fb),
	.w5(32'h3bfdc45b),
	.w6(32'hbacb1903),
	.w7(32'h3c2a2137),
	.w8(32'h3c36638c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b0655),
	.w1(32'hbad05c34),
	.w2(32'hbb47eeb6),
	.w3(32'hbbb277fb),
	.w4(32'hbb141ec0),
	.w5(32'hbb8496dc),
	.w6(32'hbb98089c),
	.w7(32'hbbfca166),
	.w8(32'hbbcf0990),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4e9d9),
	.w1(32'hbb059131),
	.w2(32'hbc01c465),
	.w3(32'h39d1d942),
	.w4(32'hbb1843a6),
	.w5(32'hbc433a8b),
	.w6(32'hbbd44723),
	.w7(32'hbbe875b7),
	.w8(32'hbc367e9c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb3051),
	.w1(32'hb85218ba),
	.w2(32'hb98c3baf),
	.w3(32'hbb48317d),
	.w4(32'h3ae7e558),
	.w5(32'hbb024b33),
	.w6(32'h3a5ef92d),
	.w7(32'hbb6301cc),
	.w8(32'hbb406608),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8b124),
	.w1(32'hbb00b997),
	.w2(32'h3b1a4c90),
	.w3(32'h3b005e57),
	.w4(32'h3abe7a78),
	.w5(32'h3a5ed43d),
	.w6(32'hbbcc1aa2),
	.w7(32'hbb068239),
	.w8(32'hbb1e164f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfca3f0),
	.w1(32'h3c3fbfd5),
	.w2(32'h3c3d6cb3),
	.w3(32'h3b6218b0),
	.w4(32'h3c13a107),
	.w5(32'h3c6eee8d),
	.w6(32'h3b896d79),
	.w7(32'h3b4a1a1e),
	.w8(32'h3c029b06),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51c726),
	.w1(32'hbb5160c8),
	.w2(32'hbaddea94),
	.w3(32'hbb3aa2e9),
	.w4(32'hba9f05b0),
	.w5(32'hbb078b33),
	.w6(32'hba8153e7),
	.w7(32'h3a03efa2),
	.w8(32'hb9ff5459),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb52dad),
	.w1(32'h3b2e94ea),
	.w2(32'hbc1ca52e),
	.w3(32'h3bf1c6e2),
	.w4(32'h3b62861f),
	.w5(32'hbb584ae1),
	.w6(32'h3bc6f66a),
	.w7(32'h3a4902f8),
	.w8(32'h39ca046a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0ddd),
	.w1(32'h3b1363ee),
	.w2(32'h3b4c998c),
	.w3(32'hb8c47f93),
	.w4(32'h3b3a0bee),
	.w5(32'h3a6a68d8),
	.w6(32'hba9cd780),
	.w7(32'h3b0f550e),
	.w8(32'h3b00a918),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a460f44),
	.w1(32'hbb4fb951),
	.w2(32'hbb0420cc),
	.w3(32'h3b005fb8),
	.w4(32'h3a1db78a),
	.w5(32'hbb86a5b3),
	.w6(32'h393ed00f),
	.w7(32'hba8f2937),
	.w8(32'hbb2ea120),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a901bb0),
	.w1(32'h3a201b4c),
	.w2(32'h3bd3c5a5),
	.w3(32'hbb01dce1),
	.w4(32'h376e1833),
	.w5(32'hbb0452da),
	.w6(32'hbb3643c6),
	.w7(32'h3b72d736),
	.w8(32'h3bd1f921),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ce9c),
	.w1(32'hbb754f24),
	.w2(32'hbbcd5cd4),
	.w3(32'hb9d28a82),
	.w4(32'hbb8969a8),
	.w5(32'hbbdcef15),
	.w6(32'hbaedc1e2),
	.w7(32'hba012e39),
	.w8(32'hbb01c821),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e71a),
	.w1(32'h3af463fc),
	.w2(32'h3acdb457),
	.w3(32'hbb141aeb),
	.w4(32'h3a8d1677),
	.w5(32'hbb279dcc),
	.w6(32'h39dcb0c7),
	.w7(32'h3b0db51e),
	.w8(32'h3b6de2cb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f366d8),
	.w1(32'hb9e6306d),
	.w2(32'h3b8fc911),
	.w3(32'h3b3a5b2e),
	.w4(32'hb92709ec),
	.w5(32'h3b680d1b),
	.w6(32'hbaad36aa),
	.w7(32'h3ad2a5b6),
	.w8(32'h3b73f9d0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4f2d8),
	.w1(32'hbc92dd01),
	.w2(32'h3c07181a),
	.w3(32'hbc22b969),
	.w4(32'hbccc0cd9),
	.w5(32'h3c574895),
	.w6(32'hbbee4537),
	.w7(32'hbc4a9629),
	.w8(32'h3c1494d4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd78416),
	.w1(32'h38d71ace),
	.w2(32'hbc03ed57),
	.w3(32'h3b14791f),
	.w4(32'h3abcbc87),
	.w5(32'hbc1f4c4d),
	.w6(32'h3c0b8717),
	.w7(32'hbb22e892),
	.w8(32'hbbddad88),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8400f9),
	.w1(32'h3ca23e59),
	.w2(32'h3c2dc7b3),
	.w3(32'h3c626382),
	.w4(32'h3c97c188),
	.w5(32'h3c65b700),
	.w6(32'h3baca119),
	.w7(32'h3bc2dca8),
	.w8(32'hbae5efd6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40f543),
	.w1(32'hb9f61a47),
	.w2(32'hbaf4a055),
	.w3(32'h3b52fc72),
	.w4(32'h3ad3ecd8),
	.w5(32'hba99f3cc),
	.w6(32'h3b4028ce),
	.w7(32'h3a8ee778),
	.w8(32'hbb273f6c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b36e4),
	.w1(32'h3bec9833),
	.w2(32'hbafb6f2a),
	.w3(32'h3ab1cb21),
	.w4(32'hb9045115),
	.w5(32'hbba9b19a),
	.w6(32'hba681215),
	.w7(32'h3ae8f6bb),
	.w8(32'h3be51442),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba388df7),
	.w1(32'h39d52205),
	.w2(32'h3a8fbc07),
	.w3(32'hba1e1a63),
	.w4(32'hbb83309e),
	.w5(32'h3c0a279e),
	.w6(32'h393cd268),
	.w7(32'hbaec1aec),
	.w8(32'hbb8d9ffb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1df36),
	.w1(32'hbaa81c01),
	.w2(32'h39c31afc),
	.w3(32'hb8574c25),
	.w4(32'hbb837f22),
	.w5(32'h3b5326bb),
	.w6(32'h3a052d47),
	.w7(32'hba57c02e),
	.w8(32'h3a8ce57b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57f8b3),
	.w1(32'h3c01ca5c),
	.w2(32'h3c181381),
	.w3(32'h3b9f6b57),
	.w4(32'h3c188d0c),
	.w5(32'h3c697741),
	.w6(32'h3b39cd0d),
	.w7(32'h3b9ecbf9),
	.w8(32'h3b89038a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41cbd1),
	.w1(32'h3a4770dc),
	.w2(32'h3a336150),
	.w3(32'hba3195c8),
	.w4(32'hbac81771),
	.w5(32'hb9200987),
	.w6(32'hbb2f34f7),
	.w7(32'hbba4eb90),
	.w8(32'hbb993b60),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09432d),
	.w1(32'hbb023693),
	.w2(32'h3a8d2bdc),
	.w3(32'hbbf93ac5),
	.w4(32'hbb4a92e7),
	.w5(32'hb932e490),
	.w6(32'hbbfb0d72),
	.w7(32'hbb44d792),
	.w8(32'h3b07300f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34f12),
	.w1(32'hb95025d9),
	.w2(32'hbad147e9),
	.w3(32'hbabb7111),
	.w4(32'h39ce2ff0),
	.w5(32'hbba5defd),
	.w6(32'hba2ea7e4),
	.w7(32'hbaf5d4bf),
	.w8(32'h3a3c055f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d85e6),
	.w1(32'h3bce17f9),
	.w2(32'h3c9428c9),
	.w3(32'hba087191),
	.w4(32'h3c14cca6),
	.w5(32'h3c812607),
	.w6(32'h3b6d96bf),
	.w7(32'h3c6900ca),
	.w8(32'h3c5786fc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae920d0),
	.w1(32'hba97d570),
	.w2(32'h3ae04d65),
	.w3(32'hba48a86a),
	.w4(32'hb8037fa1),
	.w5(32'h39cfc114),
	.w6(32'hbacb01ef),
	.w7(32'h3b7f7bea),
	.w8(32'h3bb8042c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bbf87),
	.w1(32'h3a39ce44),
	.w2(32'hbb7b453d),
	.w3(32'h3afa092b),
	.w4(32'h3a8de8a3),
	.w5(32'hbb463052),
	.w6(32'h3b960ded),
	.w7(32'h3bb95209),
	.w8(32'h3b30ab33),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fafef),
	.w1(32'hbb06a64e),
	.w2(32'hbb1426ee),
	.w3(32'h3ae81caa),
	.w4(32'h3a010cf0),
	.w5(32'h3ab5126d),
	.w6(32'h3a9d739b),
	.w7(32'h3a155663),
	.w8(32'h3ad67fea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4a439),
	.w1(32'h3bdc67f2),
	.w2(32'h3bdcd32f),
	.w3(32'h3b6b9df9),
	.w4(32'hbb45a56b),
	.w5(32'hbb830c0c),
	.w6(32'h3b0777e5),
	.w7(32'h3a9f6aea),
	.w8(32'h3aa37f82),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2ac7e),
	.w1(32'hbb4f6eae),
	.w2(32'hb917446c),
	.w3(32'hba6396ec),
	.w4(32'h3b048d89),
	.w5(32'hb9d8568b),
	.w6(32'h3a9bee75),
	.w7(32'h3a6be1d9),
	.w8(32'h3a93e5dd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c9287),
	.w1(32'hbb690777),
	.w2(32'h3c166a50),
	.w3(32'h37ba3388),
	.w4(32'h3bfd13e8),
	.w5(32'h3baa0334),
	.w6(32'hba928dac),
	.w7(32'h3c07d6b4),
	.w8(32'h3c100118),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba41fcd),
	.w1(32'hbac0b5fd),
	.w2(32'h3aa2c96e),
	.w3(32'h3b22493e),
	.w4(32'h3acf8968),
	.w5(32'h3a6237fa),
	.w6(32'h3ad1bde9),
	.w7(32'h3add5744),
	.w8(32'h3a34339b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1542d5),
	.w1(32'hbb326e1d),
	.w2(32'h3b0ff74b),
	.w3(32'hbab616b4),
	.w4(32'h3a25cace),
	.w5(32'hb9253739),
	.w6(32'h3a33c71a),
	.w7(32'hbb3a1516),
	.w8(32'hb9cd42c0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22709a),
	.w1(32'h395dd6ef),
	.w2(32'hbb123c9a),
	.w3(32'h38bc34ca),
	.w4(32'h3a1fad20),
	.w5(32'h3a71880e),
	.w6(32'hba3e68a9),
	.w7(32'hbaad740c),
	.w8(32'hba1e7674),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f8b80),
	.w1(32'h3a8cb618),
	.w2(32'h3a53355d),
	.w3(32'hba25d3ea),
	.w4(32'hba0cb525),
	.w5(32'h3b0e7ed2),
	.w6(32'h3ab1da8f),
	.w7(32'h39850f98),
	.w8(32'h3a7f6715),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a3acf),
	.w1(32'h3a364808),
	.w2(32'h3abde535),
	.w3(32'h397ebf2d),
	.w4(32'hba9cd8b1),
	.w5(32'h3b2c3af8),
	.w6(32'hbac2cef8),
	.w7(32'hbb7e0595),
	.w8(32'hbb8e8477),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5b8fb),
	.w1(32'h3a016082),
	.w2(32'h3b9f3e25),
	.w3(32'h3ac63eab),
	.w4(32'h3bf97b62),
	.w5(32'h3a9cfcb8),
	.w6(32'h3a97e068),
	.w7(32'h3b10fb61),
	.w8(32'h3aec0022),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c2686),
	.w1(32'h3abc1364),
	.w2(32'h3b417de4),
	.w3(32'hba87a64d),
	.w4(32'h3b66ae04),
	.w5(32'h3b4f1f46),
	.w6(32'h3abddf0d),
	.w7(32'h3b88d9d3),
	.w8(32'h3a3c8e8d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12c5cf),
	.w1(32'h3a56d652),
	.w2(32'h3ba75e75),
	.w3(32'h39ca05df),
	.w4(32'hb9aa037e),
	.w5(32'h3c0c2e6d),
	.w6(32'h3baa27c8),
	.w7(32'hb907350a),
	.w8(32'hbbc48a89),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a900184),
	.w1(32'hba2935ca),
	.w2(32'hb927afbd),
	.w3(32'hba9d737c),
	.w4(32'hbb8dc151),
	.w5(32'hba7324bd),
	.w6(32'h3972f5d6),
	.w7(32'hbb34ace7),
	.w8(32'hb9b98111),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb069c),
	.w1(32'h39b7337e),
	.w2(32'hba76394a),
	.w3(32'h3b5cc3ed),
	.w4(32'h3b5ebf5a),
	.w5(32'h3b194511),
	.w6(32'hb9a2c42b),
	.w7(32'hbaa80840),
	.w8(32'h39b6eecd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d145),
	.w1(32'h3b55b4a2),
	.w2(32'hb9b47e57),
	.w3(32'h3a81bd81),
	.w4(32'h3b99e03b),
	.w5(32'hbab8242b),
	.w6(32'hbad5108a),
	.w7(32'h3b81016b),
	.w8(32'h3b49ef7c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b10f5),
	.w1(32'h398319d2),
	.w2(32'h3b97c42e),
	.w3(32'h3b0846fd),
	.w4(32'h3959e405),
	.w5(32'h3c01e236),
	.w6(32'h3ae94058),
	.w7(32'h3ad0e1df),
	.w8(32'hba870564),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8122fe),
	.w1(32'hbb73c02d),
	.w2(32'h3c070f60),
	.w3(32'hba26878f),
	.w4(32'hb9f27462),
	.w5(32'hbab34d7a),
	.w6(32'h39c679ad),
	.w7(32'h3c377ed8),
	.w8(32'h3c1ab982),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fe8cd),
	.w1(32'hbb0836af),
	.w2(32'hbb2cee37),
	.w3(32'hbb01bf80),
	.w4(32'hb92bb465),
	.w5(32'h3bc6bb4c),
	.w6(32'hba8fc25a),
	.w7(32'hbc19858c),
	.w8(32'hbb576d01),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e7a4d),
	.w1(32'hb74dac38),
	.w2(32'h3c128b1b),
	.w3(32'h3b3ff888),
	.w4(32'hbabe791e),
	.w5(32'h3c108c72),
	.w6(32'h3b096162),
	.w7(32'h3aabd3bf),
	.w8(32'h3b2aa313),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284ae0),
	.w1(32'h3aeb9784),
	.w2(32'hbbdab4cd),
	.w3(32'h3aeaa76e),
	.w4(32'h3a284a61),
	.w5(32'hbc12f7d0),
	.w6(32'hbb393364),
	.w7(32'hbb9dc592),
	.w8(32'hbc0553c5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b22246),
	.w1(32'h37cb76c5),
	.w2(32'hb560f693),
	.w3(32'h36173afb),
	.w4(32'hb6f88cfd),
	.w5(32'h388574cc),
	.w6(32'hb5924967),
	.w7(32'h37b915df),
	.w8(32'h3845f6cf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f8fb9),
	.w1(32'hb8309db0),
	.w2(32'hb9094e91),
	.w3(32'h37a680b7),
	.w4(32'hb89b94de),
	.w5(32'hb90b81c6),
	.w6(32'hb6b2b13a),
	.w7(32'hb8b108a0),
	.w8(32'hb8edb276),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380cfef2),
	.w1(32'h37fc3bfa),
	.w2(32'hb782f574),
	.w3(32'h36f8a04e),
	.w4(32'h3794d18a),
	.w5(32'hb86e37c1),
	.w6(32'h38a7c3ce),
	.w7(32'h38980f9c),
	.w8(32'hb8846a01),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42ca4c),
	.w1(32'h3a0199a3),
	.w2(32'h3b54e5a2),
	.w3(32'hba3a6dc1),
	.w4(32'h3a857fce),
	.w5(32'h3b3e77a3),
	.w6(32'h3ab6db97),
	.w7(32'h3b19d67f),
	.w8(32'h3ae08af0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d72359),
	.w1(32'hb80a4782),
	.w2(32'hb81f7188),
	.w3(32'hb763bfc5),
	.w4(32'hb7b7d005),
	.w5(32'hb7dd04ca),
	.w6(32'h36c0c8b6),
	.w7(32'h37738b26),
	.w8(32'hb7fc91f5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb529e45),
	.w1(32'h3a68a13e),
	.w2(32'h3c06b8f6),
	.w3(32'hb9f5bac4),
	.w4(32'h3b269f2f),
	.w5(32'h3b7845a9),
	.w6(32'hb873abdf),
	.w7(32'h3ba3c647),
	.w8(32'h3bcffa3a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa748b),
	.w1(32'hba1f0d68),
	.w2(32'h3b630af6),
	.w3(32'hbada3e9a),
	.w4(32'h3b808d8b),
	.w5(32'h3ba73b07),
	.w6(32'hbb2a247b),
	.w7(32'h3b13d9cd),
	.w8(32'h3bb059b0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20fd4d),
	.w1(32'hb9def321),
	.w2(32'hbb736fc5),
	.w3(32'hbb0cbd27),
	.w4(32'hbb262453),
	.w5(32'hbb8b631b),
	.w6(32'hbb562f8c),
	.w7(32'hbb21ac6c),
	.w8(32'hbb35bbbb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba889694),
	.w1(32'hbadf4fe1),
	.w2(32'hb9df0967),
	.w3(32'hbac1148b),
	.w4(32'hba5e59a4),
	.w5(32'hb9605646),
	.w6(32'hba425588),
	.w7(32'h3a1b033d),
	.w8(32'hba75b0fc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a507933),
	.w1(32'h3b1dac01),
	.w2(32'h3bbfb352),
	.w3(32'h3ab48cc9),
	.w4(32'h39a957a4),
	.w5(32'h3b8aa482),
	.w6(32'h3a196bda),
	.w7(32'h3bbeea06),
	.w8(32'h3bbf64e3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab166c7),
	.w1(32'h3ae25fab),
	.w2(32'hb94b313b),
	.w3(32'h3901a52a),
	.w4(32'hb9ced644),
	.w5(32'h39164cd4),
	.w6(32'hbaba7248),
	.w7(32'hba876dd0),
	.w8(32'h385494f6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf86ffe),
	.w1(32'h3b1a4052),
	.w2(32'h3bf8b9aa),
	.w3(32'hba9d82c0),
	.w4(32'h3b3d5166),
	.w5(32'h3bd5e7a5),
	.w6(32'h3a869790),
	.w7(32'h3baadcb2),
	.w8(32'h3bbe2f86),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37608214),
	.w1(32'hb7861620),
	.w2(32'hb7361a87),
	.w3(32'h368b313c),
	.w4(32'hb7909316),
	.w5(32'hb7749241),
	.w6(32'hb6526e0e),
	.w7(32'hb6fcbe8c),
	.w8(32'hb74dcec3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bfd264),
	.w1(32'hb8d5f6c3),
	.w2(32'hb8a52538),
	.w3(32'hb7f919a0),
	.w4(32'hb90b0708),
	.w5(32'hb8836f2e),
	.w6(32'hb7ba1838),
	.w7(32'hb9197521),
	.w8(32'hb8c7262e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c4e04),
	.w1(32'hb855aaff),
	.w2(32'hb983a42c),
	.w3(32'hb88e36ae),
	.w4(32'hb873f959),
	.w5(32'hb94a1557),
	.w6(32'hb9444188),
	.w7(32'hb95b9428),
	.w8(32'hb9aa75da),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a567b1f),
	.w1(32'h3aaacf77),
	.w2(32'h38fee6d8),
	.w3(32'h3ad4ff40),
	.w4(32'h3af59d58),
	.w5(32'h39a6016c),
	.w6(32'h3a3077e0),
	.w7(32'h3a9183ec),
	.w8(32'h39019ea8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f1e60),
	.w1(32'hbb35e616),
	.w2(32'hbb8f70c6),
	.w3(32'h3a399fd4),
	.w4(32'hbba41443),
	.w5(32'hbb84b2ac),
	.w6(32'hba95a9cf),
	.w7(32'hbb431303),
	.w8(32'hba7b72f8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b10193),
	.w1(32'hba326207),
	.w2(32'hb9e66be4),
	.w3(32'h38ea1dfd),
	.w4(32'hba0c8bea),
	.w5(32'hb993c0a0),
	.w6(32'h38378ee1),
	.w7(32'hba1369cf),
	.w8(32'hba2b875a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f0e582),
	.w1(32'hbb6b6c10),
	.w2(32'hbbb3be7b),
	.w3(32'hbb6c4ec7),
	.w4(32'hbb8f736f),
	.w5(32'hbb284226),
	.w6(32'hbb5d5230),
	.w7(32'hbb7bbbab),
	.w8(32'hbb5bb5eb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c48ea),
	.w1(32'h3b293763),
	.w2(32'h3c2d2ca8),
	.w3(32'hbab11ae4),
	.w4(32'h3c0680e1),
	.w5(32'h3bde05bd),
	.w6(32'h3b44a6d1),
	.w7(32'h3bfce70a),
	.w8(32'h3bfed022),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b699fca),
	.w1(32'h3ba22d9d),
	.w2(32'h3b9d1121),
	.w3(32'h3b89d8a7),
	.w4(32'h3b85edb0),
	.w5(32'h3b3d4d63),
	.w6(32'h3aadbc7c),
	.w7(32'h3b00deb1),
	.w8(32'h3b5ecd62),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd7f8c),
	.w1(32'hbb8e923e),
	.w2(32'h3c0cee4c),
	.w3(32'hbbbfd5b7),
	.w4(32'hbb4b0fe8),
	.w5(32'h3c050114),
	.w6(32'hbb08862a),
	.w7(32'h3bf106f5),
	.w8(32'h3c212d8c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bfabb),
	.w1(32'h3b922445),
	.w2(32'h3aa70558),
	.w3(32'h3bb5e62e),
	.w4(32'h3bcc953f),
	.w5(32'h3a93ccfc),
	.w6(32'h3bad5ec9),
	.w7(32'h3b606c42),
	.w8(32'hbb24fe75),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c725),
	.w1(32'hbb82b9fa),
	.w2(32'hbb8c1330),
	.w3(32'hbbafd4ca),
	.w4(32'hbb86e631),
	.w5(32'hbb3060a4),
	.w6(32'hbb5247a3),
	.w7(32'hbaba6d23),
	.w8(32'hbb3e9009),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46c10a),
	.w1(32'h3a7b311a),
	.w2(32'hba864a82),
	.w3(32'hbaf0db5f),
	.w4(32'hbb853015),
	.w5(32'hba79a3e2),
	.w6(32'hba10d60a),
	.w7(32'hba3b9deb),
	.w8(32'hbb3c2dc0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3729),
	.w1(32'h3b4b0df8),
	.w2(32'hbb92262b),
	.w3(32'h3b814250),
	.w4(32'h3a5cd350),
	.w5(32'hbb8fb020),
	.w6(32'h3aba523a),
	.w7(32'h3993d7da),
	.w8(32'hbb09220d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b17cd6),
	.w1(32'h38732802),
	.w2(32'hb6410515),
	.w3(32'h392c0abb),
	.w4(32'h38c3cf06),
	.w5(32'hb8f47973),
	.w6(32'h3936ba6c),
	.w7(32'h39076bb0),
	.w8(32'hb90f2d35),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fce7b),
	.w1(32'h3777deac),
	.w2(32'h3bb35964),
	.w3(32'hbb167069),
	.w4(32'h3aeb6e0d),
	.w5(32'h3bb0e9f2),
	.w6(32'hbab98036),
	.w7(32'h3b2bfdb8),
	.w8(32'h3b2d8fd1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a359b),
	.w1(32'hb8b991c5),
	.w2(32'h3c421c92),
	.w3(32'h3a0af629),
	.w4(32'h3917e7b7),
	.w5(32'h3bbe89d2),
	.w6(32'hbb29e0d4),
	.w7(32'h3be3c9a8),
	.w8(32'h3c397353),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944614),
	.w1(32'hbc89b375),
	.w2(32'hbac3aa06),
	.w3(32'hbb950ffb),
	.w4(32'hbca4f3d0),
	.w5(32'hbb9b5380),
	.w6(32'hbb24978b),
	.w7(32'hbc7781ed),
	.w8(32'hbbe68ff8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9f05),
	.w1(32'hbbc72d2c),
	.w2(32'hbc136b1c),
	.w3(32'h3b9611e5),
	.w4(32'hbbc221f9),
	.w5(32'hbbea5a7d),
	.w6(32'h3aa433e3),
	.w7(32'hbbc4590e),
	.w8(32'hbb8bcf84),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d8e85),
	.w1(32'hbaa7efe7),
	.w2(32'hbbeb70c3),
	.w3(32'hb98292bb),
	.w4(32'hbb1161fd),
	.w5(32'hbbf6dbe4),
	.w6(32'hbb6f1893),
	.w7(32'hbb85eb0e),
	.w8(32'hbbc5c45a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93df3d),
	.w1(32'hbb9e5867),
	.w2(32'h3bc96874),
	.w3(32'hbac9cae9),
	.w4(32'hbb20572a),
	.w5(32'h3bc69d86),
	.w6(32'hbaae5876),
	.w7(32'h3ab364a5),
	.w8(32'h3c0a3ab4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a9794),
	.w1(32'h382ef3e3),
	.w2(32'h36fb3bd3),
	.w3(32'h385e4658),
	.w4(32'h3845c8df),
	.w5(32'hb6591a1a),
	.w6(32'h3865c6a2),
	.w7(32'h383539b6),
	.w8(32'hb708d1ac),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba45908),
	.w1(32'hbc45b185),
	.w2(32'hba88be6e),
	.w3(32'h3a71b2ad),
	.w4(32'hbc56fbd9),
	.w5(32'hbb50ae7e),
	.w6(32'hbb8ff720),
	.w7(32'hbb98ae5e),
	.w8(32'h3bb81d63),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432163),
	.w1(32'h3b45a15c),
	.w2(32'h3c324e94),
	.w3(32'h3b8051ca),
	.w4(32'h3b8cb249),
	.w5(32'h3c2aca46),
	.w6(32'h39724854),
	.w7(32'h3ae93c76),
	.w8(32'h3c0c4014),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bd7719),
	.w1(32'hb496f9f7),
	.w2(32'hb921a1a9),
	.w3(32'hb74c6ed5),
	.w4(32'hb8989034),
	.w5(32'hb95615d5),
	.w6(32'hb84d1105),
	.w7(32'hb9143f46),
	.w8(32'hb98c109c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8ac51),
	.w1(32'hb9c6cb33),
	.w2(32'hb8770fc2),
	.w3(32'hb89eba4f),
	.w4(32'hbb74953d),
	.w5(32'hbb29844e),
	.w6(32'hbac03faf),
	.w7(32'hbad9dc7a),
	.w8(32'hba98cbff),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb784095),
	.w1(32'h3ad321d0),
	.w2(32'h3b7a32fc),
	.w3(32'hbb31711a),
	.w4(32'h3b2dbaca),
	.w5(32'h3ba376c8),
	.w6(32'hbae08f5c),
	.w7(32'h3b33f17b),
	.w8(32'h3b73d8b8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afad6ca),
	.w1(32'h3adbacbb),
	.w2(32'hbb65ea25),
	.w3(32'h3a59dcec),
	.w4(32'h3a85e313),
	.w5(32'hbb95fe21),
	.w6(32'hbb566b11),
	.w7(32'hbabdf4c3),
	.w8(32'hbb8a0d41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb12c6f),
	.w1(32'h3c4beaf9),
	.w2(32'h3bce680f),
	.w3(32'h3b8d97f4),
	.w4(32'h3c11f082),
	.w5(32'h3bb8adf2),
	.w6(32'h3af991a6),
	.w7(32'h3be9492e),
	.w8(32'h3b0fd699),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80dd2ce),
	.w1(32'hbb0cab16),
	.w2(32'hbba9c8e0),
	.w3(32'hba9af034),
	.w4(32'hbb6a8a97),
	.w5(32'hbb8ce3de),
	.w6(32'hba118968),
	.w7(32'hba8b62cd),
	.w8(32'hba7ade16),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5d68b),
	.w1(32'hbba180ca),
	.w2(32'hbaf30374),
	.w3(32'hbb9c6086),
	.w4(32'hbc0e74d9),
	.w5(32'h3b1c4134),
	.w6(32'hbb893354),
	.w7(32'hbc30cc39),
	.w8(32'hbbd3c4d0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e0637),
	.w1(32'hbae207ce),
	.w2(32'hbb83143e),
	.w3(32'hb9eda7eb),
	.w4(32'hbba8a83c),
	.w5(32'hbb2a439d),
	.w6(32'h395eefba),
	.w7(32'hbb029cb4),
	.w8(32'hbb6de3b3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7afeb9),
	.w1(32'hb899dcce),
	.w2(32'hbaacd5af),
	.w3(32'hba9d62ee),
	.w4(32'hb766f28e),
	.w5(32'hba85f548),
	.w6(32'hbb2c9488),
	.w7(32'hbab15ac5),
	.w8(32'hba9d29b2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad1266),
	.w1(32'h373c4ea7),
	.w2(32'h36af8823),
	.w3(32'h3710ccde),
	.w4(32'hb89edf5e),
	.w5(32'hb877c540),
	.w6(32'h380470d1),
	.w7(32'hb866c5e1),
	.w8(32'hb89550b0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978d42b),
	.w1(32'hba8017cb),
	.w2(32'hba6561ec),
	.w3(32'hba32b091),
	.w4(32'hbac328bd),
	.w5(32'hb9a52acf),
	.w6(32'hb9ba954a),
	.w7(32'hba4c8b64),
	.w8(32'h37d25511),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b0d7de),
	.w1(32'hb5b379cc),
	.w2(32'h37a3b3e9),
	.w3(32'h3881ec8b),
	.w4(32'h351c7f42),
	.w5(32'hb8a88d26),
	.w6(32'h37f97627),
	.w7(32'hb7be873c),
	.w8(32'h35b5ec89),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6cc76),
	.w1(32'hb82f64e2),
	.w2(32'hb6a0c4a5),
	.w3(32'hb8ce53ac),
	.w4(32'hb8cc3d5c),
	.w5(32'hb9054351),
	.w6(32'h37c1dc87),
	.w7(32'h3885f277),
	.w8(32'hb97203c9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c258b),
	.w1(32'hba7219d2),
	.w2(32'hbaef7eff),
	.w3(32'hbae1110f),
	.w4(32'hbad322d3),
	.w5(32'hba93ddc5),
	.w6(32'hbb44ab21),
	.w7(32'hbb0838fa),
	.w8(32'hbaeefa69),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cf851),
	.w1(32'h383c428e),
	.w2(32'h3963b01d),
	.w3(32'h389c13a5),
	.w4(32'hb884bbd2),
	.w5(32'h3944be17),
	.w6(32'h396e9d5c),
	.w7(32'h39e1e8f4),
	.w8(32'h3a187fa9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d1bc5),
	.w1(32'h3a8a52bf),
	.w2(32'h3ba76266),
	.w3(32'hba59868e),
	.w4(32'h39202893),
	.w5(32'h3b585479),
	.w6(32'hb8c320b1),
	.w7(32'h3a6a3d13),
	.w8(32'h3b59a5e5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a776866),
	.w1(32'hbb0ad0af),
	.w2(32'hbc0be1ff),
	.w3(32'hbaa1a425),
	.w4(32'hbb844ce7),
	.w5(32'hbbf2ca30),
	.w6(32'hbb1636d2),
	.w7(32'hbb5370f1),
	.w8(32'hbbbeac40),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c1ac40),
	.w1(32'hb93acded),
	.w2(32'hb8b50152),
	.w3(32'hb8770c0e),
	.w4(32'hb9799662),
	.w5(32'hb85c2b2b),
	.w6(32'hb904fa8d),
	.w7(32'hb9396507),
	.w8(32'hb8a3421d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c9878),
	.w1(32'hb9bbefc0),
	.w2(32'hb8072df3),
	.w3(32'hb9108bf6),
	.w4(32'hb98cb95f),
	.w5(32'h38032941),
	.w6(32'h3681efd0),
	.w7(32'hb9049d4b),
	.w8(32'h38e0717e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb778140d),
	.w1(32'hb79ebf3c),
	.w2(32'hb7bba0f6),
	.w3(32'hb6a85f0e),
	.w4(32'hb74a3f61),
	.w5(32'hb786933e),
	.w6(32'h36a96e99),
	.w7(32'hb6ee6907),
	.w8(32'hb79b6b63),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01852e),
	.w1(32'hb993b669),
	.w2(32'hba014810),
	.w3(32'hb9f75b7c),
	.w4(32'hb95a08f2),
	.w5(32'hb9dd4172),
	.w6(32'hb9a318ba),
	.w7(32'hb896562a),
	.w8(32'hb8d3d2a0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb879859c),
	.w1(32'h3be9d3a7),
	.w2(32'h3b400e0b),
	.w3(32'h396ec275),
	.w4(32'h3b4e1fa7),
	.w5(32'h3c5297a7),
	.w6(32'hbb828336),
	.w7(32'hbb1edb87),
	.w8(32'hba68478e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0edd5),
	.w1(32'h383db16a),
	.w2(32'h3b997900),
	.w3(32'h39692081),
	.w4(32'h3b914e8c),
	.w5(32'h3bd45f99),
	.w6(32'hb938dea0),
	.w7(32'h3bc0db15),
	.w8(32'h3ba117e0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d6033),
	.w1(32'hb9c19437),
	.w2(32'h3aa226a8),
	.w3(32'hba8dbcf7),
	.w4(32'h38f82bd0),
	.w5(32'h3ab382ba),
	.w6(32'hba444ee9),
	.w7(32'h3a561b37),
	.w8(32'h3aae64c0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15d02c),
	.w1(32'hbaacf19a),
	.w2(32'hba0889f0),
	.w3(32'h39ac676a),
	.w4(32'h399f2c7e),
	.w5(32'h3a850509),
	.w6(32'h3a610857),
	.w7(32'h3a86b77a),
	.w8(32'h39cbcfec),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c3a75),
	.w1(32'hb9b13aaa),
	.w2(32'hb8e6fecb),
	.w3(32'hb986bfca),
	.w4(32'hba83cc9a),
	.w5(32'hb801612f),
	.w6(32'hba793745),
	.w7(32'hba892a26),
	.w8(32'h3937744b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba630bb2),
	.w1(32'hbac3fbde),
	.w2(32'hba2a1f36),
	.w3(32'hbb0f2357),
	.w4(32'hba89213b),
	.w5(32'hba6389a5),
	.w6(32'hbb022ef1),
	.w7(32'hbab6f2e1),
	.w8(32'hba8367dd),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6a2da),
	.w1(32'h3a7a6fe1),
	.w2(32'hbbcb716f),
	.w3(32'h399ca0cc),
	.w4(32'hbb0fef33),
	.w5(32'hbb5a4a5e),
	.w6(32'hbb3331ba),
	.w7(32'hbb8bf4c4),
	.w8(32'hbb2fe80a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16de0),
	.w1(32'h3b5782ae),
	.w2(32'h3c77bad0),
	.w3(32'h39506ab6),
	.w4(32'h3b832ea1),
	.w5(32'h3c273694),
	.w6(32'h3b55ee26),
	.w7(32'h3c23a00c),
	.w8(32'h3c1d4141),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e2da5),
	.w1(32'hbad6d23b),
	.w2(32'hbba89c26),
	.w3(32'hb9c5c027),
	.w4(32'hbb1fee63),
	.w5(32'hbb75dd8e),
	.w6(32'hbacfb249),
	.w7(32'hbb4097a5),
	.w8(32'hbb3bcf4a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae03cdf),
	.w1(32'h39851a45),
	.w2(32'h3b628587),
	.w3(32'hbb280772),
	.w4(32'hbb2a9bc9),
	.w5(32'h3b15ecd1),
	.w6(32'hb9b8c425),
	.w7(32'h394331da),
	.w8(32'h3b26bd85),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88731f),
	.w1(32'h3a502b45),
	.w2(32'h3c28b6c9),
	.w3(32'hbb7720a6),
	.w4(32'h3af3d951),
	.w5(32'h3be070b6),
	.w6(32'hbb0e1e0d),
	.w7(32'h3b1a867b),
	.w8(32'h3bbc78d9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f9fd4),
	.w1(32'hbb8acf54),
	.w2(32'hbb86067a),
	.w3(32'hbb42f373),
	.w4(32'hbbd043a6),
	.w5(32'hbb144302),
	.w6(32'hbb89bb37),
	.w7(32'hbbefb829),
	.w8(32'hbb8c5a12),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38191d),
	.w1(32'hbab40a5f),
	.w2(32'h3a8b94fe),
	.w3(32'hbae3b258),
	.w4(32'hb94e4590),
	.w5(32'h3b1b61c0),
	.w6(32'hba1f27a8),
	.w7(32'h3b24ce78),
	.w8(32'h3b684fa0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3969da),
	.w1(32'hb9f197c2),
	.w2(32'hb9a1b153),
	.w3(32'hba3409d9),
	.w4(32'hb9bddd6b),
	.w5(32'hb85daa63),
	.w6(32'hba3f9aa1),
	.w7(32'hb957f106),
	.w8(32'h349f6ced),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba808d),
	.w1(32'h3bc8b225),
	.w2(32'hbb88ccff),
	.w3(32'h3b7ed1fe),
	.w4(32'h3bdbb539),
	.w5(32'hb98e2825),
	.w6(32'h3aaad4cd),
	.w7(32'h3b33b8fe),
	.w8(32'hbae0fca7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9e492),
	.w1(32'hb98b4b6d),
	.w2(32'h3b116f41),
	.w3(32'h389f8522),
	.w4(32'h391c1338),
	.w5(32'h3abc2443),
	.w6(32'h396cb628),
	.w7(32'h3823353d),
	.w8(32'h3a6136c1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b44d41),
	.w1(32'h38b7714c),
	.w2(32'h395b7f41),
	.w3(32'hb87d7305),
	.w4(32'h38dbb360),
	.w5(32'h38a633e5),
	.w6(32'h37692780),
	.w7(32'h37d67eae),
	.w8(32'h361f6e40),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38550900),
	.w1(32'h3803da25),
	.w2(32'h39002506),
	.w3(32'h36977a53),
	.w4(32'hb866bec7),
	.w5(32'h3894ce3d),
	.w6(32'h389f518f),
	.w7(32'hb8dc8510),
	.w8(32'h3862a612),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99602c3),
	.w1(32'hbb038f56),
	.w2(32'h3635968a),
	.w3(32'hb958512b),
	.w4(32'hb9f17c56),
	.w5(32'h39ccf9ec),
	.w6(32'hba7a2050),
	.w7(32'hba169517),
	.w8(32'h3a5190c9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc790a),
	.w1(32'hbb42ec04),
	.w2(32'hbac2bf3c),
	.w3(32'h3afa270e),
	.w4(32'hbb8e504d),
	.w5(32'hbb23c762),
	.w6(32'hb81fef30),
	.w7(32'hbb612626),
	.w8(32'h3a42aa60),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39e9a9),
	.w1(32'h3a4027cb),
	.w2(32'h3ab9d9dd),
	.w3(32'hbb115989),
	.w4(32'h3ad3d7e0),
	.w5(32'h3a903c09),
	.w6(32'hbb15e5f7),
	.w7(32'h3aff80bb),
	.w8(32'h3a9d8577),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3824f429),
	.w1(32'h3747655c),
	.w2(32'hb80d1cfd),
	.w3(32'h3716a958),
	.w4(32'hb7f63406),
	.w5(32'hb8491613),
	.w6(32'h37fba15a),
	.w7(32'hb7d0dc5a),
	.w8(32'hb85cc9a4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1f67),
	.w1(32'h39316d34),
	.w2(32'h3ac4205f),
	.w3(32'hbaad2387),
	.w4(32'h3a350c55),
	.w5(32'h3b440376),
	.w6(32'hb9f42602),
	.w7(32'h3b1ea7c5),
	.w8(32'h3b601865),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8bae1),
	.w1(32'hba3080ac),
	.w2(32'hbb0cd13a),
	.w3(32'hba9123e6),
	.w4(32'hba02bce6),
	.w5(32'hbae622fa),
	.w6(32'hbb139d3a),
	.w7(32'hbabf29d2),
	.w8(32'hbaadda44),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8a351),
	.w1(32'h3ac710cc),
	.w2(32'h3bf88b99),
	.w3(32'hbbdaf7a4),
	.w4(32'hbb0f8da9),
	.w5(32'h3b2e21cb),
	.w6(32'hbb635c32),
	.w7(32'h3b30033f),
	.w8(32'h3b9fc9ca),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35d988),
	.w1(32'h3c73bb59),
	.w2(32'h3bd12d84),
	.w3(32'h3ab245a3),
	.w4(32'h3c1dc3fa),
	.w5(32'h3c0ae567),
	.w6(32'h3b3cc684),
	.w7(32'h3be562e9),
	.w8(32'h3c0eec29),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af044c2),
	.w1(32'hbac2a7bf),
	.w2(32'hbb2ba73d),
	.w3(32'hb9d4b19f),
	.w4(32'hbae389a6),
	.w5(32'hbb46ab73),
	.w6(32'hba3a9a21),
	.w7(32'hbabef54a),
	.w8(32'hbb1943d9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d59f94),
	.w1(32'hb9d9fa48),
	.w2(32'hb9292e41),
	.w3(32'hb66f3aaf),
	.w4(32'hb9e82a2c),
	.w5(32'hb89207ae),
	.w6(32'hb8413101),
	.w7(32'hb9dd3f31),
	.w8(32'hb956e0c2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae767f7),
	.w1(32'hbb0769b6),
	.w2(32'hbb19b0d3),
	.w3(32'hbaafa1a9),
	.w4(32'hbadcf0a1),
	.w5(32'hbaa376c6),
	.w6(32'hbb1e0afa),
	.w7(32'hbb281393),
	.w8(32'hbac8430e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1289e3),
	.w1(32'hbaaac02e),
	.w2(32'hb8c11815),
	.w3(32'h39b4724c),
	.w4(32'hbb0161aa),
	.w5(32'hba86eba4),
	.w6(32'h3a087806),
	.w7(32'hbb1ec1af),
	.w8(32'hb99d83a6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d485d),
	.w1(32'hbae1cfb7),
	.w2(32'hbb62f3e6),
	.w3(32'h393bd27f),
	.w4(32'hbb10211a),
	.w5(32'hbb6fed72),
	.w6(32'h37e08c2d),
	.w7(32'hbb043bed),
	.w8(32'hbb21870a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17c53d),
	.w1(32'h3a7b5812),
	.w2(32'h3b325cdc),
	.w3(32'hb9ad452f),
	.w4(32'h3a87ac08),
	.w5(32'h3b047f55),
	.w6(32'h3a1fa656),
	.w7(32'h3b0cb92e),
	.w8(32'h3b24b077),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9b54c),
	.w1(32'hb98b2427),
	.w2(32'hba00119b),
	.w3(32'hb968a8e2),
	.w4(32'hb9d2a3b0),
	.w5(32'hba23df93),
	.w6(32'hb9871f00),
	.w7(32'hb99b217c),
	.w8(32'hb9f8a321),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ad97),
	.w1(32'h39a56ce5),
	.w2(32'h3b6e6af4),
	.w3(32'hbb108f78),
	.w4(32'h39a6aa0a),
	.w5(32'h3b899b14),
	.w6(32'hbb332c30),
	.w7(32'h3b11c8a1),
	.w8(32'h3b5b3789),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1099c),
	.w1(32'h3b1a8267),
	.w2(32'h3b534c8a),
	.w3(32'hb7f83ada),
	.w4(32'h3b2254c6),
	.w5(32'h3affd633),
	.w6(32'hbad24431),
	.w7(32'h3a85f3ae),
	.w8(32'h3ad86a5d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4de8c),
	.w1(32'h38a6c2a2),
	.w2(32'hba91da78),
	.w3(32'h3a30f595),
	.w4(32'hb8541f4d),
	.w5(32'h3984ff6d),
	.w6(32'h3a013c2c),
	.w7(32'hba07a59d),
	.w8(32'hbac8ff5c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe438e),
	.w1(32'hb9924ee9),
	.w2(32'h36b8ed9c),
	.w3(32'hb8b065ee),
	.w4(32'hb967ab27),
	.w5(32'h38bf609a),
	.w6(32'hb8c0bd72),
	.w7(32'hb9638c51),
	.w8(32'h3885895a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf613df),
	.w1(32'hb8475b3f),
	.w2(32'hba20bada),
	.w3(32'hba80cdba),
	.w4(32'h3abe71b4),
	.w5(32'h3ab9f6ab),
	.w6(32'h3921ebca),
	.w7(32'h3baaa5a4),
	.w8(32'h3b538700),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853fae8),
	.w1(32'h3833be97),
	.w2(32'hb6d60f9f),
	.w3(32'h38290ee4),
	.w4(32'h37e37aa7),
	.w5(32'hb7e8507e),
	.w6(32'h3815bba9),
	.w7(32'h374e6ccc),
	.w8(32'hb815255f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388af708),
	.w1(32'h391a7ac9),
	.w2(32'h39fe8af7),
	.w3(32'h38328b46),
	.w4(32'h392ca302),
	.w5(32'h39c847cb),
	.w6(32'h3855961d),
	.w7(32'h39be3b5a),
	.w8(32'h39bc4779),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d6b6f),
	.w1(32'h39bba109),
	.w2(32'hbb2dd5b9),
	.w3(32'hb922772c),
	.w4(32'hba91fdc7),
	.w5(32'hbb37af45),
	.w6(32'hbaa03231),
	.w7(32'hbb1e24b0),
	.w8(32'hbb38f5fe),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4a09),
	.w1(32'h3a88de99),
	.w2(32'h3bac940c),
	.w3(32'hbb65b07f),
	.w4(32'h3b89acc1),
	.w5(32'h3c190fde),
	.w6(32'hbb5e74b5),
	.w7(32'h3b048710),
	.w8(32'h3b989898),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edbc25),
	.w1(32'hbab3c867),
	.w2(32'hba2408b2),
	.w3(32'hb9856aae),
	.w4(32'hba91b06e),
	.w5(32'hb9d93272),
	.w6(32'hb981e822),
	.w7(32'hba344ee2),
	.w8(32'h3937d312),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993b3d2),
	.w1(32'hb80c457f),
	.w2(32'hbb8785c9),
	.w3(32'h39494db4),
	.w4(32'h38deb87e),
	.w5(32'hbb47069e),
	.w6(32'hbae09d9c),
	.w7(32'hbab1f2d4),
	.w8(32'hbb0a9a64),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ace7ea),
	.w1(32'h3add4af7),
	.w2(32'h3b7cbc7b),
	.w3(32'hb885c592),
	.w4(32'h3a782bd6),
	.w5(32'h3b61da45),
	.w6(32'h3aff152c),
	.w7(32'h3aa13286),
	.w8(32'h3b7f1ff9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3edb7c),
	.w1(32'h3bc38ff1),
	.w2(32'h3bf931d6),
	.w3(32'h3b4e8221),
	.w4(32'h3ba003a6),
	.w5(32'h3bfd25ea),
	.w6(32'h3ba5ea4c),
	.w7(32'h3b8231ec),
	.w8(32'h3a395575),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a31c0),
	.w1(32'h3abd0477),
	.w2(32'h3ae6666d),
	.w3(32'hb9947c7f),
	.w4(32'hb94f5edc),
	.w5(32'h3903e27c),
	.w6(32'hbb46fb57),
	.w7(32'hb997b81f),
	.w8(32'h3a258b3e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb229e64),
	.w1(32'h3b03692c),
	.w2(32'h3bb69937),
	.w3(32'hba63ca50),
	.w4(32'h3b7c16b2),
	.w5(32'h3bb97d2f),
	.w6(32'h3a981b3e),
	.w7(32'h3bc25370),
	.w8(32'h3b9d54ce),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392fff21),
	.w1(32'h3775c836),
	.w2(32'hb7aec484),
	.w3(32'hb67ae85c),
	.w4(32'hb77d5956),
	.w5(32'hb897fd5b),
	.w6(32'hb89d9a37),
	.w7(32'hb8e03f46),
	.w8(32'hb9368c93),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9a3c3),
	.w1(32'h39eee992),
	.w2(32'hba299af4),
	.w3(32'hbb1dc8c6),
	.w4(32'hbb3aa6af),
	.w5(32'hbaaa9e38),
	.w6(32'hbae12311),
	.w7(32'hbaf95d67),
	.w8(32'hba5034ec),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3701b18f),
	.w1(32'h37461876),
	.w2(32'hb812c7c3),
	.w3(32'h37b1d72f),
	.w4(32'h38206742),
	.w5(32'hb805c309),
	.w6(32'h36f62a0c),
	.w7(32'h38016d5e),
	.w8(32'hb7e0fd5e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982d1d2),
	.w1(32'h389a517d),
	.w2(32'h3a1bd290),
	.w3(32'h39750414),
	.w4(32'h3a165d1d),
	.w5(32'h39222c30),
	.w6(32'h39a8e705),
	.w7(32'h3a493a20),
	.w8(32'hb90a08f3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9954595),
	.w1(32'h371f523d),
	.w2(32'hba35f218),
	.w3(32'hb91b9dbc),
	.w4(32'hb902fab9),
	.w5(32'hba820cd4),
	.w6(32'h39384014),
	.w7(32'h39b394a6),
	.w8(32'hba48df2c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4855c6),
	.w1(32'hba2210f0),
	.w2(32'hbacc4fbf),
	.w3(32'hbac27a8c),
	.w4(32'hbb681845),
	.w5(32'hba0287c2),
	.w6(32'h3a0867db),
	.w7(32'hbac1cfe4),
	.w8(32'hbb3c745e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716a3cd),
	.w1(32'hb7da401c),
	.w2(32'hb81ab026),
	.w3(32'hb6b84d13),
	.w4(32'hb80fffc1),
	.w5(32'hb8284c0f),
	.w6(32'h36ac997d),
	.w7(32'hb7e3a828),
	.w8(32'hb7d024fc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e9897c),
	.w1(32'hb7c1ce61),
	.w2(32'hb8022cd7),
	.w3(32'hb79616f1),
	.w4(32'h3742ab41),
	.w5(32'h381416c1),
	.w6(32'h370e0f17),
	.w7(32'h37647a55),
	.w8(32'h37a1df36),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0da00),
	.w1(32'h3980aafc),
	.w2(32'hba9b36e6),
	.w3(32'hba1aaadf),
	.w4(32'h39a7be7d),
	.w5(32'hba8d7357),
	.w6(32'hba048d50),
	.w7(32'h3a57e2e9),
	.w8(32'hba4384eb),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b6c9b),
	.w1(32'hbadfa1d3),
	.w2(32'h3b8b841d),
	.w3(32'h3b0b343e),
	.w4(32'hbb4c800e),
	.w5(32'h3b95ed86),
	.w6(32'hba49437c),
	.w7(32'h3b5d9549),
	.w8(32'h3bac247b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800e18),
	.w1(32'hbbb7bf64),
	.w2(32'h3ae404ab),
	.w3(32'h3b00e595),
	.w4(32'hbbc1b5c9),
	.w5(32'h3b099227),
	.w6(32'h3af473fa),
	.w7(32'hba80cb4d),
	.w8(32'h3bbc5d78),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a158f4d),
	.w1(32'h3a8ad2b6),
	.w2(32'h3a58fbb8),
	.w3(32'h3a622bdd),
	.w4(32'h3a84de96),
	.w5(32'h3a177fe2),
	.w6(32'h3aae895f),
	.w7(32'h3ab2cca2),
	.w8(32'h3a83f366),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185296),
	.w1(32'h3bd9d56d),
	.w2(32'h3c56ea67),
	.w3(32'hb8c1f15d),
	.w4(32'h3c13a63c),
	.w5(32'h3c4a18c1),
	.w6(32'h3b8d3f7e),
	.w7(32'h3c497062),
	.w8(32'h3b9e62d1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b097cc0),
	.w1(32'h3b1ead10),
	.w2(32'hb9a08a3a),
	.w3(32'hbb4ca57e),
	.w4(32'hbb459150),
	.w5(32'h3b1ddea0),
	.w6(32'hbb8f8d4d),
	.w7(32'hbb6898a8),
	.w8(32'h39f5a958),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2c3d5),
	.w1(32'h3a72c067),
	.w2(32'h3ba6626e),
	.w3(32'hb9ad01ac),
	.w4(32'h3b04f37b),
	.w5(32'h3b74d3ca),
	.w6(32'hba7bc40c),
	.w7(32'h3b3941f9),
	.w8(32'h3b87abf7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3848c228),
	.w1(32'h375201a7),
	.w2(32'h36442e70),
	.w3(32'h3884a8b4),
	.w4(32'h379962b1),
	.w5(32'h371473e3),
	.w6(32'h3880abbe),
	.w7(32'h383d4c6c),
	.w8(32'h37a8b9b0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c5fd8),
	.w1(32'hb86aee56),
	.w2(32'hb8a99650),
	.w3(32'h3833e8ff),
	.w4(32'hb897a761),
	.w5(32'hb889547c),
	.w6(32'h3805c34b),
	.w7(32'hb88d6be2),
	.w8(32'hb8408061),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35930c99),
	.w1(32'h35b1bf63),
	.w2(32'hb717064e),
	.w3(32'h371d0539),
	.w4(32'h36fa2358),
	.w5(32'hb716b7f4),
	.w6(32'h3780f61f),
	.w7(32'h374a02cf),
	.w8(32'hb71685d1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cd259),
	.w1(32'h388a40ef),
	.w2(32'h3b955da4),
	.w3(32'h38e0ed86),
	.w4(32'h3a275695),
	.w5(32'h3ba55d03),
	.w6(32'hba5dd8e3),
	.w7(32'h3a8baef0),
	.w8(32'h3b945947),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a9e0f),
	.w1(32'hba29c611),
	.w2(32'h3b2cf004),
	.w3(32'hbb204b99),
	.w4(32'hb9b81221),
	.w5(32'h3b13da1b),
	.w6(32'hbab5b82b),
	.w7(32'hb81a37d2),
	.w8(32'h3b16b65e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fcfa6),
	.w1(32'hbb565efd),
	.w2(32'hbc06284e),
	.w3(32'hbabb4610),
	.w4(32'hbba7a35e),
	.w5(32'hbbf46b57),
	.w6(32'hbb38f1b6),
	.w7(32'hbb822b79),
	.w8(32'hbbaba28f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c372ab),
	.w1(32'hb9fd3dec),
	.w2(32'hba81eeb1),
	.w3(32'h3872d669),
	.w4(32'hb9693758),
	.w5(32'hba41065f),
	.w6(32'hb956ae70),
	.w7(32'hb8dcf5c3),
	.w8(32'hba0ed05c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79831c),
	.w1(32'h3ba651c2),
	.w2(32'h3c2de583),
	.w3(32'hbb0d9ca4),
	.w4(32'h3bb51d7c),
	.w5(32'h3ca6146d),
	.w6(32'hba7061b6),
	.w7(32'h3c7c9c88),
	.w8(32'h3c286c78),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ccb40),
	.w1(32'h3b5ad443),
	.w2(32'h3c146def),
	.w3(32'h3bd23f03),
	.w4(32'h3c1a3348),
	.w5(32'h3ba13df7),
	.w6(32'h3bf060d8),
	.w7(32'h3af9d883),
	.w8(32'hba413f5e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a354cb1),
	.w1(32'h3bef8be0),
	.w2(32'h3c1084f1),
	.w3(32'hbb8ddbda),
	.w4(32'h3c0ac356),
	.w5(32'h3a85c859),
	.w6(32'hbbeff3a1),
	.w7(32'h3ba039f0),
	.w8(32'h3a9da832),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff07c),
	.w1(32'hbac02c9d),
	.w2(32'h3aa35fb1),
	.w3(32'h3b7421d6),
	.w4(32'h3c13f8df),
	.w5(32'h3b41758a),
	.w6(32'hbb65f17f),
	.w7(32'h3b8f4b89),
	.w8(32'h3afd4087),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5168b9),
	.w1(32'hba285626),
	.w2(32'h3a652fe0),
	.w3(32'h3b025135),
	.w4(32'hbbe4a54f),
	.w5(32'hbc4037a7),
	.w6(32'h3beb4f5d),
	.w7(32'hbb80b225),
	.w8(32'hbc2b92d6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97cd9d),
	.w1(32'hbbb9e7e1),
	.w2(32'h3a8bcd52),
	.w3(32'hbbcdc6ee),
	.w4(32'hbad2edf5),
	.w5(32'h3bfc246c),
	.w6(32'hbc1c99a2),
	.w7(32'h3b38a033),
	.w8(32'h3bdfb46a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0349),
	.w1(32'hbc7c8b3f),
	.w2(32'hbcba8a61),
	.w3(32'h3afc9641),
	.w4(32'hbb2658f4),
	.w5(32'hbc5b5a2c),
	.w6(32'hbb991576),
	.w7(32'h3be278cd),
	.w8(32'h3c072125),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc794dea),
	.w1(32'h3c88ddcf),
	.w2(32'h3bec9980),
	.w3(32'hbbfccaf3),
	.w4(32'h3c2d4c7a),
	.w5(32'h3b862d8d),
	.w6(32'hbb2c902b),
	.w7(32'h3c0acdd1),
	.w8(32'h3bf06be4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d925b),
	.w1(32'hbbd4d6f8),
	.w2(32'h3c87fb9e),
	.w3(32'h3b475743),
	.w4(32'hbbb71714),
	.w5(32'h3c5675b3),
	.w6(32'h3bf17b9a),
	.w7(32'hbc0f5b79),
	.w8(32'hbba24c0d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73d527),
	.w1(32'hbbfc7042),
	.w2(32'hba34020e),
	.w3(32'h3c9d665a),
	.w4(32'hbc8d0e2a),
	.w5(32'h3c478b25),
	.w6(32'h3b5f033f),
	.w7(32'hbc821e1d),
	.w8(32'h3afe625d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d04b4),
	.w1(32'hbabef911),
	.w2(32'hbbb224dd),
	.w3(32'h3c326cfb),
	.w4(32'h3ba17d57),
	.w5(32'h39b18f4d),
	.w6(32'h3bbc81c8),
	.w7(32'hbb069b75),
	.w8(32'h3b02ae57),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1fafe),
	.w1(32'hb9e21e12),
	.w2(32'h3b19b6ec),
	.w3(32'h3bcce702),
	.w4(32'hbc6cc02c),
	.w5(32'h3b836581),
	.w6(32'hbae12da3),
	.w7(32'hbbe95493),
	.w8(32'hbb67c25f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6337f5),
	.w1(32'h3b7d4c30),
	.w2(32'hbb86f16e),
	.w3(32'h39732bf2),
	.w4(32'h3bed7d84),
	.w5(32'hbc024973),
	.w6(32'h3aef753c),
	.w7(32'h3bdfee01),
	.w8(32'hbacdfc2b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad49279),
	.w1(32'hbb13c835),
	.w2(32'hbbccc6b1),
	.w3(32'hbb886fd5),
	.w4(32'hbb9c21be),
	.w5(32'hbc50711b),
	.w6(32'hbb54fe2c),
	.w7(32'hbbabcaee),
	.w8(32'hbc775dd9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe62f6),
	.w1(32'h3c09e8c5),
	.w2(32'h3c5cd4db),
	.w3(32'hbc8081c0),
	.w4(32'h3bb68f26),
	.w5(32'h3bdd6c5a),
	.w6(32'hbc9553fa),
	.w7(32'h3b9dad9a),
	.w8(32'h3c0d94dd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9465bb),
	.w1(32'hba3cc028),
	.w2(32'h3c313de9),
	.w3(32'h3c1d8b71),
	.w4(32'h3c61715b),
	.w5(32'h3c24fdf0),
	.w6(32'h3c3241a3),
	.w7(32'h39ee29a2),
	.w8(32'h3c33e0f2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0770f),
	.w1(32'h3b2da885),
	.w2(32'hbbb47aeb),
	.w3(32'h3be0c41e),
	.w4(32'hbbf2547c),
	.w5(32'hbc81d6c3),
	.w6(32'h3b28c76b),
	.w7(32'hbc74cc3e),
	.w8(32'hbc4ae8e9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda8470),
	.w1(32'hbc312f05),
	.w2(32'h3bc529b2),
	.w3(32'hbc1ee631),
	.w4(32'hbc84c06d),
	.w5(32'h3aaa77d3),
	.w6(32'hbc225477),
	.w7(32'hbc480333),
	.w8(32'hbc23a421),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae68ba7),
	.w1(32'h3c16ac74),
	.w2(32'h3bb689f4),
	.w3(32'h3af9742a),
	.w4(32'h3bb28f8a),
	.w5(32'h3b56ed5d),
	.w6(32'hbbbbe309),
	.w7(32'hbc4650bf),
	.w8(32'hbc59564b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d9552),
	.w1(32'h3c2411b8),
	.w2(32'h3bd9011e),
	.w3(32'hbb919ba1),
	.w4(32'h3b45b9f9),
	.w5(32'hbba85738),
	.w6(32'hbc3589eb),
	.w7(32'hbac64789),
	.w8(32'hbb4cc88f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4e097),
	.w1(32'hbb14b5e2),
	.w2(32'h3c883ff7),
	.w3(32'h38e95d9b),
	.w4(32'hbb11db0b),
	.w5(32'h3cb38400),
	.w6(32'h3aea4f59),
	.w7(32'h3b053d90),
	.w8(32'h3c8a29ab),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6edee6),
	.w1(32'h3a3f239c),
	.w2(32'h3b6aaa0f),
	.w3(32'hba9796f0),
	.w4(32'h3c4f6f6f),
	.w5(32'hbac4c533),
	.w6(32'hbb8274db),
	.w7(32'h3c2447e1),
	.w8(32'hba9e68f5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd43f6),
	.w1(32'h3c2b6248),
	.w2(32'h3bceb007),
	.w3(32'hbc8e99b6),
	.w4(32'hbb418534),
	.w5(32'h3c070a7e),
	.w6(32'hbc5b149a),
	.w7(32'hbb2b0855),
	.w8(32'h3b383e5b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a2bd),
	.w1(32'hbc02ebe0),
	.w2(32'hbbbe8baa),
	.w3(32'h3c365af7),
	.w4(32'hbb2b816b),
	.w5(32'h3a980824),
	.w6(32'h3b2cbf62),
	.w7(32'hb82c8349),
	.w8(32'h3c0f2591),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52891b),
	.w1(32'h3a79eead),
	.w2(32'hbc2c0f04),
	.w3(32'h3b642b55),
	.w4(32'hbb336de9),
	.w5(32'h3b17ca7d),
	.w6(32'h3bda592c),
	.w7(32'h3b98b05b),
	.w8(32'h3c1693d3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1192cc),
	.w1(32'h3cd15071),
	.w2(32'h3cc57585),
	.w3(32'hb8793963),
	.w4(32'h3b79b2d4),
	.w5(32'hbc17290d),
	.w6(32'h3c128073),
	.w7(32'hbbcfe4d2),
	.w8(32'hbbbbdbdb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90c422),
	.w1(32'h3bf3f699),
	.w2(32'h3bbc57cd),
	.w3(32'hbb3cfd9a),
	.w4(32'h3c87e01c),
	.w5(32'h3bae0333),
	.w6(32'hba7255fb),
	.w7(32'h3b555910),
	.w8(32'hbb50d273),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c104),
	.w1(32'h3b736c8d),
	.w2(32'h3b430165),
	.w3(32'h39f91ac9),
	.w4(32'h3c1deaaa),
	.w5(32'hbb89a341),
	.w6(32'hbb8b9178),
	.w7(32'h3b842b7a),
	.w8(32'hbab2f431),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cdb16),
	.w1(32'h3bfe18fe),
	.w2(32'hb9f4fa1f),
	.w3(32'hb9cd28e8),
	.w4(32'h3b68a6bc),
	.w5(32'hbb9ed871),
	.w6(32'hbc0f783c),
	.w7(32'h3b3434a7),
	.w8(32'h3bae45af),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaba4d),
	.w1(32'hbb83f806),
	.w2(32'hbb12d4b8),
	.w3(32'h3be537da),
	.w4(32'hbbb57ab1),
	.w5(32'hbb4815ed),
	.w6(32'h3be7c2c0),
	.w7(32'h3c4b7771),
	.w8(32'h3c3f5ed5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7261),
	.w1(32'hbc7ae739),
	.w2(32'hbc3c2ea3),
	.w3(32'hbba3c3b2),
	.w4(32'hbba86f33),
	.w5(32'h3a9ba7e9),
	.w6(32'hb9409606),
	.w7(32'h3c60da49),
	.w8(32'h3b909091),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82f846),
	.w1(32'h3b73b2b0),
	.w2(32'h3c30bb01),
	.w3(32'h3b6eb06a),
	.w4(32'h3c04f54a),
	.w5(32'h3bd50e58),
	.w6(32'h3afb81e9),
	.w7(32'h3b529d8d),
	.w8(32'h3be26086),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846848),
	.w1(32'hbbd8acb5),
	.w2(32'hbc074317),
	.w3(32'h3b308077),
	.w4(32'h3b19d8b3),
	.w5(32'hbc328e24),
	.w6(32'h3b000836),
	.w7(32'hb98b6dd9),
	.w8(32'hbc0a6e3b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc670697),
	.w1(32'h3c81230e),
	.w2(32'h3d0f4b14),
	.w3(32'hbc5f15c3),
	.w4(32'h3cc913c0),
	.w5(32'h3d104f85),
	.w6(32'hbc926617),
	.w7(32'h3c501bea),
	.w8(32'h3c316634),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49798a),
	.w1(32'h3b5c697c),
	.w2(32'h3cded89b),
	.w3(32'hbbb3e784),
	.w4(32'hb9bca41c),
	.w5(32'h3d1736e2),
	.w6(32'hbc2ebd78),
	.w7(32'hbc047b99),
	.w8(32'h3c38ceaa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b715cfc),
	.w1(32'hbbdf6d4f),
	.w2(32'hbc356c3a),
	.w3(32'h3c29944d),
	.w4(32'hbb476eb7),
	.w5(32'h3b5b24c0),
	.w6(32'hba022b75),
	.w7(32'hbb532ec9),
	.w8(32'h3c0832a6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dea80),
	.w1(32'hbc1ec8e8),
	.w2(32'h3b13dbf0),
	.w3(32'hbb459248),
	.w4(32'hbbb1bde1),
	.w5(32'h3c0f6e80),
	.w6(32'h3b88de3a),
	.w7(32'h3b6eaaff),
	.w8(32'h3c701611),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bade98d),
	.w1(32'h3c8ce17e),
	.w2(32'hbb7c00a6),
	.w3(32'h3bcc38ef),
	.w4(32'h3c32fcd7),
	.w5(32'hbc35aa46),
	.w6(32'h3be68463),
	.w7(32'h3b9202ec),
	.w8(32'hbc22c2f9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4048),
	.w1(32'hbbe3e507),
	.w2(32'h3b9b4912),
	.w3(32'hbc591b6b),
	.w4(32'hbc868e0c),
	.w5(32'h3ba2ffbf),
	.w6(32'hbc69187c),
	.w7(32'hbc662466),
	.w8(32'h3a98153c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11fe87),
	.w1(32'hbbe61c4f),
	.w2(32'hbbdd7ee6),
	.w3(32'h3bdad88c),
	.w4(32'hbb233754),
	.w5(32'hbc20fce5),
	.w6(32'h3b872d71),
	.w7(32'hbb8c7792),
	.w8(32'hbbf10ad2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4c58f),
	.w1(32'hbb9f13cb),
	.w2(32'hbc7d4f87),
	.w3(32'hbb9ef482),
	.w4(32'h3c8f133e),
	.w5(32'h3c41d2b5),
	.w6(32'hbc193f6a),
	.w7(32'h3c094940),
	.w8(32'h3cb3350b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc7cfb),
	.w1(32'h3c23c1b2),
	.w2(32'h3b2044fd),
	.w3(32'h3955e2a6),
	.w4(32'hbb062990),
	.w5(32'hbb179a43),
	.w6(32'h3bef4d63),
	.w7(32'hbbb230fb),
	.w8(32'hbb344d2c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6320d),
	.w1(32'hbb4beff7),
	.w2(32'h3c081d4f),
	.w3(32'h3a3e67e2),
	.w4(32'hbb5872f1),
	.w5(32'h3bbf6ee7),
	.w6(32'hbacf259f),
	.w7(32'h3ba4181f),
	.w8(32'h3baa042c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f5c26),
	.w1(32'h3b071683),
	.w2(32'hbb37a426),
	.w3(32'hb8c5e6eb),
	.w4(32'h3b98966a),
	.w5(32'hbc62e251),
	.w6(32'hbb62974b),
	.w7(32'h3b8ec021),
	.w8(32'hbc16bcb6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc410376),
	.w1(32'h3b84e02b),
	.w2(32'h3afffac5),
	.w3(32'hbc52f74a),
	.w4(32'hbab2e65a),
	.w5(32'hba2b74f5),
	.w6(32'hbac96dd7),
	.w7(32'h3bb776cc),
	.w8(32'hbaa53948),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3acc3),
	.w1(32'hbbfa8166),
	.w2(32'hbb919d15),
	.w3(32'hbbfee4cb),
	.w4(32'hbc49eba7),
	.w5(32'hbb8ab2eb),
	.w6(32'hbc8d4e6b),
	.w7(32'hbc27013e),
	.w8(32'hbb18c80f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2639c),
	.w1(32'hbbad7fb9),
	.w2(32'h3c298fe8),
	.w3(32'h3bdaf9a7),
	.w4(32'hb9e388e0),
	.w5(32'h3c8e591c),
	.w6(32'h3ba58863),
	.w7(32'h3b0b908e),
	.w8(32'h3c637140),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bc90a),
	.w1(32'h3c95ca56),
	.w2(32'hb91e5766),
	.w3(32'h3be01ac6),
	.w4(32'h3d141401),
	.w5(32'hba976f73),
	.w6(32'h3bd9e3d6),
	.w7(32'h3cd1e8d1),
	.w8(32'h3c8757e0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ffd8),
	.w1(32'hbc8b8a23),
	.w2(32'hbcc97b1a),
	.w3(32'hbc53bf06),
	.w4(32'h3a9683f9),
	.w5(32'hb9fa1a67),
	.w6(32'hbc07119d),
	.w7(32'h3c34671d),
	.w8(32'h3c98d20b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82ae29),
	.w1(32'hbbc4c50a),
	.w2(32'h3bca00d7),
	.w3(32'hbbbe0be3),
	.w4(32'hbb916670),
	.w5(32'hbaf117ca),
	.w6(32'h3baf28a4),
	.w7(32'hbc62f3c3),
	.w8(32'hbc88649c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc93f55),
	.w1(32'h3bd69f0e),
	.w2(32'h3bee7863),
	.w3(32'hbb367e8f),
	.w4(32'h3cb333b2),
	.w5(32'h3c92f097),
	.w6(32'hbc41a285),
	.w7(32'h3a71df62),
	.w8(32'h3baba197),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8a9a5),
	.w1(32'h3b672054),
	.w2(32'h3b82c1d2),
	.w3(32'hba2bdef1),
	.w4(32'hbb8b9e0f),
	.w5(32'h3b2b2275),
	.w6(32'hbbf556a7),
	.w7(32'hbb619712),
	.w8(32'h3ba74e2d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fd5eb),
	.w1(32'hbc7f4f31),
	.w2(32'hbc10753c),
	.w3(32'h3bb36b79),
	.w4(32'hbc0f66a7),
	.w5(32'h3bdd5128),
	.w6(32'h3ba0360e),
	.w7(32'h38859e4c),
	.w8(32'h3c2961cb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b35d),
	.w1(32'h3cb7352c),
	.w2(32'h3bcb5aac),
	.w3(32'h3b75aa30),
	.w4(32'h3c4dad50),
	.w5(32'hbc167c00),
	.w6(32'hb9f8cffb),
	.w7(32'h3ab3d88c),
	.w8(32'hbc780630),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c995),
	.w1(32'hbb989217),
	.w2(32'h3a2272af),
	.w3(32'hbc79d97c),
	.w4(32'hbc751a63),
	.w5(32'hbc2b6b6b),
	.w6(32'hbc404147),
	.w7(32'hbbc9bb85),
	.w8(32'hbbb59b08),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17e831),
	.w1(32'hbbfc1063),
	.w2(32'hbc20f0fe),
	.w3(32'hbb5e3ccc),
	.w4(32'h3c3c7dd8),
	.w5(32'hbc5475f0),
	.w6(32'hbbe77cd3),
	.w7(32'h3bde1346),
	.w8(32'hb9f6e8f9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae6693),
	.w1(32'hbbbd109a),
	.w2(32'hbc07a383),
	.w3(32'hbca470af),
	.w4(32'hbbc3c6ad),
	.w5(32'h3c82cd8f),
	.w6(32'hbc3b2b68),
	.w7(32'h3b0237e9),
	.w8(32'h3cb5964e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48c3c),
	.w1(32'h3b26cb76),
	.w2(32'h3bed5aeb),
	.w3(32'h3bc4673e),
	.w4(32'h3b93f86d),
	.w5(32'hba44e95a),
	.w6(32'h3c3f51f9),
	.w7(32'hbadcca08),
	.w8(32'hb9444342),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cc898),
	.w1(32'h3ca058e7),
	.w2(32'h3c040b1d),
	.w3(32'hbb8096f5),
	.w4(32'h3c19e2b3),
	.w5(32'hbbd56ab8),
	.w6(32'hbc46dec4),
	.w7(32'hba85b0da),
	.w8(32'hbbe2f4c3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule