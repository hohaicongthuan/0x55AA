module layer_10_featuremap_469(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d628b),
	.w1(32'h3a2ad646),
	.w2(32'hba9bc1a7),
	.w3(32'h3a44920a),
	.w4(32'hba9cdd39),
	.w5(32'hbb8825d7),
	.w6(32'h3ad62f32),
	.w7(32'hba870ed8),
	.w8(32'hbae0a3d5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9019109),
	.w1(32'h3b61ad91),
	.w2(32'hb97a33f6),
	.w3(32'hba941e0c),
	.w4(32'h3bd3b0ca),
	.w5(32'hb9f891e5),
	.w6(32'h3a162761),
	.w7(32'h3baa21fb),
	.w8(32'hbaeee4cc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6ed22),
	.w1(32'h3bccd2a4),
	.w2(32'hbb1a9c1b),
	.w3(32'hb91b2759),
	.w4(32'h3b27154e),
	.w5(32'hbb303343),
	.w6(32'hba50e0e1),
	.w7(32'h3b8d5349),
	.w8(32'h3a53f7bf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6a136),
	.w1(32'hbaaff7ad),
	.w2(32'hba6d194b),
	.w3(32'hbaa0a044),
	.w4(32'h39c797b8),
	.w5(32'hbb765f1a),
	.w6(32'h3b00fc85),
	.w7(32'h3b0025cd),
	.w8(32'hbb2aecbb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef61f2),
	.w1(32'hba29fbc3),
	.w2(32'hba49e663),
	.w3(32'h39ad3343),
	.w4(32'hba5cb18c),
	.w5(32'hbaffc4a4),
	.w6(32'h390b524f),
	.w7(32'hb98811ed),
	.w8(32'hbac853a9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4718f),
	.w1(32'hbaaaf8b3),
	.w2(32'h3a17e00c),
	.w3(32'hba4986d7),
	.w4(32'h3b4ae3e8),
	.w5(32'h3b6324bb),
	.w6(32'hb92882c6),
	.w7(32'h3ad427f8),
	.w8(32'h3b2dda09),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76f8be),
	.w1(32'hba4cb0f5),
	.w2(32'h3ae95a2f),
	.w3(32'hba8e322c),
	.w4(32'hba182e0e),
	.w5(32'hbb42b351),
	.w6(32'h3a253424),
	.w7(32'hbb185056),
	.w8(32'hbb13b0fb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d145ac),
	.w1(32'h3ad3d53e),
	.w2(32'hbb8b664e),
	.w3(32'hba7b675b),
	.w4(32'h3b4a1da1),
	.w5(32'hbadad033),
	.w6(32'h3b11ebfa),
	.w7(32'h3b265efd),
	.w8(32'h3a7b97ba),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfb19e),
	.w1(32'hba398580),
	.w2(32'h3ac05564),
	.w3(32'hba264663),
	.w4(32'h3a819e64),
	.w5(32'h3a8b7f04),
	.w6(32'h3b86f876),
	.w7(32'h3b5f04da),
	.w8(32'h39c8289a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9973a7),
	.w1(32'h3a9dda16),
	.w2(32'h3b562532),
	.w3(32'h3bbe2906),
	.w4(32'h3b44ce04),
	.w5(32'h3bf595d3),
	.w6(32'h3be51c89),
	.w7(32'h3b8c9818),
	.w8(32'h3b7311c1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696887),
	.w1(32'hb9df4437),
	.w2(32'hbb4dcb00),
	.w3(32'h3bae4711),
	.w4(32'hb8aec5c3),
	.w5(32'h3a0f848a),
	.w6(32'h3b98e4f4),
	.w7(32'h3b51a7c9),
	.w8(32'h3b192e16),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80277f),
	.w1(32'h3a8f5e78),
	.w2(32'hba9743ca),
	.w3(32'hb9127d03),
	.w4(32'hb9eb4a1b),
	.w5(32'h3a01e2e7),
	.w6(32'h3a34bef9),
	.w7(32'h3a62df3e),
	.w8(32'hba2b9db6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab19c69),
	.w1(32'h3ad13c6e),
	.w2(32'h39fb5723),
	.w3(32'hbaeded02),
	.w4(32'h3b1c0754),
	.w5(32'h3b0631c6),
	.w6(32'hbafe8f22),
	.w7(32'h3b1917ab),
	.w8(32'h3a629ba5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae10c15),
	.w1(32'h3b061b0a),
	.w2(32'h3a049698),
	.w3(32'h3aaa2955),
	.w4(32'h3a1fac21),
	.w5(32'h3bc18ed0),
	.w6(32'h3a39e836),
	.w7(32'hbadc1a8f),
	.w8(32'h3b48a740),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0183ef),
	.w1(32'h3b358b4f),
	.w2(32'hbb3050e5),
	.w3(32'h3ba5b46d),
	.w4(32'h3bbdd5e1),
	.w5(32'h3b492a32),
	.w6(32'h3b58a98a),
	.w7(32'h3b5c75cf),
	.w8(32'hbb04f1e6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7152e7),
	.w1(32'h3ab9e3b9),
	.w2(32'hba6bca5f),
	.w3(32'hbb9884be),
	.w4(32'h3b037500),
	.w5(32'h3ab9d279),
	.w6(32'hbbeb7a0c),
	.w7(32'h3b3cc5ab),
	.w8(32'h39546bf9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba075524),
	.w1(32'hbb28f616),
	.w2(32'hba83888c),
	.w3(32'hba92ff21),
	.w4(32'hbb71bde1),
	.w5(32'hbb662a12),
	.w6(32'hbab981a8),
	.w7(32'hbb4a77de),
	.w8(32'hbb246318),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e9453),
	.w1(32'hba6b9b14),
	.w2(32'h37daa880),
	.w3(32'hbb819de3),
	.w4(32'hbb172228),
	.w5(32'hba93ba8e),
	.w6(32'hbb074c06),
	.w7(32'hbb051f4b),
	.w8(32'hbab1d153),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa132a),
	.w1(32'h3b66c4ca),
	.w2(32'h3a38f993),
	.w3(32'hba310add),
	.w4(32'h3b470ddf),
	.w5(32'h3ae70c49),
	.w6(32'h3aa8c393),
	.w7(32'h3b3043b4),
	.w8(32'h371fb8a0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f755a),
	.w1(32'h3b1bffe6),
	.w2(32'h39170c91),
	.w3(32'hb94988a1),
	.w4(32'h3b3f9a77),
	.w5(32'hbb322f2d),
	.w6(32'hb8c32ddc),
	.w7(32'h3b392534),
	.w8(32'hbb160040),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b33e52),
	.w1(32'h3b3e5309),
	.w2(32'hba2fb930),
	.w3(32'hbac8ba6e),
	.w4(32'h3ba99d7c),
	.w5(32'h3b36c8d5),
	.w6(32'hbad40fd6),
	.w7(32'h3b6d3b69),
	.w8(32'hb9fd90b7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719cfb),
	.w1(32'h3c35b3a5),
	.w2(32'hba6b57a0),
	.w3(32'hbb162a25),
	.w4(32'h3c261483),
	.w5(32'hba8a8b96),
	.w6(32'hbb69aacd),
	.w7(32'h3c370055),
	.w8(32'h398bf489),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af79f64),
	.w1(32'h372a8203),
	.w2(32'h3abbf610),
	.w3(32'h3a80dcb4),
	.w4(32'h3b8d03e5),
	.w5(32'h3c2b3c35),
	.w6(32'h3a00ee13),
	.w7(32'h3a9efb1d),
	.w8(32'h3b95b8e1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba759711),
	.w1(32'h3b5bdb07),
	.w2(32'h3b274983),
	.w3(32'h3a70dd52),
	.w4(32'h3a9f72a7),
	.w5(32'h3ab7a9eb),
	.w6(32'hbaa5e4b9),
	.w7(32'h3b40e50c),
	.w8(32'h3afcefec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05c361),
	.w1(32'hb9528bd9),
	.w2(32'h3acb1eeb),
	.w3(32'h3a36ba37),
	.w4(32'hb4d3fc92),
	.w5(32'h3c12546e),
	.w6(32'h3a17f2ed),
	.w7(32'h3b197c6f),
	.w8(32'h3bc4f2aa),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2a8a3),
	.w1(32'h3aba24ce),
	.w2(32'h3a456a84),
	.w3(32'h3abd9f7e),
	.w4(32'h3b3c2d89),
	.w5(32'h3bae8f6f),
	.w6(32'h3b1be6b6),
	.w7(32'h3b1bbfd1),
	.w8(32'h3b800ae7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7636f),
	.w1(32'h3c034cb0),
	.w2(32'h3a872680),
	.w3(32'h3aed76f9),
	.w4(32'h3baec05a),
	.w5(32'h3ac925ad),
	.w6(32'hbae385e9),
	.w7(32'h3b2776a6),
	.w8(32'h3bc2dce5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae78000),
	.w1(32'h3a146708),
	.w2(32'h3996186b),
	.w3(32'h3b62a520),
	.w4(32'h3aa2f1a7),
	.w5(32'h3a431627),
	.w6(32'h3b760cb0),
	.w7(32'h3af0756e),
	.w8(32'h3b4e69a5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd168f),
	.w1(32'hba3a96fc),
	.w2(32'hba9546e2),
	.w3(32'h3bae5f62),
	.w4(32'h3954e004),
	.w5(32'h3ac4a7d0),
	.w6(32'h3bf3e24c),
	.w7(32'hbb67158b),
	.w8(32'hb9128930),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba979fe4),
	.w1(32'h3b007397),
	.w2(32'hba15d310),
	.w3(32'h3962a9b1),
	.w4(32'h3b3a1aa9),
	.w5(32'h3aebb118),
	.w6(32'h3a67a9a2),
	.w7(32'h3b0e1935),
	.w8(32'h3a9ccafd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d45d),
	.w1(32'h39457319),
	.w2(32'h3aa6d0da),
	.w3(32'hbb342edf),
	.w4(32'h3a757c6d),
	.w5(32'h394de2a2),
	.w6(32'hbb01742a),
	.w7(32'hb92811eb),
	.w8(32'hb97bda5a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adedf21),
	.w1(32'h39da3a36),
	.w2(32'h3aa57d1a),
	.w3(32'h3b059e8c),
	.w4(32'h3b2920d5),
	.w5(32'h3b542479),
	.w6(32'h3b240f57),
	.w7(32'h3b6c0709),
	.w8(32'h3b4ba5f3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32661a),
	.w1(32'hbb6def6e),
	.w2(32'hba916b12),
	.w3(32'h3aec1224),
	.w4(32'hbb097e39),
	.w5(32'hbb4d7446),
	.w6(32'h396610a3),
	.w7(32'h3a3dbc57),
	.w8(32'h3bdead6e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac94779),
	.w1(32'h3a0852f9),
	.w2(32'h3ae46d46),
	.w3(32'hba7ce522),
	.w4(32'hb9674016),
	.w5(32'h39cde7a1),
	.w6(32'h3b8e265b),
	.w7(32'hba9c11f0),
	.w8(32'h3b3256a1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d29ebc),
	.w1(32'h392663be),
	.w2(32'hbb3b3cbe),
	.w3(32'h3a6cdce8),
	.w4(32'hbab009bc),
	.w5(32'h3a531c0e),
	.w6(32'h3abe60b1),
	.w7(32'hbb6fb271),
	.w8(32'hbb268fad),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14f543),
	.w1(32'h3a8a105f),
	.w2(32'h3b4608eb),
	.w3(32'h3990f156),
	.w4(32'hb8908998),
	.w5(32'h3b33dd63),
	.w6(32'hb9f41fcd),
	.w7(32'h3ab5286b),
	.w8(32'h3abe16a3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae96f0),
	.w1(32'h3b6b0ffe),
	.w2(32'h3be3479e),
	.w3(32'h39d57ea6),
	.w4(32'h3b859e7f),
	.w5(32'h3ba2910a),
	.w6(32'h3ae68b40),
	.w7(32'h3b1d443c),
	.w8(32'h3b9a945f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab31674),
	.w1(32'hb89db6a8),
	.w2(32'h3b3bada1),
	.w3(32'h3a54b038),
	.w4(32'h3ac98ca4),
	.w5(32'h3b583edb),
	.w6(32'h3acebb75),
	.w7(32'h3aaf9153),
	.w8(32'h3b74a989),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ce9c0),
	.w1(32'hbb1a8bdc),
	.w2(32'hba8cb603),
	.w3(32'h3b2a6291),
	.w4(32'hbb45fc11),
	.w5(32'hbb013520),
	.w6(32'h3b244fcd),
	.w7(32'hbb10cc03),
	.w8(32'hb9b3e8a2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57f5c4),
	.w1(32'hba5b6fbf),
	.w2(32'hb94e4de4),
	.w3(32'h3b517b00),
	.w4(32'hbaa3537f),
	.w5(32'hbae1d44f),
	.w6(32'h3b2ce90c),
	.w7(32'hba84e001),
	.w8(32'h3a70bcc3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a776b),
	.w1(32'h3b14c64f),
	.w2(32'hbba60093),
	.w3(32'h3b94d769),
	.w4(32'h3bc33045),
	.w5(32'hba3b140a),
	.w6(32'h3b5fd051),
	.w7(32'h3b0fe214),
	.w8(32'hbb11ab46),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c837b),
	.w1(32'h3b8c49de),
	.w2(32'h3a13c4db),
	.w3(32'h3b5c4cf0),
	.w4(32'h3bb4b896),
	.w5(32'h3adea906),
	.w6(32'hba1444bb),
	.w7(32'h3b83a6b1),
	.w8(32'h3aa34d74),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a78d),
	.w1(32'h3b5a8d3e),
	.w2(32'h3b651cd2),
	.w3(32'h3b253564),
	.w4(32'h3ba7f255),
	.w5(32'h3b86b5b3),
	.w6(32'h3919d59d),
	.w7(32'h3b86a5c0),
	.w8(32'h3b22f7f8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a87cc6),
	.w1(32'h3accdee4),
	.w2(32'hba36db53),
	.w3(32'h3ac790fe),
	.w4(32'h392fc292),
	.w5(32'hbbc87550),
	.w6(32'h3aae2f92),
	.w7(32'hb9bb3008),
	.w8(32'hbb4edc99),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c1701),
	.w1(32'h3a4f55bc),
	.w2(32'h3a40c5c4),
	.w3(32'hba92fcd4),
	.w4(32'h3adf25f2),
	.w5(32'h3b4900bb),
	.w6(32'hbb0beb6b),
	.w7(32'h3b080008),
	.w8(32'h3b2bb077),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74d4cf1),
	.w1(32'hba8494a8),
	.w2(32'hbafb6b3c),
	.w3(32'h3a1b2e9b),
	.w4(32'h3a8a8bae),
	.w5(32'h3990ec80),
	.w6(32'h3ab90ba2),
	.w7(32'h3b90cb3e),
	.w8(32'hbab653b8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c24eb),
	.w1(32'h3c07b1e3),
	.w2(32'h3b013aed),
	.w3(32'hba5183f2),
	.w4(32'h3b705e3c),
	.w5(32'h3aa41263),
	.w6(32'hbac8ff62),
	.w7(32'h3b4bc56e),
	.w8(32'h39a4a48b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee896),
	.w1(32'hbb161539),
	.w2(32'hbae69788),
	.w3(32'h3b5ffcb3),
	.w4(32'hbb1fc958),
	.w5(32'hbb1db634),
	.w6(32'h3ac3d420),
	.w7(32'hbb282382),
	.w8(32'hbaef4ab5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a94c9),
	.w1(32'h3a53df28),
	.w2(32'h3afa48fb),
	.w3(32'h3ad42284),
	.w4(32'hbb0bae6e),
	.w5(32'h3b3787b3),
	.w6(32'h3adb4706),
	.w7(32'h399d1b47),
	.w8(32'h3a885c96),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5764d6),
	.w1(32'hb9a54821),
	.w2(32'h3b1dd0f2),
	.w3(32'hbaa7b1e5),
	.w4(32'h3b2d2ef3),
	.w5(32'h3b50a301),
	.w6(32'hba4d66bb),
	.w7(32'h3b39dd1b),
	.w8(32'h3ad532e2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f8965),
	.w1(32'hba76b6b5),
	.w2(32'h3a2678a5),
	.w3(32'hbaeb7727),
	.w4(32'hba42a858),
	.w5(32'h3b76fdc1),
	.w6(32'hba829251),
	.w7(32'hbae715e1),
	.w8(32'h3a98c709),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a4d72),
	.w1(32'h3bb27b9d),
	.w2(32'h3b493609),
	.w3(32'h3a665d33),
	.w4(32'h3bc808ea),
	.w5(32'h3b08b113),
	.w6(32'h38d06f9e),
	.w7(32'h3be77991),
	.w8(32'h3a7af631),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02b781),
	.w1(32'hba1e48ce),
	.w2(32'h3a2af2b7),
	.w3(32'hba155ff4),
	.w4(32'hb9205a09),
	.w5(32'h3ae0c7ff),
	.w6(32'hb90d04fe),
	.w7(32'h3987eb93),
	.w8(32'h3b2c657b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c7a39),
	.w1(32'h3ace8db2),
	.w2(32'hba2baf77),
	.w3(32'hbab0de94),
	.w4(32'h3afb034e),
	.w5(32'h3b171ff3),
	.w6(32'h3a5bde94),
	.w7(32'hbaa8b12c),
	.w8(32'h3a486bf9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4fce4),
	.w1(32'hb9f7891b),
	.w2(32'h3b3281e8),
	.w3(32'h3a5f9289),
	.w4(32'h3a545483),
	.w5(32'h3a9ac190),
	.w6(32'h3b329054),
	.w7(32'hba2a4b75),
	.w8(32'h3ab48216),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d14e),
	.w1(32'h3a9d5e8e),
	.w2(32'h3a885643),
	.w3(32'h3a3a4141),
	.w4(32'h398d4ba1),
	.w5(32'hbaa09005),
	.w6(32'h3b4793b6),
	.w7(32'hbb2cd75b),
	.w8(32'hbaa14322),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80b216),
	.w1(32'hb9b738b1),
	.w2(32'hba3b2009),
	.w3(32'hb9fd0ab4),
	.w4(32'hb96bc6db),
	.w5(32'h3a74f4fa),
	.w6(32'h3a1fcdcd),
	.w7(32'hba51720b),
	.w8(32'h3a05400a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab20d46),
	.w1(32'hbb244146),
	.w2(32'hbbd3a6c7),
	.w3(32'hbae1240e),
	.w4(32'hbb526d15),
	.w5(32'hbbebbfed),
	.w6(32'hba5ca868),
	.w7(32'h3ae1a26f),
	.w8(32'hbba56f81),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e266f),
	.w1(32'hbb0ae29d),
	.w2(32'hbb2d393b),
	.w3(32'hbb165982),
	.w4(32'hbb708d7c),
	.w5(32'hbb0fddb3),
	.w6(32'hbb2d54ff),
	.w7(32'hbb800477),
	.w8(32'hba94cd5b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b33e),
	.w1(32'hbacf4820),
	.w2(32'h3b00af03),
	.w3(32'hbadb22f6),
	.w4(32'h3ac64ddb),
	.w5(32'h3bb36d96),
	.w6(32'hbb0f8899),
	.w7(32'h3a3b361b),
	.w8(32'h3afa6549),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0825f),
	.w1(32'h3bd4e8e8),
	.w2(32'h3be53201),
	.w3(32'h3b0ad459),
	.w4(32'h3ab6704a),
	.w5(32'h3ac72b57),
	.w6(32'h39e8ab97),
	.w7(32'h3b2834fc),
	.w8(32'h3ba12701),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d889e),
	.w1(32'hb92d4625),
	.w2(32'hba5c0a90),
	.w3(32'h3ada3809),
	.w4(32'hba8d1979),
	.w5(32'hba6e191f),
	.w6(32'h3b4e042a),
	.w7(32'hbab2a93e),
	.w8(32'hbad1509c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4be0b8),
	.w1(32'h3a55813d),
	.w2(32'h3b425537),
	.w3(32'h3aad08a0),
	.w4(32'h3adbbc59),
	.w5(32'h3bb3d2fb),
	.w6(32'hb9c6815c),
	.w7(32'h3abc915f),
	.w8(32'h3b355fb1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d2608),
	.w1(32'hba58c4c3),
	.w2(32'hbaf6966c),
	.w3(32'h3b08c8a1),
	.w4(32'hbae48307),
	.w5(32'hbb0b46d8),
	.w6(32'h3afb33f0),
	.w7(32'hbab6f368),
	.w8(32'hbb31989a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9431a5),
	.w1(32'h3a086496),
	.w2(32'hbb439746),
	.w3(32'hbaf9359d),
	.w4(32'hbb4e7228),
	.w5(32'hbbdde229),
	.w6(32'hbab84e23),
	.w7(32'hba94cb2b),
	.w8(32'hbb7bb230),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13be37),
	.w1(32'hba12b551),
	.w2(32'h3acb0faa),
	.w3(32'h3a30f063),
	.w4(32'hbb297acf),
	.w5(32'h3b03fd64),
	.w6(32'h3ada36f8),
	.w7(32'hbb0638e5),
	.w8(32'h3aa41c56),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cd4f5),
	.w1(32'hbb85f8c7),
	.w2(32'hbbd81cf6),
	.w3(32'hb981bc1b),
	.w4(32'hbbcf36f7),
	.w5(32'hbb89f0d1),
	.w6(32'h396704af),
	.w7(32'hbbab00d8),
	.w8(32'hbb7cbc4f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2adb4),
	.w1(32'h3b5a173f),
	.w2(32'h3b8ae6c5),
	.w3(32'hba70bf9b),
	.w4(32'h3b463be0),
	.w5(32'h3b8ae05c),
	.w6(32'hb92c3879),
	.w7(32'h3b2ab0d9),
	.w8(32'h3908cb89),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0acf),
	.w1(32'h3b5f5623),
	.w2(32'h392a3784),
	.w3(32'h396300b1),
	.w4(32'h3c0954e2),
	.w5(32'hbb1e5a38),
	.w6(32'h3a4f7969),
	.w7(32'h3b52c25e),
	.w8(32'hbb96ea81),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a449a),
	.w1(32'h3b91c495),
	.w2(32'hbbd871d4),
	.w3(32'hbb590159),
	.w4(32'h3c74311b),
	.w5(32'hba448a97),
	.w6(32'hbb94975e),
	.w7(32'h3c467ccc),
	.w8(32'hbba451ac),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b6ba4),
	.w1(32'hbb8e2777),
	.w2(32'hbb22d966),
	.w3(32'hbbdd693e),
	.w4(32'h3c171096),
	.w5(32'h3c445821),
	.w6(32'hbbc17ebb),
	.w7(32'h3ba9acd3),
	.w8(32'h3b5985b8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafca6f7),
	.w1(32'h3a5d5690),
	.w2(32'hbbe8d34a),
	.w3(32'h3bc5c70d),
	.w4(32'hbace6d11),
	.w5(32'h3a8cf86b),
	.w6(32'h3b164981),
	.w7(32'hbbb31cfc),
	.w8(32'h3b1e6173),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac13f94),
	.w1(32'hbb0d4f83),
	.w2(32'hbb7e9bcc),
	.w3(32'h3b9f2426),
	.w4(32'h379d8128),
	.w5(32'hbc03f46e),
	.w6(32'hbb05fe84),
	.w7(32'h3af5a2ad),
	.w8(32'hbb61a140),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4dcea),
	.w1(32'h3bf99967),
	.w2(32'h3c2aad17),
	.w3(32'hbc095a4b),
	.w4(32'h3b58fb60),
	.w5(32'h3b6ab65c),
	.w6(32'hbb1cf72a),
	.w7(32'h3ae83d6c),
	.w8(32'hbb7dec18),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0020a2),
	.w1(32'hbb3ada25),
	.w2(32'hbb106e23),
	.w3(32'hbb91198e),
	.w4(32'h3be01d94),
	.w5(32'h3c967f3f),
	.w6(32'hb8b2d969),
	.w7(32'hbc2c3868),
	.w8(32'h3b8f12a7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea8e68),
	.w1(32'h3bc352f5),
	.w2(32'h3bd3cd0b),
	.w3(32'h3c0c7df0),
	.w4(32'h3b867ee7),
	.w5(32'h3c2e8e91),
	.w6(32'h3b9bee9f),
	.w7(32'hba0add44),
	.w8(32'hbaa74e5e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c145e60),
	.w1(32'hbb72393b),
	.w2(32'hbb0f7cff),
	.w3(32'h3b9c2145),
	.w4(32'h3bc58dfb),
	.w5(32'h3a4256f4),
	.w6(32'h3b052393),
	.w7(32'h3ba7e07c),
	.w8(32'hbb09fa4e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaf7e3),
	.w1(32'h3b1c0a76),
	.w2(32'h3b052cba),
	.w3(32'hbaf16d86),
	.w4(32'h3aec0c14),
	.w5(32'h3bacdc8c),
	.w6(32'hbbc33153),
	.w7(32'hbbe17ca0),
	.w8(32'hbc713d17),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93612b),
	.w1(32'hbb430afb),
	.w2(32'hbb101f63),
	.w3(32'h3bf54631),
	.w4(32'hbb6043ee),
	.w5(32'hbaa4e393),
	.w6(32'hbc11b799),
	.w7(32'hbba66fbb),
	.w8(32'h3a912593),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b8fc),
	.w1(32'h39536991),
	.w2(32'hbbb6d147),
	.w3(32'hbb6ad79c),
	.w4(32'h3bdf27f3),
	.w5(32'h3a03db7e),
	.w6(32'hbbc2c6ba),
	.w7(32'h3b2821fd),
	.w8(32'hba943301),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cfcb1),
	.w1(32'hbb99d1fe),
	.w2(32'hbbf008d5),
	.w3(32'hbb2f5c0e),
	.w4(32'hbb6e04c0),
	.w5(32'hbae6cc34),
	.w6(32'hb8ba36b2),
	.w7(32'hbc181a82),
	.w8(32'hbc3057d2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb26359),
	.w1(32'hbb75ccc2),
	.w2(32'h3a4a5c12),
	.w3(32'hbb8fb0bd),
	.w4(32'hbb4b75d1),
	.w5(32'h3b95f595),
	.w6(32'hbc36727e),
	.w7(32'hbbf42ec3),
	.w8(32'hbb1937e9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eb617),
	.w1(32'hbb795626),
	.w2(32'hbc362f98),
	.w3(32'h3c0f16a3),
	.w4(32'hbb36492c),
	.w5(32'hbb9cff0f),
	.w6(32'h3b5892ae),
	.w7(32'hba9ef7e3),
	.w8(32'h3b7be4c1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d6a0d),
	.w1(32'hbb830c49),
	.w2(32'hb9b1e709),
	.w3(32'hbafdb2f1),
	.w4(32'hbba235c9),
	.w5(32'h3b43a636),
	.w6(32'h3a9c2768),
	.w7(32'hba8a8951),
	.w8(32'h3b586d12),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b105817),
	.w1(32'hbbc9d1aa),
	.w2(32'hbb5c3366),
	.w3(32'h3bcc9887),
	.w4(32'h3b257a6f),
	.w5(32'h3b2d74b8),
	.w6(32'h3bb56de0),
	.w7(32'h396438de),
	.w8(32'h3b607663),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4192),
	.w1(32'hbb640ed6),
	.w2(32'hbb49466b),
	.w3(32'h3ae33460),
	.w4(32'hbb38b5d3),
	.w5(32'h3b00679b),
	.w6(32'hbb6bef93),
	.w7(32'hb9daabed),
	.w8(32'h3c005786),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943bb2c),
	.w1(32'hba8ef736),
	.w2(32'h3bdf3b9a),
	.w3(32'h3991504c),
	.w4(32'hbace358b),
	.w5(32'h3cb45aaf),
	.w6(32'h39a32bfc),
	.w7(32'hbb29e7c2),
	.w8(32'h3b288e5e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc680c),
	.w1(32'hba18a513),
	.w2(32'h3c1664f3),
	.w3(32'h3c578e87),
	.w4(32'h3b57266f),
	.w5(32'h3c834670),
	.w6(32'h3c06ce69),
	.w7(32'hbc0a1479),
	.w8(32'hbb8c33f4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2eef2),
	.w1(32'hbc08f213),
	.w2(32'hbb5a9247),
	.w3(32'h3bdd0a20),
	.w4(32'hbbd92395),
	.w5(32'hba847fda),
	.w6(32'h3b6cf5fc),
	.w7(32'hba7611de),
	.w8(32'hba8db4c4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbff6dc),
	.w1(32'hbbff1e1f),
	.w2(32'hbb8d1c48),
	.w3(32'hba97525c),
	.w4(32'hbc192b5d),
	.w5(32'h3aa6701f),
	.w6(32'hbb66a12a),
	.w7(32'hbbfd6e4d),
	.w8(32'hbb7d4da2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed6bb5),
	.w1(32'h39d6e1e8),
	.w2(32'h3b819684),
	.w3(32'h3bfbbd63),
	.w4(32'hbb52bad9),
	.w5(32'hbbe51b2b),
	.w6(32'hbb68690c),
	.w7(32'hbab3b6aa),
	.w8(32'hbb965843),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1adc5),
	.w1(32'hbbb3d9af),
	.w2(32'hbb497dbd),
	.w3(32'h3b192d33),
	.w4(32'hbae91373),
	.w5(32'h3b5627c2),
	.w6(32'hbb056bdb),
	.w7(32'hbc137a8d),
	.w8(32'h3b676515),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20eb0c),
	.w1(32'hbb9e0fe4),
	.w2(32'hbbfb4199),
	.w3(32'h3bce47c4),
	.w4(32'hbba408a9),
	.w5(32'hbbc67137),
	.w6(32'h3b1b58b2),
	.w7(32'hbbb614f8),
	.w8(32'h3ba4e86d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5d98d),
	.w1(32'h395663d6),
	.w2(32'hbb12fefe),
	.w3(32'hbc080a3a),
	.w4(32'hbb7b566a),
	.w5(32'hbbd139af),
	.w6(32'hbbad2983),
	.w7(32'h3b319b66),
	.w8(32'hbb7fbac1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6795ed),
	.w1(32'hbbad2625),
	.w2(32'hbc3a68f3),
	.w3(32'hbb7b2f7b),
	.w4(32'h3abfe1d0),
	.w5(32'h399fe110),
	.w6(32'h3aa7c511),
	.w7(32'hbb1a9b92),
	.w8(32'h3b8b118f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf38e7d),
	.w1(32'h3bdc4586),
	.w2(32'h3b453e56),
	.w3(32'h3a3bf0b4),
	.w4(32'h3c7d0a0f),
	.w5(32'hbc398a1e),
	.w6(32'hb8fa06c6),
	.w7(32'h3bb0ce6c),
	.w8(32'hbc46489f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857549),
	.w1(32'hb88c4c4d),
	.w2(32'h3b997b91),
	.w3(32'hbbbe751d),
	.w4(32'h3c2bb3b5),
	.w5(32'h3c955645),
	.w6(32'hbc4f91fc),
	.w7(32'h3bbc8ab9),
	.w8(32'h3c0ba678),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7e1c),
	.w1(32'hbada3114),
	.w2(32'hbb03e2a7),
	.w3(32'h3b62928b),
	.w4(32'hbb845ba9),
	.w5(32'hbbb569ec),
	.w6(32'h3abf76b6),
	.w7(32'h3aa5bfff),
	.w8(32'h3b0e6cd5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18acaa),
	.w1(32'hbb538a59),
	.w2(32'h39a8107f),
	.w3(32'hbb492ad6),
	.w4(32'hbbce99aa),
	.w5(32'hbc315d90),
	.w6(32'h39d936ba),
	.w7(32'hb93823c1),
	.w8(32'hbb23ef0f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95d8b),
	.w1(32'h3b9e2480),
	.w2(32'h3c29fa4d),
	.w3(32'h3b6c683e),
	.w4(32'hbbae9bc2),
	.w5(32'h3724dcca),
	.w6(32'h3a3ea5df),
	.w7(32'hbb1e96a9),
	.w8(32'hbab4657a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f2e54),
	.w1(32'h3ba04f15),
	.w2(32'h3c1c9b17),
	.w3(32'h3b4b4436),
	.w4(32'h3aa94328),
	.w5(32'h3c5911b1),
	.w6(32'h3a886561),
	.w7(32'h3c067580),
	.w8(32'h3b7edc0b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf8675),
	.w1(32'hbb0594d2),
	.w2(32'hbbd20ba6),
	.w3(32'hb9d8a278),
	.w4(32'h3c977b12),
	.w5(32'h3b5f64e2),
	.w6(32'h3ba7d387),
	.w7(32'h3c54a5de),
	.w8(32'h3c411fc3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178f43),
	.w1(32'hbb2370b9),
	.w2(32'hbb50c890),
	.w3(32'hbbbb85cc),
	.w4(32'h3c2fd600),
	.w5(32'h3c0ae219),
	.w6(32'hbb9711aa),
	.w7(32'h3b6b73ad),
	.w8(32'h3bed8c28),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f7fba),
	.w1(32'hbadc8813),
	.w2(32'h3b421966),
	.w3(32'h3b69ac9e),
	.w4(32'h3c875acf),
	.w5(32'h3c6bdb3b),
	.w6(32'hbb95b632),
	.w7(32'h3c09e431),
	.w8(32'h3c1bf6b2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8633),
	.w1(32'hbb5202dc),
	.w2(32'hbb59f892),
	.w3(32'h3b916507),
	.w4(32'hbb9d0983),
	.w5(32'hbac9ed1f),
	.w6(32'hbbbb5696),
	.w7(32'h3b8c600b),
	.w8(32'h3c41f7fc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8e4f),
	.w1(32'h3a8e7815),
	.w2(32'h3b32a10c),
	.w3(32'hbba8b144),
	.w4(32'hba1bc1d6),
	.w5(32'hbade21ea),
	.w6(32'h3ba7b1db),
	.w7(32'h3bafd2d7),
	.w8(32'h3be69a1a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1a3d2),
	.w1(32'hba6870ca),
	.w2(32'hbb5d557e),
	.w3(32'h3bb9db70),
	.w4(32'h3c3ec253),
	.w5(32'h3c933975),
	.w6(32'h3bbac38b),
	.w7(32'h3a7e4d24),
	.w8(32'h3b1c54e3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a449b),
	.w1(32'h3adcb38b),
	.w2(32'hbc00c0bf),
	.w3(32'hbb64ac75),
	.w4(32'h3b6e92a7),
	.w5(32'hbc437a50),
	.w6(32'hbc0605ed),
	.w7(32'h3bc8f13e),
	.w8(32'hbb074db6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a390),
	.w1(32'hbbd9474a),
	.w2(32'h3b0c920b),
	.w3(32'hbbc3a63e),
	.w4(32'hbb0a5fae),
	.w5(32'h3c2be724),
	.w6(32'hba50740a),
	.w7(32'hbba31fa5),
	.w8(32'h3bcc0ad2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a3ae),
	.w1(32'h3ad07ae1),
	.w2(32'hbbf09a1a),
	.w3(32'hb8845898),
	.w4(32'h3bac47c3),
	.w5(32'hbbee6ee8),
	.w6(32'hbbb8b188),
	.w7(32'h3cada3cb),
	.w8(32'h3c4c871b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf4358),
	.w1(32'hbb85a907),
	.w2(32'hbc033874),
	.w3(32'hbc0d3212),
	.w4(32'hbc4317ea),
	.w5(32'hbbf10672),
	.w6(32'h3b6785d4),
	.w7(32'hbbf45591),
	.w8(32'h3bcf6918),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04b12d),
	.w1(32'h3a44571f),
	.w2(32'h3a29013b),
	.w3(32'hbb0a05b8),
	.w4(32'hbb91a058),
	.w5(32'h3b8983cf),
	.w6(32'h3bfd3832),
	.w7(32'hbb88748c),
	.w8(32'hb99e0ada),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a846501),
	.w1(32'hbaf721ea),
	.w2(32'hba8f7860),
	.w3(32'h3ba32192),
	.w4(32'hbb8b1567),
	.w5(32'hbc28f490),
	.w6(32'hbb515a84),
	.w7(32'hbb30d634),
	.w8(32'hbb973a31),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6ebf),
	.w1(32'hba122c31),
	.w2(32'h3ab85be1),
	.w3(32'hbbb67b34),
	.w4(32'hbb2eeb99),
	.w5(32'h3cc20cec),
	.w6(32'hbb20220d),
	.w7(32'hba9174b1),
	.w8(32'hba32305f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c94e8),
	.w1(32'hba5ccc38),
	.w2(32'hbb701f2d),
	.w3(32'hbc661e36),
	.w4(32'hbbd7be1f),
	.w5(32'h3a9ca10f),
	.w6(32'hbc04fd2e),
	.w7(32'hbb9672a8),
	.w8(32'h3b95fb78),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d01211),
	.w1(32'h399f92cd),
	.w2(32'hbacdd1cf),
	.w3(32'h3bc0d5a0),
	.w4(32'h3abb2987),
	.w5(32'h3b035ae9),
	.w6(32'h3b3b455b),
	.w7(32'h3b77f190),
	.w8(32'h39036dec),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40860f),
	.w1(32'h3b9d8d93),
	.w2(32'hb957efdd),
	.w3(32'hbaf571f3),
	.w4(32'h3bbad0dc),
	.w5(32'hba961fbd),
	.w6(32'hbb3425c4),
	.w7(32'h3b9ce043),
	.w8(32'h3b1f999f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f985b),
	.w1(32'hbb8fa131),
	.w2(32'hbc55b795),
	.w3(32'h386bd275),
	.w4(32'hbb3fdec0),
	.w5(32'hbc58c965),
	.w6(32'hbade46f8),
	.w7(32'h3b58bf03),
	.w8(32'hba454f76),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb02e96),
	.w1(32'hbb770457),
	.w2(32'h3c14fa58),
	.w3(32'hbbee3a4d),
	.w4(32'h39aea09f),
	.w5(32'h3c0607d5),
	.w6(32'hbb31fa6b),
	.w7(32'hbc55575d),
	.w8(32'hbb98415f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df78a),
	.w1(32'hbb534707),
	.w2(32'h3aafee60),
	.w3(32'h3b3ceaa3),
	.w4(32'hbb687dc2),
	.w5(32'h3bd116a5),
	.w6(32'hbb6bd48d),
	.w7(32'hbac6dfa3),
	.w8(32'h3bffd89f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b472b92),
	.w1(32'h3a5824fe),
	.w2(32'h38966b56),
	.w3(32'h3c843682),
	.w4(32'h3b6b0fd7),
	.w5(32'h3bc20330),
	.w6(32'h3c07c3b0),
	.w7(32'h39f9bc1a),
	.w8(32'hb89ccd0f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd543bd),
	.w1(32'h3b541b46),
	.w2(32'h3c01ae29),
	.w3(32'hba939d9f),
	.w4(32'h3baf9a92),
	.w5(32'h3c126b50),
	.w6(32'hbbe7d26b),
	.w7(32'hbb367827),
	.w8(32'hbba91467),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae78456),
	.w1(32'hbbd675cb),
	.w2(32'hbbdd6203),
	.w3(32'hb9315a6b),
	.w4(32'h3bac71df),
	.w5(32'h3c00e7ba),
	.w6(32'hbc0e16f5),
	.w7(32'hba5c27c2),
	.w8(32'h39986df4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d820d),
	.w1(32'hbb7982f2),
	.w2(32'hbbe035ca),
	.w3(32'h3aaebf73),
	.w4(32'h3a867ab7),
	.w5(32'hbbc26e1d),
	.w6(32'hbb852353),
	.w7(32'hbbb0329a),
	.w8(32'hbbb91a94),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800e17),
	.w1(32'h3aa851d1),
	.w2(32'hbbd876f4),
	.w3(32'hbafb2f6b),
	.w4(32'h3b844f95),
	.w5(32'h3b890276),
	.w6(32'hbbaff857),
	.w7(32'h39561e9f),
	.w8(32'h3c146e93),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5665ab),
	.w1(32'h3b24d723),
	.w2(32'h3b14a12f),
	.w3(32'hbb247204),
	.w4(32'hbb184131),
	.w5(32'h3b002477),
	.w6(32'hbaa3f1b6),
	.w7(32'hbaf0534c),
	.w8(32'h3bc5086e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98fbd7),
	.w1(32'hbb09a3a4),
	.w2(32'hbb1a9f74),
	.w3(32'hbb93c1d3),
	.w4(32'hbb9cda0e),
	.w5(32'hbb8e6bd4),
	.w6(32'h3a841b48),
	.w7(32'hb9f456ae),
	.w8(32'h3a3ee7c4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32d5f2),
	.w1(32'hbc00258c),
	.w2(32'h3b52d19e),
	.w3(32'h39a33c59),
	.w4(32'hbb8443f4),
	.w5(32'h3c4a5303),
	.w6(32'h3a0b9eaa),
	.w7(32'hbadff769),
	.w8(32'h3c37a003),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90a674),
	.w1(32'hbb1580aa),
	.w2(32'h39cf13e1),
	.w3(32'h3c173f4e),
	.w4(32'hbb725665),
	.w5(32'h39950c5c),
	.w6(32'h3c1154eb),
	.w7(32'hbb990276),
	.w8(32'h3a09e2c5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c9ff7),
	.w1(32'hb8e0f903),
	.w2(32'hbbc82bb2),
	.w3(32'h3a89b371),
	.w4(32'hbb82b09e),
	.w5(32'hbbe1136c),
	.w6(32'h3b3ab5d8),
	.w7(32'hbbe50321),
	.w8(32'hbbe5eb63),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5358c4),
	.w1(32'h3c1e0474),
	.w2(32'h3c218178),
	.w3(32'h3c13c6ed),
	.w4(32'h3b45b758),
	.w5(32'h3c8e69e6),
	.w6(32'h3a822a04),
	.w7(32'h3c36f365),
	.w8(32'h3be9c684),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ce46),
	.w1(32'hba917c4c),
	.w2(32'hb948aa75),
	.w3(32'hbb629cbe),
	.w4(32'hbc19d0c9),
	.w5(32'h3bca7aba),
	.w6(32'hba2c8a08),
	.w7(32'hbc123546),
	.w8(32'h3bd860ea),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba549d3),
	.w1(32'hbb3f0b57),
	.w2(32'hbb2f0a29),
	.w3(32'h3bc69311),
	.w4(32'h3afd6cfa),
	.w5(32'hbb01754f),
	.w6(32'h3b34f7e2),
	.w7(32'h3afd1f28),
	.w8(32'h3b568c7a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931d59),
	.w1(32'h3a8b1b03),
	.w2(32'hbab3d8a8),
	.w3(32'hb9b6ab03),
	.w4(32'h3b39642b),
	.w5(32'h3b6f72a9),
	.w6(32'hb99e7ce0),
	.w7(32'hbb0a3d7e),
	.w8(32'h3a6a24c3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a8534),
	.w1(32'h3be10e6d),
	.w2(32'h3c94fc0d),
	.w3(32'h3b526d30),
	.w4(32'h3bd25874),
	.w5(32'h3bfb68ea),
	.w6(32'hbbc6445b),
	.w7(32'hbbd11b2b),
	.w8(32'hbc145609),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba66dda),
	.w1(32'h3bedfd0e),
	.w2(32'h3bf0b1db),
	.w3(32'h3abfb673),
	.w4(32'hbc05623a),
	.w5(32'hbc2b783c),
	.w6(32'hbbc0cc8e),
	.w7(32'hbba92bee),
	.w8(32'hbc83d7ba),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2acb7),
	.w1(32'hbab003da),
	.w2(32'h3bb408e9),
	.w3(32'hbb60fe11),
	.w4(32'h3bf59e66),
	.w5(32'h3be40d12),
	.w6(32'hbc289474),
	.w7(32'h3b72b2a2),
	.w8(32'h3a3fa3a8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dd5cc),
	.w1(32'hbbc86c86),
	.w2(32'hba6f16d8),
	.w3(32'hbbad9318),
	.w4(32'hbba8ad4a),
	.w5(32'h3bc1ee5b),
	.w6(32'hbba5ecac),
	.w7(32'h3ae3a068),
	.w8(32'h3c0ae398),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1b84),
	.w1(32'hbb2abb5c),
	.w2(32'hb8be3d5c),
	.w3(32'h3c070285),
	.w4(32'h3babc47c),
	.w5(32'h3bfeaac5),
	.w6(32'h38040d17),
	.w7(32'h3b55df94),
	.w8(32'h3be88632),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fea38),
	.w1(32'h3b37c1e2),
	.w2(32'h3b40c36d),
	.w3(32'h3b44c0df),
	.w4(32'h3bd54027),
	.w5(32'h3bc087c9),
	.w6(32'h3b3f9c12),
	.w7(32'h3a4e0234),
	.w8(32'hbb4adbae),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4ff58),
	.w1(32'hbbda9638),
	.w2(32'hbc716571),
	.w3(32'h3b77d182),
	.w4(32'hbbe30811),
	.w5(32'hbc15e273),
	.w6(32'hba1fc62a),
	.w7(32'hbbc6b2c8),
	.w8(32'hbc0294c3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb23509),
	.w1(32'hbbf79748),
	.w2(32'hbc3a490a),
	.w3(32'hbb4235d8),
	.w4(32'h397bbcb9),
	.w5(32'hbc5e3392),
	.w6(32'hbb40a67e),
	.w7(32'h3b43f01c),
	.w8(32'hbb88358b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6cd9e),
	.w1(32'hba916e0c),
	.w2(32'hbb2b707a),
	.w3(32'hbc093d32),
	.w4(32'h3b99dd5c),
	.w5(32'h3c100e7e),
	.w6(32'hbbe6f244),
	.w7(32'hbb413277),
	.w8(32'hb888547d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0163),
	.w1(32'h3be44805),
	.w2(32'hbad9a1f7),
	.w3(32'hba7ce695),
	.w4(32'h3cbb250f),
	.w5(32'h3c5c3697),
	.w6(32'hbba5df5a),
	.w7(32'h3c00ac3a),
	.w8(32'hb939b618),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc239381),
	.w1(32'h3c23cf96),
	.w2(32'h3b070b57),
	.w3(32'hbbb87099),
	.w4(32'h3b8a2d19),
	.w5(32'h3a9881bd),
	.w6(32'hbbfdf08d),
	.w7(32'hbb100a6b),
	.w8(32'hbb4990e6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5fac8),
	.w1(32'h3bbab808),
	.w2(32'h3bebcdc4),
	.w3(32'h3b0ff93d),
	.w4(32'h3b6f028d),
	.w5(32'hbb1bbf0c),
	.w6(32'h3b36201a),
	.w7(32'h3ba4668b),
	.w8(32'h3aeb60a1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3780806c),
	.w1(32'hb95a14b2),
	.w2(32'hbb46ad5d),
	.w3(32'hbb574e0e),
	.w4(32'h3c04e850),
	.w5(32'h3c7525fa),
	.w6(32'hb9fd1888),
	.w7(32'h3bd08662),
	.w8(32'h3b938f36),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a12b),
	.w1(32'hbb17e76b),
	.w2(32'h3bec6c80),
	.w3(32'h3b98288b),
	.w4(32'hbc354f08),
	.w5(32'hbb811117),
	.w6(32'h3a1c3e18),
	.w7(32'hbc06eee7),
	.w8(32'hbb4f6dd3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcf9d1),
	.w1(32'h3af9b2f4),
	.w2(32'h39fcb08c),
	.w3(32'h3bde33d0),
	.w4(32'h3c4d7a92),
	.w5(32'h3c6c9232),
	.w6(32'h3adfa388),
	.w7(32'h3b9b7f69),
	.w8(32'h3ba639e1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c904),
	.w1(32'hbc01d664),
	.w2(32'hbba0efa9),
	.w3(32'hbb2c8aa4),
	.w4(32'hbc3d6d22),
	.w5(32'hbaae2310),
	.w6(32'hbbc6a692),
	.w7(32'hbb344c47),
	.w8(32'h3b2ca8c5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818e9b),
	.w1(32'hbb8f911e),
	.w2(32'h3b75ff39),
	.w3(32'hba88f53f),
	.w4(32'hbb64a8d7),
	.w5(32'hbb47951d),
	.w6(32'hba3317fd),
	.w7(32'h3a3318d9),
	.w8(32'hbab1e4cb),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38626333),
	.w1(32'h3bd1b831),
	.w2(32'h3b10e806),
	.w3(32'hbc056388),
	.w4(32'h3ccaa2cd),
	.w5(32'h3cc6f3ef),
	.w6(32'h3aa20d96),
	.w7(32'h3bccf1f9),
	.w8(32'h3b1a405d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04cbcb),
	.w1(32'h3b6219c2),
	.w2(32'h3b2651e0),
	.w3(32'h3c7acea4),
	.w4(32'h3ba720eb),
	.w5(32'hbb7214cd),
	.w6(32'hbb9c5c5f),
	.w7(32'h3c5e45f1),
	.w8(32'h3ba738cf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57691d),
	.w1(32'h3c0a2719),
	.w2(32'hba5a52f3),
	.w3(32'hbba8ac07),
	.w4(32'h3c050817),
	.w5(32'h3aea1df0),
	.w6(32'hbb1c93db),
	.w7(32'h3bc3cf7f),
	.w8(32'h3b8814b6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6a5b),
	.w1(32'h3bae57e4),
	.w2(32'h3a466520),
	.w3(32'h3afc912b),
	.w4(32'h389aa178),
	.w5(32'h3999228b),
	.w6(32'hb9b86969),
	.w7(32'hb9a7b954),
	.w8(32'hbb02d077),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43b2f5),
	.w1(32'h3b1c2b72),
	.w2(32'h3be3060d),
	.w3(32'h3b3b5d22),
	.w4(32'h3c14f492),
	.w5(32'h3aa4c2ab),
	.w6(32'hbb8e4650),
	.w7(32'h3b62a6d5),
	.w8(32'hbb1e6264),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57ab68),
	.w1(32'h3bd107ae),
	.w2(32'h3c8661e8),
	.w3(32'hbb710ab7),
	.w4(32'h3c3c06b0),
	.w5(32'h3b187dbe),
	.w6(32'hbc0669b9),
	.w7(32'h3a9bf33a),
	.w8(32'hbbe4dbe9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817e9c),
	.w1(32'hbb257b40),
	.w2(32'hbb2ff945),
	.w3(32'hbb885fe4),
	.w4(32'h38233f99),
	.w5(32'hbb1a01f4),
	.w6(32'hbbfb7399),
	.w7(32'hbb9589ae),
	.w8(32'hbb33d564),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac91980),
	.w1(32'h3b97dbaf),
	.w2(32'h3b554284),
	.w3(32'hba6440fb),
	.w4(32'h3b08fdd4),
	.w5(32'h3a658a24),
	.w6(32'hbb9a985b),
	.w7(32'hbbaf4674),
	.w8(32'hbb82e677),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f9e3),
	.w1(32'hbb697303),
	.w2(32'h3aaaf508),
	.w3(32'h3ba5a608),
	.w4(32'hbbd65799),
	.w5(32'h3b42b0e0),
	.w6(32'hb9374a09),
	.w7(32'hbbba2dfb),
	.w8(32'hbaaebc99),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae90582),
	.w1(32'hbb8f80e6),
	.w2(32'h3ba5e35a),
	.w3(32'h3c6c87d0),
	.w4(32'hbc03ccb0),
	.w5(32'hbb9d860f),
	.w6(32'h3af3410b),
	.w7(32'hbb3a4d86),
	.w8(32'hbc38051c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1744d2),
	.w1(32'h3b617ac2),
	.w2(32'h3b84107e),
	.w3(32'hbb2b1f54),
	.w4(32'hb8e3eb81),
	.w5(32'hbc1e6173),
	.w6(32'hbb9ae70f),
	.w7(32'h3a9d919e),
	.w8(32'hbc0cefb7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74bb44),
	.w1(32'hba62950d),
	.w2(32'hbc6a798d),
	.w3(32'hbbabae15),
	.w4(32'h3c18a68d),
	.w5(32'hb9910a62),
	.w6(32'hbb8aeac6),
	.w7(32'h3c1e2370),
	.w8(32'h3bd63cd0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43b0d8),
	.w1(32'hbbac4b61),
	.w2(32'hbbb17379),
	.w3(32'hba413a48),
	.w4(32'hbba31221),
	.w5(32'hbb3b4d77),
	.w6(32'hba1e53e7),
	.w7(32'hbc106250),
	.w8(32'hbc11a845),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c1992),
	.w1(32'h3b3a6203),
	.w2(32'h3c24d3c4),
	.w3(32'hbabde002),
	.w4(32'h3c8df13b),
	.w5(32'h3ca8af39),
	.w6(32'hbbcc5d24),
	.w7(32'h3ae004d0),
	.w8(32'h3c3aee93),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17bcac),
	.w1(32'hba4c4264),
	.w2(32'h3ae18688),
	.w3(32'h3c29264f),
	.w4(32'hbb4ffe06),
	.w5(32'h3ab8aab9),
	.w6(32'h3b720e2d),
	.w7(32'hbb8ce37e),
	.w8(32'hbbe188ba),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c068e86),
	.w1(32'hbc265335),
	.w2(32'hbc185d7b),
	.w3(32'h3c7aa295),
	.w4(32'h3923cfbe),
	.w5(32'hbbb044a9),
	.w6(32'h38e1a0a7),
	.w7(32'h3a1e75d2),
	.w8(32'hbbaba07e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f1911),
	.w1(32'hbb458d50),
	.w2(32'h3a7c731f),
	.w3(32'hb9d5d7a1),
	.w4(32'hbada0ddf),
	.w5(32'h3c5e6099),
	.w6(32'hbb7644ab),
	.w7(32'hbaa11c2e),
	.w8(32'h3bc6e6c5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5de677),
	.w1(32'h3c1f6788),
	.w2(32'h3a9142a4),
	.w3(32'h3bbd408d),
	.w4(32'h3c376848),
	.w5(32'hbb07edfa),
	.w6(32'h3b78450c),
	.w7(32'hbc07f6d6),
	.w8(32'hbbb47ca0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbea125),
	.w1(32'hbbd7b598),
	.w2(32'hbb704165),
	.w3(32'hbad7208c),
	.w4(32'h3bb834cd),
	.w5(32'h3b4ceeb8),
	.w6(32'hbbfbadd4),
	.w7(32'h3a914c87),
	.w8(32'h3b6420fc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd88683),
	.w1(32'hbbe11e24),
	.w2(32'hbc0c9114),
	.w3(32'h3bc1e390),
	.w4(32'hbc050a82),
	.w5(32'h3a66975d),
	.w6(32'h3b86912b),
	.w7(32'hbc5efb9c),
	.w8(32'h3b1d199d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5d31),
	.w1(32'h39c76b4f),
	.w2(32'h3b848e36),
	.w3(32'h3bab979e),
	.w4(32'hbbba561d),
	.w5(32'h3bd66fab),
	.w6(32'h3b285dcf),
	.w7(32'hbb574d5f),
	.w8(32'h3bbe3905),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32e232),
	.w1(32'h3ba8410a),
	.w2(32'hb9b26f95),
	.w3(32'h3ab4fba9),
	.w4(32'h3c0a4ac5),
	.w5(32'hbac78c4e),
	.w6(32'hba9ed335),
	.w7(32'h3b20d331),
	.w8(32'hba9a3075),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3020ce),
	.w1(32'h3b926f91),
	.w2(32'h3b846792),
	.w3(32'h3a8e7d4d),
	.w4(32'h3cbbb099),
	.w5(32'h3c6f09d7),
	.w6(32'h3bb94fed),
	.w7(32'h3b3f7ad6),
	.w8(32'hbb02dee0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd3ba7),
	.w1(32'hbb5ae04b),
	.w2(32'hbbe1dcad),
	.w3(32'h3bb9cd91),
	.w4(32'hbbf0e19f),
	.w5(32'hbc2556fd),
	.w6(32'hbb87a96b),
	.w7(32'hbbb18759),
	.w8(32'hba16c5a3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbedf4),
	.w1(32'h3b017ee0),
	.w2(32'h396f506d),
	.w3(32'hbc3113f9),
	.w4(32'h3c74305b),
	.w5(32'h3a2382e5),
	.w6(32'h3b09231e),
	.w7(32'h3bc811c6),
	.w8(32'hbbccc991),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0f9b),
	.w1(32'h3b8ac30c),
	.w2(32'h3b510bc2),
	.w3(32'hbb2d8118),
	.w4(32'h3b4dfb58),
	.w5(32'hb8c15b9e),
	.w6(32'hbbfe9cc1),
	.w7(32'h3a9cd89a),
	.w8(32'hbb0d858d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60521f),
	.w1(32'hbbe708cc),
	.w2(32'hbb3ac575),
	.w3(32'hbb9f27af),
	.w4(32'hbbf5cd9e),
	.w5(32'hbaba6788),
	.w6(32'hbc2ed0ab),
	.w7(32'hbc78c678),
	.w8(32'hbb9d41cb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aafed),
	.w1(32'h39959f9e),
	.w2(32'hba6bd686),
	.w3(32'h3c1f94b1),
	.w4(32'h3baa39a9),
	.w5(32'h3bfc58ba),
	.w6(32'h3b3124a7),
	.w7(32'h3a9cdc00),
	.w8(32'h3b8d065f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07422),
	.w1(32'h3bec0fbe),
	.w2(32'h3b640146),
	.w3(32'h3b644f28),
	.w4(32'h3c6202c2),
	.w5(32'h3bf59e9a),
	.w6(32'hbb1bb19a),
	.w7(32'h3c22e773),
	.w8(32'h395f7378),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf60da4),
	.w1(32'hbb7ac6d5),
	.w2(32'h39f5da40),
	.w3(32'h3a1193c1),
	.w4(32'h37c89952),
	.w5(32'hbaed8f63),
	.w6(32'h3abfd617),
	.w7(32'hbbb567a7),
	.w8(32'hbc13785d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa49dcc),
	.w1(32'hbc146438),
	.w2(32'hbba28436),
	.w3(32'h3b0b427b),
	.w4(32'hbb90dd2a),
	.w5(32'hbb142039),
	.w6(32'hbbc0ef96),
	.w7(32'hb8fafdf1),
	.w8(32'hbbd2a128),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb964d40),
	.w1(32'h3b05f24e),
	.w2(32'h3c1dec45),
	.w3(32'hbba14bb0),
	.w4(32'h3b4ac147),
	.w5(32'h3c869e29),
	.w6(32'hbb830932),
	.w7(32'hba36802b),
	.w8(32'h3c0452d6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2473d),
	.w1(32'hbb67b0a6),
	.w2(32'hb9f78231),
	.w3(32'h3c5d0eef),
	.w4(32'h3a66545e),
	.w5(32'h3b9abda1),
	.w6(32'h3ba44d13),
	.w7(32'hb766396f),
	.w8(32'hbafff6af),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9ab99),
	.w1(32'hbbcbfaeb),
	.w2(32'hbae5e815),
	.w3(32'h3b9edd6e),
	.w4(32'hbb59ea00),
	.w5(32'h3bd36304),
	.w6(32'hbaff02cb),
	.w7(32'hbc086e90),
	.w8(32'hbb1d2516),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3b1d),
	.w1(32'h3ae5a3ab),
	.w2(32'h3a9561f4),
	.w3(32'h3b8082e0),
	.w4(32'hbb066e01),
	.w5(32'h3b883415),
	.w6(32'hbb1a3597),
	.w7(32'hbb12df8e),
	.w8(32'h3b4c4f7e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940847),
	.w1(32'hbb36ad64),
	.w2(32'h3b06ae5f),
	.w3(32'h3af79c1a),
	.w4(32'hba34152f),
	.w5(32'h3c0baefb),
	.w6(32'hbb289ca1),
	.w7(32'hba0075f0),
	.w8(32'h3b6f1200),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3bec4),
	.w1(32'hbb62a7d5),
	.w2(32'hbbfd1a92),
	.w3(32'hba70d2ca),
	.w4(32'h3a8feda8),
	.w5(32'hbb347b6a),
	.w6(32'hbb13940b),
	.w7(32'h3b5dbb96),
	.w8(32'hb8621dfd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae85418),
	.w1(32'h3a48c27e),
	.w2(32'hb97270c0),
	.w3(32'hbb21bf7b),
	.w4(32'h3bc479ed),
	.w5(32'h3c09dec4),
	.w6(32'h3b6138bb),
	.w7(32'h3bad33c5),
	.w8(32'h3c032b0e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66b9f),
	.w1(32'hb9a3c22a),
	.w2(32'h3ba7d2ba),
	.w3(32'h3bee76e1),
	.w4(32'hbadaa7c2),
	.w5(32'hba846a0c),
	.w6(32'h3bb6c1dc),
	.w7(32'hbb8da61a),
	.w8(32'h3a1f78c7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcacd02),
	.w1(32'h3ad75952),
	.w2(32'h3b9c82fc),
	.w3(32'h3b87c6d6),
	.w4(32'h3a537a5c),
	.w5(32'h3c0f63b1),
	.w6(32'h3ab362dc),
	.w7(32'h38cf2c68),
	.w8(32'h3c0f4f26),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ef896),
	.w1(32'h3891b08a),
	.w2(32'hba5f0098),
	.w3(32'h3c66e50c),
	.w4(32'hbaa1f4d7),
	.w5(32'h3b0b576a),
	.w6(32'h3c80c99f),
	.w7(32'h3ab9348e),
	.w8(32'hba84e680),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb361c27),
	.w1(32'hbc2b6ff6),
	.w2(32'hbc365903),
	.w3(32'hba5d50c1),
	.w4(32'hbc15d9ac),
	.w5(32'hbb680143),
	.w6(32'hbb496c86),
	.w7(32'hbc89d696),
	.w8(32'hbc4729bc),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc653dde),
	.w1(32'hbadf7b8e),
	.w2(32'h3b23a4ec),
	.w3(32'hbc1401ca),
	.w4(32'h3bfd53b4),
	.w5(32'h3ad97b16),
	.w6(32'hbc82adbd),
	.w7(32'hba7cb530),
	.w8(32'hbb63214f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8bf2e),
	.w1(32'h3b641e44),
	.w2(32'hbb02accd),
	.w3(32'hb63617e2),
	.w4(32'hbaeab9ef),
	.w5(32'hbc80db2d),
	.w6(32'hbbd68d5f),
	.w7(32'h3c16df28),
	.w8(32'hbace8438),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40f9fa),
	.w1(32'h3badc933),
	.w2(32'h3b8cafa8),
	.w3(32'h3b0fa922),
	.w4(32'h3bf33719),
	.w5(32'hba2f6b46),
	.w6(32'h3c155e57),
	.w7(32'h3c1f27d6),
	.w8(32'h3babcb37),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c9f26),
	.w1(32'hb8f8496f),
	.w2(32'hbaa02ab4),
	.w3(32'hbb106758),
	.w4(32'h3be891c0),
	.w5(32'h3a82a97f),
	.w6(32'hbb9db2aa),
	.w7(32'hb9f7dcb1),
	.w8(32'h38c637a9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc661eed),
	.w1(32'hba0d8551),
	.w2(32'hbaf1c338),
	.w3(32'hbc128659),
	.w4(32'h36d7afbd),
	.w5(32'hb98aa801),
	.w6(32'hbc316f97),
	.w7(32'hba00b679),
	.w8(32'h39b95142),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1672c),
	.w1(32'hb6dbe429),
	.w2(32'hb9aab98c),
	.w3(32'hbaa0cdde),
	.w4(32'hba221ede),
	.w5(32'hba0c8292),
	.w6(32'hba078ca3),
	.w7(32'hbaa76441),
	.w8(32'hba3e6cfd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba370f13),
	.w1(32'h3a3476b4),
	.w2(32'h3a667ec8),
	.w3(32'hba5a7b42),
	.w4(32'hbac26420),
	.w5(32'hba8ebb3c),
	.w6(32'hb98ea62b),
	.w7(32'hba1c0479),
	.w8(32'h3aadf119),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69fc16),
	.w1(32'hb9c36b5e),
	.w2(32'hbac43cc1),
	.w3(32'h3aa43140),
	.w4(32'h3a7d0ca5),
	.w5(32'hba34e14a),
	.w6(32'h3acae2a5),
	.w7(32'hb95de9ab),
	.w8(32'hba264388),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba924f58),
	.w1(32'hba5ce1f0),
	.w2(32'h3948ef81),
	.w3(32'hbae22952),
	.w4(32'hba23ae37),
	.w5(32'hba84d250),
	.w6(32'hba986f67),
	.w7(32'hba800733),
	.w8(32'hba4e1fce),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb2524),
	.w1(32'hb9fd20e5),
	.w2(32'hba18976c),
	.w3(32'hb987efa1),
	.w4(32'h399cda1b),
	.w5(32'hb92c1935),
	.w6(32'hba7b6d8b),
	.w7(32'hbad9e8fa),
	.w8(32'hba8c97a3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81b764),
	.w1(32'h3948f461),
	.w2(32'h3a397141),
	.w3(32'h390bc0ff),
	.w4(32'hb8510f59),
	.w5(32'hba8876a7),
	.w6(32'hbace8751),
	.w7(32'hbaa29b2e),
	.w8(32'hb9b600a5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b96b94),
	.w1(32'hbb1a7175),
	.w2(32'hbb577608),
	.w3(32'hb9640021),
	.w4(32'hbb5a9033),
	.w5(32'hbb3f521c),
	.w6(32'hba512b57),
	.w7(32'hbb33ea3c),
	.w8(32'hbb5bede1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bf8b1),
	.w1(32'hba925d9d),
	.w2(32'hb85c63da),
	.w3(32'hba8f9631),
	.w4(32'hb91c600c),
	.w5(32'h3a8d9346),
	.w6(32'hba7f5faa),
	.w7(32'hb9888870),
	.w8(32'h3ad8f1f9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a932bbb),
	.w1(32'h3ab81ccb),
	.w2(32'h3aa0637b),
	.w3(32'h39ae2ebc),
	.w4(32'h3afc72e4),
	.w5(32'h3b13db3e),
	.w6(32'hb8a02681),
	.w7(32'h3a5696a8),
	.w8(32'h3ad005b0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4974c),
	.w1(32'hbac24c6a),
	.w2(32'hba8b490f),
	.w3(32'h3aae9a81),
	.w4(32'hbad009d0),
	.w5(32'hbaf5348d),
	.w6(32'h3a20da47),
	.w7(32'hbab2016b),
	.w8(32'hbb28f1e2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ad276),
	.w1(32'h3ad6260c),
	.w2(32'h3adb35ef),
	.w3(32'hba92adfa),
	.w4(32'h3ac23f69),
	.w5(32'h3a673efb),
	.w6(32'hba96ce2c),
	.w7(32'h3b398488),
	.w8(32'h3b656b62),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a049643),
	.w1(32'h3a008231),
	.w2(32'h3a302bca),
	.w3(32'h3a839b09),
	.w4(32'hb9e96f7a),
	.w5(32'h38d51c8c),
	.w6(32'h3b098a86),
	.w7(32'hb949dbe7),
	.w8(32'hba259630),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10bd3c),
	.w1(32'h383ffe7e),
	.w2(32'h3a315cdd),
	.w3(32'hbab87522),
	.w4(32'hba4a9bb7),
	.w5(32'h39a8b5ba),
	.w6(32'hbaa37331),
	.w7(32'hb988b8e3),
	.w8(32'h3a7d37b5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c672e8),
	.w1(32'h3a415dae),
	.w2(32'hbab68670),
	.w3(32'hb9dacd57),
	.w4(32'h3a7ca935),
	.w5(32'hb78843c6),
	.w6(32'h3a0f4611),
	.w7(32'hba5a76ab),
	.w8(32'hbaa815ab),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92aeef),
	.w1(32'hba7a1391),
	.w2(32'hb9bcac47),
	.w3(32'hbaf25861),
	.w4(32'hbabd42b6),
	.w5(32'hba009d00),
	.w6(32'hbb20428b),
	.w7(32'hba3f9ebf),
	.w8(32'hb8256672),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa8b9a),
	.w1(32'hbabd69aa),
	.w2(32'h3a1f033f),
	.w3(32'hbae7df1c),
	.w4(32'hbb1f956e),
	.w5(32'h3a49d0b3),
	.w6(32'hba0fdd16),
	.w7(32'hbadf95ae),
	.w8(32'hb8cc2f84),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37b956),
	.w1(32'hba63610d),
	.w2(32'hba81c111),
	.w3(32'h3949da1b),
	.w4(32'h3917ecfd),
	.w5(32'hb8fe563a),
	.w6(32'h3a6b5c34),
	.w7(32'h3abe4bc2),
	.w8(32'h3a850dc6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6a327),
	.w1(32'hba13be7b),
	.w2(32'hbab4d2cc),
	.w3(32'hb9e84cc7),
	.w4(32'hb9f18606),
	.w5(32'hbb51a898),
	.w6(32'hb9d39e1d),
	.w7(32'h3a054d83),
	.w8(32'hba0dc69f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cb473),
	.w1(32'h38ed55b7),
	.w2(32'hbac94261),
	.w3(32'hba8abea4),
	.w4(32'h392ed2f5),
	.w5(32'hba8c9747),
	.w6(32'hba957a13),
	.w7(32'hbab99f0c),
	.w8(32'hbb00587f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba443a),
	.w1(32'h3b0eff04),
	.w2(32'h3a8991ce),
	.w3(32'hba316602),
	.w4(32'h3b1ea1a0),
	.w5(32'h3a9ca70d),
	.w6(32'hba35ae13),
	.w7(32'h3ad5b7a3),
	.w8(32'h3a0ec2e8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeba2d3),
	.w1(32'hbac003b0),
	.w2(32'hba86d5d1),
	.w3(32'h3a6da693),
	.w4(32'hbaace37e),
	.w5(32'hba07fa7f),
	.w6(32'hb8c8f2f7),
	.w7(32'hbaa75fe3),
	.w8(32'hbaa12e3f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba877f06),
	.w1(32'h3aa3bb1b),
	.w2(32'h3a00d8cc),
	.w3(32'hbaf24f8a),
	.w4(32'h3adf575b),
	.w5(32'h3b0e9308),
	.w6(32'hbafd848a),
	.w7(32'h3a1687ad),
	.w8(32'h3a045c82),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb844262b),
	.w1(32'h3b0917b5),
	.w2(32'h3b1e0721),
	.w3(32'h3a80cd9f),
	.w4(32'h3ad2b653),
	.w5(32'h3a92a172),
	.w6(32'hb8d03b6b),
	.w7(32'h3ad68355),
	.w8(32'h3afec782),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a413775),
	.w1(32'h38e239e1),
	.w2(32'h3a1b660f),
	.w3(32'h3a4c0c76),
	.w4(32'h3a826cf1),
	.w5(32'h3a953335),
	.w6(32'h3af91630),
	.w7(32'h39a1d559),
	.w8(32'h39e51005),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a2db0),
	.w1(32'hba5937ab),
	.w2(32'h38237e78),
	.w3(32'hb9874d9a),
	.w4(32'hb98cca43),
	.w5(32'h39941a52),
	.w6(32'hb70c59fa),
	.w7(32'hb8d5202d),
	.w8(32'h39848600),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39184030),
	.w1(32'hb9fcc042),
	.w2(32'hbaf69dfc),
	.w3(32'hbaa8c09b),
	.w4(32'hba875892),
	.w5(32'hba0ca6cb),
	.w6(32'hb9f62bc1),
	.w7(32'hb9c31a3b),
	.w8(32'hba73f64c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa089ca),
	.w1(32'hb97af77d),
	.w2(32'h3a268870),
	.w3(32'hb93ac0fa),
	.w4(32'hba225b94),
	.w5(32'h3aa9ba68),
	.w6(32'h3a0a4871),
	.w7(32'hb963965b),
	.w8(32'hb9ed0db3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a823310),
	.w1(32'hb8436b14),
	.w2(32'h3a1ecadd),
	.w3(32'h3a1c6029),
	.w4(32'hbabc21f7),
	.w5(32'h39b23afd),
	.w6(32'h3a3d765e),
	.w7(32'hba78429b),
	.w8(32'h3a113cac),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961e699),
	.w1(32'h3adad111),
	.w2(32'h399936b8),
	.w3(32'h394bb81f),
	.w4(32'h3b0cde19),
	.w5(32'h3a7a74ff),
	.w6(32'h38fb1bb5),
	.w7(32'h3af902f7),
	.w8(32'hb9eea2e5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab7d5e),
	.w1(32'h3aa21232),
	.w2(32'h3a7b0aa8),
	.w3(32'h3922267d),
	.w4(32'h3a98666c),
	.w5(32'h3aaac974),
	.w6(32'hba0c1244),
	.w7(32'hba7763a7),
	.w8(32'h375a3063),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92bd95),
	.w1(32'h381b46ba),
	.w2(32'h39bad58f),
	.w3(32'h3ad1e690),
	.w4(32'h3a5c65ea),
	.w5(32'hb9a5babc),
	.w6(32'hb8e80fa6),
	.w7(32'h3a332e31),
	.w8(32'hb8f32554),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8196c4),
	.w1(32'hba5e74df),
	.w2(32'hba0a0438),
	.w3(32'h39d579ae),
	.w4(32'hbaccbdd7),
	.w5(32'h3a460e01),
	.w6(32'h3a5fe626),
	.w7(32'hbaef12e7),
	.w8(32'hba49ae31),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7455e5),
	.w1(32'hb9a61037),
	.w2(32'hbaa4649b),
	.w3(32'hba9b5293),
	.w4(32'hbab845eb),
	.w5(32'hbb0c4c3b),
	.w6(32'h394a98a9),
	.w7(32'hb9a2f5a2),
	.w8(32'hb8fe04e1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b2dbb),
	.w1(32'h3a556975),
	.w2(32'h399ccea9),
	.w3(32'h3a0ed08b),
	.w4(32'hba162ec2),
	.w5(32'hba038dd8),
	.w6(32'h3a75fdcc),
	.w7(32'hb885f10b),
	.w8(32'hb9987ddc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb051bbc),
	.w1(32'h39f93cbe),
	.w2(32'h39f0e565),
	.w3(32'hbb482472),
	.w4(32'h394748fd),
	.w5(32'hb8f8178d),
	.w6(32'hba6482b2),
	.w7(32'hb985e747),
	.w8(32'h3a875e95),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82ad643),
	.w1(32'hb9526212),
	.w2(32'h39f4f828),
	.w3(32'h3a30cc55),
	.w4(32'hba662174),
	.w5(32'h37ccb38c),
	.w6(32'h3acc7113),
	.w7(32'hba4f132c),
	.w8(32'hb9d76604),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d319b),
	.w1(32'h3ab4b85d),
	.w2(32'h3ab814c7),
	.w3(32'hb930853e),
	.w4(32'h3a289f5b),
	.w5(32'h392e783e),
	.w6(32'hb952b875),
	.w7(32'h384d5c17),
	.w8(32'h399003d3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a842521),
	.w1(32'h39aa93c4),
	.w2(32'h39753cf7),
	.w3(32'hb91f3276),
	.w4(32'h3a48866a),
	.w5(32'h3b0697e5),
	.w6(32'hb9833667),
	.w7(32'h39af7d38),
	.w8(32'h3a81777b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba720ebb),
	.w1(32'hba002e16),
	.w2(32'h3979c12f),
	.w3(32'hb922bee9),
	.w4(32'hb9c62ab1),
	.w5(32'hba44e432),
	.w6(32'hba043c8a),
	.w7(32'hb9999e7f),
	.w8(32'h3a479b22),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e2b3d),
	.w1(32'hba9cb0e9),
	.w2(32'hbac93164),
	.w3(32'hb91b7a25),
	.w4(32'hba036e17),
	.w5(32'hba63871d),
	.w6(32'h3a987365),
	.w7(32'hba408386),
	.w8(32'hba8ad552),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891aeb),
	.w1(32'hb9eb22a7),
	.w2(32'h3ab732e8),
	.w3(32'hbaf062f4),
	.w4(32'h394c47e9),
	.w5(32'h3aa353a9),
	.w6(32'hbaa7973b),
	.w7(32'hb9f6fa53),
	.w8(32'hb9657d72),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1122a2),
	.w1(32'hb98f7154),
	.w2(32'h3a9d6081),
	.w3(32'h3a5ae970),
	.w4(32'hba8080f9),
	.w5(32'h3aa9cbe1),
	.w6(32'hb8199630),
	.w7(32'hbab2773f),
	.w8(32'h39d8d975),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae45f71),
	.w1(32'hbabc44e0),
	.w2(32'hba966862),
	.w3(32'h3a56afb9),
	.w4(32'hbad3aeb4),
	.w5(32'hba26d2d7),
	.w6(32'h3a9dc68c),
	.w7(32'hba4c4ccc),
	.w8(32'hba6d86b7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcabaa),
	.w1(32'hbaf9f478),
	.w2(32'h3a9c82fc),
	.w3(32'hb76e6ed4),
	.w4(32'hbb0d70d9),
	.w5(32'hba867784),
	.w6(32'h39ca0e05),
	.w7(32'hbb1e2995),
	.w8(32'hba5eb769),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39667d79),
	.w1(32'h381a54c1),
	.w2(32'h3aa1319f),
	.w3(32'hb98125f0),
	.w4(32'h3a806513),
	.w5(32'h3b394c65),
	.w6(32'hbaa545cc),
	.w7(32'h3aa97df1),
	.w8(32'h3b2ea1a4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965d865),
	.w1(32'hb9b38190),
	.w2(32'h396698cb),
	.w3(32'h3a966785),
	.w4(32'hba4e8598),
	.w5(32'h3a2007d0),
	.w6(32'h3a92aa9b),
	.w7(32'hbaa9a9a4),
	.w8(32'hb91977de),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabc3c2),
	.w1(32'hbaa8f946),
	.w2(32'hba466faf),
	.w3(32'h3a7a60e7),
	.w4(32'hba04b77c),
	.w5(32'h3a1d6a1c),
	.w6(32'h3a9f2b10),
	.w7(32'hbaf63fb6),
	.w8(32'hbaa1a6f3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42d36),
	.w1(32'h3af2d2b9),
	.w2(32'h3b84d27d),
	.w3(32'hba925d44),
	.w4(32'h3aca02ec),
	.w5(32'h3ad30440),
	.w6(32'hba8750aa),
	.w7(32'h3a428fb4),
	.w8(32'h3a3733e2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc8bf),
	.w1(32'h38fff1c8),
	.w2(32'h3a1ed237),
	.w3(32'h39f93aa8),
	.w4(32'hb9fea822),
	.w5(32'hbb08ef82),
	.w6(32'hb6b753fc),
	.w7(32'h38cd716f),
	.w8(32'hb919e944),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f07cc),
	.w1(32'hbae96b71),
	.w2(32'hbaaebb8d),
	.w3(32'h39c494ba),
	.w4(32'hbb3d836a),
	.w5(32'hba8c1bd6),
	.w6(32'h395e6b4c),
	.w7(32'hbb023dcb),
	.w8(32'hba831424),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384272c4),
	.w1(32'hb9fcbd78),
	.w2(32'hbaccb8d0),
	.w3(32'hba96b8ea),
	.w4(32'hb9795c37),
	.w5(32'hba948078),
	.w6(32'hb6f56cc2),
	.w7(32'hba10272d),
	.w8(32'hbaec0223),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b310d),
	.w1(32'h3a79895c),
	.w2(32'hb898a80e),
	.w3(32'hbaa577fa),
	.w4(32'h3ae5a3e6),
	.w5(32'hb9a0f13c),
	.w6(32'hba5d1fd1),
	.w7(32'h3a066793),
	.w8(32'h3a764938),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972b29f),
	.w1(32'hba1bad80),
	.w2(32'hba7a9dfe),
	.w3(32'h39964a27),
	.w4(32'hba80530e),
	.w5(32'hba87ffd1),
	.w6(32'h39a5619d),
	.w7(32'hba136b45),
	.w8(32'hbaa95f55),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bf298),
	.w1(32'h39d6416a),
	.w2(32'h3a18c3b4),
	.w3(32'hba7481d4),
	.w4(32'hb906831e),
	.w5(32'h3ae0598e),
	.w6(32'hb879a3b6),
	.w7(32'hb9bc7781),
	.w8(32'h3a03af58),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b299d),
	.w1(32'h3b0982a1),
	.w2(32'h3b2ade1a),
	.w3(32'h3ae250fc),
	.w4(32'h399774a2),
	.w5(32'hbaa7dca3),
	.w6(32'h3af1c932),
	.w7(32'hba249a9c),
	.w8(32'h3a2c32b3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5ee67),
	.w1(32'hb78cdb26),
	.w2(32'h3ae1e5b3),
	.w3(32'h3967bc8d),
	.w4(32'hba00ce0c),
	.w5(32'h3a173b25),
	.w6(32'h3ac2f01f),
	.w7(32'hba58eb4c),
	.w8(32'h3a1eaf49),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57aac4),
	.w1(32'hbacb8dff),
	.w2(32'hbafd0fb5),
	.w3(32'h399edb8d),
	.w4(32'hbb7516e4),
	.w5(32'hbb493f36),
	.w6(32'hb8a41fbc),
	.w7(32'hbb01a505),
	.w8(32'hbb21ef41),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c53006),
	.w1(32'hba227135),
	.w2(32'hbac4aebf),
	.w3(32'hbacef0d7),
	.w4(32'hb9f4b372),
	.w5(32'hb9970917),
	.w6(32'hba90a312),
	.w7(32'hba5a1053),
	.w8(32'hba645ff4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule