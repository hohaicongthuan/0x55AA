module layer_10_featuremap_228(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106f96),
	.w1(32'h3aaed674),
	.w2(32'h3c8427db),
	.w3(32'hbad27507),
	.w4(32'hbb8a0859),
	.w5(32'h3c0b5492),
	.w6(32'h3b71f675),
	.w7(32'h3a5ded67),
	.w8(32'hbbc27efe),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf1d2b),
	.w1(32'hbac16d3c),
	.w2(32'h3cf89996),
	.w3(32'hbb5c823c),
	.w4(32'h39e5f286),
	.w5(32'hbb5bc066),
	.w6(32'hba2d2db5),
	.w7(32'h3cdb82be),
	.w8(32'h3b9945a3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ba2e),
	.w1(32'hba8eee39),
	.w2(32'hbd16bc56),
	.w3(32'h3ca0b4bd),
	.w4(32'h3ba7d0bc),
	.w5(32'hbc3bdace),
	.w6(32'h3d0a33c0),
	.w7(32'h3bfd6dbc),
	.w8(32'hbb5a5ac5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831aad),
	.w1(32'hbc0244ad),
	.w2(32'hbc7d4a15),
	.w3(32'hbc328579),
	.w4(32'hbc01a149),
	.w5(32'h39acd2a1),
	.w6(32'hbb31e020),
	.w7(32'h3c548a47),
	.w8(32'hb9dce5c8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8e405),
	.w1(32'hbc226113),
	.w2(32'h3ad1eda7),
	.w3(32'hbc2cb500),
	.w4(32'h3c1c0e6a),
	.w5(32'h3a841333),
	.w6(32'hbc3dbf30),
	.w7(32'hbba78e69),
	.w8(32'h3b0ef7f3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e1f66),
	.w1(32'hbb563abf),
	.w2(32'hbaa4474c),
	.w3(32'hbc45620a),
	.w4(32'hb997af17),
	.w5(32'h3bf4e538),
	.w6(32'h3b07fdab),
	.w7(32'hbc172cbf),
	.w8(32'hba485f30),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e89b2),
	.w1(32'h3b17e818),
	.w2(32'h3c0e14e1),
	.w3(32'hbc8c2979),
	.w4(32'hba61ea00),
	.w5(32'h3c749f2f),
	.w6(32'h3b94f79b),
	.w7(32'hbc18de9c),
	.w8(32'hbbef6fcb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16e806),
	.w1(32'hbc284acc),
	.w2(32'h3cbae23a),
	.w3(32'hbbdfcdfa),
	.w4(32'hbb8957d3),
	.w5(32'hb93950d3),
	.w6(32'hbc855c8f),
	.w7(32'hbc0b179b),
	.w8(32'h3cc39f32),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c3d0c),
	.w1(32'hbb25f183),
	.w2(32'h3c96b0c5),
	.w3(32'hbc836b08),
	.w4(32'h3b21a442),
	.w5(32'hbc493ad4),
	.w6(32'hbba9954f),
	.w7(32'hbbed117a),
	.w8(32'hba72d1a3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc646215),
	.w1(32'h382c5f36),
	.w2(32'h3c3d64bc),
	.w3(32'h3ca6f3c4),
	.w4(32'hbc643a16),
	.w5(32'hbbe1c4f4),
	.w6(32'hbc45a4d9),
	.w7(32'hbb5f62d2),
	.w8(32'hbc4d0ef1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269f1e),
	.w1(32'h3c4981a6),
	.w2(32'h39c9c8a8),
	.w3(32'hbbf865c3),
	.w4(32'hbbc10b61),
	.w5(32'h3bf7626b),
	.w6(32'hbc14cd46),
	.w7(32'hbc17127d),
	.w8(32'h3b385a9f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f162d),
	.w1(32'h3a8e9c0a),
	.w2(32'hbbd89133),
	.w3(32'hbc9df617),
	.w4(32'h3c5908f0),
	.w5(32'hb7575f22),
	.w6(32'h3b56304d),
	.w7(32'hb78d6dd1),
	.w8(32'h3b9a67c3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1688b6),
	.w1(32'hbc4e8d5b),
	.w2(32'h386d5c62),
	.w3(32'h3b6bb7a7),
	.w4(32'h3a0f2aa7),
	.w5(32'h3cf7bbac),
	.w6(32'h3c67fdaf),
	.w7(32'hbc85ea36),
	.w8(32'h3c36b8b9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92c5e4),
	.w1(32'hbc9ad018),
	.w2(32'hbcfc0ff3),
	.w3(32'hbcbc4ecd),
	.w4(32'hbc1c3b3a),
	.w5(32'h3a5faa7f),
	.w6(32'hba07d2b1),
	.w7(32'hbbf13d65),
	.w8(32'h3b97f53f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b89a4),
	.w1(32'h3ca58b50),
	.w2(32'h394de08e),
	.w3(32'hbbb14565),
	.w4(32'hbbe7a163),
	.w5(32'hba32563d),
	.w6(32'h3bfaa690),
	.w7(32'hbbecc44c),
	.w8(32'h39fc072f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6566d6),
	.w1(32'hbb36ee17),
	.w2(32'h3a1bc0f6),
	.w3(32'hbc93665b),
	.w4(32'h3a17172e),
	.w5(32'hbbf29e1a),
	.w6(32'h3c074863),
	.w7(32'h3b125014),
	.w8(32'h3bdc72f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb171e0e),
	.w1(32'h3c201032),
	.w2(32'hbc0acc8e),
	.w3(32'h3b6e0960),
	.w4(32'hb6b4731d),
	.w5(32'hbc13cd95),
	.w6(32'hb9291e66),
	.w7(32'hbb199a25),
	.w8(32'hbbf652ad),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35e310),
	.w1(32'hbb1f9d15),
	.w2(32'h3b874d2c),
	.w3(32'hbc84024c),
	.w4(32'hbba507fd),
	.w5(32'h39adb085),
	.w6(32'h3c00f5ac),
	.w7(32'hbb3032cb),
	.w8(32'hbc170c71),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c644f44),
	.w1(32'h3a239193),
	.w2(32'hbb9619cf),
	.w3(32'h3b56f53e),
	.w4(32'h3adb2820),
	.w5(32'hbbd09067),
	.w6(32'hbbbdd2f2),
	.w7(32'hbc4b30ec),
	.w8(32'h3b0c93aa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0315d),
	.w1(32'hbc43f8c8),
	.w2(32'hbba79ac7),
	.w3(32'hbbea6470),
	.w4(32'hbac0bcec),
	.w5(32'h3b32d1ca),
	.w6(32'hbc6c0bc5),
	.w7(32'hbbd0fbb1),
	.w8(32'hbb8a1f90),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c7726),
	.w1(32'hbaffcde4),
	.w2(32'hbc2ed0f4),
	.w3(32'h3b8a37f0),
	.w4(32'hbb8da5f1),
	.w5(32'hbbe0bd68),
	.w6(32'hbb8e9273),
	.w7(32'h3b0f79d1),
	.w8(32'hbbe6686e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e27f7),
	.w1(32'hbd006c4b),
	.w2(32'hba14ea8f),
	.w3(32'hbb1b6cb4),
	.w4(32'h3bb0e22e),
	.w5(32'h3ab4dc22),
	.w6(32'hbb3dd4b9),
	.w7(32'hb99ae385),
	.w8(32'hbbcf1525),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745fe3),
	.w1(32'hb8f35d3a),
	.w2(32'hbbdd5c9f),
	.w3(32'hbaa6ae59),
	.w4(32'h3a8704c6),
	.w5(32'hbc1e54b7),
	.w6(32'h3acaa222),
	.w7(32'h3b410fe6),
	.w8(32'hbc3c212a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b930d98),
	.w1(32'hbc53ab5a),
	.w2(32'h3c8a8b88),
	.w3(32'h3c197e7f),
	.w4(32'h3aa91db8),
	.w5(32'hbc19e6a3),
	.w6(32'h3c9f3d76),
	.w7(32'hb9a083d7),
	.w8(32'h38044ce8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab52f),
	.w1(32'h3bc38f31),
	.w2(32'h3c8fcd93),
	.w3(32'h3b9b1d1d),
	.w4(32'hbc2906c0),
	.w5(32'h3c7837d0),
	.w6(32'hbaad0960),
	.w7(32'h3b7d3556),
	.w8(32'hba22f3d3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb456f48),
	.w1(32'h3b30035f),
	.w2(32'h3c16da45),
	.w3(32'h3d102158),
	.w4(32'h3bf6988b),
	.w5(32'hbc939b89),
	.w6(32'hbb9f9645),
	.w7(32'h3b979735),
	.w8(32'h395cb5cf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf13ce0),
	.w1(32'h3cb5c1be),
	.w2(32'h3b091409),
	.w3(32'h3be0ff66),
	.w4(32'hb9daf0c1),
	.w5(32'hbb09124d),
	.w6(32'hbc578129),
	.w7(32'hbc259dd9),
	.w8(32'hbc477a14),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb397b34),
	.w1(32'hbc271ca2),
	.w2(32'h3aa67c36),
	.w3(32'h3a903af9),
	.w4(32'hbbb7a55f),
	.w5(32'hbb5344a0),
	.w6(32'h3aa2563d),
	.w7(32'hbc4bf52c),
	.w8(32'hbbf93e90),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b627e3f),
	.w1(32'hbba7417d),
	.w2(32'h3c36f6aa),
	.w3(32'h3c239190),
	.w4(32'hbb67a89d),
	.w5(32'hbc037d3d),
	.w6(32'h3c2da2bd),
	.w7(32'hbb0ad0df),
	.w8(32'hbb90774f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e6234),
	.w1(32'h3cc15a44),
	.w2(32'h3c9c6fe4),
	.w3(32'hbb68480e),
	.w4(32'h3b175e36),
	.w5(32'hbca973cb),
	.w6(32'h3c82a225),
	.w7(32'hbac69e97),
	.w8(32'h3b8df3ca),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a30e9),
	.w1(32'hbc41d7ac),
	.w2(32'hbbb8b07e),
	.w3(32'hbb0ddff7),
	.w4(32'hbb7d8048),
	.w5(32'hba4344d3),
	.w6(32'h3bf2479d),
	.w7(32'h3b7dda4d),
	.w8(32'h3c64f0f9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bad26),
	.w1(32'hbbc863b1),
	.w2(32'hbbc6ae45),
	.w3(32'hbafbf3c4),
	.w4(32'h3a2ac65b),
	.w5(32'hbb972fa7),
	.w6(32'hbb258fb1),
	.w7(32'hbc2fb660),
	.w8(32'hba23548b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db5bb9),
	.w1(32'hbc7eb605),
	.w2(32'h3abd7ee0),
	.w3(32'hbc79faac),
	.w4(32'hbc2b459a),
	.w5(32'h3c1b6064),
	.w6(32'h3c836900),
	.w7(32'hbc1bb4b0),
	.w8(32'hbba9251f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c0f9e),
	.w1(32'hbccae1b9),
	.w2(32'h3c5a8835),
	.w3(32'hbc36114d),
	.w4(32'h3c68f251),
	.w5(32'h3caf60a4),
	.w6(32'h3b20665e),
	.w7(32'hbb901fd9),
	.w8(32'h3978e98a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc965fa),
	.w1(32'hbc2df0c5),
	.w2(32'hbc97203a),
	.w3(32'hb9db5bae),
	.w4(32'hbb961d03),
	.w5(32'hba4328d2),
	.w6(32'h3b22680e),
	.w7(32'hbcbb0e31),
	.w8(32'hbb4d1a4f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02b1db),
	.w1(32'h3b5a5769),
	.w2(32'hbca2b89a),
	.w3(32'hbb6f0708),
	.w4(32'hbaef5fc6),
	.w5(32'h3b85f1b6),
	.w6(32'h3c2feb74),
	.w7(32'hb9bacea6),
	.w8(32'h3a283c4c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b381e58),
	.w1(32'hbca21914),
	.w2(32'hbb91a7a9),
	.w3(32'h3c25e86e),
	.w4(32'h3bd0cddb),
	.w5(32'hb98bd3d8),
	.w6(32'hbbc72390),
	.w7(32'h3b97ef2e),
	.w8(32'hbc0923ab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b10c),
	.w1(32'h3a206201),
	.w2(32'h3b8cbea0),
	.w3(32'hbbf82b4f),
	.w4(32'hbc9d3303),
	.w5(32'hb8ea9412),
	.w6(32'hbc07ecf8),
	.w7(32'hbc8b0517),
	.w8(32'h3b329c4d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30e915),
	.w1(32'h3b0491ed),
	.w2(32'h3bd1e6b1),
	.w3(32'h3c7be440),
	.w4(32'hbc091dcc),
	.w5(32'hbb2e6caa),
	.w6(32'hbc358679),
	.w7(32'h3a57b84f),
	.w8(32'hbbd8e7c1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ce47),
	.w1(32'h3b796053),
	.w2(32'hba5f2689),
	.w3(32'h39949d17),
	.w4(32'hb8a8802a),
	.w5(32'h3c110b30),
	.w6(32'h3b94a420),
	.w7(32'h3c2862ba),
	.w8(32'hbc85e23e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35164430),
	.w1(32'h3b101078),
	.w2(32'hba48fe79),
	.w3(32'hbc2742a6),
	.w4(32'hbc128dac),
	.w5(32'h3b48ccb8),
	.w6(32'h3992ea08),
	.w7(32'hbaad2342),
	.w8(32'hbbdcbffa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c4e86),
	.w1(32'hbb4fcc1a),
	.w2(32'h3c4cf063),
	.w3(32'h3c092fd6),
	.w4(32'hb8038ba8),
	.w5(32'hbc1141f2),
	.w6(32'hbb355f07),
	.w7(32'hbc8ede6e),
	.w8(32'hb9a6fa9b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdab4bf),
	.w1(32'hbc044dbf),
	.w2(32'h3b676e07),
	.w3(32'hbc6028f4),
	.w4(32'h3b330426),
	.w5(32'hbb84f1b7),
	.w6(32'hbc67915c),
	.w7(32'hbc01eb00),
	.w8(32'h3c3e41e8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5205b5),
	.w1(32'h3b4efbc4),
	.w2(32'h3c15adf7),
	.w3(32'h3b9eef4a),
	.w4(32'h3bab6698),
	.w5(32'hbab266e9),
	.w6(32'hbc892533),
	.w7(32'h3c56b22d),
	.w8(32'hba4a0024),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee0d84),
	.w1(32'hbb78d2db),
	.w2(32'hba55c9fa),
	.w3(32'hbc014f5b),
	.w4(32'h3ba90634),
	.w5(32'hbb7b2d08),
	.w6(32'h3b8071e4),
	.w7(32'h3ab193e3),
	.w8(32'h364d908c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a498f),
	.w1(32'hbbc6b7c9),
	.w2(32'h3cb1cb4d),
	.w3(32'hbbafd242),
	.w4(32'hbc1d18f6),
	.w5(32'h3c826534),
	.w6(32'hbca612a9),
	.w7(32'h3b91eba1),
	.w8(32'hbc65b5c5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b281db3),
	.w1(32'h3c79ad1a),
	.w2(32'hbb8d35cd),
	.w3(32'hbc977065),
	.w4(32'h3c22a5b7),
	.w5(32'hbb8bc474),
	.w6(32'h3986a69b),
	.w7(32'hbabf1356),
	.w8(32'hbb9dc271),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc065994),
	.w1(32'h3c9560b2),
	.w2(32'h3c2c54a5),
	.w3(32'hbab9bbb8),
	.w4(32'hbbe44a55),
	.w5(32'hb86c9a2b),
	.w6(32'hbc93bab2),
	.w7(32'hba4c111c),
	.w8(32'h3c3fda2d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8593d),
	.w1(32'hbc26b2cf),
	.w2(32'h3c749d08),
	.w3(32'hbc712f38),
	.w4(32'h3c842713),
	.w5(32'hbba318da),
	.w6(32'h3a86fd3b),
	.w7(32'hbc1c6cc5),
	.w8(32'hbc63c69b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f5a09),
	.w1(32'h3ccf2117),
	.w2(32'hbb66bba1),
	.w3(32'h3c42a532),
	.w4(32'hbb9d2bf2),
	.w5(32'hbb73ea1f),
	.w6(32'hba9269d4),
	.w7(32'h3c21a945),
	.w8(32'h3bb598fd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ccf7e2),
	.w1(32'hbb9afbba),
	.w2(32'h3bb1814a),
	.w3(32'h3ab176e8),
	.w4(32'h39ff0258),
	.w5(32'h36da6a6b),
	.w6(32'hbbb55c22),
	.w7(32'hbc0b3aa1),
	.w8(32'hba2096e8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd9f86),
	.w1(32'hbc6a66c3),
	.w2(32'h3acc5e97),
	.w3(32'hbc150792),
	.w4(32'hbc0fe032),
	.w5(32'h3ac27341),
	.w6(32'h3bce42cd),
	.w7(32'hbb8788e2),
	.w8(32'hbb2356b8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b7e5d),
	.w1(32'hbba59229),
	.w2(32'hbaeeff45),
	.w3(32'hbc7a34f4),
	.w4(32'h3bf9ff9d),
	.w5(32'hbc924ee6),
	.w6(32'h39f5940c),
	.w7(32'hbb9cbdd5),
	.w8(32'hbcb5f514),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb894be),
	.w1(32'hbacf84f7),
	.w2(32'hbb80e73b),
	.w3(32'hbb00fe85),
	.w4(32'hbb933acc),
	.w5(32'hbc7f59ab),
	.w6(32'h3cac766b),
	.w7(32'hbc71cd7d),
	.w8(32'hbcbb997c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be715),
	.w1(32'h3afc8481),
	.w2(32'hbac3b6af),
	.w3(32'h3cfcd532),
	.w4(32'h3ad34517),
	.w5(32'h3ac8dc21),
	.w6(32'h3b117d5c),
	.w7(32'hbaa211e6),
	.w8(32'hbbe047df),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c06a4),
	.w1(32'h3b6ccda5),
	.w2(32'hbb897832),
	.w3(32'h3c7be14a),
	.w4(32'h3c17e545),
	.w5(32'hbbd41c04),
	.w6(32'hbad8b5a2),
	.w7(32'hba36be40),
	.w8(32'h3b94695b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8daaaa),
	.w1(32'h3b03d000),
	.w2(32'h3b987294),
	.w3(32'hbb800e11),
	.w4(32'hbc1e35be),
	.w5(32'hbaa050ec),
	.w6(32'hbbf1b1e7),
	.w7(32'hb8c6d6cf),
	.w8(32'hbc05cc73),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf96ef9),
	.w1(32'h3bb84cf1),
	.w2(32'hbd10cdec),
	.w3(32'hbc752ae4),
	.w4(32'h3b86225b),
	.w5(32'hbb86cdd1),
	.w6(32'h3b503227),
	.w7(32'hb9a2e041),
	.w8(32'h3b39c2ce),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b88cb),
	.w1(32'hbc2b67cb),
	.w2(32'hbbe84f7d),
	.w3(32'h3990e57e),
	.w4(32'h3be72fc8),
	.w5(32'h3b7c236e),
	.w6(32'h3c33e73e),
	.w7(32'hbbc8f446),
	.w8(32'h3b88bdcc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d7385),
	.w1(32'hba8b581f),
	.w2(32'h3be7c69c),
	.w3(32'h3c2d0b1b),
	.w4(32'h385f5af5),
	.w5(32'h3b4a0b55),
	.w6(32'hbb9a3fc2),
	.w7(32'h3c66c0ae),
	.w8(32'h3c8f2b94),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19aa32),
	.w1(32'h3afe4b97),
	.w2(32'hbb8e5dd1),
	.w3(32'h3c00afb2),
	.w4(32'hbbe9e060),
	.w5(32'hbb9f324e),
	.w6(32'h3b8067dc),
	.w7(32'h3c222151),
	.w8(32'h3b6aad4e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13dc54),
	.w1(32'hba0d11a6),
	.w2(32'hbad76729),
	.w3(32'hbb09a7e5),
	.w4(32'hbbd1a0f1),
	.w5(32'h3b283197),
	.w6(32'h3c5582f1),
	.w7(32'h3af29fe7),
	.w8(32'h3be10f64),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205dec),
	.w1(32'hba7cc842),
	.w2(32'hbd0c80c6),
	.w3(32'hbbe4919c),
	.w4(32'h3b838e92),
	.w5(32'h3c02c3bf),
	.w6(32'hb89b69c8),
	.w7(32'hbbf0e2bf),
	.w8(32'h3b811a63),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9c2c9),
	.w1(32'hbc33c3fc),
	.w2(32'h3ae6970b),
	.w3(32'h3c368496),
	.w4(32'hbb7e7654),
	.w5(32'hbba6b3f7),
	.w6(32'h3bdd4ebd),
	.w7(32'hbb04d40f),
	.w8(32'hb9aac15f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a7791),
	.w1(32'h3a558363),
	.w2(32'hba6c7be4),
	.w3(32'hbbafe799),
	.w4(32'h391283fd),
	.w5(32'h3c219acb),
	.w6(32'h3bdb0a19),
	.w7(32'h3ace25f7),
	.w8(32'hbbea6890),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2414a8),
	.w1(32'h39955116),
	.w2(32'h3c0b9996),
	.w3(32'h3c9124c6),
	.w4(32'h3bd46a0e),
	.w5(32'hba611517),
	.w6(32'h3bd38bde),
	.w7(32'h3c5c713f),
	.w8(32'h3b8786b0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd4ac7),
	.w1(32'h3c004570),
	.w2(32'h38dff6b7),
	.w3(32'h3c4cea6a),
	.w4(32'h3b8c019b),
	.w5(32'h3c70224f),
	.w6(32'h3875a313),
	.w7(32'hbbe1eb06),
	.w8(32'h3ba330f5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b130c66),
	.w1(32'h3cb1141e),
	.w2(32'h3b026fc7),
	.w3(32'h3a2bebe2),
	.w4(32'h3a18514d),
	.w5(32'h3cb8d165),
	.w6(32'h3b916a67),
	.w7(32'h3b6dcd3a),
	.w8(32'h3b27849d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdada58),
	.w1(32'h3b86af78),
	.w2(32'h396ba054),
	.w3(32'hbb845ab2),
	.w4(32'hb49795a7),
	.w5(32'hba844ad0),
	.w6(32'h3ae92085),
	.w7(32'h3b13f642),
	.w8(32'h3cb91185),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefda3e),
	.w1(32'hbb8f6825),
	.w2(32'hbc809698),
	.w3(32'hbc81e4f9),
	.w4(32'hbac00199),
	.w5(32'hba6994e0),
	.w6(32'h3aa51f7e),
	.w7(32'h3a883ada),
	.w8(32'hbaecb5fe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06f62),
	.w1(32'h3bfa0700),
	.w2(32'h3b88fc7b),
	.w3(32'hbb4bda54),
	.w4(32'h3b3a7870),
	.w5(32'hb956dbc9),
	.w6(32'h3b05d5a0),
	.w7(32'h3c98f593),
	.w8(32'h3bd2d37b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e226b),
	.w1(32'hbc50898f),
	.w2(32'hbba79f0c),
	.w3(32'h3cc7c602),
	.w4(32'h3bb412a7),
	.w5(32'hbaf424bf),
	.w6(32'hbbdc43de),
	.w7(32'hbc024eb0),
	.w8(32'hbc03e3a8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff9846),
	.w1(32'hbbc6bc8b),
	.w2(32'hb9e77108),
	.w3(32'hbac972d2),
	.w4(32'h3c031061),
	.w5(32'hbbe3ba99),
	.w6(32'hba919ac3),
	.w7(32'hbc3b683a),
	.w8(32'hbbd36c1b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66df19),
	.w1(32'h35a45af3),
	.w2(32'h3c91332b),
	.w3(32'hbbc7c795),
	.w4(32'hb8584602),
	.w5(32'h3b27210b),
	.w6(32'h3b6d48f8),
	.w7(32'hbb0c22bf),
	.w8(32'h3bac21c0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b60b8),
	.w1(32'hbae57fa3),
	.w2(32'hb97fd64c),
	.w3(32'hbc1058cc),
	.w4(32'hba243880),
	.w5(32'hbb9339d8),
	.w6(32'h3bab8957),
	.w7(32'hbaab5d28),
	.w8(32'h3bd57832),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8440b),
	.w1(32'h3c352a66),
	.w2(32'h396060bf),
	.w3(32'h3b7d7b76),
	.w4(32'h3be87c65),
	.w5(32'hbbafba20),
	.w6(32'hbb1cf2f2),
	.w7(32'h392d1bd6),
	.w8(32'h3b0eb1e5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65303c),
	.w1(32'hbc30ebee),
	.w2(32'hbc2db81f),
	.w3(32'h3bf4ffdf),
	.w4(32'h3a87ae59),
	.w5(32'h3a9afe45),
	.w6(32'h3c3143b2),
	.w7(32'h3b1a874a),
	.w8(32'h3c012749),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eef00),
	.w1(32'hbad3ea3e),
	.w2(32'h3ce8e277),
	.w3(32'h3c23022a),
	.w4(32'h3bad70dd),
	.w5(32'hbb223303),
	.w6(32'hbb846dd1),
	.w7(32'hbc6f6631),
	.w8(32'h3cad7266),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba824fed),
	.w1(32'h3a34d9d9),
	.w2(32'h3a5dc657),
	.w3(32'hbc4c7b61),
	.w4(32'hb94d8e3e),
	.w5(32'hbc15876d),
	.w6(32'h3b960607),
	.w7(32'h3b660227),
	.w8(32'hbb94590b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86aa6f),
	.w1(32'h3c0e1da1),
	.w2(32'hbc99ace2),
	.w3(32'hba50a6fd),
	.w4(32'hbc190147),
	.w5(32'h3c0cf26d),
	.w6(32'h3a6642c5),
	.w7(32'h3bd73383),
	.w8(32'hb97723fc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909d1a6),
	.w1(32'h3bbfd825),
	.w2(32'h3b9a408f),
	.w3(32'hbaad6732),
	.w4(32'h3beca99b),
	.w5(32'h3ae848a3),
	.w6(32'hbb8527d5),
	.w7(32'h3c9cb41d),
	.w8(32'hbae1523b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77331),
	.w1(32'h3a13fb89),
	.w2(32'hbb2279a2),
	.w3(32'h3b592d96),
	.w4(32'hbb0987af),
	.w5(32'h3be782c1),
	.w6(32'hbb055938),
	.w7(32'hba94332d),
	.w8(32'h3d01356e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb586f90),
	.w1(32'h3ccde08d),
	.w2(32'h3b3cff1f),
	.w3(32'hb907d6e9),
	.w4(32'h3aa7cfd1),
	.w5(32'hbbaacc25),
	.w6(32'hbabb470f),
	.w7(32'hbb2cf9af),
	.w8(32'hbbd2e66f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2cba),
	.w1(32'h3bb8951d),
	.w2(32'hbb17de7d),
	.w3(32'hbb14fa76),
	.w4(32'hb9678df6),
	.w5(32'hbbacf1c6),
	.w6(32'hbb2c70b3),
	.w7(32'hbb6135c3),
	.w8(32'hbb559a0f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42f04),
	.w1(32'hba85dd6e),
	.w2(32'hbc85c3c5),
	.w3(32'h3b9f0862),
	.w4(32'hbd025d57),
	.w5(32'h3aa6718c),
	.w6(32'hbc01c3d0),
	.w7(32'hbb65ac45),
	.w8(32'hbbd8c4d4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5067dd),
	.w1(32'h3b255be9),
	.w2(32'hbb91c43a),
	.w3(32'h3a6eea33),
	.w4(32'hbb906468),
	.w5(32'hbb9d037b),
	.w6(32'hba749df0),
	.w7(32'h3bb35dfc),
	.w8(32'h398086e2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7bb6d),
	.w1(32'h3ca691d8),
	.w2(32'h3c0ca31c),
	.w3(32'h3c55ecb6),
	.w4(32'h3b6a8ab8),
	.w5(32'hba799874),
	.w6(32'hbc26c5a9),
	.w7(32'hbb46bb86),
	.w8(32'hbc00e476),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4164a4),
	.w1(32'h3bddce42),
	.w2(32'hbb942b52),
	.w3(32'hbb82b34d),
	.w4(32'h3aeb64f4),
	.w5(32'hbc6d2d6f),
	.w6(32'hbb29e857),
	.w7(32'hbb5d9ed9),
	.w8(32'hba9dc674),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b252c),
	.w1(32'hba4390d0),
	.w2(32'hbbfd63f7),
	.w3(32'h3b4fefee),
	.w4(32'hbb6f3d09),
	.w5(32'h3c7e0c99),
	.w6(32'hbbfccb63),
	.w7(32'hbb578f02),
	.w8(32'hbbc2b1bb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda5811),
	.w1(32'hbab47752),
	.w2(32'h3b3d62dc),
	.w3(32'hbbb8861c),
	.w4(32'hbbab1163),
	.w5(32'h39d1fdd5),
	.w6(32'hb9264360),
	.w7(32'hbaceeae9),
	.w8(32'h3a68d0cd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ec5a0),
	.w1(32'h3ac80e7e),
	.w2(32'hbc96e205),
	.w3(32'hba3e08d3),
	.w4(32'h3bca4b3a),
	.w5(32'hba491e84),
	.w6(32'hbc1382d2),
	.w7(32'hbb1adfb9),
	.w8(32'h3b8999c1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a4dd3),
	.w1(32'hbbadf685),
	.w2(32'h3bb112fa),
	.w3(32'hbb87a1ad),
	.w4(32'hbb8e5b30),
	.w5(32'hbc75d5ea),
	.w6(32'h3b89e142),
	.w7(32'h3bac943c),
	.w8(32'hbaca29f9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69e5a9),
	.w1(32'hba3f578f),
	.w2(32'hbb3254a6),
	.w3(32'h3ce30748),
	.w4(32'h3b508783),
	.w5(32'h3a2f53a9),
	.w6(32'hba16eb49),
	.w7(32'hbc5da4f8),
	.w8(32'hbb9e3d58),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898416),
	.w1(32'hbcbc14b5),
	.w2(32'h3c159786),
	.w3(32'h3affe878),
	.w4(32'h39c48d86),
	.w5(32'hbb9aa02d),
	.w6(32'hbb904eb2),
	.w7(32'hbbe5017f),
	.w8(32'hba945fae),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa09ef),
	.w1(32'hbbddcc49),
	.w2(32'h37eadbeb),
	.w3(32'hbc28cef9),
	.w4(32'hbaa21f8d),
	.w5(32'h39a7af7d),
	.w6(32'h3a22d369),
	.w7(32'h390d85a7),
	.w8(32'hbbb5e693),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397775d3),
	.w1(32'hbc09bf62),
	.w2(32'hbba0d8c5),
	.w3(32'hbb7df2c8),
	.w4(32'hbb771c4b),
	.w5(32'hbc35ddf1),
	.w6(32'hbb79a58f),
	.w7(32'hba642798),
	.w8(32'hbac2c748),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bdae6),
	.w1(32'hb9ad9482),
	.w2(32'h37ad9376),
	.w3(32'hbd894214),
	.w4(32'h37903bc2),
	.w5(32'hbc1edd34),
	.w6(32'hbbbe6935),
	.w7(32'hbbba32db),
	.w8(32'hb276bf70),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc304b04),
	.w1(32'hbc560295),
	.w2(32'hbbe1e956),
	.w3(32'h3897fca4),
	.w4(32'h39063abb),
	.w5(32'hbc1ac6b9),
	.w6(32'hbbda0925),
	.w7(32'h3c37e7c2),
	.w8(32'hbbb92e29),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994cf39),
	.w1(32'hbcbc9b46),
	.w2(32'hba67fa24),
	.w3(32'h3bc4a755),
	.w4(32'hbbe270b1),
	.w5(32'h3c78b251),
	.w6(32'hbb26d99b),
	.w7(32'hbc18ec50),
	.w8(32'hbc4bbff3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f1207),
	.w1(32'hbc20cfb8),
	.w2(32'h3bde8196),
	.w3(32'h3aa03fb1),
	.w4(32'hbb0b30f7),
	.w5(32'hbbe12e2b),
	.w6(32'h3a803fbb),
	.w7(32'hbc038ca7),
	.w8(32'hbb0089cd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8d95),
	.w1(32'hbc0e7d66),
	.w2(32'h3a970f68),
	.w3(32'hbaf277a1),
	.w4(32'hbb814f99),
	.w5(32'hbbd61f63),
	.w6(32'h3a6309de),
	.w7(32'hbbb6d09f),
	.w8(32'hbc247e1e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f6ba),
	.w1(32'hbb97cf98),
	.w2(32'h3c35b56e),
	.w3(32'hbb3a42b8),
	.w4(32'hbbb9e9a0),
	.w5(32'h35ea9c84),
	.w6(32'h3d048c6c),
	.w7(32'h3b9bcf64),
	.w8(32'hbbc91890),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153d82),
	.w1(32'hbbbf6b3a),
	.w2(32'hbce6e793),
	.w3(32'hbc5e2c8b),
	.w4(32'h3a998036),
	.w5(32'h3b055aa8),
	.w6(32'hb92d88e8),
	.w7(32'hbc1d75c0),
	.w8(32'h3bf6520a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab1615),
	.w1(32'h3b87a856),
	.w2(32'hbb872b86),
	.w3(32'h3a2a031c),
	.w4(32'hbb7734f9),
	.w5(32'h3aba17e0),
	.w6(32'hbb9c04ec),
	.w7(32'hbb926417),
	.w8(32'hbbed7c99),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04ec5),
	.w1(32'hbd1c7119),
	.w2(32'h3a246fc4),
	.w3(32'h3ad2f23f),
	.w4(32'hbbf40fee),
	.w5(32'hbc50c63c),
	.w6(32'h39d08e28),
	.w7(32'hbc19ffa2),
	.w8(32'hbba156bc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5466ba),
	.w1(32'hbb49fa2b),
	.w2(32'hbb9317c7),
	.w3(32'h3c03e9ef),
	.w4(32'hbbc8d824),
	.w5(32'hbaa52fd7),
	.w6(32'hbbec6ed0),
	.w7(32'hbb36d1b2),
	.w8(32'h3a190581),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0579d4),
	.w1(32'h3962b250),
	.w2(32'h3b6ecad0),
	.w3(32'hbb8f7a2a),
	.w4(32'hbb0ff813),
	.w5(32'hbb8cc558),
	.w6(32'hbba6b76d),
	.w7(32'hbc848052),
	.w8(32'h380e0385),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21824d),
	.w1(32'hbba415fc),
	.w2(32'hb8b03913),
	.w3(32'h3ab9fe40),
	.w4(32'hb98be944),
	.w5(32'h3b2eac23),
	.w6(32'h39681fff),
	.w7(32'h39cf8c75),
	.w8(32'h39b2b0e5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d92f132),
	.w1(32'h3c2f3473),
	.w2(32'h3ba99e96),
	.w3(32'hbc789e14),
	.w4(32'hbb29637d),
	.w5(32'hbaa590e1),
	.w6(32'hbcab8d04),
	.w7(32'h3a606537),
	.w8(32'h3cc5cc65),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148d95),
	.w1(32'hbb7e1dab),
	.w2(32'hbbf84e7b),
	.w3(32'hbc0e77c8),
	.w4(32'hbb605dae),
	.w5(32'hbce77257),
	.w6(32'hba824c47),
	.w7(32'h3a3ec440),
	.w8(32'h3bc530ee),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc44691),
	.w1(32'h3c063d42),
	.w2(32'hbbbec63d),
	.w3(32'hbb20a7e4),
	.w4(32'hbb8f4203),
	.w5(32'hbc1fe606),
	.w6(32'hbc6fb9d2),
	.w7(32'hbb8e3dd6),
	.w8(32'h3acf5dbc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c5ed4),
	.w1(32'h3b37393d),
	.w2(32'hba8e96f9),
	.w3(32'hba923751),
	.w4(32'hbc1c2b9a),
	.w5(32'hbba1d9de),
	.w6(32'hbba6bc3f),
	.w7(32'h3a9bbd37),
	.w8(32'hbb8c685e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6810ef),
	.w1(32'h3ac55dfa),
	.w2(32'hbbc3bcdd),
	.w3(32'h3af5645f),
	.w4(32'hba9ec0dc),
	.w5(32'hbb6bde37),
	.w6(32'h399e03ae),
	.w7(32'hbc0f09e5),
	.w8(32'h3c1dcb8a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f08f8),
	.w1(32'hbbd73a2c),
	.w2(32'hbab27abd),
	.w3(32'h3b74d588),
	.w4(32'h39271d90),
	.w5(32'hbb63be3b),
	.w6(32'h39dd4ef7),
	.w7(32'hbc12623f),
	.w8(32'hbb2f8b61),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaff16),
	.w1(32'hba04eb25),
	.w2(32'hbbc87fec),
	.w3(32'hbbad20e2),
	.w4(32'hbb88cb73),
	.w5(32'hbc3e15df),
	.w6(32'h3b8c0793),
	.w7(32'hbc8989f9),
	.w8(32'hbc3426a5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c311217),
	.w1(32'hbbda49a2),
	.w2(32'hbb9a2f65),
	.w3(32'h3b2153f8),
	.w4(32'hbbe9489f),
	.w5(32'h3b2d04c0),
	.w6(32'hbbd0e1c6),
	.w7(32'h3b4a9bb7),
	.w8(32'h3b17e560),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc36b),
	.w1(32'h3b20175e),
	.w2(32'h3b0ff2b8),
	.w3(32'hba9dd3a8),
	.w4(32'h3ca00800),
	.w5(32'h3c3d0be2),
	.w6(32'h3c97632f),
	.w7(32'hbba9872f),
	.w8(32'h3a5147c3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14f703),
	.w1(32'hbc0e7bfa),
	.w2(32'h3ba312bd),
	.w3(32'hbc008cb5),
	.w4(32'hbbaeb373),
	.w5(32'hb9cd6907),
	.w6(32'hbb95ded0),
	.w7(32'h3bd5829f),
	.w8(32'h3c8dcd6e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd713bc),
	.w1(32'hbc18839d),
	.w2(32'hbc688de6),
	.w3(32'h3cdf2ecc),
	.w4(32'h3b2c3a53),
	.w5(32'h3bf7de50),
	.w6(32'hbb23cb60),
	.w7(32'hbb1a54e7),
	.w8(32'hba557555),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b4a44),
	.w1(32'h3b5db8bb),
	.w2(32'hba992277),
	.w3(32'hbc924b27),
	.w4(32'h3bb1d0bc),
	.w5(32'hba41672f),
	.w6(32'h3b66345e),
	.w7(32'hbca811e6),
	.w8(32'hbc891c8f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122dcc),
	.w1(32'h39c529bf),
	.w2(32'hbb99971e),
	.w3(32'hbbd06496),
	.w4(32'hbc422e99),
	.w5(32'hba183ea2),
	.w6(32'h3c9ef45c),
	.w7(32'hba9c08cf),
	.w8(32'h3c4e3a00),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba001e3),
	.w1(32'hbc2beb55),
	.w2(32'hbc2c84d1),
	.w3(32'h3bb34d17),
	.w4(32'hba61d596),
	.w5(32'h39111f9e),
	.w6(32'hbbbded61),
	.w7(32'hbb679cca),
	.w8(32'h3c358940),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d7d90),
	.w1(32'hbbbda4e2),
	.w2(32'h3a3cbd1f),
	.w3(32'hbb47308f),
	.w4(32'h39bcd9e2),
	.w5(32'hbc513062),
	.w6(32'h3aefab2b),
	.w7(32'hbb48572b),
	.w8(32'hbbe7a382),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d97c),
	.w1(32'h3c428c72),
	.w2(32'h3cc56b09),
	.w3(32'h396211a8),
	.w4(32'h3cc54793),
	.w5(32'h3b481d30),
	.w6(32'h3aae07aa),
	.w7(32'h3b889d7a),
	.w8(32'h3c67be9e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb685c54),
	.w1(32'h3bd5fb6b),
	.w2(32'hb9c30083),
	.w3(32'h3b3d7611),
	.w4(32'h3ad1db83),
	.w5(32'h3a843c5d),
	.w6(32'h3b001787),
	.w7(32'h3a9a1b6f),
	.w8(32'h3ab270c5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81cdd3),
	.w1(32'hb509834d),
	.w2(32'hba89af35),
	.w3(32'hbc123629),
	.w4(32'hbca59503),
	.w5(32'hbc9dafc5),
	.w6(32'hbaeb2db7),
	.w7(32'hbaec96f6),
	.w8(32'hbc018795),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8440a6),
	.w1(32'h3b963fcf),
	.w2(32'h3c325f6f),
	.w3(32'h3b077ae5),
	.w4(32'hbb4ec5d9),
	.w5(32'hbabe7535),
	.w6(32'hbb91304e),
	.w7(32'h3c783bfa),
	.w8(32'hbb12b970),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa9604),
	.w1(32'h3b036c3f),
	.w2(32'h3ca170ae),
	.w3(32'hbcc324ed),
	.w4(32'hbcd211c7),
	.w5(32'hbbbcf43e),
	.w6(32'h3c1ea32b),
	.w7(32'h3beb04cc),
	.w8(32'hb985201e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9aa46f),
	.w1(32'hbb93dbbc),
	.w2(32'h3ad8cf28),
	.w3(32'hbbad513d),
	.w4(32'hbbe49340),
	.w5(32'h3abd7c04),
	.w6(32'hbbba7c84),
	.w7(32'hbb7a578b),
	.w8(32'hbbbfa878),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd27d30),
	.w1(32'h3b297070),
	.w2(32'h3b3c93b2),
	.w3(32'hbb19826e),
	.w4(32'h3c1c5be7),
	.w5(32'hbb91db13),
	.w6(32'hbb9223ce),
	.w7(32'hbc5b5ae4),
	.w8(32'hbc167571),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc4d22),
	.w1(32'hbc1a74ba),
	.w2(32'hbacb81f8),
	.w3(32'h3ca5934a),
	.w4(32'hba695353),
	.w5(32'h3bf98a6c),
	.w6(32'hb52a2ee2),
	.w7(32'h3b15dcfb),
	.w8(32'hbb01de03),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fad5a),
	.w1(32'hbcc39ced),
	.w2(32'hbb9919a3),
	.w3(32'hbca0b4b0),
	.w4(32'h3b4b4370),
	.w5(32'h3bc86815),
	.w6(32'hba53773e),
	.w7(32'h389cd16a),
	.w8(32'hbbfed4a7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf384e),
	.w1(32'h3c8309ab),
	.w2(32'hbb022106),
	.w3(32'h3c7bde1b),
	.w4(32'h3b1c72c7),
	.w5(32'hbbb8ec3d),
	.w6(32'hb8b9c1ec),
	.w7(32'hbc267007),
	.w8(32'h3b9e91cf),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5ec9f),
	.w1(32'h3bc2845a),
	.w2(32'hbbfe723b),
	.w3(32'h3b9f6d2c),
	.w4(32'hbbb2ac7a),
	.w5(32'hbc212ac9),
	.w6(32'h3c8a36a1),
	.w7(32'hbc160dd7),
	.w8(32'h3c15ab66),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba572a65),
	.w1(32'hb9ca678e),
	.w2(32'hba58a2a9),
	.w3(32'hba5d91e2),
	.w4(32'h3c9c6ac9),
	.w5(32'h3cd44107),
	.w6(32'h3bdcbe19),
	.w7(32'h3c3b91cb),
	.w8(32'h3a8aa4fb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49fc0d),
	.w1(32'hb9d05d0d),
	.w2(32'hba7b43d5),
	.w3(32'h3c21a9a0),
	.w4(32'h3aaa1038),
	.w5(32'hbc3e5de4),
	.w6(32'hbb25e7ef),
	.w7(32'hbae54798),
	.w8(32'h3abba0f9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1254ac),
	.w1(32'hbb984505),
	.w2(32'h3bc7b16f),
	.w3(32'h3a01bf9e),
	.w4(32'h3a831623),
	.w5(32'hbb550eb7),
	.w6(32'hbc094a07),
	.w7(32'hbca1e5e4),
	.w8(32'hbb6ba438),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccdc78),
	.w1(32'hbc3055ea),
	.w2(32'hbb861b67),
	.w3(32'hbba522c3),
	.w4(32'hbbaadf86),
	.w5(32'h395aeaca),
	.w6(32'hbbbb0d13),
	.w7(32'hbbbcdbc7),
	.w8(32'hbad5e9ff),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ec1a),
	.w1(32'hbb127c9d),
	.w2(32'hbca63f9f),
	.w3(32'hbba5f6cf),
	.w4(32'hbbc0aa91),
	.w5(32'hbb325892),
	.w6(32'hbc349a95),
	.w7(32'hbb88cbf7),
	.w8(32'hbbf478ed),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8223b6),
	.w1(32'h3b7cb228),
	.w2(32'hbb0fec8e),
	.w3(32'h3a047fe4),
	.w4(32'hbb6ab397),
	.w5(32'h3bbd04d7),
	.w6(32'h3ad683bf),
	.w7(32'hbb611ef0),
	.w8(32'h3b6a7b7d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf3b04),
	.w1(32'hbaeb6a84),
	.w2(32'hbc26d194),
	.w3(32'h3ba78263),
	.w4(32'h3c9f0699),
	.w5(32'h3baaba98),
	.w6(32'h3b4e2480),
	.w7(32'hbb5583e1),
	.w8(32'hbb950cf0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb809a2ec),
	.w1(32'hbc0c752d),
	.w2(32'hbb8ca206),
	.w3(32'hbc49bbd6),
	.w4(32'h3b36bf01),
	.w5(32'hbc12e908),
	.w6(32'hbad9dbcb),
	.w7(32'hbc466121),
	.w8(32'hba05f9d3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8e42),
	.w1(32'hbb01db73),
	.w2(32'hbbf5d2be),
	.w3(32'hbc5a532a),
	.w4(32'hbb238849),
	.w5(32'hbb674de0),
	.w6(32'hbb152ae6),
	.w7(32'hbba128cd),
	.w8(32'hba3c5c19),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5618a6),
	.w1(32'hbc01dfe4),
	.w2(32'h39e38fea),
	.w3(32'h3ad76dd7),
	.w4(32'hbb33eb42),
	.w5(32'hbcc09ad7),
	.w6(32'h3bd41a4d),
	.w7(32'hbc570f4d),
	.w8(32'h3c2a7dce),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e19d1),
	.w1(32'hbb2e1722),
	.w2(32'h3ca604b0),
	.w3(32'h3bddd61a),
	.w4(32'hbbcea8c7),
	.w5(32'h3c290a70),
	.w6(32'h3b33f0f8),
	.w7(32'h3b4fb173),
	.w8(32'h3cbfb8d3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb30aac),
	.w1(32'hbc8ee93e),
	.w2(32'hbc05a1aa),
	.w3(32'hbaf50721),
	.w4(32'h3b2b1912),
	.w5(32'hbc6cb089),
	.w6(32'h3c90177c),
	.w7(32'h3b3a6716),
	.w8(32'hbc32566a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b491),
	.w1(32'hbc183a08),
	.w2(32'h3c8f1399),
	.w3(32'hbaa3579b),
	.w4(32'h3c86d697),
	.w5(32'hbaae2950),
	.w6(32'h3bf36e32),
	.w7(32'h3bc93196),
	.w8(32'h3ac5a0f6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cadf6),
	.w1(32'h3cb770d5),
	.w2(32'hb809dd1a),
	.w3(32'hbc05aeab),
	.w4(32'hbc03dd01),
	.w5(32'h3b833db3),
	.w6(32'h3c28ef04),
	.w7(32'hbaae25aa),
	.w8(32'h3abc78a7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9fa81),
	.w1(32'hbb693565),
	.w2(32'hbc203efd),
	.w3(32'hbc33580c),
	.w4(32'hbbb4acad),
	.w5(32'hbbbb6d13),
	.w6(32'hb7c684d3),
	.w7(32'h3c0fde85),
	.w8(32'h3c156ccc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b560ad6),
	.w1(32'h3b3e425d),
	.w2(32'hbb4bc8d2),
	.w3(32'hbaca8797),
	.w4(32'hbd1906d4),
	.w5(32'h3b0f96bb),
	.w6(32'hbb835dc8),
	.w7(32'hbc1cfeee),
	.w8(32'h3bf3e740),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07124a),
	.w1(32'hbb8f8bb3),
	.w2(32'h3b25bc02),
	.w3(32'hbc6d8ce9),
	.w4(32'hbbc6b4d8),
	.w5(32'h3ae7c587),
	.w6(32'h3a7cbd19),
	.w7(32'hbb945eb0),
	.w8(32'h3b997ffb),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41f90a),
	.w1(32'hbc7983d4),
	.w2(32'hbc193a12),
	.w3(32'h39eedacf),
	.w4(32'hbc4e3c4f),
	.w5(32'hbb11fa71),
	.w6(32'hbc0296be),
	.w7(32'hb70aec0d),
	.w8(32'h3afc37e6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc228dbd),
	.w1(32'hba8be227),
	.w2(32'hba0d62fa),
	.w3(32'hbc105340),
	.w4(32'h3bf9e989),
	.w5(32'h3bb662be),
	.w6(32'hbb6780d5),
	.w7(32'hbb1b9b7d),
	.w8(32'h3c27f8df),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b264455),
	.w1(32'h3b0348ce),
	.w2(32'hbc64c471),
	.w3(32'h3b88878a),
	.w4(32'hbb2c8db2),
	.w5(32'h35d35e38),
	.w6(32'hbb4301e2),
	.w7(32'hbb8106de),
	.w8(32'h3beb5fee),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf584b4),
	.w1(32'hbc310af0),
	.w2(32'h3c0a0e01),
	.w3(32'h3ab175fe),
	.w4(32'hbbb57579),
	.w5(32'hba97fe63),
	.w6(32'hbc9908b8),
	.w7(32'hbbc5acd0),
	.w8(32'h3c4e28e2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0060f1),
	.w1(32'hbc8947a8),
	.w2(32'h3c9ee86e),
	.w3(32'hbb5c60fb),
	.w4(32'h3ba58ffc),
	.w5(32'hbb8200f3),
	.w6(32'h3bcaf9ca),
	.w7(32'h3c0e7d96),
	.w8(32'h3d0988bd),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c8e61),
	.w1(32'hbc6d565e),
	.w2(32'hbb8eaf7f),
	.w3(32'hbb9e7e11),
	.w4(32'h3b22c0d5),
	.w5(32'h3a5f5a72),
	.w6(32'hbbf5d4fd),
	.w7(32'h3b77f69f),
	.w8(32'hbc34366c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4db20),
	.w1(32'h3b78e06e),
	.w2(32'hbbf17110),
	.w3(32'h3acfe37c),
	.w4(32'h3b8f88cb),
	.w5(32'h3b214c77),
	.w6(32'hbc5823d9),
	.w7(32'h3b65bfeb),
	.w8(32'hba5c0387),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcf61a),
	.w1(32'hbb36b603),
	.w2(32'h35a76e1f),
	.w3(32'hba70ca05),
	.w4(32'h3a390310),
	.w5(32'hbb88c11f),
	.w6(32'h3b39c7f1),
	.w7(32'hba98a505),
	.w8(32'hbc0903d6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe387f8),
	.w1(32'hbc01cbac),
	.w2(32'h3811a2f0),
	.w3(32'h3b8a15fd),
	.w4(32'hbb8f49a6),
	.w5(32'h3b99f81c),
	.w6(32'hbc64c604),
	.w7(32'hbaa2e29f),
	.w8(32'h3b5fce7e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983fef3),
	.w1(32'hbbf292b9),
	.w2(32'h3b4e8897),
	.w3(32'h3bb84af9),
	.w4(32'hbbe3ed07),
	.w5(32'hbb07f2f4),
	.w6(32'h3b2cc286),
	.w7(32'hbb0889c0),
	.w8(32'h3b648ef2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc213f25),
	.w1(32'hbbd969b3),
	.w2(32'hbbef9ed3),
	.w3(32'hbc21fa49),
	.w4(32'h3abe1b83),
	.w5(32'h3a6d7721),
	.w6(32'hbc01c713),
	.w7(32'h3c76086b),
	.w8(32'hbbfd21d7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96110d),
	.w1(32'hba636a1a),
	.w2(32'h3b1422e0),
	.w3(32'hbc450591),
	.w4(32'h3bc7b8ee),
	.w5(32'hbbe0fc4c),
	.w6(32'h3cb6157b),
	.w7(32'hbb903d7d),
	.w8(32'h3b1805e5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85fb35),
	.w1(32'h3b8314cf),
	.w2(32'hbb5c9da9),
	.w3(32'h3bf3318b),
	.w4(32'hbbee5a89),
	.w5(32'h3630a915),
	.w6(32'hbbb137d7),
	.w7(32'h3c58d1b5),
	.w8(32'h3b893712),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d2300),
	.w1(32'hbb28fb0a),
	.w2(32'h3ae32264),
	.w3(32'hbb8e30b4),
	.w4(32'hbb28ca15),
	.w5(32'hbbf01ffc),
	.w6(32'h3c296479),
	.w7(32'hb9ff02fd),
	.w8(32'h3bcb8a73),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65cebf),
	.w1(32'hbb061ca8),
	.w2(32'h3ce47d26),
	.w3(32'hbc96b810),
	.w4(32'hbbe1037e),
	.w5(32'h3bd8ca2a),
	.w6(32'hbad59e7f),
	.w7(32'h3c334be5),
	.w8(32'h3b13f51c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa3ce),
	.w1(32'hbb8c7fc4),
	.w2(32'hbc386824),
	.w3(32'hbad76f6e),
	.w4(32'hbade4b85),
	.w5(32'hbbdd73e3),
	.w6(32'hba9263ba),
	.w7(32'hbbac7628),
	.w8(32'hb8d791a5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a900cc0),
	.w1(32'hbca3edd2),
	.w2(32'h3c0a599f),
	.w3(32'hbbe8b78a),
	.w4(32'hbae515b0),
	.w5(32'h3c304cf0),
	.w6(32'hba14b280),
	.w7(32'hbb8f6ef7),
	.w8(32'h3cd8adf7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829c17),
	.w1(32'hbbe0df65),
	.w2(32'h3ae8057d),
	.w3(32'h3b44da60),
	.w4(32'hbc3c7d55),
	.w5(32'hbb3e9272),
	.w6(32'hbbbeaf64),
	.w7(32'h3c52a038),
	.w8(32'hbb0e16a9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3e97d),
	.w1(32'h3bb1bb4b),
	.w2(32'h3c28f1c0),
	.w3(32'h3c0776a0),
	.w4(32'h3ba07e4a),
	.w5(32'h3c4a6c12),
	.w6(32'h3bc86ff1),
	.w7(32'hb95ae15e),
	.w8(32'h3b83b6a4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc244e5f),
	.w1(32'h3bdce570),
	.w2(32'hbbba7514),
	.w3(32'h3b473062),
	.w4(32'h3af81680),
	.w5(32'hbaf30c85),
	.w6(32'hbbc89414),
	.w7(32'h3c1ad28b),
	.w8(32'hbbda38d6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ce50e),
	.w1(32'hbaaaba3f),
	.w2(32'hbacfd873),
	.w3(32'h3b92ef85),
	.w4(32'h3c48d2dd),
	.w5(32'h3c17ad32),
	.w6(32'h3af12d0e),
	.w7(32'h3be0acbc),
	.w8(32'hbb441750),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130203),
	.w1(32'hba8f83e1),
	.w2(32'h3c43f88a),
	.w3(32'h3cc59c72),
	.w4(32'hbaf7b36e),
	.w5(32'h3a120538),
	.w6(32'h3aab37b2),
	.w7(32'hbbabf4dd),
	.w8(32'hbb9d2cc7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04d16f),
	.w1(32'hbc0c3834),
	.w2(32'hbbef1fdf),
	.w3(32'hbcfdbf91),
	.w4(32'h3bbe0564),
	.w5(32'hbbc48dac),
	.w6(32'h3ba2ad67),
	.w7(32'hbada95f3),
	.w8(32'hbab443db),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8619cd),
	.w1(32'h3c1a9c3e),
	.w2(32'h3c0d335d),
	.w3(32'h3b5e4c65),
	.w4(32'hbbb45bc9),
	.w5(32'h3bd896d6),
	.w6(32'hb89eb545),
	.w7(32'h3b94324a),
	.w8(32'h3c4ad774),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cd158),
	.w1(32'hb9a4ac90),
	.w2(32'h3c37570a),
	.w3(32'hbc860f52),
	.w4(32'h3956ac4b),
	.w5(32'hb96c8e3b),
	.w6(32'hbba817d8),
	.w7(32'hbbb12ab4),
	.w8(32'hba9a5c40),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada8b19),
	.w1(32'h3c0be12a),
	.w2(32'h3b0b147f),
	.w3(32'h3b74db69),
	.w4(32'h3b123678),
	.w5(32'h3b57bddb),
	.w6(32'h3abbbf39),
	.w7(32'h3c69b407),
	.w8(32'hbbcefe58),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87fdcc),
	.w1(32'hbbfee0f6),
	.w2(32'h3d032bc9),
	.w3(32'hbbed0ac5),
	.w4(32'h3ae25228),
	.w5(32'h3a4f59e4),
	.w6(32'hbb99c18a),
	.w7(32'hbaff7e1b),
	.w8(32'hbc9b0739),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ead62),
	.w1(32'hbb9cc73e),
	.w2(32'hbbad344d),
	.w3(32'hbb83a9ae),
	.w4(32'h39f0acda),
	.w5(32'h3cab753f),
	.w6(32'h3c1f35a9),
	.w7(32'h3b6d63f4),
	.w8(32'hbab432eb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45fec4),
	.w1(32'hbc54518c),
	.w2(32'h3b413c9b),
	.w3(32'hbc477905),
	.w4(32'hbc0b89d7),
	.w5(32'h3be5c80a),
	.w6(32'h3bc21b3b),
	.w7(32'h399d65f5),
	.w8(32'h3ba13569),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ab97eb),
	.w1(32'hbc46da44),
	.w2(32'hbbd3bb13),
	.w3(32'h3b0f472a),
	.w4(32'h3a9c4397),
	.w5(32'h3d5b08a6),
	.w6(32'hbc755c4b),
	.w7(32'h3b9dbfa0),
	.w8(32'hbc05cea1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bb1fa4),
	.w1(32'h3c0356ed),
	.w2(32'h3ac10d1f),
	.w3(32'hbb9a1f71),
	.w4(32'hbb879688),
	.w5(32'hbb5b2906),
	.w6(32'hbc1b8e14),
	.w7(32'hbba22f47),
	.w8(32'h3b531d67),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd62dc3),
	.w1(32'h39e045f5),
	.w2(32'hbc38bd7c),
	.w3(32'h3a779227),
	.w4(32'hb9c589be),
	.w5(32'h3c106a37),
	.w6(32'h32384e2f),
	.w7(32'hbb247c0d),
	.w8(32'hbb55ab2e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1be52),
	.w1(32'hbb122aa0),
	.w2(32'h3b44d706),
	.w3(32'h3bf4850e),
	.w4(32'hbb42aa94),
	.w5(32'h3b9437cf),
	.w6(32'h3c29df03),
	.w7(32'h3c09ca7a),
	.w8(32'hbc3968a4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e76f),
	.w1(32'h3c7f5f8d),
	.w2(32'hbc45e001),
	.w3(32'hba7552c6),
	.w4(32'h3b60718d),
	.w5(32'hbb26872a),
	.w6(32'h3bfa2e71),
	.w7(32'hbb9b50c5),
	.w8(32'h3af5f58f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74d7bf),
	.w1(32'h37ebd63e),
	.w2(32'h3bda7040),
	.w3(32'hbb5d2edd),
	.w4(32'h3c2a9e38),
	.w5(32'h3bcc8fa6),
	.w6(32'h3cb9398e),
	.w7(32'h3a2fc5f7),
	.w8(32'h3c6c35ae),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a149d09),
	.w1(32'hbc0fc034),
	.w2(32'h3b268588),
	.w3(32'h3bb6836f),
	.w4(32'h3bc67ffb),
	.w5(32'hba295bd4),
	.w6(32'hba059fc7),
	.w7(32'hbb02f663),
	.w8(32'h3bb57ec0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d5416),
	.w1(32'h3c1eefb5),
	.w2(32'hbae37c21),
	.w3(32'hb78e6c96),
	.w4(32'h3b3397b6),
	.w5(32'h3b08a1d2),
	.w6(32'hbb9cc9df),
	.w7(32'h3a6117f9),
	.w8(32'hba669919),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1c597),
	.w1(32'hbb7e9f98),
	.w2(32'h3c01a33d),
	.w3(32'h3b2bd0cb),
	.w4(32'hb9fdc01f),
	.w5(32'h372a194a),
	.w6(32'h3b549643),
	.w7(32'h3b347b9b),
	.w8(32'h3bd424c2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68910c),
	.w1(32'h3a4b0439),
	.w2(32'hbba52840),
	.w3(32'h3b86bfef),
	.w4(32'hbac6943d),
	.w5(32'h3a9c82f6),
	.w6(32'h3b06b723),
	.w7(32'h3b537403),
	.w8(32'h3a8b2957),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8d387),
	.w1(32'h3c3e4bd0),
	.w2(32'hbc52328c),
	.w3(32'hbc59af87),
	.w4(32'hbbca2be9),
	.w5(32'hbb4be329),
	.w6(32'hbbc7ade4),
	.w7(32'hba8765e0),
	.w8(32'h38feefe0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0500),
	.w1(32'h3c3509c3),
	.w2(32'hbc3ff0f4),
	.w3(32'h3a06d7a8),
	.w4(32'h39969200),
	.w5(32'hbb021aa9),
	.w6(32'h3c2d162f),
	.w7(32'h3ab1d649),
	.w8(32'h3c31bb47),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00255),
	.w1(32'h3b84f8a1),
	.w2(32'hbb8961e9),
	.w3(32'h3b8fb519),
	.w4(32'h3a381345),
	.w5(32'hbbb527f1),
	.w6(32'h39508590),
	.w7(32'hbbf798d5),
	.w8(32'hba872d82),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e8538),
	.w1(32'h39649f80),
	.w2(32'h3ae3e1d8),
	.w3(32'h3b7cd1c3),
	.w4(32'h3a1ae7f3),
	.w5(32'h3b23ea14),
	.w6(32'h3a104389),
	.w7(32'h3c1b2a54),
	.w8(32'h3a3171aa),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c613e),
	.w1(32'h3a7e2feb),
	.w2(32'hbb0b0efe),
	.w3(32'h3c319eeb),
	.w4(32'hbb4daac9),
	.w5(32'hbba1905c),
	.w6(32'hba872a97),
	.w7(32'h3bb4ae9f),
	.w8(32'hba3591d2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf380ca),
	.w1(32'h3b44b7cf),
	.w2(32'hbc38bbc3),
	.w3(32'hbae9598a),
	.w4(32'hbc1f045f),
	.w5(32'h3b4b1216),
	.w6(32'h3c88f409),
	.w7(32'h3bab808b),
	.w8(32'h3c01541b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41ffa4),
	.w1(32'h3b860ba7),
	.w2(32'hbc4b5a28),
	.w3(32'hbbf03282),
	.w4(32'h3c0b4b1b),
	.w5(32'hbb77bcac),
	.w6(32'h3c3e773d),
	.w7(32'h3bebd4ef),
	.w8(32'h3b86bf86),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb944),
	.w1(32'hbbe02f1a),
	.w2(32'hbc460cdc),
	.w3(32'h3c481639),
	.w4(32'hb9a5e7ee),
	.w5(32'h3a46d335),
	.w6(32'hbaf8c741),
	.w7(32'h3ab098dc),
	.w8(32'hbb5faf0d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba713586),
	.w1(32'hbb8d0258),
	.w2(32'h3c22e5de),
	.w3(32'h3bc84b63),
	.w4(32'h3ac39dfd),
	.w5(32'hba821b2b),
	.w6(32'hbb963a21),
	.w7(32'h3befa487),
	.w8(32'h3a840e4c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe94bee),
	.w1(32'hbb344d80),
	.w2(32'h3cdb7736),
	.w3(32'h3ab8b96a),
	.w4(32'hbbee0074),
	.w5(32'hbb825640),
	.w6(32'hbb36b461),
	.w7(32'hbbce8d9d),
	.w8(32'hbc19fa35),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdbb41),
	.w1(32'h3b07fac3),
	.w2(32'h3a4f56f5),
	.w3(32'hbb6f2fdf),
	.w4(32'hbb57d74f),
	.w5(32'hbbd9f1f3),
	.w6(32'hbc6b5fce),
	.w7(32'hbbc36687),
	.w8(32'hbbae9c67),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea8500),
	.w1(32'hbc27bebf),
	.w2(32'h3be0583b),
	.w3(32'h3c90b662),
	.w4(32'hba7b94ad),
	.w5(32'h3c2f3e69),
	.w6(32'hba50bc37),
	.w7(32'hbaddafb7),
	.w8(32'hbb08c396),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac689df),
	.w1(32'hba94deed),
	.w2(32'hbba42c74),
	.w3(32'h39e18a2f),
	.w4(32'hbba04fea),
	.w5(32'hbaba6541),
	.w6(32'h3cceead3),
	.w7(32'h3c4e0f95),
	.w8(32'hba5c2874),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f390e),
	.w1(32'hbbe1ff02),
	.w2(32'hbb18c234),
	.w3(32'hbc76aa84),
	.w4(32'hbbab087c),
	.w5(32'h3bfc52d8),
	.w6(32'hb999da3a),
	.w7(32'hbb93421c),
	.w8(32'hbad7aa3c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebcb29),
	.w1(32'h3bb9824b),
	.w2(32'h3bdcbb92),
	.w3(32'h3c359b2b),
	.w4(32'h3ba48a7b),
	.w5(32'hbbde8007),
	.w6(32'h3b59116d),
	.w7(32'h39d77ab0),
	.w8(32'h3beef38b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94df630),
	.w1(32'h3b891ab7),
	.w2(32'h3bb23262),
	.w3(32'h3a820216),
	.w4(32'hbc99de92),
	.w5(32'h3a836e67),
	.w6(32'h3bca2b23),
	.w7(32'h3c3e88e6),
	.w8(32'hbc5c7a31),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefe746),
	.w1(32'h3bb01891),
	.w2(32'hbba1099c),
	.w3(32'hbb0b534b),
	.w4(32'hbb5e5dd6),
	.w5(32'h3b9a4a71),
	.w6(32'hbc5ef45f),
	.w7(32'hbb9014ab),
	.w8(32'hbb59a11e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72e7e),
	.w1(32'h3b5206fa),
	.w2(32'hbb8b6e39),
	.w3(32'hbb839814),
	.w4(32'h3b3fee38),
	.w5(32'hbc16599b),
	.w6(32'hbc004712),
	.w7(32'hbc4d6489),
	.w8(32'hbbcb60eb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadca9ba),
	.w1(32'hbc1b386c),
	.w2(32'h3a9df4ab),
	.w3(32'hbc1264d6),
	.w4(32'h38a33a58),
	.w5(32'hbb947a71),
	.w6(32'hbc601593),
	.w7(32'h3b3f3805),
	.w8(32'hbbc8ccdf),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccda17),
	.w1(32'h3b43fafb),
	.w2(32'hb983f8a6),
	.w3(32'hbb175a9c),
	.w4(32'h3af51312),
	.w5(32'hbbe1fd41),
	.w6(32'hbc29864a),
	.w7(32'hbac71b33),
	.w8(32'hbbe31b23),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc190),
	.w1(32'hbbf63d20),
	.w2(32'hb54bc9c6),
	.w3(32'hbb50ee90),
	.w4(32'hbb84b11e),
	.w5(32'h3bb33c48),
	.w6(32'hbbb7e348),
	.w7(32'hbb989ff6),
	.w8(32'hb9b71b21),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4819e),
	.w1(32'hbb0b276b),
	.w2(32'hbc3ff5f0),
	.w3(32'hba5c25d3),
	.w4(32'h3b280b5f),
	.w5(32'h3bb8ff24),
	.w6(32'hbc502057),
	.w7(32'hb733d223),
	.w8(32'hbb257c08),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90de50),
	.w1(32'h3c96b04c),
	.w2(32'h3bb1687d),
	.w3(32'h3b16fa9e),
	.w4(32'h3b220b18),
	.w5(32'hbbeba25a),
	.w6(32'h3b42e7d6),
	.w7(32'h3aa4f8b0),
	.w8(32'hbba647f9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146f4b),
	.w1(32'hbb7c7ccc),
	.w2(32'h3a1919fb),
	.w3(32'h3bcd418c),
	.w4(32'hbaee78ba),
	.w5(32'hbbccb2d9),
	.w6(32'hbba15262),
	.w7(32'h3a94f0de),
	.w8(32'h3b5280d9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a2661),
	.w1(32'hbbe91b73),
	.w2(32'h3b962926),
	.w3(32'h3b3118e2),
	.w4(32'hb92843c5),
	.w5(32'h3bc8a3d5),
	.w6(32'h3b3d9b90),
	.w7(32'hba3d5a81),
	.w8(32'h3b84754f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fd88),
	.w1(32'hbbca8d1e),
	.w2(32'h39bb4b2f),
	.w3(32'h3bd67123),
	.w4(32'h3abad017),
	.w5(32'hbb76d4be),
	.w6(32'hbb188f44),
	.w7(32'hb51e11a1),
	.w8(32'h3b53dad0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dbd5d),
	.w1(32'hbc2d5ffd),
	.w2(32'hbb64b488),
	.w3(32'h3c4c464e),
	.w4(32'hbb8bd6af),
	.w5(32'hbb826cc8),
	.w6(32'h3c4cbc9a),
	.w7(32'h3b71ee0f),
	.w8(32'hb79566a1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4d3d9),
	.w1(32'h3ac9ec08),
	.w2(32'h3a88fb84),
	.w3(32'hbb044249),
	.w4(32'hb9d70cd4),
	.w5(32'hbaba0625),
	.w6(32'hbbc149cf),
	.w7(32'hba94ecbe),
	.w8(32'hbc8fb59c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b890dc6),
	.w1(32'hbb869753),
	.w2(32'h3ba56725),
	.w3(32'hbb3e7703),
	.w4(32'h3d05c3d9),
	.w5(32'h3afffc8d),
	.w6(32'h38757a04),
	.w7(32'hbc17e190),
	.w8(32'hbc2e0adb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10424b),
	.w1(32'h3b64f514),
	.w2(32'h3c01bbd1),
	.w3(32'hbb8ced22),
	.w4(32'h3b48aa95),
	.w5(32'h3bb20171),
	.w6(32'hbb298e3a),
	.w7(32'h3bb0a68f),
	.w8(32'h3aadb894),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dcf6d),
	.w1(32'h3c211831),
	.w2(32'hb8b148a7),
	.w3(32'hbb9dd604),
	.w4(32'h3cb4882e),
	.w5(32'hbb2cd2cb),
	.w6(32'hb96eb1eb),
	.w7(32'hbbab52b6),
	.w8(32'h3a982705),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd4a67),
	.w1(32'hbad9b363),
	.w2(32'h3c315a8a),
	.w3(32'hbb9a696b),
	.w4(32'hb79534fc),
	.w5(32'h3b38c4b0),
	.w6(32'hbaa7ef93),
	.w7(32'hbbe54764),
	.w8(32'h3c1a1d5e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c656b3e),
	.w1(32'h3b7ab190),
	.w2(32'hbb1992f4),
	.w3(32'hbb9b9cdb),
	.w4(32'h3abfa9e6),
	.w5(32'h3c170212),
	.w6(32'h3c054388),
	.w7(32'hbbd19658),
	.w8(32'hbbc6b351),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c2ae8),
	.w1(32'hbb42caf2),
	.w2(32'h39cdb3b5),
	.w3(32'hba3bf45f),
	.w4(32'h3c23ff83),
	.w5(32'hbba62903),
	.w6(32'hbc03946d),
	.w7(32'hbc71d5c9),
	.w8(32'h3b38e29a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c3c9),
	.w1(32'hb9e0d9a9),
	.w2(32'h39f929c6),
	.w3(32'h3b79d8fe),
	.w4(32'h3b41a1e8),
	.w5(32'hbc230b57),
	.w6(32'hbbc3b570),
	.w7(32'h3c1a8888),
	.w8(32'hbb6918e8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb720a1f),
	.w1(32'hbb8b52eb),
	.w2(32'hbbd9ffb6),
	.w3(32'h3b842690),
	.w4(32'hbc24fa43),
	.w5(32'hbc863215),
	.w6(32'hbc94f65d),
	.w7(32'h3a0d6ceb),
	.w8(32'hba9653e6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe16e0),
	.w1(32'hbb6e5c54),
	.w2(32'h3c8736be),
	.w3(32'hbc54671c),
	.w4(32'hbc05b91e),
	.w5(32'hbcb573a9),
	.w6(32'hbc84fd57),
	.w7(32'hbbf5cbc1),
	.w8(32'h3ca9f702),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf461ce),
	.w1(32'hbcc4b2cb),
	.w2(32'hbbd2d509),
	.w3(32'hbb9ee081),
	.w4(32'hbc435c90),
	.w5(32'hbb62d314),
	.w6(32'hbbda9df4),
	.w7(32'hbbcf821a),
	.w8(32'hbc53afb6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c371d59),
	.w1(32'h3d138a39),
	.w2(32'hbc448924),
	.w3(32'hbc2a5e61),
	.w4(32'hbc789a80),
	.w5(32'h3bcfb040),
	.w6(32'hbbd869ac),
	.w7(32'h3c174cd2),
	.w8(32'h3ca590e2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeef42),
	.w1(32'hbc8c221c),
	.w2(32'h3c10e946),
	.w3(32'h39aec19f),
	.w4(32'hbc6bf712),
	.w5(32'h3c925de8),
	.w6(32'hbc890780),
	.w7(32'h3c596bf5),
	.w8(32'h3ad3c0fe),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968113),
	.w1(32'h3b70a27c),
	.w2(32'hbbf94ea9),
	.w3(32'hb88fc2e4),
	.w4(32'hbb1244e3),
	.w5(32'h3c5ef0ef),
	.w6(32'hbd0dbaaa),
	.w7(32'h3c85108b),
	.w8(32'hbc7de1b7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d1801),
	.w1(32'hbbe8486e),
	.w2(32'h3c1c7a03),
	.w3(32'hbc949fa9),
	.w4(32'hbd08f95f),
	.w5(32'hbb5f75e4),
	.w6(32'h3b8732d5),
	.w7(32'h3c476a07),
	.w8(32'hba830079),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2a36),
	.w1(32'hba59d63f),
	.w2(32'hba89d9eb),
	.w3(32'h3be7599c),
	.w4(32'h3af4beed),
	.w5(32'h3b8be0ed),
	.w6(32'hbb491c34),
	.w7(32'hbc03cb06),
	.w8(32'hbc841af4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbe645),
	.w1(32'h3ad20140),
	.w2(32'hbc9de6cd),
	.w3(32'hbc5554a8),
	.w4(32'h3c86a61c),
	.w5(32'h3cd3098d),
	.w6(32'hbca6c953),
	.w7(32'hbb8835c4),
	.w8(32'h3cc12f0a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb9e8),
	.w1(32'h3c231a21),
	.w2(32'hbc04678f),
	.w3(32'hbb996505),
	.w4(32'h3bc26eef),
	.w5(32'hbca807b3),
	.w6(32'h3bf0326c),
	.w7(32'h3b3cfb6c),
	.w8(32'hbbe2296f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb94b37),
	.w1(32'h3bbd8fcc),
	.w2(32'h3c08f05d),
	.w3(32'h3c08a404),
	.w4(32'hbc9a87fa),
	.w5(32'h3beb48b3),
	.w6(32'hba92b817),
	.w7(32'hbbd4dc44),
	.w8(32'hbc090fad),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35ab71),
	.w1(32'h3c0721df),
	.w2(32'hbc14849a),
	.w3(32'hbc88d070),
	.w4(32'hbb94ab8f),
	.w5(32'hbaa6a850),
	.w6(32'h3cb285c4),
	.w7(32'h3cb8b8b4),
	.w8(32'hba08eb8f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2efe1),
	.w1(32'hbc60e70c),
	.w2(32'hbca09f85),
	.w3(32'hbb2ee104),
	.w4(32'hbb3c6f20),
	.w5(32'hbb82398e),
	.w6(32'h3c918ce4),
	.w7(32'h3baf24cc),
	.w8(32'hbc3035a1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078d67),
	.w1(32'hbc111f27),
	.w2(32'hbc0644db),
	.w3(32'hbbd04093),
	.w4(32'h3b5b0113),
	.w5(32'hbc363fb4),
	.w6(32'hbac2ecb4),
	.w7(32'hbb08b88b),
	.w8(32'hbbabbfb7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb720a08),
	.w1(32'hba9bba84),
	.w2(32'hbc05e586),
	.w3(32'h361faa6c),
	.w4(32'hbc1432e6),
	.w5(32'h3ca0b6fa),
	.w6(32'hbc5f62d7),
	.w7(32'hbc1e3f23),
	.w8(32'hbc663084),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65a67c),
	.w1(32'hbc155d28),
	.w2(32'hbc09be0a),
	.w3(32'hbbf5d826),
	.w4(32'hbc897d40),
	.w5(32'h3a7a13ff),
	.w6(32'hbc953127),
	.w7(32'h3c117114),
	.w8(32'hbb1e32f7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390513ee),
	.w1(32'hbad02461),
	.w2(32'h3b09fda6),
	.w3(32'h3bdbd646),
	.w4(32'hbc3d7907),
	.w5(32'hbce3cdd3),
	.w6(32'h3d13b1ba),
	.w7(32'hbcd40927),
	.w8(32'hbb2e65c0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60c9bb),
	.w1(32'hbc089945),
	.w2(32'h3c4c71d3),
	.w3(32'h3b534b5d),
	.w4(32'hbb9b8e7c),
	.w5(32'h3b874843),
	.w6(32'hbc816814),
	.w7(32'hbc571dab),
	.w8(32'hbb185f6a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c6625),
	.w1(32'hbbb9aa44),
	.w2(32'h3a14b54e),
	.w3(32'h3b515199),
	.w4(32'h3b19c63d),
	.w5(32'h3bfbfad3),
	.w6(32'h3c0dfeb8),
	.w7(32'hbbf7985b),
	.w8(32'h3aa00e96),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4608b91),
	.w1(32'h3c1a74b6),
	.w2(32'hbc000285),
	.w3(32'hbc848643),
	.w4(32'h3c661301),
	.w5(32'hbce689f2),
	.w6(32'hbaf05c97),
	.w7(32'hbc95d94e),
	.w8(32'h3b491a66),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb706ac),
	.w1(32'hba4b86dd),
	.w2(32'h37154061),
	.w3(32'h3b029765),
	.w4(32'hbc27f6a3),
	.w5(32'hbab98411),
	.w6(32'hbb14cf30),
	.w7(32'h3af4448d),
	.w8(32'hbc95597a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7182a),
	.w1(32'hbc95d42e),
	.w2(32'hbc40a179),
	.w3(32'h3cc71eb0),
	.w4(32'hbb9976a4),
	.w5(32'hbc551c0e),
	.w6(32'hb922a378),
	.w7(32'h3bca1932),
	.w8(32'hbc5df62b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11e88b),
	.w1(32'hbc4ac8a8),
	.w2(32'h3c2c5cac),
	.w3(32'hbc271cfc),
	.w4(32'h39b8fade),
	.w5(32'h3babb8ff),
	.w6(32'h3c4fd9e4),
	.w7(32'hbc502a03),
	.w8(32'hbbf6dde9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a48c5),
	.w1(32'h3a93279b),
	.w2(32'h3a8146fd),
	.w3(32'hbbe1d83f),
	.w4(32'hbc58af62),
	.w5(32'hbb6aa444),
	.w6(32'hbb8a5e3f),
	.w7(32'hbc51c9ef),
	.w8(32'h3c505505),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a6651),
	.w1(32'hbc140f70),
	.w2(32'hbc1e294a),
	.w3(32'h3a3e9ef8),
	.w4(32'h3b4a4558),
	.w5(32'h3b8d08d1),
	.w6(32'hbbe0401c),
	.w7(32'hbcafa391),
	.w8(32'hba22dabf),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc245d52),
	.w1(32'h3c7391c5),
	.w2(32'hbbe1174b),
	.w3(32'hbcc26e99),
	.w4(32'h3c139581),
	.w5(32'hbcade927),
	.w6(32'hbbc58bf5),
	.w7(32'h3b1d1b2c),
	.w8(32'hbd0235ca),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6004eb),
	.w1(32'hbc215d6e),
	.w2(32'hbc7f1dbd),
	.w3(32'hbca61f26),
	.w4(32'h3a04a809),
	.w5(32'h3c6a7339),
	.w6(32'h3c5f658b),
	.w7(32'hbc93610e),
	.w8(32'h3c48e623),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0152e8),
	.w1(32'hbc99a569),
	.w2(32'hbb2abce8),
	.w3(32'hbc329041),
	.w4(32'hbb05d2b1),
	.w5(32'h3be093ea),
	.w6(32'hbb5e11f0),
	.w7(32'h3c2401b9),
	.w8(32'hbcf32e06),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c962937),
	.w1(32'h3c376cc1),
	.w2(32'hbca0fb8b),
	.w3(32'h3bdef46d),
	.w4(32'hbbcc6c68),
	.w5(32'hbaf0efdf),
	.w6(32'h3c5ead4f),
	.w7(32'hbd3c7629),
	.w8(32'hbb7eb9e9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f8967),
	.w1(32'h3a65ba54),
	.w2(32'h3a5d85cd),
	.w3(32'hbc36068b),
	.w4(32'hbbded954),
	.w5(32'hbb49d703),
	.w6(32'h3c068996),
	.w7(32'hbb0f68cb),
	.w8(32'hba9e841e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba092c0),
	.w1(32'h3c7dc5e7),
	.w2(32'hba7192dc),
	.w3(32'hbc942fa1),
	.w4(32'hbb93a630),
	.w5(32'hbb85958e),
	.w6(32'h3b639ebe),
	.w7(32'hbb1b8d8c),
	.w8(32'hbc076c13),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule