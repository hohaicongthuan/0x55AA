module layer_8_featuremap_238(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad01f3c),
	.w1(32'hbc485f5d),
	.w2(32'hbccd2b00),
	.w3(32'h3c074957),
	.w4(32'hbbe7490d),
	.w5(32'hbb4d6091),
	.w6(32'hbc0d4fbc),
	.w7(32'hbc888999),
	.w8(32'h3c2679fa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0f981),
	.w1(32'hbb8d887a),
	.w2(32'hbbba890b),
	.w3(32'h3bdbb953),
	.w4(32'hbb0c613a),
	.w5(32'h3a942932),
	.w6(32'hbb9d8c23),
	.w7(32'hbbb86796),
	.w8(32'hba6c4db6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c1b9),
	.w1(32'h3b2bdec7),
	.w2(32'h3c8968da),
	.w3(32'hbb6225dd),
	.w4(32'h3c108337),
	.w5(32'h3c1542b9),
	.w6(32'hbbb6f10c),
	.w7(32'hba7c51d6),
	.w8(32'h3b7a4bd4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2afeaf),
	.w1(32'hba6837cc),
	.w2(32'h3cd0e05e),
	.w3(32'hbc167ac4),
	.w4(32'h3ca41909),
	.w5(32'h3cf198b7),
	.w6(32'hbca8b98b),
	.w7(32'hbc873dd5),
	.w8(32'hba5f5c30),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d16f1a6),
	.w1(32'h3b694276),
	.w2(32'hbb068b6b),
	.w3(32'h3bcb6013),
	.w4(32'h3adf3c04),
	.w5(32'h3a9917f8),
	.w6(32'h3bfce95b),
	.w7(32'h3bb61d89),
	.w8(32'h3b111da3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a784f),
	.w1(32'hbc8481c6),
	.w2(32'hbcea6ec9),
	.w3(32'hba76d4a8),
	.w4(32'hbceb25e0),
	.w5(32'hbd0170ae),
	.w6(32'h3ba1c09e),
	.w7(32'hbc0db725),
	.w8(32'hbcc8e249),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ca2bc),
	.w1(32'h3b9ee64e),
	.w2(32'h3bb4c0c6),
	.w3(32'hbcd0b40e),
	.w4(32'h3a9965ea),
	.w5(32'h3b15e0d0),
	.w6(32'h3be0dddd),
	.w7(32'h3b5b2840),
	.w8(32'h3ace34c2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb9994),
	.w1(32'h39829cac),
	.w2(32'hbc0530bf),
	.w3(32'hba60d747),
	.w4(32'h3b9f6b13),
	.w5(32'h39afdecc),
	.w6(32'hbb30ac0e),
	.w7(32'hbbcc88a3),
	.w8(32'h3b8b87cc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46c213),
	.w1(32'hbbc9352e),
	.w2(32'hbb3f4605),
	.w3(32'h3981a919),
	.w4(32'h3b928a47),
	.w5(32'h3bda603f),
	.w6(32'hbb5a8785),
	.w7(32'hbc718780),
	.w8(32'h394b4cf1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4a5fb),
	.w1(32'h399b92de),
	.w2(32'hbc816f94),
	.w3(32'hb857bd60),
	.w4(32'h3b857441),
	.w5(32'h3c8cf7f4),
	.w6(32'hbbb5dcbc),
	.w7(32'hbb968903),
	.w8(32'hbbee248c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35aeaf),
	.w1(32'h3bed1034),
	.w2(32'hbb6fbc4f),
	.w3(32'h3c923720),
	.w4(32'h3ac5e729),
	.w5(32'hbc3ca3e2),
	.w6(32'h3c9ebad2),
	.w7(32'h3c64de33),
	.w8(32'h3c351ec0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb669a98),
	.w1(32'h3bbd60c9),
	.w2(32'h3c5d68b2),
	.w3(32'hbb8d783a),
	.w4(32'h3be51643),
	.w5(32'h3bf706a7),
	.w6(32'h3b9ccacb),
	.w7(32'h3c603c7b),
	.w8(32'h3c0a890d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4c93d),
	.w1(32'hbb2cc6a2),
	.w2(32'hba42ec4c),
	.w3(32'h3a4024f0),
	.w4(32'h3c0f2f36),
	.w5(32'h3c4d3354),
	.w6(32'hba40eddc),
	.w7(32'h3b91de8c),
	.w8(32'hbb2c8181),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944c9f),
	.w1(32'hbaecf458),
	.w2(32'hbc05aa3d),
	.w3(32'h3c094f2b),
	.w4(32'hbb0cd829),
	.w5(32'hbad84439),
	.w6(32'hbc1fc134),
	.w7(32'hbbb5c001),
	.w8(32'h3b4c74de),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9fcde),
	.w1(32'hbace08d6),
	.w2(32'h3a84f66b),
	.w3(32'hbb7988d8),
	.w4(32'h3b25b4f9),
	.w5(32'hba0a806b),
	.w6(32'h3b13893b),
	.w7(32'hbb8946a9),
	.w8(32'hbb43776b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7d133),
	.w1(32'hbc855d16),
	.w2(32'hbbb09874),
	.w3(32'hbc1f23a2),
	.w4(32'hbc59b1ac),
	.w5(32'h3c199423),
	.w6(32'hbb670a4f),
	.w7(32'hbc4366ea),
	.w8(32'h3b718862),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b859b3d),
	.w1(32'h3bfbbcf3),
	.w2(32'hbb463858),
	.w3(32'hbb9b7c4d),
	.w4(32'h3ac84958),
	.w5(32'h3b9dd5e8),
	.w6(32'hbb6fa23f),
	.w7(32'h3c135467),
	.w8(32'h3c188f73),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42d610),
	.w1(32'h3bf0f237),
	.w2(32'h3c254f53),
	.w3(32'h3bdf01d9),
	.w4(32'h3c086fcf),
	.w5(32'h3bb4cd85),
	.w6(32'hbb366463),
	.w7(32'h38e05042),
	.w8(32'h3bc00536),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31b518),
	.w1(32'h3bde6738),
	.w2(32'h3c36b5b9),
	.w3(32'h3bb88743),
	.w4(32'hbb1257ad),
	.w5(32'h3bfe4b2a),
	.w6(32'h3a719a6c),
	.w7(32'h3bebd5eb),
	.w8(32'h3c7e6760),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabec91),
	.w1(32'h3c24cb7c),
	.w2(32'h3adfe699),
	.w3(32'h3938f97e),
	.w4(32'h3b48650d),
	.w5(32'hbbb642e5),
	.w6(32'h3c08eac5),
	.w7(32'h3b90abb0),
	.w8(32'h39e42d6e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a082b),
	.w1(32'h3c6110e6),
	.w2(32'hbc90940d),
	.w3(32'hbc5221ce),
	.w4(32'hbc48e3ae),
	.w5(32'hbcfe174b),
	.w6(32'h3c43cc82),
	.w7(32'h3c611fb7),
	.w8(32'hbb7e341d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbeb7e2),
	.w1(32'h3be69055),
	.w2(32'h3ca62e65),
	.w3(32'hbc6d835f),
	.w4(32'h3c35248a),
	.w5(32'h3bc68ab9),
	.w6(32'hbc091864),
	.w7(32'hbb730990),
	.w8(32'h3bb4cc24),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97e2e2),
	.w1(32'h3cee68d2),
	.w2(32'h3d1f30b5),
	.w3(32'hbc2a5a3a),
	.w4(32'h3d09b3fb),
	.w5(32'h3c7ec2ee),
	.w6(32'hbc952388),
	.w7(32'h3cc91e72),
	.w8(32'h3c2f7ec4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6633f),
	.w1(32'h3c4268b4),
	.w2(32'h3bb1da8f),
	.w3(32'hbc020141),
	.w4(32'h3c058802),
	.w5(32'h39916a47),
	.w6(32'h3be3ebdd),
	.w7(32'h3b41b160),
	.w8(32'h3b9f557d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97623b),
	.w1(32'h3bc99069),
	.w2(32'h3c4dee89),
	.w3(32'h3a926d4b),
	.w4(32'h3b57f049),
	.w5(32'hbc462f2f),
	.w6(32'hbc824e54),
	.w7(32'h3b4e2cc4),
	.w8(32'h3a676c4c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba99c1b),
	.w1(32'h3cbf6bc2),
	.w2(32'h3cb153b8),
	.w3(32'hbcbb81b4),
	.w4(32'h3b354203),
	.w5(32'hbb5c0995),
	.w6(32'h3bfcae71),
	.w7(32'h3cb09061),
	.w8(32'h3cd742b8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c5d87),
	.w1(32'hbab017c4),
	.w2(32'h3cf4cae9),
	.w3(32'h3b0ad8b3),
	.w4(32'h3bceae05),
	.w5(32'h3cae6865),
	.w6(32'hbb501db1),
	.w7(32'hbbd57117),
	.w8(32'h3bbdefe6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd23100),
	.w1(32'h3c18ed5d),
	.w2(32'h3b1058b1),
	.w3(32'hbc9ace38),
	.w4(32'hbbdac3d1),
	.w5(32'hbc7a73fa),
	.w6(32'h3c1cb55c),
	.w7(32'hbb421b47),
	.w8(32'h3b3b3aa7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8f18),
	.w1(32'h3a3782a7),
	.w2(32'h3b723adb),
	.w3(32'h3c771a84),
	.w4(32'h3be4e1ea),
	.w5(32'h3cb7bcf7),
	.w6(32'h3c43282d),
	.w7(32'h3bd60873),
	.w8(32'h3b85b066),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92bcc7),
	.w1(32'h3ac264ee),
	.w2(32'h3b2d410c),
	.w3(32'h3d02f960),
	.w4(32'hbb6fcc24),
	.w5(32'hbab00932),
	.w6(32'h3b82990a),
	.w7(32'hbb0d665b),
	.w8(32'h3ad6ead6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e3a8a),
	.w1(32'h3bc36cc4),
	.w2(32'hbcb3ed9a),
	.w3(32'hbb97ee5f),
	.w4(32'hbb085274),
	.w5(32'hbb9db25f),
	.w6(32'h3c5e90d8),
	.w7(32'h3a57bcd0),
	.w8(32'hbba71487),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd0b38),
	.w1(32'hbc2b5e50),
	.w2(32'hbc803ba5),
	.w3(32'h3c6cc8f1),
	.w4(32'hbbd0c231),
	.w5(32'hba0a5ee3),
	.w6(32'h3a41f3c0),
	.w7(32'hbc14eb6a),
	.w8(32'hbb7163f7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f2a47),
	.w1(32'h3c17a0bc),
	.w2(32'h3cc3106d),
	.w3(32'h3c713f2c),
	.w4(32'h3c12eb28),
	.w5(32'h3c862118),
	.w6(32'hbb355eb1),
	.w7(32'h3bbd9b1a),
	.w8(32'h3c6868f0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62554),
	.w1(32'hba144f35),
	.w2(32'h3bb9a123),
	.w3(32'hbbc78fd3),
	.w4(32'h3b67d946),
	.w5(32'h3c4c20d6),
	.w6(32'hbb289e2a),
	.w7(32'h3b1c0a33),
	.w8(32'h3b87a0d1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b715e),
	.w1(32'hbcd1b134),
	.w2(32'hbcb9666a),
	.w3(32'h3b577b0b),
	.w4(32'hbb0de95b),
	.w5(32'hbba9c102),
	.w6(32'hbb2128de),
	.w7(32'hbc4bb606),
	.w8(32'hbc0608bb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc6ea9),
	.w1(32'h3b2ae0f9),
	.w2(32'h3c0f109b),
	.w3(32'h3b5ea5da),
	.w4(32'h3b9bf4fe),
	.w5(32'hb9ae0856),
	.w6(32'h3c632ffe),
	.w7(32'h3b302d9d),
	.w8(32'h3b53a5cc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52537),
	.w1(32'h393c4a8d),
	.w2(32'h3acfb2e4),
	.w3(32'hbb315372),
	.w4(32'h3a7dced9),
	.w5(32'hbac7e0f1),
	.w6(32'hbb21184f),
	.w7(32'h39facdad),
	.w8(32'hbb4cee26),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf00657),
	.w1(32'hbbe49366),
	.w2(32'hbb6378e3),
	.w3(32'hbbbdcd78),
	.w4(32'h3b2c80be),
	.w5(32'h3b963ab6),
	.w6(32'hbb6e1537),
	.w7(32'hbc0b7fce),
	.w8(32'h39e60def),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c4dd4),
	.w1(32'hbbd00f6f),
	.w2(32'h3ba60805),
	.w3(32'hbb8e25cf),
	.w4(32'h3a81beb6),
	.w5(32'hbb28f248),
	.w6(32'hbb6fdd19),
	.w7(32'hb96462ad),
	.w8(32'hbb1e047b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfde1c6),
	.w1(32'hbb4d7638),
	.w2(32'hbb165505),
	.w3(32'hbc4b509f),
	.w4(32'hbb6a4f2b),
	.w5(32'hbb958477),
	.w6(32'hba2b0331),
	.w7(32'hbb17b839),
	.w8(32'hbb45ce3e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87589c),
	.w1(32'hba950a23),
	.w2(32'hbc2d1579),
	.w3(32'h3a85d03b),
	.w4(32'h3a3cd970),
	.w5(32'hbc1f6f95),
	.w6(32'h3b865123),
	.w7(32'hbc332c84),
	.w8(32'hbb38dd8a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeac1a),
	.w1(32'h3adbae8f),
	.w2(32'h3a15c477),
	.w3(32'hbb0c3ed9),
	.w4(32'hbc39baac),
	.w5(32'hbcc4d69e),
	.w6(32'hba39c5d9),
	.w7(32'h3b4c31e0),
	.w8(32'hba71867e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c1a86),
	.w1(32'hbac15463),
	.w2(32'hbb2478bb),
	.w3(32'hbcca6779),
	.w4(32'hbadd8d75),
	.w5(32'hbc5bddca),
	.w6(32'h3b57e423),
	.w7(32'h3b81e652),
	.w8(32'h3b19aec6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2649da),
	.w1(32'hbb908ed9),
	.w2(32'h3bec1ae8),
	.w3(32'hbb8e0495),
	.w4(32'h3c3da1ed),
	.w5(32'h3c5d3cb2),
	.w6(32'h39b74377),
	.w7(32'h3b94d3d4),
	.w8(32'h3bcd9b15),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b823c),
	.w1(32'hb7a92295),
	.w2(32'h3ae85934),
	.w3(32'hbb26072a),
	.w4(32'hbbb81338),
	.w5(32'hbbaa9a92),
	.w6(32'h3b95327b),
	.w7(32'h3bbc0730),
	.w8(32'h3ae1d715),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16e3e),
	.w1(32'h3b97a0b9),
	.w2(32'h395a7527),
	.w3(32'hbbfdf87a),
	.w4(32'hbb84dfe5),
	.w5(32'hbc4e7921),
	.w6(32'h3bda1df6),
	.w7(32'hbad8325b),
	.w8(32'hbbd11baa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf23f0),
	.w1(32'h3c64f292),
	.w2(32'h3b86033f),
	.w3(32'hbc72a91e),
	.w4(32'h3ab79808),
	.w5(32'hbc1ebd4b),
	.w6(32'h3c6cfe7a),
	.w7(32'h3c49f0aa),
	.w8(32'h3aaf91c2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18f3c2),
	.w1(32'h3b260bf2),
	.w2(32'h3c9259da),
	.w3(32'hbbb9cfcf),
	.w4(32'h3c6b5891),
	.w5(32'h3c0d1e41),
	.w6(32'h38858a9e),
	.w7(32'h3b30a71c),
	.w8(32'h3b488428),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56c4d6),
	.w1(32'h3bae559a),
	.w2(32'h3bca1736),
	.w3(32'hb9c4379b),
	.w4(32'h3ba628c9),
	.w5(32'h3bf1a20f),
	.w6(32'hbbb21381),
	.w7(32'hbbd1c7a9),
	.w8(32'h3ba5c998),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9097bb),
	.w1(32'h3c07e80f),
	.w2(32'hbcbcd906),
	.w3(32'h3adbd399),
	.w4(32'hbbd3c552),
	.w5(32'hbcad4e57),
	.w6(32'h3c694957),
	.w7(32'hbc423e57),
	.w8(32'hbc26eb3f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc028308),
	.w1(32'h3b2ed20a),
	.w2(32'h3c5791d7),
	.w3(32'hbc855370),
	.w4(32'hba36a4f4),
	.w5(32'h3bec64e2),
	.w6(32'hbc5c3e31),
	.w7(32'hbb2d528d),
	.w8(32'h3b5c0175),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35772c),
	.w1(32'h3ba1c486),
	.w2(32'h3bb4106e),
	.w3(32'h3b40a8e3),
	.w4(32'hbbae0097),
	.w5(32'hbbbac42c),
	.w6(32'hbc535c20),
	.w7(32'hbbd8df31),
	.w8(32'hbac3f887),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d85df),
	.w1(32'hb8ecb1d2),
	.w2(32'hbc0b5a95),
	.w3(32'hbbd1826a),
	.w4(32'h3c136f6c),
	.w5(32'h3b7b691d),
	.w6(32'h3a1a1539),
	.w7(32'hbbf36020),
	.w8(32'h3ba1cb6c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00bcbc),
	.w1(32'hbba19c6a),
	.w2(32'hbc0601fb),
	.w3(32'h3bc6d105),
	.w4(32'hbbb0fa1e),
	.w5(32'hbc1227f0),
	.w6(32'h3c1d622c),
	.w7(32'hbb8e11e8),
	.w8(32'h3b78be8e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e515a),
	.w1(32'hbb9b0365),
	.w2(32'h3c64db37),
	.w3(32'hb78a25fa),
	.w4(32'h3c1105f0),
	.w5(32'h3be5deae),
	.w6(32'hbc8e8a1e),
	.w7(32'h3c14074e),
	.w8(32'h3c25e88c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380874),
	.w1(32'h3b0b3aa0),
	.w2(32'hbae74dec),
	.w3(32'h3b487195),
	.w4(32'h3c14438c),
	.w5(32'h3ba2bccf),
	.w6(32'hba5b5c2b),
	.w7(32'h3b8f6d79),
	.w8(32'h3b7771fe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52acb8),
	.w1(32'hbca8cae2),
	.w2(32'hbd22fdbc),
	.w3(32'hba8bd33e),
	.w4(32'hbca5e6a1),
	.w5(32'hbc7fe6af),
	.w6(32'h3b2bf4fb),
	.w7(32'hbc963f48),
	.w8(32'hbd008247),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f74b7),
	.w1(32'hbc1c0917),
	.w2(32'hbc7bf44a),
	.w3(32'h3c408cba),
	.w4(32'hbc5b2202),
	.w5(32'hbc32ed9f),
	.w6(32'h39d7f257),
	.w7(32'hbc6603bc),
	.w8(32'hbc1a5945),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c68b),
	.w1(32'hba89905e),
	.w2(32'h3a1f9430),
	.w3(32'hbb44c6e9),
	.w4(32'h3b41a8b7),
	.w5(32'hbaa7d990),
	.w6(32'hbb1066c1),
	.w7(32'h3aa86858),
	.w8(32'h3a9e66b7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96beda2),
	.w1(32'h3bad7245),
	.w2(32'h3cd73f29),
	.w3(32'h3a96ac67),
	.w4(32'h3c50c880),
	.w5(32'h3c81c797),
	.w6(32'hbb8e9abd),
	.w7(32'h3b97b15f),
	.w8(32'h3af17c35),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a46ae),
	.w1(32'hbc0f7be9),
	.w2(32'hbc9f73b2),
	.w3(32'h3bffbc9b),
	.w4(32'hbc9d305a),
	.w5(32'hbc2bad89),
	.w6(32'h3bc2a7b1),
	.w7(32'hbbba3857),
	.w8(32'hbb8b2875),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a5859),
	.w1(32'hbc4e3815),
	.w2(32'h3ae8c1ce),
	.w3(32'hbc862cdb),
	.w4(32'hb9ec7fa0),
	.w5(32'hbb521a52),
	.w6(32'hbc4e46af),
	.w7(32'hbc64c15d),
	.w8(32'hba92d3d9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bb709),
	.w1(32'h3bda3b9d),
	.w2(32'hbbc35096),
	.w3(32'hbc77eb67),
	.w4(32'h3c0f5829),
	.w5(32'h3b46ca76),
	.w6(32'h3c9bad61),
	.w7(32'h3b14f9e6),
	.w8(32'h3c36431d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35218b),
	.w1(32'h3b78d188),
	.w2(32'h3c1c9360),
	.w3(32'h3cabe8fc),
	.w4(32'h3be1a41a),
	.w5(32'h3c08b4b9),
	.w6(32'h3bdf3d20),
	.w7(32'h3bcd8606),
	.w8(32'h3ae5b91b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c6286),
	.w1(32'h3b07a244),
	.w2(32'h3ad4cc7f),
	.w3(32'h39caae18),
	.w4(32'h3be4e259),
	.w5(32'h3bc06e30),
	.w6(32'h3946dae6),
	.w7(32'h3a97ae17),
	.w8(32'h3b6536d7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9710863),
	.w1(32'hba068f86),
	.w2(32'h3b662365),
	.w3(32'h3b291d1c),
	.w4(32'hbbc28a5e),
	.w5(32'h3bc74ea4),
	.w6(32'h3afbaa5c),
	.w7(32'h3b8eb9a6),
	.w8(32'hbac708f3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13de95),
	.w1(32'hbc62eadc),
	.w2(32'h3b47c0aa),
	.w3(32'hbbbca94e),
	.w4(32'h3cbf1ba0),
	.w5(32'h3ccadbb6),
	.w6(32'hbc93f2b6),
	.w7(32'hbb9fa5e8),
	.w8(32'h3c1d8b9f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4985d1),
	.w1(32'h3cb22abc),
	.w2(32'h3c5893ff),
	.w3(32'h3b73e903),
	.w4(32'hbb2ede77),
	.w5(32'hbc8f04ad),
	.w6(32'h3ca9562a),
	.w7(32'h3c687d1a),
	.w8(32'hba81b8cd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06d2bc),
	.w1(32'h3bfd1762),
	.w2(32'h3c1e0e94),
	.w3(32'hbc4a89ca),
	.w4(32'h3c0a5d9b),
	.w5(32'h3c9338e9),
	.w6(32'hbb3883a6),
	.w7(32'hbbc7130c),
	.w8(32'h3b2d76db),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8178a),
	.w1(32'hba1b3dc0),
	.w2(32'h3bcf7273),
	.w3(32'h3aaec7f5),
	.w4(32'h3b0b1fba),
	.w5(32'h3b2ced35),
	.w6(32'h3c196d03),
	.w7(32'h3c03c545),
	.w8(32'hbc1fdc80),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c5d7),
	.w1(32'hbc352e6b),
	.w2(32'hbb9a1315),
	.w3(32'h3ba3a195),
	.w4(32'hbc00955c),
	.w5(32'hbb653db7),
	.w6(32'hbc21386c),
	.w7(32'hbc2b5779),
	.w8(32'hba390c81),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ff43),
	.w1(32'h3c43a74f),
	.w2(32'h3c12b2e2),
	.w3(32'hbc3c353f),
	.w4(32'hb9847626),
	.w5(32'h3a9fcba2),
	.w6(32'hbb404a6d),
	.w7(32'h3b91525d),
	.w8(32'h3b9cb700),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c099b54),
	.w1(32'h3bf0c40d),
	.w2(32'h3c95c389),
	.w3(32'hbaa3dadc),
	.w4(32'h3ab65b81),
	.w5(32'h3c0221c3),
	.w6(32'hbb7ade97),
	.w7(32'h3ad86589),
	.w8(32'hbaabe634),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e1c98),
	.w1(32'hbbf8c585),
	.w2(32'hbd22264b),
	.w3(32'hbc0c4424),
	.w4(32'hbc610682),
	.w5(32'hbbcf0bb3),
	.w6(32'h3c807607),
	.w7(32'hbca36135),
	.w8(32'hbc342ddb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3407cc),
	.w1(32'hbc8c3163),
	.w2(32'h39861766),
	.w3(32'h3c7ec8b7),
	.w4(32'hbc4be312),
	.w5(32'hbb65b942),
	.w6(32'hbcefacd6),
	.w7(32'hbc849fc3),
	.w8(32'hbc608043),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89a155),
	.w1(32'hbc8c5490),
	.w2(32'hbcaffca4),
	.w3(32'hbc878bbe),
	.w4(32'hbc0094af),
	.w5(32'hbc1a3c6b),
	.w6(32'hbc945f57),
	.w7(32'hbcca4586),
	.w8(32'hbc51b9ca),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8e21),
	.w1(32'hbb8a829e),
	.w2(32'hbc8b5263),
	.w3(32'h3c55148b),
	.w4(32'hbc8b60f0),
	.w5(32'hbc3c8bc5),
	.w6(32'h3b9e01f6),
	.w7(32'hba085c50),
	.w8(32'hbc18def9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8306e),
	.w1(32'hbba454b0),
	.w2(32'hbc4006dd),
	.w3(32'h3bbd457f),
	.w4(32'hbc0df773),
	.w5(32'hbc394b27),
	.w6(32'hbbcb3975),
	.w7(32'hbc305be2),
	.w8(32'hbb07a856),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b834740),
	.w1(32'hbb95be23),
	.w2(32'hbab5eb62),
	.w3(32'hbb3838aa),
	.w4(32'hbba92015),
	.w5(32'hbb3262c6),
	.w6(32'hbc1d7a75),
	.w7(32'hba80dcff),
	.w8(32'h3bf4da26),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83d96c),
	.w1(32'hbb828e56),
	.w2(32'h3c5b9790),
	.w3(32'h3b28170a),
	.w4(32'hb7a03ee7),
	.w5(32'h3c40d911),
	.w6(32'h39832a67),
	.w7(32'h3ae3a061),
	.w8(32'h3c04481e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bee0f),
	.w1(32'h3b339795),
	.w2(32'h3c47765e),
	.w3(32'hbb7243fd),
	.w4(32'hbbfd1a87),
	.w5(32'hbc4c58f0),
	.w6(32'hbb993c09),
	.w7(32'h3be226d7),
	.w8(32'h3b516f79),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbb6c2),
	.w1(32'h39870882),
	.w2(32'h3c345a0e),
	.w3(32'hbca74189),
	.w4(32'h3c25f527),
	.w5(32'h3c36692d),
	.w6(32'hba987c2f),
	.w7(32'h3ba10a52),
	.w8(32'h3b8b610d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba30c5),
	.w1(32'h3c2daf37),
	.w2(32'hba92cfe0),
	.w3(32'h3c5e266b),
	.w4(32'h3ba40ca3),
	.w5(32'hbbdfb972),
	.w6(32'h3b220270),
	.w7(32'h3b8b858a),
	.w8(32'hbb100371),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f986),
	.w1(32'h3c1e2b2a),
	.w2(32'h3d5fb9a8),
	.w3(32'hbbadafea),
	.w4(32'h3ce09d09),
	.w5(32'h3d4bca1b),
	.w6(32'hbbb7ba56),
	.w7(32'h3b15b956),
	.w8(32'h3d0ac9af),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7c8e5b),
	.w1(32'h3bf001dc),
	.w2(32'h3b849153),
	.w3(32'h3c87b00f),
	.w4(32'h3b83d7a3),
	.w5(32'h3b8c4e14),
	.w6(32'h39a71db2),
	.w7(32'h3b61b32e),
	.w8(32'h3bd7229f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b0d24),
	.w1(32'hbbbf9b19),
	.w2(32'hbc960799),
	.w3(32'hbc3eb7f4),
	.w4(32'hbb7cbd13),
	.w5(32'hbc0c17b4),
	.w6(32'h3bfc75bb),
	.w7(32'h3b885d0e),
	.w8(32'hbbaca9ba),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60396b),
	.w1(32'hbc4cc574),
	.w2(32'hbc8a3d53),
	.w3(32'hbb2ba892),
	.w4(32'hbb77a3ae),
	.w5(32'hbb753a84),
	.w6(32'hbaebb60b),
	.w7(32'hbb6935be),
	.w8(32'hbbbe7441),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f298f),
	.w1(32'h3a82dd0b),
	.w2(32'hbbc76c16),
	.w3(32'hba902b9e),
	.w4(32'hbc7c9a80),
	.w5(32'hbcf64c9d),
	.w6(32'hbb814719),
	.w7(32'h3ab01b52),
	.w8(32'hbb92bad0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd065a8),
	.w1(32'hbc8f0855),
	.w2(32'hbcbd6864),
	.w3(32'hbcebcdff),
	.w4(32'hba4fd489),
	.w5(32'h3aed5f0a),
	.w6(32'hbb92a724),
	.w7(32'hbc2a15c2),
	.w8(32'hbc8dba0a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64f787),
	.w1(32'hba6df5a0),
	.w2(32'h3caec275),
	.w3(32'h3b93f3be),
	.w4(32'h3bf52d2b),
	.w5(32'h3cc11b0c),
	.w6(32'hbb88fd36),
	.w7(32'h3b006db5),
	.w8(32'h3c3282c8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c562d95),
	.w1(32'h3b0b60e2),
	.w2(32'h3817aeda),
	.w3(32'h3c029c1a),
	.w4(32'h3baaab8d),
	.w5(32'h3b570965),
	.w6(32'h3a7c7091),
	.w7(32'hba44a350),
	.w8(32'h3b3e8962),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a3144),
	.w1(32'h3a8c3975),
	.w2(32'h3c50ae2e),
	.w3(32'h39f1d5a7),
	.w4(32'h3c2fecec),
	.w5(32'h3c5f6a41),
	.w6(32'h3b3b32b8),
	.w7(32'h3b4d891b),
	.w8(32'h3a9edfb6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9dab9),
	.w1(32'h3afb93d6),
	.w2(32'h3b4eec56),
	.w3(32'h3abb3ea0),
	.w4(32'hbb8a0f4e),
	.w5(32'hb9b2f2e7),
	.w6(32'hbadb1bae),
	.w7(32'h3adbc3f4),
	.w8(32'h3b4db289),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be429a2),
	.w1(32'h3c4576f2),
	.w2(32'h3c261f35),
	.w3(32'h3b74d199),
	.w4(32'h3bee5751),
	.w5(32'h3af91813),
	.w6(32'h3bec15b5),
	.w7(32'h3c43b789),
	.w8(32'h3bbdfc40),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba817749),
	.w1(32'h3c09f153),
	.w2(32'hbc7abcf0),
	.w3(32'hbb5d1ca9),
	.w4(32'h3b41b2d6),
	.w5(32'h3bac39a3),
	.w6(32'h3bff4d0e),
	.w7(32'hbc5ac00c),
	.w8(32'hbc23a31c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1008b),
	.w1(32'hbc5d903e),
	.w2(32'hbcb5f518),
	.w3(32'hbb1727d0),
	.w4(32'hbc34944e),
	.w5(32'hbc537742),
	.w6(32'h39835fbd),
	.w7(32'hbc0d8077),
	.w8(32'hbc107e35),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd81974),
	.w1(32'h3cc97018),
	.w2(32'h3d5629d2),
	.w3(32'hbad041fd),
	.w4(32'h3cd98fa8),
	.w5(32'h3c865256),
	.w6(32'hbb64b681),
	.w7(32'h3c4c0632),
	.w8(32'h3c670583),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac023f),
	.w1(32'hbb967a83),
	.w2(32'h3cd0cfce),
	.w3(32'hbbbf52ab),
	.w4(32'h3c0bb5e9),
	.w5(32'h3cacfd88),
	.w6(32'hbb701b70),
	.w7(32'hbb38202c),
	.w8(32'h3be0ec96),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75f92c),
	.w1(32'h374d6a71),
	.w2(32'h3aec66fe),
	.w3(32'hbc2781a2),
	.w4(32'hbb5f1c2a),
	.w5(32'hbbc39183),
	.w6(32'hbb2894d3),
	.w7(32'h3baff7f0),
	.w8(32'hbb5f6d82),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938d858),
	.w1(32'hbb832623),
	.w2(32'hbb4ea0bb),
	.w3(32'hbc0aaef9),
	.w4(32'hb9a7d1b6),
	.w5(32'hbb87caee),
	.w6(32'hbc118060),
	.w7(32'hbb91ff4d),
	.w8(32'hbb6fd801),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8121c99),
	.w1(32'hbbc9ac4a),
	.w2(32'hbc04f78f),
	.w3(32'h3b1771a1),
	.w4(32'h3c2a5558),
	.w5(32'hba12c493),
	.w6(32'h3aec2db3),
	.w7(32'hbb687beb),
	.w8(32'hbc39e2ec),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce0034),
	.w1(32'hbb0e8706),
	.w2(32'hbbc338bb),
	.w3(32'hbc2f72ae),
	.w4(32'h3b89e644),
	.w5(32'h3c83f0d4),
	.w6(32'h3be22c3c),
	.w7(32'hba37d6f1),
	.w8(32'hba3f5be4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59c4e6),
	.w1(32'h3bcdadb3),
	.w2(32'h3bbc5191),
	.w3(32'h3c34bc4a),
	.w4(32'h3b49d060),
	.w5(32'h3c28de01),
	.w6(32'hbb46284b),
	.w7(32'hbb65c103),
	.w8(32'h3ab50b6d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c0e79),
	.w1(32'hbd3f1ff5),
	.w2(32'hbd1b0367),
	.w3(32'h3b7c367f),
	.w4(32'hbc892082),
	.w5(32'hbb661718),
	.w6(32'hbc0a9001),
	.w7(32'hbd06fc4f),
	.w8(32'hbc9f6f01),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93563e),
	.w1(32'hbbd4779a),
	.w2(32'h3c60ebab),
	.w3(32'hb90fdcda),
	.w4(32'hbb6e9d4c),
	.w5(32'hbc0ee4a0),
	.w6(32'hbc3bafb5),
	.w7(32'h3c5cde3f),
	.w8(32'h3be4fc02),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa10ef2),
	.w1(32'h3c6af68c),
	.w2(32'h3c323e65),
	.w3(32'hbad00ea2),
	.w4(32'h3c75b40b),
	.w5(32'h3c0156ac),
	.w6(32'h3c351997),
	.w7(32'h3c00e56c),
	.w8(32'h3c4b18ed),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f0bc3),
	.w1(32'hbc037897),
	.w2(32'hbd15a89f),
	.w3(32'h3bb8d8d7),
	.w4(32'hbbb40935),
	.w5(32'hbc5dce58),
	.w6(32'h3bb49c6e),
	.w7(32'hbc091bb3),
	.w8(32'hbc996fa3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9d7b8),
	.w1(32'hba6697fe),
	.w2(32'hbb70dca4),
	.w3(32'h3b276ee1),
	.w4(32'h3ba907fb),
	.w5(32'hbbf1f28f),
	.w6(32'hbc8f77b0),
	.w7(32'hbbdbadd6),
	.w8(32'hbbb511e1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f078),
	.w1(32'h3bfa1c71),
	.w2(32'h3b8c4d61),
	.w3(32'hbb94d1a4),
	.w4(32'h3b8a645b),
	.w5(32'h3a4b56f6),
	.w6(32'h3c939da5),
	.w7(32'h3c6b9d5e),
	.w8(32'h3c27575a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef8fa),
	.w1(32'h3b27def6),
	.w2(32'hba9020e1),
	.w3(32'h3b2e5c93),
	.w4(32'h3bc6caf6),
	.w5(32'h3bce7e2e),
	.w6(32'h3961b558),
	.w7(32'h3a64306e),
	.w8(32'h3bbfa4fa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee24bf),
	.w1(32'h3ba2c8b1),
	.w2(32'h3c1ba0e6),
	.w3(32'h3bebeae6),
	.w4(32'h3b1cf904),
	.w5(32'h3be0af7f),
	.w6(32'hbbb1d141),
	.w7(32'h39d5415b),
	.w8(32'h3c17a51d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dab16),
	.w1(32'h3bb7bee4),
	.w2(32'h3bbb8130),
	.w3(32'hbb079f80),
	.w4(32'h3b23ccc2),
	.w5(32'hbb78ce0f),
	.w6(32'h3af0bc7a),
	.w7(32'h3aa898c7),
	.w8(32'hba1b1e53),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9300a82),
	.w1(32'hbb889ea0),
	.w2(32'h3abd7f60),
	.w3(32'hbbd50256),
	.w4(32'hbbabef52),
	.w5(32'h3c14075e),
	.w6(32'hbb685400),
	.w7(32'hbbb3c94a),
	.w8(32'h3b64102a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb445a55),
	.w1(32'h3d30e87c),
	.w2(32'h3d782ee4),
	.w3(32'h3adc3504),
	.w4(32'h3c9d231e),
	.w5(32'h3bbc7b4d),
	.w6(32'h3b6139ce),
	.w7(32'h3cdac216),
	.w8(32'h3ccd7408),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c907655),
	.w1(32'hbbdd5f71),
	.w2(32'hbc05e192),
	.w3(32'h3ac51822),
	.w4(32'hbb29a893),
	.w5(32'h3ad2d02d),
	.w6(32'h3b4b235c),
	.w7(32'h3ae111b7),
	.w8(32'h39b0a48b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f467),
	.w1(32'hb8f1e0be),
	.w2(32'hbb413e4b),
	.w3(32'h3adf7dd6),
	.w4(32'h3b81918d),
	.w5(32'h3b8c5d1c),
	.w6(32'h38e61de5),
	.w7(32'hb985a8a8),
	.w8(32'h3b89fbe9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadabbb0),
	.w1(32'hba1c172f),
	.w2(32'h3c289093),
	.w3(32'h3be0909a),
	.w4(32'hbbaa80b7),
	.w5(32'hbb385540),
	.w6(32'hbb55be7d),
	.w7(32'h3ac3996a),
	.w8(32'h3a838c88),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab02b7),
	.w1(32'hbb192213),
	.w2(32'h3c02fb69),
	.w3(32'hbbe71086),
	.w4(32'h3bb38abb),
	.w5(32'h3c057317),
	.w6(32'hbaf9bfd3),
	.w7(32'h3aaa2e82),
	.w8(32'h3bd596a5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfde7cd),
	.w1(32'h3b2ac8f4),
	.w2(32'h3c9106d7),
	.w3(32'h3b1a428b),
	.w4(32'h3ab78af3),
	.w5(32'h3b021673),
	.w6(32'hbc690e01),
	.w7(32'hbc44792b),
	.w8(32'h3bbb05cd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd43ddc),
	.w1(32'hbacbe526),
	.w2(32'h3bf0d5f7),
	.w3(32'h3abdbca8),
	.w4(32'h3982a016),
	.w5(32'hbb89d03a),
	.w6(32'hbc47eb8e),
	.w7(32'hbacdd2bb),
	.w8(32'hba98daa5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc61869),
	.w1(32'h3c17afb7),
	.w2(32'h3c63acdf),
	.w3(32'hbc9db121),
	.w4(32'hbae63ed8),
	.w5(32'hbb22476c),
	.w6(32'h3c1eb5fd),
	.w7(32'h3bb42eb5),
	.w8(32'hb9707543),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7092fb7),
	.w1(32'hbca8ed09),
	.w2(32'hbc72474c),
	.w3(32'h3b665553),
	.w4(32'hbbd555f4),
	.w5(32'hbbf93085),
	.w6(32'hbb78840c),
	.w7(32'hbc527479),
	.w8(32'hbc4c2836),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9afb2a),
	.w1(32'h3b65ec70),
	.w2(32'h3a960436),
	.w3(32'hbc76e661),
	.w4(32'h38933d9d),
	.w5(32'hbb6bfe40),
	.w6(32'h3b4c3b2d),
	.w7(32'hb835417e),
	.w8(32'h3a9baf9c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f2a0),
	.w1(32'hbc1443e3),
	.w2(32'hbbd85d5b),
	.w3(32'hbb4bfd88),
	.w4(32'hbb6a9645),
	.w5(32'hbba0ef80),
	.w6(32'h39d5e752),
	.w7(32'hbb4a806a),
	.w8(32'hbbd3723a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c665c),
	.w1(32'hbc9386af),
	.w2(32'hbc5db3de),
	.w3(32'h38b56942),
	.w4(32'hbc322a2c),
	.w5(32'hbc67d5be),
	.w6(32'hbcd23ce5),
	.w7(32'hbd0ad6b0),
	.w8(32'hbc455d37),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba911093),
	.w1(32'h3c1f81d5),
	.w2(32'h3d06235a),
	.w3(32'hbad1eeb6),
	.w4(32'h3c9d57f2),
	.w5(32'h3ccdb596),
	.w6(32'h39d124ed),
	.w7(32'h3c8d98e5),
	.w8(32'h3cc89242),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51659b),
	.w1(32'hba7cd67f),
	.w2(32'hbb97b6e0),
	.w3(32'h3bfc0ee3),
	.w4(32'hbb3afd0f),
	.w5(32'hbbd02c6c),
	.w6(32'hbb6f63c0),
	.w7(32'hbbc31fa3),
	.w8(32'hb9dca0cd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe4270),
	.w1(32'hbb7f6c6a),
	.w2(32'h3b1eca40),
	.w3(32'hb9a18f7c),
	.w4(32'h3b4aadeb),
	.w5(32'h3b8f949e),
	.w6(32'hbb9b8358),
	.w7(32'hb9395a65),
	.w8(32'hbacbcf8e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule