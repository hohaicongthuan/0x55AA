module layer_8_featuremap_208(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fd4ca),
	.w1(32'h3c9b5b84),
	.w2(32'h3c786a8a),
	.w3(32'hbb004671),
	.w4(32'h3b8fe451),
	.w5(32'h3b2a259a),
	.w6(32'h3bde1e94),
	.w7(32'h3c2b30ab),
	.w8(32'h3c9ec52d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f0359),
	.w1(32'h3c0360a2),
	.w2(32'h3abdd59b),
	.w3(32'hbcbfd51c),
	.w4(32'h3aa77bfb),
	.w5(32'h3ad7bea5),
	.w6(32'h3ae07ff5),
	.w7(32'h3a676174),
	.w8(32'hbb431b2c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2449b5),
	.w1(32'h3bb99638),
	.w2(32'hbb98033c),
	.w3(32'hbc308622),
	.w4(32'hbbd60e40),
	.w5(32'hbc1f9ef8),
	.w6(32'hbbf90957),
	.w7(32'hbb47d624),
	.w8(32'hbb1c5ba8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5afd7c),
	.w1(32'h3a86047b),
	.w2(32'h3b5b592c),
	.w3(32'hbadc9df3),
	.w4(32'hb9998071),
	.w5(32'h3b1b4003),
	.w6(32'h3a569ada),
	.w7(32'h3b98f0cd),
	.w8(32'hb99102af),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cab45),
	.w1(32'hbb86d83b),
	.w2(32'h3bd9563a),
	.w3(32'h3b63f0eb),
	.w4(32'h3a1f9d8b),
	.w5(32'h3bfad991),
	.w6(32'hba22074a),
	.w7(32'hba48e600),
	.w8(32'h3b907791),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24d804),
	.w1(32'h3c63571c),
	.w2(32'hbb088a20),
	.w3(32'hbb8d0587),
	.w4(32'h3b30c9de),
	.w5(32'hbb741c57),
	.w6(32'h3c778434),
	.w7(32'h3b8ba854),
	.w8(32'hbc2e74a3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6110e2),
	.w1(32'hbc25a169),
	.w2(32'h3abc41ad),
	.w3(32'h3c857c4d),
	.w4(32'hbbd43335),
	.w5(32'hb9ab9b91),
	.w6(32'hbc018bfb),
	.w7(32'hbb883c47),
	.w8(32'h39dcc618),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93cbdd),
	.w1(32'h3c6abacc),
	.w2(32'hbc7165f4),
	.w3(32'hbbc3f433),
	.w4(32'h3b24517d),
	.w5(32'hbbf95d74),
	.w6(32'h3c4a7581),
	.w7(32'hbba4d1d6),
	.w8(32'h3ba80e10),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3040),
	.w1(32'hbb2f143f),
	.w2(32'h3c618bba),
	.w3(32'hbbe71568),
	.w4(32'h3b07012a),
	.w5(32'h3c4687b0),
	.w6(32'hbb3627a0),
	.w7(32'h3b80db32),
	.w8(32'h3bdbf71b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf93b7a),
	.w1(32'hbbb7b9ec),
	.w2(32'hbce88858),
	.w3(32'hbc3071fc),
	.w4(32'hbad56b2d),
	.w5(32'hbc4a9bac),
	.w6(32'h3b809dda),
	.w7(32'hbc5735ff),
	.w8(32'hbbf43c95),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc953531),
	.w1(32'h3c5ac0eb),
	.w2(32'hba5dbf7a),
	.w3(32'hbbd27450),
	.w4(32'h3a7de85f),
	.w5(32'hbbb59d97),
	.w6(32'h39ee6b2a),
	.w7(32'h3af5b365),
	.w8(32'h3bf0b79e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15c157),
	.w1(32'h3a517fab),
	.w2(32'h3bb480a2),
	.w3(32'hbc122fb1),
	.w4(32'h3523df9c),
	.w5(32'h3bc7ec76),
	.w6(32'h3aafc089),
	.w7(32'hba961461),
	.w8(32'h39de863c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71bf4f),
	.w1(32'hbb704e99),
	.w2(32'hbc689cc0),
	.w3(32'h3c71d370),
	.w4(32'h3b0e457c),
	.w5(32'hbbe325f6),
	.w6(32'hbaf52b95),
	.w7(32'hbb8b6a7b),
	.w8(32'hbbc4a855),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3a006),
	.w1(32'h3c3b3975),
	.w2(32'h3b3c22bc),
	.w3(32'hbacaab12),
	.w4(32'hbab20bc5),
	.w5(32'hbb4ba7f5),
	.w6(32'h3c2ced84),
	.w7(32'h3b5e7ada),
	.w8(32'h3c00029a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dfefb),
	.w1(32'hbb5f1654),
	.w2(32'h38350b8a),
	.w3(32'hbc22746c),
	.w4(32'hba9fa78c),
	.w5(32'hbac1262a),
	.w6(32'hbab0f522),
	.w7(32'hbaf5c298),
	.w8(32'h3ac5a32e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1f3da),
	.w1(32'hbbe3662e),
	.w2(32'h3bb684eb),
	.w3(32'hbb00b853),
	.w4(32'hbc8dcc4b),
	.w5(32'h3af152b9),
	.w6(32'hbc75cadb),
	.w7(32'h3a2c5efe),
	.w8(32'hbba42cf6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0074c9),
	.w1(32'h3c19404e),
	.w2(32'h3c30c267),
	.w3(32'hbb615976),
	.w4(32'h3a8fd33b),
	.w5(32'h3b2c1f8c),
	.w6(32'h3bb0c5fc),
	.w7(32'h3cb35c77),
	.w8(32'h3b518e90),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabbe52),
	.w1(32'hbb92068d),
	.w2(32'h3c5247a8),
	.w3(32'hbc4466d8),
	.w4(32'hbbad893a),
	.w5(32'h3aae81ea),
	.w6(32'hbc562682),
	.w7(32'hbb84f055),
	.w8(32'hb98ed77f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ba9f6),
	.w1(32'h3d10a730),
	.w2(32'h3cb6e524),
	.w3(32'h3a73a359),
	.w4(32'h3cbde35b),
	.w5(32'h3b79f964),
	.w6(32'h3a5f9552),
	.w7(32'hbbde13aa),
	.w8(32'hbbe3e4d7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02a75d),
	.w1(32'h3bef5e93),
	.w2(32'h3c4a0f3e),
	.w3(32'hbc38b66b),
	.w4(32'h3b9a414e),
	.w5(32'h3c6f7cfb),
	.w6(32'h3b58ee1b),
	.w7(32'h3b8017a3),
	.w8(32'h3c28dd6f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf638a),
	.w1(32'hbb52496d),
	.w2(32'hbc59c638),
	.w3(32'hb919f3cb),
	.w4(32'hbc3be247),
	.w5(32'hbbbb1aac),
	.w6(32'hbabfbb7b),
	.w7(32'hbbf6b554),
	.w8(32'h3b0a0bdf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b888bca),
	.w1(32'hbc96b03b),
	.w2(32'hbccf42c4),
	.w3(32'h3b9cfee4),
	.w4(32'hbcbf5b3e),
	.w5(32'hbc9b5ec5),
	.w6(32'hbbbd03a0),
	.w7(32'hbccecdac),
	.w8(32'hbbed7604),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacc3f7),
	.w1(32'h3cf3bbf6),
	.w2(32'h3c8b12df),
	.w3(32'hbc27bf59),
	.w4(32'hbab9b68c),
	.w5(32'hbc05a1dd),
	.w6(32'h3c519c84),
	.w7(32'h3c80f7b8),
	.w8(32'h3c870609),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0b38),
	.w1(32'h3b4cca38),
	.w2(32'h3c95723b),
	.w3(32'hbc45e619),
	.w4(32'h3afe098e),
	.w5(32'h3c0f19b6),
	.w6(32'h3c1a2f05),
	.w7(32'hba8e9d97),
	.w8(32'h3be5ca92),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2272f2),
	.w1(32'h3b7170b0),
	.w2(32'h3c09463f),
	.w3(32'h3aeb94e5),
	.w4(32'h3be835ca),
	.w5(32'h3bb0f035),
	.w6(32'h3b775fc5),
	.w7(32'h39beec6c),
	.w8(32'hb8a26bf5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3cd8),
	.w1(32'h3c1cc79c),
	.w2(32'h3c2559af),
	.w3(32'h3c8e73c4),
	.w4(32'hbb1f6aff),
	.w5(32'h3c8929b5),
	.w6(32'h3c1efad1),
	.w7(32'h3c1d20e8),
	.w8(32'h3cea568e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00b3ce),
	.w1(32'h3bbff280),
	.w2(32'hbb4035ae),
	.w3(32'h3ae9080b),
	.w4(32'hbc10961d),
	.w5(32'hbb830aa8),
	.w6(32'hba0180cb),
	.w7(32'hb79fee52),
	.w8(32'h39d4504c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc76fb0),
	.w1(32'h3d6aa6a7),
	.w2(32'h3da077ed),
	.w3(32'h3d029c25),
	.w4(32'h3d59081e),
	.w5(32'h3d909e5b),
	.w6(32'h3de97eca),
	.w7(32'h3de905ed),
	.w8(32'h3d4ba4a4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122375),
	.w1(32'hbbc4fd4e),
	.w2(32'hbc522165),
	.w3(32'hba010da0),
	.w4(32'hbc2da5ea),
	.w5(32'hbba8d969),
	.w6(32'h3b08b84f),
	.w7(32'hbc250fe1),
	.w8(32'hb910ca09),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d733),
	.w1(32'hbba45a5c),
	.w2(32'hbc1d3b17),
	.w3(32'hb9d33fd1),
	.w4(32'h3bb6a52c),
	.w5(32'h3b0297c1),
	.w6(32'hbb1746b2),
	.w7(32'hbbc02f01),
	.w8(32'hbc0966de),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc420b5d),
	.w1(32'hbc812671),
	.w2(32'hbc5f5ac7),
	.w3(32'hb90226de),
	.w4(32'hbcd146a5),
	.w5(32'hbc4e5c94),
	.w6(32'hbb5b57a9),
	.w7(32'hbc43388a),
	.w8(32'hbae877fd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba31a31),
	.w1(32'h3ce6bba4),
	.w2(32'hbc9f4c09),
	.w3(32'hbaa87742),
	.w4(32'h3c9147c4),
	.w5(32'hbc345a84),
	.w6(32'h3ca3ed1b),
	.w7(32'hbb61c7a3),
	.w8(32'hbb8cf594),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabc739),
	.w1(32'hbce019a0),
	.w2(32'hbcdcfff8),
	.w3(32'hbc2d0208),
	.w4(32'hbcc7ceee),
	.w5(32'hbcb28c42),
	.w6(32'hbc91aadd),
	.w7(32'hbcb581a0),
	.w8(32'hbb1cb82b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b07e),
	.w1(32'h3bae6e89),
	.w2(32'h3bd09c92),
	.w3(32'hbb6c96e6),
	.w4(32'h3be45b07),
	.w5(32'h3a3431d5),
	.w6(32'h3b2bedcf),
	.w7(32'h3bddc0a5),
	.w8(32'h3b8a182e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc3e64),
	.w1(32'hbcd6444b),
	.w2(32'hbc25ae37),
	.w3(32'hbbbd737c),
	.w4(32'hbc4db42e),
	.w5(32'h3b0aff6f),
	.w6(32'hbc8a8ede),
	.w7(32'hbc93c8dd),
	.w8(32'h387074fa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7576f),
	.w1(32'h3bfd359d),
	.w2(32'h3c225c5f),
	.w3(32'h3cdeb399),
	.w4(32'h3aec8cc9),
	.w5(32'h3c1ab620),
	.w6(32'hb9e2cc4d),
	.w7(32'h3c0e7090),
	.w8(32'h3c27cb62),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c394a01),
	.w1(32'hbbdccb99),
	.w2(32'hbbe0be06),
	.w3(32'h3c21c680),
	.w4(32'hbbb977e6),
	.w5(32'hbb0a50a2),
	.w6(32'hb9806872),
	.w7(32'hbb964432),
	.w8(32'hbb4cda0c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7bc50),
	.w1(32'hb9c4b4f4),
	.w2(32'hb9d9c1db),
	.w3(32'hbb058243),
	.w4(32'hbad3737c),
	.w5(32'hba800fc1),
	.w6(32'h3ba77404),
	.w7(32'hbaad6621),
	.w8(32'h3b7346f9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6496f),
	.w1(32'hbc52ed63),
	.w2(32'h3af124b6),
	.w3(32'hbb199c68),
	.w4(32'hbc9ac939),
	.w5(32'h3b2b8da1),
	.w6(32'hbc223fc0),
	.w7(32'hbc07d0fc),
	.w8(32'h3c16570a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f4045),
	.w1(32'h3ae89c7a),
	.w2(32'hbbace056),
	.w3(32'h3bcc028b),
	.w4(32'h3b65332a),
	.w5(32'hbad94a68),
	.w6(32'h3c10f814),
	.w7(32'h3b0f4780),
	.w8(32'h3aa4ce14),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8accac),
	.w1(32'h3b918430),
	.w2(32'h3b3c76d9),
	.w3(32'h3c1542fe),
	.w4(32'h3afb8588),
	.w5(32'h3b5493de),
	.w6(32'hb98ff0bb),
	.w7(32'h3acb5f27),
	.w8(32'h3ba3e025),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad0dce),
	.w1(32'h3c25ddc5),
	.w2(32'h3b6f3803),
	.w3(32'hbba869fb),
	.w4(32'h3be0bbf3),
	.w5(32'hbbf3d8ca),
	.w6(32'hbc18da77),
	.w7(32'h3a236742),
	.w8(32'hbc52090c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39bdd2),
	.w1(32'hbc517edf),
	.w2(32'hbc31c021),
	.w3(32'hbb54c15a),
	.w4(32'hbb9a57ff),
	.w5(32'hba652a4b),
	.w6(32'hbbf1f5bc),
	.w7(32'hbc28a0b1),
	.w8(32'hbb400b67),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b5efa),
	.w1(32'h3bc75876),
	.w2(32'h3a3d8d70),
	.w3(32'h3c58b945),
	.w4(32'h3bba1691),
	.w5(32'h3b55c491),
	.w6(32'hbb52162d),
	.w7(32'hbb149ac5),
	.w8(32'h3bf5568f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1968ec),
	.w1(32'h3a0340ea),
	.w2(32'h3c46a10b),
	.w3(32'h3b24b18d),
	.w4(32'hb9a004a4),
	.w5(32'h3c4edfb4),
	.w6(32'hbae7e992),
	.w7(32'h3bef2c7d),
	.w8(32'h3babba19),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24a62b),
	.w1(32'h3ad25a00),
	.w2(32'h3be7c610),
	.w3(32'hba333a78),
	.w4(32'h3ad986f7),
	.w5(32'h3bc631f7),
	.w6(32'hb98c9eb9),
	.w7(32'h3baf4e9a),
	.w8(32'hbac4245a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab188be),
	.w1(32'hbb5cb3e2),
	.w2(32'h3c1ef5f1),
	.w3(32'hbb060ddd),
	.w4(32'h39a616e0),
	.w5(32'h3be44f6d),
	.w6(32'hba4e668d),
	.w7(32'h3b167fd8),
	.w8(32'h3bf8a153),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c770c79),
	.w1(32'hbb4eb2b6),
	.w2(32'h3c6ffd04),
	.w3(32'h3c280d45),
	.w4(32'h3a07a8e3),
	.w5(32'h3c801cdd),
	.w6(32'h3ab7b44d),
	.w7(32'h3bb3d981),
	.w8(32'h3c636aae),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f2736),
	.w1(32'hbb705b2c),
	.w2(32'hbc035d1a),
	.w3(32'h3c365967),
	.w4(32'h3b6a293b),
	.w5(32'hbafa8489),
	.w6(32'hbc6c3fec),
	.w7(32'hbbcf9c84),
	.w8(32'hbb719d97),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3307),
	.w1(32'h3c734b5d),
	.w2(32'h3c807573),
	.w3(32'hba6d9642),
	.w4(32'h3a87ad42),
	.w5(32'h3b80f8e6),
	.w6(32'h3c3d3da8),
	.w7(32'h3c4c0764),
	.w8(32'h3c70de95),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c881acc),
	.w1(32'hbb5f8f3a),
	.w2(32'hbb977bcc),
	.w3(32'hbbf1f420),
	.w4(32'hbbeb9f25),
	.w5(32'hbaf70cf4),
	.w6(32'hb956f0a3),
	.w7(32'hbaa76c8e),
	.w8(32'h3b3cd935),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24179),
	.w1(32'h3cbc8e7c),
	.w2(32'h3c49d32e),
	.w3(32'h39779a75),
	.w4(32'h3cbaa888),
	.w5(32'h3c3f9845),
	.w6(32'h3ae817cb),
	.w7(32'hbb6c4674),
	.w8(32'hba377467),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f5df),
	.w1(32'h3cb330b1),
	.w2(32'h3c00af90),
	.w3(32'hba947c18),
	.w4(32'h3ca24d76),
	.w5(32'h3c3a0880),
	.w6(32'h3c8d4190),
	.w7(32'h3c1c3c43),
	.w8(32'h3bb79fcc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2956a5),
	.w1(32'hbaefbddf),
	.w2(32'hbca167fd),
	.w3(32'hbbc573ce),
	.w4(32'hbc09de42),
	.w5(32'hbc8e7ab8),
	.w6(32'hbb8bf4c0),
	.w7(32'hbbaa7e6c),
	.w8(32'hbc407d7f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c310c),
	.w1(32'hbc5bfadc),
	.w2(32'hbc5db817),
	.w3(32'hbc2f92c2),
	.w4(32'hbc9e6aff),
	.w5(32'hbc808f71),
	.w6(32'hbb7c5fb1),
	.w7(32'hbc124dd9),
	.w8(32'hb9c3c2b8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22c1de),
	.w1(32'hb8c23e06),
	.w2(32'h3beb83a1),
	.w3(32'hb9be752b),
	.w4(32'hbc0e2ee6),
	.w5(32'hba338ed1),
	.w6(32'hbbae09a6),
	.w7(32'hbb0b8b5a),
	.w8(32'h3c033d1c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc25f08),
	.w1(32'hbbd17210),
	.w2(32'h3d476aa6),
	.w3(32'hbc0f032a),
	.w4(32'h3aa03d22),
	.w5(32'h3cbf835f),
	.w6(32'hbc854842),
	.w7(32'h3c65d4d2),
	.w8(32'h3c1072aa),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8071f9),
	.w1(32'hbc94d2f4),
	.w2(32'hbc9db789),
	.w3(32'hbb106c24),
	.w4(32'hbc471933),
	.w5(32'hbc0a0c54),
	.w6(32'hbbcd9a4d),
	.w7(32'hbc8a80f2),
	.w8(32'hbb273232),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384fc54b),
	.w1(32'hbaf16ef5),
	.w2(32'h3b0ee4ad),
	.w3(32'h3bdecd5b),
	.w4(32'h3b35527a),
	.w5(32'h3b924645),
	.w6(32'h3a237962),
	.w7(32'h3b05a65f),
	.w8(32'h3acda078),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0668f),
	.w1(32'h3bc03ac9),
	.w2(32'h3ac77756),
	.w3(32'hb9ada773),
	.w4(32'hbc03e562),
	.w5(32'h3c347dbc),
	.w6(32'h3bac874e),
	.w7(32'hbca2b377),
	.w8(32'h3bb6798c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e696),
	.w1(32'h3c97a18f),
	.w2(32'h3c8e400e),
	.w3(32'h3b16d9ba),
	.w4(32'h3c8f684b),
	.w5(32'h3b60fa96),
	.w6(32'hbb44996f),
	.w7(32'h3c512536),
	.w8(32'h3c1b3491),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393233a7),
	.w1(32'hb9d3cdf6),
	.w2(32'hba29944d),
	.w3(32'hbc8aa4b1),
	.w4(32'h3ace6d96),
	.w5(32'hbbe09121),
	.w6(32'hbb2122a8),
	.w7(32'h3bfe5a2c),
	.w8(32'hbb7eaf95),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a747e),
	.w1(32'h3c89ca6a),
	.w2(32'hbc4254d8),
	.w3(32'hbc103764),
	.w4(32'h3c8d9fe9),
	.w5(32'h39b537d4),
	.w6(32'h3c4be065),
	.w7(32'hba104c7b),
	.w8(32'hba96a14a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fe207),
	.w1(32'h393e8ff7),
	.w2(32'h3bb5dc3c),
	.w3(32'h3b505f38),
	.w4(32'h3b79a643),
	.w5(32'h3bfdef30),
	.w6(32'hbc0a3550),
	.w7(32'hbb2a07df),
	.w8(32'h3b1b1065),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0079ff),
	.w1(32'h3c7e55d7),
	.w2(32'h392203cd),
	.w3(32'h3bf0dcce),
	.w4(32'h3c522167),
	.w5(32'h3adca9e9),
	.w6(32'h3c4fd6ac),
	.w7(32'h3b930613),
	.w8(32'h3a8180c8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc72ce5),
	.w1(32'hbba991a6),
	.w2(32'hbbbb955b),
	.w3(32'h3b113e4b),
	.w4(32'h3a970999),
	.w5(32'h3b074526),
	.w6(32'h3be3d6d1),
	.w7(32'hba8ca050),
	.w8(32'hba171e8d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1419),
	.w1(32'hbbf0c927),
	.w2(32'hbc373f2b),
	.w3(32'hbb44b413),
	.w4(32'hbbe80dbe),
	.w5(32'h3b74f65b),
	.w6(32'hbc1ed196),
	.w7(32'hbb6acd01),
	.w8(32'hbc2ee883),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b022e0e),
	.w1(32'hbad29925),
	.w2(32'h3c1330a8),
	.w3(32'h3c4f88f9),
	.w4(32'h3bd54b74),
	.w5(32'h3c2dbddf),
	.w6(32'hbbd2885f),
	.w7(32'hba8faca9),
	.w8(32'h3c6a1667),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1170e8),
	.w1(32'h3c03020e),
	.w2(32'hbb6a46e3),
	.w3(32'hbbedc1db),
	.w4(32'hba701460),
	.w5(32'hbbcaffa4),
	.w6(32'h3c9278fb),
	.w7(32'h3c36d2b1),
	.w8(32'h3b993ec6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819861),
	.w1(32'h3c1251c8),
	.w2(32'h3ceba924),
	.w3(32'h3b32a674),
	.w4(32'h3c4c1854),
	.w5(32'h3d061c40),
	.w6(32'h3c0797d9),
	.w7(32'h3b8affd5),
	.w8(32'h3c42cf73),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f68f8),
	.w1(32'h3b3d3f72),
	.w2(32'hb88ac773),
	.w3(32'h3bb68bad),
	.w4(32'h3aafe333),
	.w5(32'hbbf3a1d7),
	.w6(32'hbc3fe93b),
	.w7(32'hbbfac39e),
	.w8(32'hbc0ffc5a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40fb18),
	.w1(32'h3c630b67),
	.w2(32'h3cdaec42),
	.w3(32'hbbd835fc),
	.w4(32'h3c362082),
	.w5(32'h3c98e9fa),
	.w6(32'h3ca0c784),
	.w7(32'h3c92572d),
	.w8(32'h3c731057),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fbe6b),
	.w1(32'h3c1674e7),
	.w2(32'h3c49f5e7),
	.w3(32'h3bbd9134),
	.w4(32'h3c568759),
	.w5(32'h3c511c9e),
	.w6(32'hba6fce0e),
	.w7(32'h3a87d160),
	.w8(32'h3a6c421a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af96cb7),
	.w1(32'hbc477d0c),
	.w2(32'hbb281cac),
	.w3(32'h3b780b98),
	.w4(32'hbc4d8e4f),
	.w5(32'h3ba9c1ed),
	.w6(32'hbc0a4e4c),
	.w7(32'hbc1c998f),
	.w8(32'h3b4e3ab8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0814fc),
	.w1(32'h3b824cfb),
	.w2(32'h3b3292dd),
	.w3(32'h3b47cc50),
	.w4(32'hbbd36b5e),
	.w5(32'hbc666486),
	.w6(32'h393d1ffc),
	.w7(32'hbb6cd381),
	.w8(32'hbc390ccd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92713d),
	.w1(32'h3c915c9e),
	.w2(32'h3d290208),
	.w3(32'hbc8d395a),
	.w4(32'hba864060),
	.w5(32'h3c890754),
	.w6(32'hbb0da9ba),
	.w7(32'h3cdca25d),
	.w8(32'h3c1ac6dc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468254),
	.w1(32'hbcb59ca0),
	.w2(32'hbbc8046f),
	.w3(32'hbc314468),
	.w4(32'hbc8527ca),
	.w5(32'hba80732f),
	.w6(32'hbca31ce0),
	.w7(32'hbc540481),
	.w8(32'hbb1f1897),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6135ba),
	.w1(32'hbc2d76c9),
	.w2(32'h3c0d3366),
	.w3(32'h3c15f102),
	.w4(32'hbbeed131),
	.w5(32'h3c1f038d),
	.w6(32'hbb86efca),
	.w7(32'hba7edc69),
	.w8(32'h3bdab46a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b27f),
	.w1(32'h3bacd6c0),
	.w2(32'h3bbfcb83),
	.w3(32'hbb74702c),
	.w4(32'h3b82dac0),
	.w5(32'hbbd893d0),
	.w6(32'h3bf48325),
	.w7(32'h3c0f0962),
	.w8(32'h3b82fe78),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea279),
	.w1(32'hbc1394c6),
	.w2(32'hbb6756bc),
	.w3(32'hbc25a8e1),
	.w4(32'hbb69461c),
	.w5(32'hbbce9216),
	.w6(32'hbb06c565),
	.w7(32'h3bdd3e16),
	.w8(32'h39ad2f0c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075602),
	.w1(32'hbb9927fe),
	.w2(32'hbb4ed567),
	.w3(32'h3b280cc4),
	.w4(32'hbc079804),
	.w5(32'hbc1d4052),
	.w6(32'hbb038421),
	.w7(32'hba567eef),
	.w8(32'hbb293919),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a736),
	.w1(32'hbbaf20d0),
	.w2(32'hbb8e4dca),
	.w3(32'hbbf30142),
	.w4(32'h3ad79f18),
	.w5(32'hbbf9c842),
	.w6(32'hbb002360),
	.w7(32'h3c08ca15),
	.w8(32'h3ac82f62),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388fcf53),
	.w1(32'h3ce730ed),
	.w2(32'h3d16518f),
	.w3(32'hbc1ec49f),
	.w4(32'h3cabf010),
	.w5(32'h3c7c683c),
	.w6(32'h3c377d87),
	.w7(32'h3c6afccf),
	.w8(32'h3b8f8675),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8804f),
	.w1(32'hbba4c9c6),
	.w2(32'hbb1c0934),
	.w3(32'hbbb8c5ef),
	.w4(32'hbc4d873c),
	.w5(32'hbb488d88),
	.w6(32'hba2c7d8f),
	.w7(32'hbc25fdbf),
	.w8(32'hbb7addb5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2210bd),
	.w1(32'h3c9ed946),
	.w2(32'h3bd8c3d0),
	.w3(32'h3cbbedb9),
	.w4(32'h3c04545f),
	.w5(32'h3c5edc27),
	.w6(32'h3c6a65a5),
	.w7(32'h3c151c34),
	.w8(32'h3c8e3e38),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7c86),
	.w1(32'h3c0ef7e2),
	.w2(32'h3b319bc2),
	.w3(32'hbc399892),
	.w4(32'h3a9a11e9),
	.w5(32'h3bd9027b),
	.w6(32'h3b7a1223),
	.w7(32'hbb88a37d),
	.w8(32'h3c355573),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4df95b),
	.w1(32'hbaea3042),
	.w2(32'hbab9f179),
	.w3(32'h3c15d7c2),
	.w4(32'hbbdc8e00),
	.w5(32'hbbf5d79d),
	.w6(32'h3a6ae8fd),
	.w7(32'h3a97dad2),
	.w8(32'h3b909fb0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71eec7),
	.w1(32'h3bbda31a),
	.w2(32'hbbb84239),
	.w3(32'hbb436240),
	.w4(32'h3bd551b9),
	.w5(32'hbb660f85),
	.w6(32'h3b14b851),
	.w7(32'h3beeef95),
	.w8(32'h3b8b6abf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3b877),
	.w1(32'hbc12d878),
	.w2(32'hbb5d39ab),
	.w3(32'h3c04bf47),
	.w4(32'hbc27df26),
	.w5(32'hbbd59dae),
	.w6(32'h39ed1741),
	.w7(32'hbb6fafe0),
	.w8(32'h3b0485cc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43cf95),
	.w1(32'h3bd8e0ce),
	.w2(32'h3bbb8a2b),
	.w3(32'h3b6eed2c),
	.w4(32'hbb5ed1b9),
	.w5(32'h3bd25014),
	.w6(32'hbb5e1ff5),
	.w7(32'h3ae31931),
	.w8(32'h3adefd84),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc583e9),
	.w1(32'h3c445ece),
	.w2(32'h3cb8b30e),
	.w3(32'hb9d3c543),
	.w4(32'h3c668053),
	.w5(32'h3c3279d2),
	.w6(32'h3be92845),
	.w7(32'h3c2a12af),
	.w8(32'h3c3b981d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fad5a),
	.w1(32'h3b8a09a0),
	.w2(32'h3bea6993),
	.w3(32'h3a7121fc),
	.w4(32'hba4dd9e8),
	.w5(32'h3ab69944),
	.w6(32'h3a1c3968),
	.w7(32'h3bcbbe3e),
	.w8(32'h39c798c0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fed52),
	.w1(32'hbae76397),
	.w2(32'h3b108ff2),
	.w3(32'hbbe8fd48),
	.w4(32'hbb69d64a),
	.w5(32'h3aa8339f),
	.w6(32'hb9b04ffd),
	.w7(32'h3921bc6a),
	.w8(32'hbbbb838b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0430cb),
	.w1(32'h3bf568ac),
	.w2(32'h3b82b550),
	.w3(32'h3b0d9e08),
	.w4(32'h3b3de476),
	.w5(32'h3be64ca3),
	.w6(32'h3b851ee8),
	.w7(32'h3a70f975),
	.w8(32'h3bb089c0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accdd6b),
	.w1(32'hbc0b3c81),
	.w2(32'hbd226406),
	.w3(32'h3b378da6),
	.w4(32'hbccd6b30),
	.w5(32'hbce53f60),
	.w6(32'h3b9f7d75),
	.w7(32'hbc94ecc7),
	.w8(32'h3bfd5e8a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce17a08),
	.w1(32'hbbe7d15a),
	.w2(32'h3bb78e8a),
	.w3(32'h3cf4e487),
	.w4(32'hbb1e17b4),
	.w5(32'h3c0ccaed),
	.w6(32'hbab4a88f),
	.w7(32'h3b25c536),
	.w8(32'h3c06e4a1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31ab76),
	.w1(32'hb8970853),
	.w2(32'h3ca1e215),
	.w3(32'h3bed589f),
	.w4(32'hbc050960),
	.w5(32'h3cb9bdcf),
	.w6(32'hbbe15e37),
	.w7(32'h3c2593a2),
	.w8(32'h3ce841db),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d7624),
	.w1(32'hbc21120c),
	.w2(32'hbb0ecfae),
	.w3(32'h3cf2ca87),
	.w4(32'hbcb627fb),
	.w5(32'hbb837174),
	.w6(32'hbc39146d),
	.w7(32'hbc9cad92),
	.w8(32'hba47dce5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c568039),
	.w1(32'hbb49b6a1),
	.w2(32'h3c916b14),
	.w3(32'h3c103f57),
	.w4(32'hbc01fc14),
	.w5(32'h3c18d71b),
	.w6(32'hbbf0ad79),
	.w7(32'h3b1913c3),
	.w8(32'h3ba2150b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b684e),
	.w1(32'hbc3aa6a4),
	.w2(32'hbcc8107b),
	.w3(32'h3b43951f),
	.w4(32'hbc4b0d70),
	.w5(32'hbcba78c2),
	.w6(32'hbb273ef0),
	.w7(32'hbca53a80),
	.w8(32'hbc7dd804),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a49b2),
	.w1(32'hba1114ef),
	.w2(32'h3b366fea),
	.w3(32'hbc55033c),
	.w4(32'h3c2b7e26),
	.w5(32'h3b3fb9a5),
	.w6(32'h3b9c619a),
	.w7(32'h3c0bf218),
	.w8(32'hb92e0f9b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980c636),
	.w1(32'h3c4f6b19),
	.w2(32'hba803cfb),
	.w3(32'hbc487f6d),
	.w4(32'h3b92c247),
	.w5(32'hbc11f1d7),
	.w6(32'h3c804f09),
	.w7(32'h3c2d5010),
	.w8(32'hbbe6fdc6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9757c3),
	.w1(32'h3c04950c),
	.w2(32'h3c3ecc4c),
	.w3(32'hbc04626a),
	.w4(32'h3b88dc7b),
	.w5(32'hbbd9afdd),
	.w6(32'h3c20cd32),
	.w7(32'h3c4b7b8c),
	.w8(32'h39d3a762),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cad60),
	.w1(32'h3c97703e),
	.w2(32'h3d2570b4),
	.w3(32'hbafb2a5e),
	.w4(32'h3c86a953),
	.w5(32'h3c66f8f5),
	.w6(32'hbb965f69),
	.w7(32'h3cc30934),
	.w8(32'h3c514526),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63b37a),
	.w1(32'h3bc1eeb8),
	.w2(32'h3ce02282),
	.w3(32'hbc8a8432),
	.w4(32'h3bd7321c),
	.w5(32'h3beda931),
	.w6(32'hbc30587b),
	.w7(32'h3cb764d6),
	.w8(32'h38d16687),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb772f66),
	.w1(32'h3cc1c3db),
	.w2(32'h3c7be084),
	.w3(32'h3a66dfae),
	.w4(32'h3c8dd3fd),
	.w5(32'h3c3f725c),
	.w6(32'h3c91c540),
	.w7(32'h3c509acd),
	.w8(32'h3b97c3f5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed1684),
	.w1(32'hbc050043),
	.w2(32'h3c4b01d1),
	.w3(32'h3a858af8),
	.w4(32'h3a54d7db),
	.w5(32'h3c7f5b20),
	.w6(32'h3bcd8477),
	.w7(32'h3aa52884),
	.w8(32'h3c9f57d9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c738cbc),
	.w1(32'hbada9627),
	.w2(32'h3b1ab35d),
	.w3(32'hba3bd2ea),
	.w4(32'h39a7358d),
	.w5(32'h3bfa4ebc),
	.w6(32'h3a941726),
	.w7(32'h3b60caf0),
	.w8(32'hbaeabd39),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0d9d2),
	.w1(32'hbb91562d),
	.w2(32'hbc6c1061),
	.w3(32'hbbaf807a),
	.w4(32'h3b205e69),
	.w5(32'hbc008d0d),
	.w6(32'h3a4b561c),
	.w7(32'hbb804605),
	.w8(32'h3b34fbb2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3239d),
	.w1(32'h3c71309e),
	.w2(32'h3b633e6c),
	.w3(32'hbc22638b),
	.w4(32'h3c1b3f37),
	.w5(32'h3b554091),
	.w6(32'h3c6fcad2),
	.w7(32'h3bf65358),
	.w8(32'h3b926b85),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1add),
	.w1(32'h3c06cce6),
	.w2(32'h3c8a341f),
	.w3(32'hbaacfcbd),
	.w4(32'h3c064af5),
	.w5(32'h3b7d20e5),
	.w6(32'h3c886ed1),
	.w7(32'h3c3cdf99),
	.w8(32'h3c73f3aa),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8caf0a),
	.w1(32'h3b9b5a96),
	.w2(32'h3996d4bd),
	.w3(32'hbb905d22),
	.w4(32'h3a640e5b),
	.w5(32'h3ab4022e),
	.w6(32'h39cfd0e8),
	.w7(32'h3b04d3a2),
	.w8(32'hba58a53c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d7ce),
	.w1(32'hbb84c667),
	.w2(32'h3b0a0308),
	.w3(32'hba8a7dca),
	.w4(32'hbb36e5e6),
	.w5(32'h3ad61d94),
	.w6(32'hbc33d298),
	.w7(32'hba572ba9),
	.w8(32'hbaa4ce9c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3d789),
	.w1(32'hbbc62bce),
	.w2(32'hb830d824),
	.w3(32'h3c2ede0c),
	.w4(32'hbacb4668),
	.w5(32'h3aa16c1b),
	.w6(32'h3a915da5),
	.w7(32'hba309e0d),
	.w8(32'hbbdf1ace),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41da8b),
	.w1(32'h38f7c50d),
	.w2(32'h3b08fe2e),
	.w3(32'h3c0f23a9),
	.w4(32'h3a42e81b),
	.w5(32'hbb3d2436),
	.w6(32'hbaa5b1e6),
	.w7(32'hbaf043d1),
	.w8(32'hb9e191f6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926295),
	.w1(32'h3c369a28),
	.w2(32'hbb95e1da),
	.w3(32'hbb980cfb),
	.w4(32'h3bd6f5e2),
	.w5(32'hbb777b33),
	.w6(32'h3c5d37f8),
	.w7(32'h3af2cdba),
	.w8(32'hbb7c0259),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f70b8),
	.w1(32'h3c1b656e),
	.w2(32'h3be9a5e2),
	.w3(32'hbb8f28d2),
	.w4(32'h3c53961d),
	.w5(32'h3c34138a),
	.w6(32'h3bca827e),
	.w7(32'h3baa3d47),
	.w8(32'hbc1b4191),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ad841),
	.w1(32'h3b85b227),
	.w2(32'h3b510aaf),
	.w3(32'hbcb2de55),
	.w4(32'h3c0ec7a8),
	.w5(32'h3bbdd273),
	.w6(32'h38e9ac7f),
	.w7(32'h3c26172e),
	.w8(32'h3bde2695),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd3355),
	.w1(32'h3a56cac5),
	.w2(32'hbbf894d9),
	.w3(32'h3b1a6697),
	.w4(32'h3b8b8b21),
	.w5(32'hbce00dbe),
	.w6(32'h3b0ef1f2),
	.w7(32'h3b62970b),
	.w8(32'hb9bb5506),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc333587),
	.w1(32'h3c4efe5d),
	.w2(32'h3c48aaff),
	.w3(32'hbc8dcf63),
	.w4(32'h3b8853c3),
	.w5(32'h3a1c6f3a),
	.w6(32'h3bc0721d),
	.w7(32'h3be147ef),
	.w8(32'hbaea3da8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb675c07),
	.w1(32'h3bd423f3),
	.w2(32'h3baef6b4),
	.w3(32'hbc248de0),
	.w4(32'h3af80b7a),
	.w5(32'h3b98a949),
	.w6(32'h3b90f67d),
	.w7(32'h3bba1a52),
	.w8(32'h3af0fefa),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a4553),
	.w1(32'h3b40de78),
	.w2(32'hbb2480f0),
	.w3(32'h3b6e9220),
	.w4(32'hbb262ab3),
	.w5(32'hbbf0598c),
	.w6(32'hbb9de547),
	.w7(32'hbbeab260),
	.w8(32'h3ae0b45d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9332d0),
	.w1(32'h3b94f795),
	.w2(32'h3b3330df),
	.w3(32'hbc10fe3a),
	.w4(32'h3b808be4),
	.w5(32'h3b35cfca),
	.w6(32'h3b53f2b4),
	.w7(32'h3a46aa35),
	.w8(32'h3aae5179),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f641),
	.w1(32'hbac4591b),
	.w2(32'hbbf5881f),
	.w3(32'hbb0f79e7),
	.w4(32'h3921214a),
	.w5(32'hbbca7b71),
	.w6(32'hbb6dd034),
	.w7(32'hbaf5da14),
	.w8(32'hbbce4fde),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb10da),
	.w1(32'h3c5e0ada),
	.w2(32'h3c5a5fc1),
	.w3(32'hbabafec8),
	.w4(32'h3c764d2a),
	.w5(32'h3c80df27),
	.w6(32'h3c1f56b5),
	.w7(32'h3cb05244),
	.w8(32'h38f9a7d0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26f6e3),
	.w1(32'hbcbcbc3d),
	.w2(32'hbc109db5),
	.w3(32'h3b3c8582),
	.w4(32'hbc394e1a),
	.w5(32'h3a34ec37),
	.w6(32'hbab4b7bc),
	.w7(32'hbc16cb16),
	.w8(32'hba2035c1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ecf4e),
	.w1(32'h3bdf2526),
	.w2(32'h3b7923e5),
	.w3(32'hbb73fb06),
	.w4(32'hba4bef30),
	.w5(32'h3a116a65),
	.w6(32'h3b8d21db),
	.w7(32'h3b79901d),
	.w8(32'h3b6dd748),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8302b3),
	.w1(32'h3c4e09f9),
	.w2(32'h3b2252d9),
	.w3(32'hb9bebd4f),
	.w4(32'h3c28fab7),
	.w5(32'hbb198ccf),
	.w6(32'h3b820dd4),
	.w7(32'hbb32eeab),
	.w8(32'hbae7e818),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule