module layer_10_featuremap_450(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b5fd),
	.w1(32'hbbb0a7f5),
	.w2(32'hbbae4abb),
	.w3(32'h39b35b0f),
	.w4(32'hbb63170a),
	.w5(32'hbb542bd2),
	.w6(32'h3c05feb9),
	.w7(32'h3b3966ec),
	.w8(32'h3b693625),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfc4fc),
	.w1(32'hbb37d2a2),
	.w2(32'hbb8d88f6),
	.w3(32'hbad56ee6),
	.w4(32'hb9351f9b),
	.w5(32'hba9e9d1b),
	.w6(32'h3b62251d),
	.w7(32'h3b9ec49b),
	.w8(32'hbb154841),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c150436),
	.w1(32'hb9e1aa64),
	.w2(32'h3bd53d3c),
	.w3(32'h3c0049f8),
	.w4(32'hbaf45e70),
	.w5(32'h3a8bffd9),
	.w6(32'hbb0c61ca),
	.w7(32'hbb2139a9),
	.w8(32'hbc078027),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18710),
	.w1(32'hbb9e842a),
	.w2(32'hba1df9d0),
	.w3(32'h3b44ca17),
	.w4(32'h3be2883f),
	.w5(32'h3c276ef8),
	.w6(32'hbbfed617),
	.w7(32'h3bceee03),
	.w8(32'h3c06af48),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46c3e4),
	.w1(32'hbb7a57cd),
	.w2(32'hbb7a302a),
	.w3(32'h399c0c79),
	.w4(32'h3b5166a5),
	.w5(32'h3ac79c18),
	.w6(32'hbb7234d0),
	.w7(32'hbb9ae2a0),
	.w8(32'hbb412a15),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6f2a3),
	.w1(32'h3a6818a3),
	.w2(32'h3ad0a091),
	.w3(32'h3bdaf2ca),
	.w4(32'h3bd31594),
	.w5(32'h3b43c2cf),
	.w6(32'h3b1234d2),
	.w7(32'hbb093357),
	.w8(32'h3982e96c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c274d12),
	.w1(32'h3b892eb7),
	.w2(32'hbcb00a2f),
	.w3(32'h3bd03e39),
	.w4(32'hbc5991df),
	.w5(32'hbcb83242),
	.w6(32'h3bbf2d2c),
	.w7(32'hbc8970e7),
	.w8(32'hbd10d256),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca90bb4),
	.w1(32'hbcdd06f7),
	.w2(32'hbd1986fb),
	.w3(32'hbd029028),
	.w4(32'hbcff0237),
	.w5(32'hbd177dc8),
	.w6(32'hbcced09b),
	.w7(32'hbbb8f645),
	.w8(32'hbbef3464),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e12f2),
	.w1(32'h3b5ad933),
	.w2(32'hbb08dc87),
	.w3(32'hbce0f952),
	.w4(32'hbc0bc2c1),
	.w5(32'hbc169df1),
	.w6(32'hbc737521),
	.w7(32'hbbf76adf),
	.w8(32'hbc116d91),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfccc6),
	.w1(32'hbacab8b4),
	.w2(32'h3bc839ee),
	.w3(32'hb9aaa58e),
	.w4(32'h3a5e2a6c),
	.w5(32'h3c7e2ae3),
	.w6(32'h3ba15efd),
	.w7(32'hbb92bc11),
	.w8(32'h3c088ad8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10e2c6),
	.w1(32'h3c3b04ee),
	.w2(32'h3cea1032),
	.w3(32'h3a8e26c5),
	.w4(32'hbc1793a2),
	.w5(32'h3c193e24),
	.w6(32'h3a45b43a),
	.w7(32'hbc34e206),
	.w8(32'hbcb3077e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca62413),
	.w1(32'h3bb7f58b),
	.w2(32'h3b089334),
	.w3(32'h3c647fe1),
	.w4(32'h3c083ccd),
	.w5(32'h3afbfaab),
	.w6(32'hbb0435c2),
	.w7(32'hba85f3bf),
	.w8(32'hbac81799),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f3a2),
	.w1(32'hbc858727),
	.w2(32'hbbc83e2f),
	.w3(32'h3be32e6f),
	.w4(32'hbb672458),
	.w5(32'h3b8da82e),
	.w6(32'hbb915081),
	.w7(32'h3b2c98af),
	.w8(32'hbb7f563d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6072cf),
	.w1(32'hba9d1117),
	.w2(32'hbbbf068c),
	.w3(32'h3b676d10),
	.w4(32'h3b3a30e4),
	.w5(32'h3caf9db2),
	.w6(32'hbcb72562),
	.w7(32'hbb911765),
	.w8(32'h3c1d2331),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d98e3),
	.w1(32'h3bab85a1),
	.w2(32'h3b5c6ad7),
	.w3(32'h3c593e0a),
	.w4(32'h3a5cc082),
	.w5(32'h3aaea547),
	.w6(32'hba52a962),
	.w7(32'hbb8e0dc7),
	.w8(32'hbbda59a2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60d348),
	.w1(32'hbc6e304e),
	.w2(32'h3a93a0cc),
	.w3(32'hbba1cea5),
	.w4(32'hbbb20e99),
	.w5(32'hbad34e18),
	.w6(32'hbc2798fc),
	.w7(32'h3b6f2e0b),
	.w8(32'hbb86ebda),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080bd6),
	.w1(32'h3b9317c3),
	.w2(32'h3b83d768),
	.w3(32'hbbbe1b57),
	.w4(32'hbbb2ab9b),
	.w5(32'hba9f9d5c),
	.w6(32'hbbbd1bf3),
	.w7(32'hba722a35),
	.w8(32'h3b4c2f20),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbe63f),
	.w1(32'hbb84697f),
	.w2(32'hbb1f9bea),
	.w3(32'hbc0129ef),
	.w4(32'h3c0156e9),
	.w5(32'h39c5192c),
	.w6(32'hbb4c60c9),
	.w7(32'hbb577086),
	.w8(32'hbc47d53b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0bf47),
	.w1(32'h37d5fdfa),
	.w2(32'h3b4600e7),
	.w3(32'hbbe5778a),
	.w4(32'hbb39ffab),
	.w5(32'hbb6bfb8a),
	.w6(32'hbc2ac74d),
	.w7(32'hbbac0d25),
	.w8(32'hbb87e238),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf65c3),
	.w1(32'hbbda4a7c),
	.w2(32'hba693f2e),
	.w3(32'h3bb34486),
	.w4(32'hbc392622),
	.w5(32'hbabbdb73),
	.w6(32'h3bae034e),
	.w7(32'h36ae9379),
	.w8(32'hbb514ae3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebac18),
	.w1(32'h3bfde047),
	.w2(32'h3be277a4),
	.w3(32'hbb98494f),
	.w4(32'h3ba5b916),
	.w5(32'hba29d43b),
	.w6(32'hbbf7e5b7),
	.w7(32'hbb253ed4),
	.w8(32'hbb80b0e5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac69a9f),
	.w1(32'h3a13d7c4),
	.w2(32'h3b0c50c4),
	.w3(32'hbbc72269),
	.w4(32'h3b278041),
	.w5(32'h3baae931),
	.w6(32'h39aedeb0),
	.w7(32'h3c0a6677),
	.w8(32'h3aa9886f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf267b0),
	.w1(32'hbc8cfa94),
	.w2(32'hbc100d24),
	.w3(32'h39249b65),
	.w4(32'hbbf4eda0),
	.w5(32'hbc1e7541),
	.w6(32'hbaa54cde),
	.w7(32'h3afacb46),
	.w8(32'hbbd28f8b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b182744),
	.w1(32'h3a394a43),
	.w2(32'h3b884da8),
	.w3(32'hbb9c7670),
	.w4(32'h3c19cc90),
	.w5(32'h3c4cc72a),
	.w6(32'h3a89f0da),
	.w7(32'h3c494361),
	.w8(32'h3c799106),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b346e),
	.w1(32'hb8b8f903),
	.w2(32'h3c5fa50e),
	.w3(32'h3c622a7e),
	.w4(32'h3c0ea1bb),
	.w5(32'h3c29390d),
	.w6(32'h3ca81dd6),
	.w7(32'hbbecaa75),
	.w8(32'hbc548e49),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba310efc),
	.w1(32'h3b7559d8),
	.w2(32'h3b6ff596),
	.w3(32'h3b4c5673),
	.w4(32'h3bf93fdf),
	.w5(32'hbaa5a4fb),
	.w6(32'hbc1de575),
	.w7(32'h3ad1200d),
	.w8(32'h3a037297),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4faa1),
	.w1(32'hbb042237),
	.w2(32'h3a9b330c),
	.w3(32'hbb804ca7),
	.w4(32'hbb52647b),
	.w5(32'hbc048fb1),
	.w6(32'hbb8062d6),
	.w7(32'hbb0793ef),
	.w8(32'h39cd8295),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87c6d8),
	.w1(32'h3a991982),
	.w2(32'h3c3b0433),
	.w3(32'hbc0f3fd6),
	.w4(32'hbb4fbcc8),
	.w5(32'hbb946edb),
	.w6(32'hbb409ca0),
	.w7(32'hbb8835fb),
	.w8(32'hbc39f790),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f537b),
	.w1(32'h3b3de6f4),
	.w2(32'hbc0fc535),
	.w3(32'h39ced13e),
	.w4(32'hbb230269),
	.w5(32'hbc177997),
	.w6(32'h3bd336de),
	.w7(32'hbb4a1255),
	.w8(32'hbbc9f8fa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4cf32),
	.w1(32'h3b94bf6f),
	.w2(32'h3c188173),
	.w3(32'hbb5f90b2),
	.w4(32'h3b42695d),
	.w5(32'h3adc6527),
	.w6(32'h3aa06afc),
	.w7(32'hbb929d5c),
	.w8(32'hbbd43854),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1471a4),
	.w1(32'h3ab74aa3),
	.w2(32'hbc0083bb),
	.w3(32'h3b416f30),
	.w4(32'hbbaab9e7),
	.w5(32'h3ad24335),
	.w6(32'hbbef09e8),
	.w7(32'hba5d1c88),
	.w8(32'h3983e61b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42cb2),
	.w1(32'hbc11dbec),
	.w2(32'hbb718db6),
	.w3(32'hbbad9217),
	.w4(32'hbaaf026d),
	.w5(32'h392477d7),
	.w6(32'hbb4168e6),
	.w7(32'h3b499290),
	.w8(32'hbb022cb9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d25bf),
	.w1(32'hbb99d1c5),
	.w2(32'hbbb02a02),
	.w3(32'h3b2e78b2),
	.w4(32'hbc023052),
	.w5(32'hbc062dcd),
	.w6(32'hbc0066ed),
	.w7(32'h3b8449f1),
	.w8(32'hbb800638),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ef131),
	.w1(32'hbad6dae5),
	.w2(32'hbbdf97de),
	.w3(32'hbb8c1655),
	.w4(32'hbbd1d958),
	.w5(32'hbc736f7c),
	.w6(32'h3b82fd18),
	.w7(32'h38a1088d),
	.w8(32'hbb92d095),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a129),
	.w1(32'h3c0890e7),
	.w2(32'h3c87b16a),
	.w3(32'hbc337fc6),
	.w4(32'h3c05571f),
	.w5(32'h3c0f85f2),
	.w6(32'h3b848a1b),
	.w7(32'h3c03ca10),
	.w8(32'h3c8f848f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c809481),
	.w1(32'h3b45ec03),
	.w2(32'h3bedadd9),
	.w3(32'hb9ea8e07),
	.w4(32'hbab58fa6),
	.w5(32'h3c0cb7f0),
	.w6(32'h3bb0314d),
	.w7(32'hbaa176c6),
	.w8(32'h3be6ac68),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c151cb4),
	.w1(32'h3bb01b29),
	.w2(32'h3bb9a39a),
	.w3(32'h3c7fb0a3),
	.w4(32'hbbbc14c6),
	.w5(32'h3c8a83be),
	.w6(32'h3bb72e25),
	.w7(32'hbbaa8a6b),
	.w8(32'h3b98cdba),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8183c),
	.w1(32'hbaf4fa82),
	.w2(32'h38f0c016),
	.w3(32'hba399721),
	.w4(32'hbc90e7c3),
	.w5(32'hbc832e02),
	.w6(32'h3b986a9f),
	.w7(32'hbc416af0),
	.w8(32'hbcd187aa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f766b),
	.w1(32'h3c1c5bec),
	.w2(32'h3c6d9e14),
	.w3(32'h3b9317dc),
	.w4(32'hbb5225ab),
	.w5(32'h38b0e322),
	.w6(32'hbc0273ab),
	.w7(32'hbb9e448b),
	.w8(32'hbc136ebb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaea7f0),
	.w1(32'hba634991),
	.w2(32'hba9a5d55),
	.w3(32'h3b78889f),
	.w4(32'hba905535),
	.w5(32'hbb52e128),
	.w6(32'hbac30f54),
	.w7(32'hbb0e22e6),
	.w8(32'h3babe5ba),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbef845),
	.w1(32'hbb4b4b45),
	.w2(32'hbc82756d),
	.w3(32'hba1ab71e),
	.w4(32'h3ab6d87b),
	.w5(32'h3a3a050a),
	.w6(32'hbb1effdf),
	.w7(32'hbb8fce2e),
	.w8(32'h3bd5eb70),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe23470),
	.w1(32'hbb93dc24),
	.w2(32'hb9cc0440),
	.w3(32'h3b083444),
	.w4(32'hbb412890),
	.w5(32'hbbb79947),
	.w6(32'hbb3d9e76),
	.w7(32'hbc089374),
	.w8(32'hbc1f732f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e0789f),
	.w1(32'hbbf8cc4c),
	.w2(32'hbbe5b831),
	.w3(32'h3b0dcc6d),
	.w4(32'h3ae28e58),
	.w5(32'h3a8de600),
	.w6(32'hbaa27785),
	.w7(32'hbb01dc2c),
	.w8(32'hbb5ac33d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc158e7b),
	.w1(32'hbca11314),
	.w2(32'hbbb980f2),
	.w3(32'hbac4d285),
	.w4(32'hbb70919b),
	.w5(32'hbc245952),
	.w6(32'hbc40ad5e),
	.w7(32'h3bb10b66),
	.w8(32'hba9b4aa7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc18eda),
	.w1(32'hba4bde7f),
	.w2(32'hbc0a4679),
	.w3(32'hbb3b74f7),
	.w4(32'hbbbf7c5e),
	.w5(32'hbb39165e),
	.w6(32'h39018c40),
	.w7(32'hbc0aff06),
	.w8(32'hbbab1e26),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e261),
	.w1(32'hb9c89b83),
	.w2(32'h3b8853a6),
	.w3(32'hbb298743),
	.w4(32'hba925606),
	.w5(32'h3bfb7946),
	.w6(32'h3bbbcf1d),
	.w7(32'h3b88ebcd),
	.w8(32'h3bfae3a2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0394),
	.w1(32'h3a4771ce),
	.w2(32'h3cd17868),
	.w3(32'hbba8b3f5),
	.w4(32'hb9836d4b),
	.w5(32'h3cdd7af9),
	.w6(32'hbbd6b6f3),
	.w7(32'h3a9dd579),
	.w8(32'h3c43c704),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcacf9b),
	.w1(32'hbc19b0c6),
	.w2(32'hbc6892df),
	.w3(32'h3b3f357d),
	.w4(32'hbb90c7c3),
	.w5(32'h3abee083),
	.w6(32'hbb07273c),
	.w7(32'hba1bb25f),
	.w8(32'h3b830269),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b0ab0),
	.w1(32'h3c10b9c2),
	.w2(32'hbba1e1aa),
	.w3(32'h3b870667),
	.w4(32'hbb48fceb),
	.w5(32'hbbc79ce8),
	.w6(32'h3bb81dfc),
	.w7(32'hbbf04b8c),
	.w8(32'hbb569d2f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25135b),
	.w1(32'hb96d6f0f),
	.w2(32'h3c525f7b),
	.w3(32'hbb96874d),
	.w4(32'hbbe4873e),
	.w5(32'h39d4dfb2),
	.w6(32'h3b1b7b5d),
	.w7(32'h3b210003),
	.w8(32'h3bd41b09),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c35d8),
	.w1(32'h3a7d8379),
	.w2(32'hbb11c852),
	.w3(32'hbafebf2a),
	.w4(32'h3a94f632),
	.w5(32'hbbab4cb8),
	.w6(32'hbc1fcba9),
	.w7(32'hbbcb8991),
	.w8(32'hba184e1e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbed15),
	.w1(32'h3bcb9922),
	.w2(32'hbab0575d),
	.w3(32'hbae3e116),
	.w4(32'hbbbd7200),
	.w5(32'h3bbb692d),
	.w6(32'hbb135048),
	.w7(32'hbc3d4b82),
	.w8(32'hbb3d9723),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a61ac),
	.w1(32'hbc24698b),
	.w2(32'hbc52b10f),
	.w3(32'hbb85da7e),
	.w4(32'hbc545ffc),
	.w5(32'hbc01f666),
	.w6(32'h3ba6e11e),
	.w7(32'hbc5bc6ff),
	.w8(32'hbca19333),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1efe88),
	.w1(32'hbcb00d7f),
	.w2(32'hbcac08b6),
	.w3(32'hbc659af6),
	.w4(32'hbc89ca1c),
	.w5(32'hbcce20fb),
	.w6(32'hbc7052a0),
	.w7(32'h3b4bb76c),
	.w8(32'hbc64cea9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4340f8),
	.w1(32'hbc4549fd),
	.w2(32'hbc817d25),
	.w3(32'hbc94cfe2),
	.w4(32'hbbfe128c),
	.w5(32'hbc6733f9),
	.w6(32'hbbff4f6c),
	.w7(32'h3afcecf0),
	.w8(32'hbb6c21dc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c452665),
	.w1(32'hb8dcb026),
	.w2(32'hbbe3b326),
	.w3(32'hbb32868f),
	.w4(32'hbabe5666),
	.w5(32'hbc10b946),
	.w6(32'hbc2270c4),
	.w7(32'h3b379237),
	.w8(32'hbc26dd99),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4303e),
	.w1(32'hbba396b5),
	.w2(32'h3b7af4a1),
	.w3(32'hb765bc82),
	.w4(32'hbb3ed5da),
	.w5(32'h3ab9df33),
	.w6(32'hbb6549b0),
	.w7(32'hbb17a0d1),
	.w8(32'hbb509569),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a794),
	.w1(32'hbb8645be),
	.w2(32'h3bff470c),
	.w3(32'h3bb3dda1),
	.w4(32'h3af78f5d),
	.w5(32'h3bcddc1f),
	.w6(32'h3b56fbac),
	.w7(32'hbb8775cf),
	.w8(32'h3b66c25b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27d6cf),
	.w1(32'h3bb28fee),
	.w2(32'hb9dd2920),
	.w3(32'hbb7205c0),
	.w4(32'h3c14e4fa),
	.w5(32'hba633d63),
	.w6(32'hbb4e5b2c),
	.w7(32'h3bb6c246),
	.w8(32'h3a13c19e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fa79d),
	.w1(32'hba894ace),
	.w2(32'h3c42a31b),
	.w3(32'h3aabb596),
	.w4(32'h3a654af4),
	.w5(32'h3c479dad),
	.w6(32'hbb1152a1),
	.w7(32'h3b28db54),
	.w8(32'h3bc617a5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf472af),
	.w1(32'hbb3f8f12),
	.w2(32'h3c1db042),
	.w3(32'hba78b91e),
	.w4(32'hbb1eb1ed),
	.w5(32'h3c3e4a59),
	.w6(32'hbb4c3456),
	.w7(32'h3ba77380),
	.w8(32'h3a0e6d39),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5107),
	.w1(32'hbaa83aa0),
	.w2(32'h3ac52c4d),
	.w3(32'h3b2fa1d6),
	.w4(32'h3a21228c),
	.w5(32'hba8728ca),
	.w6(32'hbb0fcfc3),
	.w7(32'hbb0d2c3c),
	.w8(32'hbbe4fb43),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb513689),
	.w1(32'hbbade9e0),
	.w2(32'hbb2b8b6d),
	.w3(32'h3bcd57b6),
	.w4(32'h3c0bda3b),
	.w5(32'hb998ffbb),
	.w6(32'h3b838b30),
	.w7(32'h3c0c459b),
	.w8(32'h3b210555),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143f10),
	.w1(32'h3afa60ed),
	.w2(32'h3ac08fc2),
	.w3(32'hbc2f049c),
	.w4(32'hba993dbb),
	.w5(32'hbb68fc57),
	.w6(32'hbc4e0962),
	.w7(32'hb90f28a3),
	.w8(32'h3b9697b0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ab02),
	.w1(32'h3b402e56),
	.w2(32'h3c36d11d),
	.w3(32'h3a82652c),
	.w4(32'h39fa66f6),
	.w5(32'h3bd2c360),
	.w6(32'hba89214f),
	.w7(32'hba05ee84),
	.w8(32'h3c05d62a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5837c),
	.w1(32'h3b076d1f),
	.w2(32'hbbce51de),
	.w3(32'h3b0e7cd5),
	.w4(32'h3a980e52),
	.w5(32'h3a1dd86d),
	.w6(32'hbb3313a1),
	.w7(32'hbc394fd6),
	.w8(32'hbc5871f7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7783c),
	.w1(32'hbc341819),
	.w2(32'hbbde4ee0),
	.w3(32'h3c0bce48),
	.w4(32'h3be8ec51),
	.w5(32'h3bd737b6),
	.w6(32'hbc0fda24),
	.w7(32'h3c0351a4),
	.w8(32'h3c2dfbe3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237a7e),
	.w1(32'h3b5c9d77),
	.w2(32'hbc2a8e17),
	.w3(32'h3c1496de),
	.w4(32'h3bbdfd53),
	.w5(32'hbb6e91f0),
	.w6(32'h3c581a93),
	.w7(32'h3c80657f),
	.w8(32'h3ccaaebc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8de0b0),
	.w1(32'hbc0c796e),
	.w2(32'hbc4873ac),
	.w3(32'hbbe6851b),
	.w4(32'hbb2d4b89),
	.w5(32'hbc19d9d3),
	.w6(32'h3c022849),
	.w7(32'hbb7f7ace),
	.w8(32'h3afb586a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27f9eb),
	.w1(32'h3bc96615),
	.w2(32'h3c1e9792),
	.w3(32'hb9b67802),
	.w4(32'hbbbfc839),
	.w5(32'h3b28055d),
	.w6(32'h3b65e561),
	.w7(32'hbc03d3e7),
	.w8(32'hb9ac8a94),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb712082e),
	.w1(32'h361a629a),
	.w2(32'h36fe5a1b),
	.w3(32'hb68f5b78),
	.w4(32'hb7502815),
	.w5(32'h381e7b83),
	.w6(32'h3600e076),
	.w7(32'hb6c32d66),
	.w8(32'h3872f9dd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e69280),
	.w1(32'hb86e2e2c),
	.w2(32'h37fc9998),
	.w3(32'hb7b34337),
	.w4(32'hb89a91a4),
	.w5(32'h38025d62),
	.w6(32'hb6b2625b),
	.w7(32'hb803fa89),
	.w8(32'h3858d73d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85dff7d),
	.w1(32'hb8cc92c7),
	.w2(32'h37edeaa9),
	.w3(32'hb8b85122),
	.w4(32'hb85bcd41),
	.w5(32'h3798b3b7),
	.w6(32'h36aa14a3),
	.w7(32'h370300ad),
	.w8(32'h37866987),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba047e8c),
	.w1(32'hbae5a50e),
	.w2(32'hbae315f3),
	.w3(32'hb8d0365a),
	.w4(32'hb780f0f0),
	.w5(32'hba4732e6),
	.w6(32'hba34532a),
	.w7(32'h3619d88f),
	.w8(32'hba202490),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38898bad),
	.w1(32'hb6eee12c),
	.w2(32'hb82891fe),
	.w3(32'h3943d63d),
	.w4(32'hb7688925),
	.w5(32'hb8a4f634),
	.w6(32'h395f42df),
	.w7(32'h37747197),
	.w8(32'hb8420bf9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0517d8),
	.w1(32'hbbbf0eff),
	.w2(32'hbbb9c908),
	.w3(32'h39d12252),
	.w4(32'hbb0cfdb8),
	.w5(32'hba829c7f),
	.w6(32'hbb0fe999),
	.w7(32'hbaa5db93),
	.w8(32'hba0931c7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78af19),
	.w1(32'hbb9dd605),
	.w2(32'hbc2e882f),
	.w3(32'hb9d9c6f5),
	.w4(32'hbb8e7a34),
	.w5(32'hba55d470),
	.w6(32'hbb470187),
	.w7(32'hbbaf5018),
	.w8(32'h3a3a5ded),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398825d6),
	.w1(32'h3b3ffea1),
	.w2(32'h3b8da674),
	.w3(32'h3aacb6d8),
	.w4(32'h3915e7d0),
	.w5(32'h3b273fed),
	.w6(32'h3b433226),
	.w7(32'h3a8f9f2d),
	.w8(32'h3b412cd5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab93475),
	.w1(32'hbb52f654),
	.w2(32'hbb1f59ab),
	.w3(32'h3956c235),
	.w4(32'hba407dc4),
	.w5(32'hbacc140f),
	.w6(32'hba2c5fc2),
	.w7(32'h396cff99),
	.w8(32'hba7124b9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5466bf),
	.w1(32'hbb4205d9),
	.w2(32'hba119fe0),
	.w3(32'h3b942f83),
	.w4(32'hba02dc46),
	.w5(32'h3a8105d6),
	.w6(32'hb8d0940a),
	.w7(32'hba29a4f6),
	.w8(32'hba2b6679),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb540939),
	.w1(32'hbb43ab04),
	.w2(32'h39b8e573),
	.w3(32'hbaa788f4),
	.w4(32'hbabff300),
	.w5(32'hb9c87828),
	.w6(32'hba672b5d),
	.w7(32'hba446bb0),
	.w8(32'hbad6f46d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a0685),
	.w1(32'hbb204331),
	.w2(32'hbb033f9b),
	.w3(32'h3a293749),
	.w4(32'h3a6a59f2),
	.w5(32'hb9a93e58),
	.w6(32'hb9662fcd),
	.w7(32'h3a4dbb34),
	.w8(32'hb8f1ca83),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c371a),
	.w1(32'hb7e263c1),
	.w2(32'h337f1864),
	.w3(32'hb818ac7a),
	.w4(32'hb81cdfe3),
	.w5(32'hb7960fd4),
	.w6(32'hb753e5af),
	.w7(32'hb5ca765c),
	.w8(32'hb697f8d6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c77043),
	.w1(32'h381dbaeb),
	.w2(32'h38262571),
	.w3(32'h39009384),
	.w4(32'hb72c2e0b),
	.w5(32'hb802108b),
	.w6(32'h379c18f3),
	.w7(32'hb847ad49),
	.w8(32'hb808b239),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923a2c3),
	.w1(32'h39024453),
	.w2(32'h395c72e5),
	.w3(32'h38d48a9a),
	.w4(32'h3895938d),
	.w5(32'h38b09973),
	.w6(32'h394061dd),
	.w7(32'h391a5e6c),
	.w8(32'h3945cb06),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393fb6e6),
	.w1(32'h3997086c),
	.w2(32'h398b05cb),
	.w3(32'hb7d3485a),
	.w4(32'hb9e83706),
	.w5(32'hb9a8ef7b),
	.w6(32'h39529d24),
	.w7(32'hb9cba50d),
	.w8(32'hb9cea96c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e43a9e),
	.w1(32'h3adb528b),
	.w2(32'h3b619bb8),
	.w3(32'h39e0099d),
	.w4(32'hbb3a2435),
	.w5(32'h3b264637),
	.w6(32'h3a7156ff),
	.w7(32'hbaf3ae8c),
	.w8(32'h3b3a4efe),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984e1b0),
	.w1(32'h39bb7dbd),
	.w2(32'h3a2e1d11),
	.w3(32'h3917d5cd),
	.w4(32'h38d4afa7),
	.w5(32'h39cff5c1),
	.w6(32'h38afa832),
	.w7(32'h38f6850f),
	.w8(32'h3a0d87dd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3112d),
	.w1(32'h3a9c03da),
	.w2(32'h3a0e52cf),
	.w3(32'hba4262f5),
	.w4(32'hb9f05118),
	.w5(32'h3b2d4dad),
	.w6(32'h3a85eeb3),
	.w7(32'h3aa5954c),
	.w8(32'h3b983f6e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aa41e),
	.w1(32'hbba4382c),
	.w2(32'hbbcddb57),
	.w3(32'hbb0564c0),
	.w4(32'hbb3645e6),
	.w5(32'hbb5f6246),
	.w6(32'hbb3bfd3a),
	.w7(32'hbab9efa6),
	.w8(32'hbb1bf078),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2236b1),
	.w1(32'h3b13763f),
	.w2(32'h3b329949),
	.w3(32'hb9db8087),
	.w4(32'h398539db),
	.w5(32'hba1150ff),
	.w6(32'h3b35b4c3),
	.w7(32'hb9e79fea),
	.w8(32'hba53b755),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11a60e),
	.w1(32'hbb448281),
	.w2(32'hbacf5865),
	.w3(32'h3bb4191a),
	.w4(32'h3addc686),
	.w5(32'h3a767072),
	.w6(32'h3b9922fb),
	.w7(32'h3a83af0f),
	.w8(32'h3b3918b7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbaf77),
	.w1(32'h3b60652d),
	.w2(32'h3a9b9d37),
	.w3(32'h39ca1eef),
	.w4(32'h3b16bf2e),
	.w5(32'h39e2dd12),
	.w6(32'h3ab21d48),
	.w7(32'h3ac24af9),
	.w8(32'h3af5e400),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0f47c),
	.w1(32'hbc5e16f4),
	.w2(32'hbc091191),
	.w3(32'hb9bd41e6),
	.w4(32'hbbd9de06),
	.w5(32'hbb936f41),
	.w6(32'hbb60dabe),
	.w7(32'hbb463c85),
	.w8(32'hba020c78),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb729ee3),
	.w1(32'hbb18e9ef),
	.w2(32'h3a92bd50),
	.w3(32'h37e7c024),
	.w4(32'hbb3ace26),
	.w5(32'hba58f84e),
	.w6(32'hb98d5422),
	.w7(32'hba0c7d4a),
	.w8(32'h39174982),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80afa1),
	.w1(32'h3a32a971),
	.w2(32'h3b65c03b),
	.w3(32'hb975c79e),
	.w4(32'hbb8d22b0),
	.w5(32'hba2d9f74),
	.w6(32'h3a222625),
	.w7(32'hbb875242),
	.w8(32'hba8a2592),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e84b7),
	.w1(32'h3aa37a2a),
	.w2(32'h3a2b452c),
	.w3(32'h3997cd61),
	.w4(32'h3a8a1107),
	.w5(32'h39240eb0),
	.w6(32'h3a088710),
	.w7(32'h392f608c),
	.w8(32'hb8476d11),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34d5a1),
	.w1(32'hbb878e41),
	.w2(32'hbb3c06a4),
	.w3(32'hbb167a32),
	.w4(32'hba56f52f),
	.w5(32'hbb289e21),
	.w6(32'hbb227954),
	.w7(32'hba6eb437),
	.w8(32'hbb5f7209),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1c3d),
	.w1(32'hbbde8d79),
	.w2(32'hb8a7d1bf),
	.w3(32'h3b2428d9),
	.w4(32'hb9d59625),
	.w5(32'hbb169def),
	.w6(32'h393dadde),
	.w7(32'hba5fb0f3),
	.w8(32'hbae605a8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb565dbf),
	.w1(32'hbc2f22e8),
	.w2(32'hbbb1ba26),
	.w3(32'hbc05e3d5),
	.w4(32'hbc7c1ad4),
	.w5(32'h3c1a832a),
	.w6(32'hba32d6b4),
	.w7(32'hbbc74e1a),
	.w8(32'h3c8b901b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0650cb),
	.w1(32'h3a663123),
	.w2(32'h3b1ae36f),
	.w3(32'hbc03493b),
	.w4(32'hbbdf09dc),
	.w5(32'hba3d8a61),
	.w6(32'hbb574db6),
	.w7(32'hbbd2c4d2),
	.w8(32'hbaab588d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e21f8),
	.w1(32'h3b136a2f),
	.w2(32'h3b829712),
	.w3(32'hbb01ef4a),
	.w4(32'hba033b82),
	.w5(32'h3ac3e441),
	.w6(32'hb98c7f69),
	.w7(32'hbb4e7f1f),
	.w8(32'h38af76be),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1128f1),
	.w1(32'hbb69f8a3),
	.w2(32'h384f0944),
	.w3(32'h3bf49d2a),
	.w4(32'h3b9887ad),
	.w5(32'h3bc1f32e),
	.w6(32'h3b4797e7),
	.w7(32'h3a930b22),
	.w8(32'h3bd15e05),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0e99a),
	.w1(32'h3b2272d2),
	.w2(32'h3ae090a0),
	.w3(32'h39ec9927),
	.w4(32'h3b3227ac),
	.w5(32'h3ac4556b),
	.w6(32'h3abebee9),
	.w7(32'h3b01cfd8),
	.w8(32'h3aa6394d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc380cd3),
	.w1(32'hbc8a9796),
	.w2(32'hbc546430),
	.w3(32'hbbd00684),
	.w4(32'hbc54104a),
	.w5(32'h3bcee9fc),
	.w6(32'h3b2034d7),
	.w7(32'hbbd509b7),
	.w8(32'h3c6a66f3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a216aae),
	.w1(32'h3b3c3f1c),
	.w2(32'h3a37c143),
	.w3(32'h3b07af1b),
	.w4(32'h3ad2c3c9),
	.w5(32'h3b526fd4),
	.w6(32'h3b29a0ca),
	.w7(32'h3a09e3c5),
	.w8(32'h3ad66d69),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a04f44),
	.w1(32'h39053d76),
	.w2(32'h3911ae82),
	.w3(32'h39a48462),
	.w4(32'h39a3ba7e),
	.w5(32'h39194c46),
	.w6(32'h3a1a1874),
	.w7(32'h3987fb3c),
	.w8(32'h394f023f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb142ab1),
	.w1(32'hbb35950f),
	.w2(32'hbac8c636),
	.w3(32'hbaadef10),
	.w4(32'hbb1bc57c),
	.w5(32'hba198d84),
	.w6(32'hb9f72212),
	.w7(32'hbaf73868),
	.w8(32'hbadce39b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a627aa2),
	.w1(32'hb9e70fe4),
	.w2(32'h3a6f27ed),
	.w3(32'h3acb5dff),
	.w4(32'h3ac30935),
	.w5(32'hb9c000bc),
	.w6(32'h3aa0b32e),
	.w7(32'h3af65fd5),
	.w8(32'hb996e029),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16d67b),
	.w1(32'h3a03aa77),
	.w2(32'h3acfcaff),
	.w3(32'hbac80217),
	.w4(32'hbb090ed5),
	.w5(32'hba815873),
	.w6(32'hba425a75),
	.w7(32'hbb66b62b),
	.w8(32'hba7d5b95),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96a117),
	.w1(32'hbb72006a),
	.w2(32'hba1bea61),
	.w3(32'h38118f6e),
	.w4(32'hbb4a3e5c),
	.w5(32'hbba24907),
	.w6(32'h3aaeb706),
	.w7(32'hbad6ece8),
	.w8(32'hbb287dbb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12fa7c),
	.w1(32'hb9ad9738),
	.w2(32'h3af0d9e4),
	.w3(32'hbab87e3c),
	.w4(32'hbb1290a6),
	.w5(32'h3a85093f),
	.w6(32'hb9489d37),
	.w7(32'hbaaeb22f),
	.w8(32'h3a7b11e0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a795e),
	.w1(32'h3c110e8e),
	.w2(32'h3b9f7dc6),
	.w3(32'hbb45a766),
	.w4(32'h3b7624ca),
	.w5(32'h3bf9357c),
	.w6(32'h3b8a8475),
	.w7(32'h3aff6779),
	.w8(32'h3bfaa6a7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d7df),
	.w1(32'hbc43319a),
	.w2(32'hbb7c48f0),
	.w3(32'hbb8cc5e8),
	.w4(32'hbbe00d30),
	.w5(32'hba8ef0d1),
	.w6(32'hbb55a2d7),
	.w7(32'hbb0c2c82),
	.w8(32'hba16cc02),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7367b7),
	.w1(32'h3a6308a6),
	.w2(32'h3ae6a11d),
	.w3(32'hba7f3780),
	.w4(32'h39d0a13b),
	.w5(32'h3acbfa61),
	.w6(32'h3aaeaa6d),
	.w7(32'h3a34084f),
	.w8(32'h3afc7f8d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905228c),
	.w1(32'h3806a0fd),
	.w2(32'h38401661),
	.w3(32'hb87758c7),
	.w4(32'hb83d27ac),
	.w5(32'hb7ff8a75),
	.w6(32'hb8fa846f),
	.w7(32'hb91e36bb),
	.w8(32'hb913117f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a63d7),
	.w1(32'hba8c003b),
	.w2(32'hb9ea3701),
	.w3(32'hb9b8b73b),
	.w4(32'hba85cbac),
	.w5(32'h3a4e094f),
	.w6(32'hba0f022f),
	.w7(32'h39ca3d66),
	.w8(32'h3a6d7563),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e878a),
	.w1(32'hb7f97027),
	.w2(32'hb6773a11),
	.w3(32'h3709c79a),
	.w4(32'hb6852a57),
	.w5(32'h37847124),
	.w6(32'h37a0120c),
	.w7(32'h36a22875),
	.w8(32'h38208e48),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ff225),
	.w1(32'h3a8b9441),
	.w2(32'h3a91f02d),
	.w3(32'h3a45c6f6),
	.w4(32'h3a7a9b07),
	.w5(32'h3a5aadce),
	.w6(32'h3a1f0bcb),
	.w7(32'h39f90ec4),
	.w8(32'h3999eef2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec052a),
	.w1(32'h3b072245),
	.w2(32'h3b5e407e),
	.w3(32'h3a5c018c),
	.w4(32'h3b14fafb),
	.w5(32'h3b66addd),
	.w6(32'h3b308050),
	.w7(32'h3b213970),
	.w8(32'h3b7a03f1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86cde50),
	.w1(32'hb996e6ee),
	.w2(32'hb9836ad7),
	.w3(32'h39d6de1f),
	.w4(32'h3947b2fa),
	.w5(32'h3948fd54),
	.w6(32'h3a83fbce),
	.w7(32'h39fa3ae7),
	.w8(32'h395ea548),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2a1c8),
	.w1(32'hbab72681),
	.w2(32'hba6aeca1),
	.w3(32'h37c59140),
	.w4(32'h3ac65c1b),
	.w5(32'h3a8ef479),
	.w6(32'hbb0e5730),
	.w7(32'hb8aaff7d),
	.w8(32'hba212fcf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed5f5f),
	.w1(32'h3b66fbbb),
	.w2(32'h3bbf4978),
	.w3(32'h3a55ee84),
	.w4(32'hbb5da481),
	.w5(32'hbada058c),
	.w6(32'h3b1249fa),
	.w7(32'hbba2c83e),
	.w8(32'hbb2aede3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd34c9),
	.w1(32'h38a1e680),
	.w2(32'h36c58a5f),
	.w3(32'h38c19b73),
	.w4(32'hb812fcef),
	.w5(32'hb8d5380f),
	.w6(32'h388caec8),
	.w7(32'hb7e81bed),
	.w8(32'hb886502f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910f046),
	.w1(32'h3830cc60),
	.w2(32'hb8a762a6),
	.w3(32'h3913be62),
	.w4(32'hb8021eed),
	.w5(32'hb8a2757b),
	.w6(32'h392d4743),
	.w7(32'hb593eab2),
	.w8(32'hb90966db),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376c2f97),
	.w1(32'hb7a27d24),
	.w2(32'hb6890995),
	.w3(32'h380683b0),
	.w4(32'h370b2739),
	.w5(32'h3867acfb),
	.w6(32'h37c251bf),
	.w7(32'h38066a6e),
	.w8(32'h38ca754a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a61701),
	.w1(32'h39bf15e5),
	.w2(32'h39e969d2),
	.w3(32'h3a1dfb74),
	.w4(32'h3a1b7047),
	.w5(32'h39fb1040),
	.w6(32'h3a41cacc),
	.w7(32'h3a4424f5),
	.w8(32'h39d833fe),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80539f),
	.w1(32'h3c0be476),
	.w2(32'hba336606),
	.w3(32'hb9c2f93e),
	.w4(32'h3b224642),
	.w5(32'h391ced70),
	.w6(32'h3b4aae05),
	.w7(32'hb9c84b9e),
	.w8(32'h3948c3bc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5c7cb),
	.w1(32'hbb841775),
	.w2(32'hbb0e4cdf),
	.w3(32'h39a62240),
	.w4(32'hbaeb3670),
	.w5(32'hba0889d5),
	.w6(32'hbaf0a76f),
	.w7(32'h3a845f07),
	.w8(32'hba2d4a2a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d52f8e),
	.w1(32'hbac8c5ee),
	.w2(32'hba80f3dd),
	.w3(32'h39a79178),
	.w4(32'hb9eb6a9e),
	.w5(32'hb9c00f29),
	.w6(32'h37eb627d),
	.w7(32'h390ea684),
	.w8(32'h39074a76),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42a1fc),
	.w1(32'hba3ead9f),
	.w2(32'hba80a1b4),
	.w3(32'hba99404e),
	.w4(32'hbacbcbb6),
	.w5(32'h37b6e5e0),
	.w6(32'hb981cd7c),
	.w7(32'hb9430efa),
	.w8(32'h3abfc195),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63ff84),
	.w1(32'hb9a3aaa0),
	.w2(32'h3a517893),
	.w3(32'h399e569e),
	.w4(32'hb94be605),
	.w5(32'h3a97270b),
	.w6(32'h3a56e73b),
	.w7(32'h39e38c3b),
	.w8(32'h3aa1609a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba440526),
	.w1(32'hbb23fc5f),
	.w2(32'hbadea922),
	.w3(32'h384e19a4),
	.w4(32'hba78474d),
	.w5(32'hba91a538),
	.w6(32'hb8b4a065),
	.w7(32'h3a65f833),
	.w8(32'h3a22a68f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4da31),
	.w1(32'hbbb1c2e1),
	.w2(32'hbac224eb),
	.w3(32'hbad97a1c),
	.w4(32'hbb8c2a3e),
	.w5(32'hba863ea0),
	.w6(32'hba8c319a),
	.w7(32'hbae7501f),
	.w8(32'hb904e5e5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66ab2b),
	.w1(32'hbbe13693),
	.w2(32'hbbc42760),
	.w3(32'hb8641bab),
	.w4(32'h39de8b25),
	.w5(32'hbaefed65),
	.w6(32'hbbb58077),
	.w7(32'hbb02960f),
	.w8(32'hbb527473),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c6a59),
	.w1(32'h3aac15f4),
	.w2(32'h3b55c9d8),
	.w3(32'hba8c7e8a),
	.w4(32'hbb26f345),
	.w5(32'h39422383),
	.w6(32'h39b714c5),
	.w7(32'hbaff2245),
	.w8(32'h3a2a7b0b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba33308),
	.w1(32'hbb949d4c),
	.w2(32'hba94f4f1),
	.w3(32'hbadbab5d),
	.w4(32'hba19a9b1),
	.w5(32'h39b8e50f),
	.w6(32'hba93d711),
	.w7(32'hbb015e4f),
	.w8(32'hb979caae),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91f9e4),
	.w1(32'hbb4caf79),
	.w2(32'hbb765d2a),
	.w3(32'h3a8dd910),
	.w4(32'h3b38f09a),
	.w5(32'h39c48cb6),
	.w6(32'h39639235),
	.w7(32'h3b578de9),
	.w8(32'hba41cd16),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918895c),
	.w1(32'h3b4d9ca6),
	.w2(32'h3b1a914a),
	.w3(32'hba890b4b),
	.w4(32'h3a13dad0),
	.w5(32'h3b90d5ca),
	.w6(32'h3b031b78),
	.w7(32'hb9b99dd0),
	.w8(32'h3bbfa5c2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d421ee),
	.w1(32'hbb2bb65d),
	.w2(32'hba26a232),
	.w3(32'hb76d9fa5),
	.w4(32'h39e05093),
	.w5(32'h3ad806ac),
	.w6(32'h3817690d),
	.w7(32'h3a83fc2a),
	.w8(32'h39bfbbd5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f3c04),
	.w1(32'hb838b2e9),
	.w2(32'h39f27d8b),
	.w3(32'hb9a59681),
	.w4(32'hb60a8f4f),
	.w5(32'h3a094c16),
	.w6(32'hb65ece74),
	.w7(32'h38ddb5cc),
	.w8(32'h39e47b9f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c3f03),
	.w1(32'hbb48e002),
	.w2(32'h3bb0a030),
	.w3(32'hb9c5d575),
	.w4(32'hbbc4dd93),
	.w5(32'hbb9f41b1),
	.w6(32'h3b48dadf),
	.w7(32'hbb8fb6b6),
	.w8(32'hbba8ebda),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1116a9),
	.w1(32'hbaa6bfbd),
	.w2(32'hba7f18db),
	.w3(32'hba9fa110),
	.w4(32'hbac3d8eb),
	.w5(32'hb984a4bb),
	.w6(32'hbabbc493),
	.w7(32'hba5e4f04),
	.w8(32'h3953bb06),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921af3e),
	.w1(32'hb9503b38),
	.w2(32'hb8af44af),
	.w3(32'hb9874df1),
	.w4(32'hb8fe8e2b),
	.w5(32'hb99e02b1),
	.w6(32'h3828170d),
	.w7(32'hb7ab7dd7),
	.w8(32'hb8affd90),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad89f4),
	.w1(32'hb8f4f3a8),
	.w2(32'h38fb4b58),
	.w3(32'h38afad27),
	.w4(32'h3864b400),
	.w5(32'h3875a374),
	.w6(32'h36240c7c),
	.w7(32'hb781dfb5),
	.w8(32'hb7f28164),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca0fac),
	.w1(32'h39c90d63),
	.w2(32'h398a9b9f),
	.w3(32'h39a26f51),
	.w4(32'hba245a73),
	.w5(32'h3aa7e7c2),
	.w6(32'h39f78969),
	.w7(32'hba3b839f),
	.w8(32'h3a685e73),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a202771),
	.w1(32'h3b619fda),
	.w2(32'h3ad9353b),
	.w3(32'h3ac12260),
	.w4(32'hbae20abd),
	.w5(32'h3b0660e1),
	.w6(32'hb9571aed),
	.w7(32'hbb716b16),
	.w8(32'h3af789c8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39540207),
	.w1(32'hba4fa14d),
	.w2(32'h3a17fb60),
	.w3(32'h3a6d6b5b),
	.w4(32'h3a6315a6),
	.w5(32'h3a70689a),
	.w6(32'h3b0f3390),
	.w7(32'h3ae18964),
	.w8(32'h3ac7535a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b549e5),
	.w1(32'hb88e7785),
	.w2(32'hb7ce125f),
	.w3(32'hb8cfd674),
	.w4(32'hb876c48f),
	.w5(32'hb80e623c),
	.w6(32'hb855ec77),
	.w7(32'hb833fabb),
	.w8(32'hb7d97c18),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac12ea4),
	.w1(32'hbb7a7e95),
	.w2(32'hb9a31beb),
	.w3(32'h369525ab),
	.w4(32'hb857dba9),
	.w5(32'hb63b06f8),
	.w6(32'hbacf8c67),
	.w7(32'hb9037715),
	.w8(32'hba99c509),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba954aa6),
	.w1(32'hbac49dfa),
	.w2(32'h39aa99ec),
	.w3(32'hba7111ea),
	.w4(32'hbaee5a81),
	.w5(32'hba0f86ce),
	.w6(32'hba148b1c),
	.w7(32'hbaa21e65),
	.w8(32'hbaa708f5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861907),
	.w1(32'hbba07d42),
	.w2(32'hbbab1fac),
	.w3(32'h3ba2037a),
	.w4(32'h3b86f97c),
	.w5(32'h3ac50080),
	.w6(32'hbb0146c5),
	.w7(32'h37225164),
	.w8(32'h3adf8ab9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb94b3f),
	.w1(32'hbb954182),
	.w2(32'h3bdf293c),
	.w3(32'h3b0b0228),
	.w4(32'hbb83fda9),
	.w5(32'h39aa8f16),
	.w6(32'h3961034b),
	.w7(32'hbaa286c4),
	.w8(32'hbb7d6f07),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39350db5),
	.w1(32'h397367b6),
	.w2(32'hb9f88cfb),
	.w3(32'h399867b1),
	.w4(32'hbacfb4d7),
	.w5(32'hbacac764),
	.w6(32'h39c8eb57),
	.w7(32'hbae78f21),
	.w8(32'hbaf21d50),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0eec0),
	.w1(32'h3b1795d5),
	.w2(32'h3b06ff97),
	.w3(32'h39117452),
	.w4(32'h3ad212cf),
	.w5(32'h3aed617f),
	.w6(32'h3a609d49),
	.w7(32'h3aad08c8),
	.w8(32'h3a87e3d8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02608f),
	.w1(32'h3a937e3b),
	.w2(32'h3b26e3e5),
	.w3(32'hbab119f5),
	.w4(32'hbab7aa15),
	.w5(32'h3ac166a3),
	.w6(32'hb8dc2a0a),
	.w7(32'hba70350d),
	.w8(32'h3af1c68b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9356eb),
	.w1(32'hba98313e),
	.w2(32'h3a47b711),
	.w3(32'hbac7be7e),
	.w4(32'hbb40bf75),
	.w5(32'h3a882d9a),
	.w6(32'h3a3f19da),
	.w7(32'hbad45d46),
	.w8(32'h3a30bb77),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab33ec2),
	.w1(32'h3b3736b8),
	.w2(32'h3b4261c3),
	.w3(32'h3adc33bf),
	.w4(32'h3a48ed38),
	.w5(32'h3a967915),
	.w6(32'h3ae0ea85),
	.w7(32'hb91d5444),
	.w8(32'h3a4e742d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba428a),
	.w1(32'hbae9babe),
	.w2(32'hba902be4),
	.w3(32'h39fd1887),
	.w4(32'h3a4d17bb),
	.w5(32'hb9254aee),
	.w6(32'hb9fd5ad8),
	.w7(32'hb992df7e),
	.w8(32'hb95389a5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38177f2c),
	.w1(32'h3993341b),
	.w2(32'h39acbfaf),
	.w3(32'h390ed85d),
	.w4(32'h3a07dbf8),
	.w5(32'h395fbae5),
	.w6(32'h39308067),
	.w7(32'h39f329b7),
	.w8(32'h38d7b06b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995b47e),
	.w1(32'hbb6b3e8a),
	.w2(32'h39750470),
	.w3(32'hba532b4b),
	.w4(32'hb9ea4e9e),
	.w5(32'h3a4f6560),
	.w6(32'hb9d71f9e),
	.w7(32'h39a51c8c),
	.w8(32'h39aa4656),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8df17),
	.w1(32'h3a80a0b3),
	.w2(32'hb9892fb7),
	.w3(32'h3b0270ae),
	.w4(32'h3a623230),
	.w5(32'hb9fa821d),
	.w6(32'h39df99f9),
	.w7(32'hb795b345),
	.w8(32'hba08ecc0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35869c),
	.w1(32'hb8b76635),
	.w2(32'h3b98badf),
	.w3(32'hbb6a8f4c),
	.w4(32'hbafc9e2e),
	.w5(32'h3a915952),
	.w6(32'h39b657b3),
	.w7(32'hb9c862d0),
	.w8(32'h39c9c080),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ef54),
	.w1(32'h3984932a),
	.w2(32'hb8dc54d4),
	.w3(32'h3a266811),
	.w4(32'h39af3133),
	.w5(32'h3917be4c),
	.w6(32'h395d5dbc),
	.w7(32'h399df63a),
	.w8(32'h39985d87),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ba69a),
	.w1(32'h3b8dce37),
	.w2(32'h3b162bbf),
	.w3(32'h3baa4a8e),
	.w4(32'h3a06a607),
	.w5(32'hbb437bc2),
	.w6(32'h3b84b8c8),
	.w7(32'hbaf11aef),
	.w8(32'hbb719e50),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a61de4),
	.w1(32'h394eb9b1),
	.w2(32'h39bcc796),
	.w3(32'h37ef05c7),
	.w4(32'h396e9305),
	.w5(32'h39b67fe2),
	.w6(32'h39605fd5),
	.w7(32'h39bd6e86),
	.w8(32'h39b00bd9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39051bd0),
	.w1(32'h3720ef68),
	.w2(32'hba2868b8),
	.w3(32'h38f34f4e),
	.w4(32'h38883b90),
	.w5(32'hb9c2d441),
	.w6(32'h38a7273b),
	.w7(32'h389eaa89),
	.w8(32'hb9817626),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab00d0),
	.w1(32'hba462b76),
	.w2(32'h3a7d5d0a),
	.w3(32'h3a94995a),
	.w4(32'hba05672b),
	.w5(32'h3a482eff),
	.w6(32'h3a0e33fe),
	.w7(32'hba8d000a),
	.w8(32'h39fbf324),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f91e4),
	.w1(32'h3ae47694),
	.w2(32'hbb069834),
	.w3(32'hbb98089e),
	.w4(32'h3a7e1129),
	.w5(32'h3b1389c7),
	.w6(32'hbb41abf4),
	.w7(32'hbb157096),
	.w8(32'h3b23d711),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad19ef5),
	.w1(32'h3a9bfd83),
	.w2(32'h3a24ea33),
	.w3(32'h3ad79912),
	.w4(32'h3a927ead),
	.w5(32'h3a1b68a7),
	.w6(32'h3b06fef7),
	.w7(32'h3aebeae5),
	.w8(32'h3a907644),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fed4cd),
	.w1(32'h3aa4800a),
	.w2(32'h3b160474),
	.w3(32'hb93b0518),
	.w4(32'hb9f6aa69),
	.w5(32'hba5d4034),
	.w6(32'h3b25af58),
	.w7(32'h39abe1f5),
	.w8(32'h39bfc5e3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a124a90),
	.w1(32'hbaf5fc12),
	.w2(32'hba141cbc),
	.w3(32'h3abf6b82),
	.w4(32'hba997a37),
	.w5(32'hbb093d2c),
	.w6(32'hbaacbcf9),
	.w7(32'h3a4b95e7),
	.w8(32'hbad94d91),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeadad),
	.w1(32'hbbd51507),
	.w2(32'h3a9201ec),
	.w3(32'hbadecf50),
	.w4(32'hba939058),
	.w5(32'hbae1333e),
	.w6(32'hb9c81079),
	.w7(32'h3aaecda7),
	.w8(32'hbbc6d311),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5507c0),
	.w1(32'hbbd84e86),
	.w2(32'hbba3347e),
	.w3(32'h3aa70c90),
	.w4(32'hbab97ade),
	.w5(32'hb9a31888),
	.w6(32'hb9214ebc),
	.w7(32'hb962a3c8),
	.w8(32'h3a430939),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94824d),
	.w1(32'hbb9223d2),
	.w2(32'hbb2eba12),
	.w3(32'hbb397fb7),
	.w4(32'hba6be985),
	.w5(32'hbaca8798),
	.w6(32'hbb54fe09),
	.w7(32'hba5bbdb0),
	.w8(32'hbb42b6a7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947c53),
	.w1(32'h3a47e119),
	.w2(32'h3a6770c9),
	.w3(32'h3a6c5761),
	.w4(32'h3aa24dbe),
	.w5(32'h3aa2362f),
	.w6(32'h3a1c260b),
	.w7(32'h3a8b1f37),
	.w8(32'h3aba5133),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafedcaa),
	.w1(32'hbb51e01a),
	.w2(32'hb9871a30),
	.w3(32'h38cf6a03),
	.w4(32'hba9c0a2c),
	.w5(32'hba188f17),
	.w6(32'hbb1e8864),
	.w7(32'hb935b56a),
	.w8(32'hb9cb7a21),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798026b),
	.w1(32'hb65111b4),
	.w2(32'h37d37460),
	.w3(32'h3807481b),
	.w4(32'h365f739d),
	.w5(32'h370dac70),
	.w6(32'h3861be8a),
	.w7(32'h37bcd8e4),
	.w8(32'h3756b8c2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba219ea6),
	.w1(32'hba0148cb),
	.w2(32'h396e04ff),
	.w3(32'hb8e93df1),
	.w4(32'h39fe3ae7),
	.w5(32'h3a06b27b),
	.w6(32'hb92cedb7),
	.w7(32'h3a0a7a0e),
	.w8(32'h398052d7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9444edf),
	.w1(32'h39a009e2),
	.w2(32'h396c0765),
	.w3(32'h38f33159),
	.w4(32'hb9815cd2),
	.w5(32'hba067046),
	.w6(32'h38226b66),
	.w7(32'hba03c731),
	.w8(32'hba149247),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e56fe),
	.w1(32'hbbc9c9d8),
	.w2(32'hbaf2aa92),
	.w3(32'hba413018),
	.w4(32'hbb0a9b75),
	.w5(32'hbae278d1),
	.w6(32'hb9da075f),
	.w7(32'h3a8230f0),
	.w8(32'hb9a54421),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bb9217),
	.w1(32'h36a21048),
	.w2(32'h36f196fa),
	.w3(32'hb7082f2d),
	.w4(32'hb6b61a1d),
	.w5(32'h378bf45f),
	.w6(32'h36c06b19),
	.w7(32'h361cbd22),
	.w8(32'h37d5d9d9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf7fac),
	.w1(32'hb9fcf146),
	.w2(32'hb989f2ff),
	.w3(32'hb9800d22),
	.w4(32'hb98aedf2),
	.w5(32'hb9869442),
	.w6(32'hb9957740),
	.w7(32'hb99ed0c0),
	.w8(32'hb95a2a83),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e04bb),
	.w1(32'h3a2453c5),
	.w2(32'h3aa4474e),
	.w3(32'h39ca7d48),
	.w4(32'hbabbefd4),
	.w5(32'hb9dc5ba7),
	.w6(32'h39da1d55),
	.w7(32'hbacddf50),
	.w8(32'h39ef3e20),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145456),
	.w1(32'hbba44565),
	.w2(32'h3aeb85e0),
	.w3(32'h3bb89066),
	.w4(32'hb99ffb5c),
	.w5(32'h3b3bf564),
	.w6(32'h3bebe6ff),
	.w7(32'h391ce373),
	.w8(32'h3849a883),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a18c1),
	.w1(32'hbb284317),
	.w2(32'hbaead887),
	.w3(32'hbb814064),
	.w4(32'hbb5116e6),
	.w5(32'h3b9971c2),
	.w6(32'hbb26bdbe),
	.w7(32'hbb09c86c),
	.w8(32'h3c000708),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f90a0),
	.w1(32'hba72c354),
	.w2(32'hbabb78cd),
	.w3(32'hb9c549ce),
	.w4(32'hba3c5552),
	.w5(32'hbaa20652),
	.w6(32'h39bb6639),
	.w7(32'hba25649d),
	.w8(32'hba08f57f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f015c),
	.w1(32'hbbb440f5),
	.w2(32'hbb76a694),
	.w3(32'hbb0aff09),
	.w4(32'hbb0132fc),
	.w5(32'hbb93c16c),
	.w6(32'hbb3201fb),
	.w7(32'hbb452b63),
	.w8(32'hbc081e6e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16200e),
	.w1(32'hbbcfa86c),
	.w2(32'h3beb1a8b),
	.w3(32'h3a876e06),
	.w4(32'hbb8d3311),
	.w5(32'h3a228fad),
	.w6(32'hbb4d9133),
	.w7(32'hb97d857b),
	.w8(32'hbb249601),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd28a4),
	.w1(32'hba4afa03),
	.w2(32'hba8e702c),
	.w3(32'h3a9393f2),
	.w4(32'h37b2ce81),
	.w5(32'hba5e88fc),
	.w6(32'h3a3b163f),
	.w7(32'hb9ead6ee),
	.w8(32'hbab6437b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d1f54),
	.w1(32'hb89ef294),
	.w2(32'hb89c1ca7),
	.w3(32'hb8c2c170),
	.w4(32'hb8d10f0e),
	.w5(32'hb8b044f2),
	.w6(32'hb847a25b),
	.w7(32'hb87db370),
	.w8(32'hb8e4eb12),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e9d00),
	.w1(32'hba2dd873),
	.w2(32'hba1173de),
	.w3(32'hba212890),
	.w4(32'hba3b1be5),
	.w5(32'hba59e4f7),
	.w6(32'hba09a2d2),
	.w7(32'hba1eeb26),
	.w8(32'hba4d574f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38420814),
	.w1(32'h3756d1b2),
	.w2(32'hb7831384),
	.w3(32'h38263657),
	.w4(32'h36b43266),
	.w5(32'hb7d16d2b),
	.w6(32'h37a033da),
	.w7(32'hb70206be),
	.w8(32'hb7160bf3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939f48),
	.w1(32'h3b17ed7a),
	.w2(32'hb994ea75),
	.w3(32'h39c07177),
	.w4(32'h3ac9555a),
	.w5(32'hba2e9934),
	.w6(32'h3a8a5aed),
	.w7(32'hbaed14b3),
	.w8(32'hbaf37eb5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919ca0d),
	.w1(32'hba85b504),
	.w2(32'hbaa56cb2),
	.w3(32'hba88f4c1),
	.w4(32'hba02f5d8),
	.w5(32'h3a2a04b0),
	.w6(32'h3a903fdf),
	.w7(32'h3a176255),
	.w8(32'h3ac00386),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4c8c4),
	.w1(32'h3b0cf9c8),
	.w2(32'h3b5b29f8),
	.w3(32'h3b2721b7),
	.w4(32'hba314e2c),
	.w5(32'h3b3e7f81),
	.w6(32'h3a149b90),
	.w7(32'hbac338bd),
	.w8(32'h3b1965f0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38249ca5),
	.w1(32'h3992cf54),
	.w2(32'h3a388c27),
	.w3(32'hb97248eb),
	.w4(32'h39d0bde8),
	.w5(32'h3a765233),
	.w6(32'h3a2748c8),
	.w7(32'h39b4c86f),
	.w8(32'h3a820488),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d88b29),
	.w1(32'hbb9474e4),
	.w2(32'hbb876e1f),
	.w3(32'h3a8f8372),
	.w4(32'hbb2810e9),
	.w5(32'hbb7ee9ad),
	.w6(32'h3aeb2d20),
	.w7(32'hba0ff68c),
	.w8(32'hbade7c88),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3046),
	.w1(32'hbc182a05),
	.w2(32'hbbd7a293),
	.w3(32'hbb4ed906),
	.w4(32'hbbbcb6a6),
	.w5(32'hbada98e8),
	.w6(32'hbae27360),
	.w7(32'hbace34e3),
	.w8(32'h3afdd52c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae0e47),
	.w1(32'h3b347d8a),
	.w2(32'h3a0d21ec),
	.w3(32'h3b8d2702),
	.w4(32'h3b1688d1),
	.w5(32'h3a0e4e82),
	.w6(32'h3c12ece4),
	.w7(32'h3ad07c0b),
	.w8(32'h3be67305),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade60dc),
	.w1(32'h3b9a21a5),
	.w2(32'h3b00b6b7),
	.w3(32'h3b1a045b),
	.w4(32'h3c1ab768),
	.w5(32'h3bc3febb),
	.w6(32'h3be55cf7),
	.w7(32'h3c19ccdc),
	.w8(32'h3c019f8e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac560a1),
	.w1(32'hba636629),
	.w2(32'h3af3481b),
	.w3(32'h3ac48f7d),
	.w4(32'hba8426a5),
	.w5(32'h3adaeaf3),
	.w6(32'h3bb557bf),
	.w7(32'hba5417e8),
	.w8(32'h3aa8cc55),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54581f),
	.w1(32'h3af71a6c),
	.w2(32'hbb1c31be),
	.w3(32'h39a3357d),
	.w4(32'h3bdcd05d),
	.w5(32'h3b21307f),
	.w6(32'hba7e2643),
	.w7(32'hb9ef4ee1),
	.w8(32'hbb0bceea),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8830b86),
	.w1(32'hbb3c89f2),
	.w2(32'hba09c978),
	.w3(32'h3b2f7178),
	.w4(32'hb799802f),
	.w5(32'h3bc62fa4),
	.w6(32'h3a85c883),
	.w7(32'h3b421378),
	.w8(32'h3bcbf1ff),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937608f),
	.w1(32'h38b034a2),
	.w2(32'hba8af432),
	.w3(32'h3c01e2fd),
	.w4(32'h3b13b489),
	.w5(32'h3be9cd0c),
	.w6(32'h3bb370a9),
	.w7(32'hba445029),
	.w8(32'h3b049ab5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61bc30),
	.w1(32'hbb878620),
	.w2(32'hbb803975),
	.w3(32'hbb95c821),
	.w4(32'hb871af43),
	.w5(32'hbbc83dc2),
	.w6(32'hbbbd554c),
	.w7(32'h3af37972),
	.w8(32'hbb7497d1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95366c),
	.w1(32'h3b855d53),
	.w2(32'h3bba8ff5),
	.w3(32'hba9dd169),
	.w4(32'h3b993e53),
	.w5(32'h3aefd654),
	.w6(32'h3b6d642c),
	.w7(32'h3a905c1c),
	.w8(32'h3b3f55d1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaf39d),
	.w1(32'hbb9ea67c),
	.w2(32'hbbc60660),
	.w3(32'hbb812c3e),
	.w4(32'hbb89fd1e),
	.w5(32'hbb64d4b5),
	.w6(32'hbbddb8cf),
	.w7(32'hbb68681f),
	.w8(32'hbbac413c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc283bb),
	.w1(32'h3c19f42f),
	.w2(32'h3bc1af4a),
	.w3(32'hbb907f61),
	.w4(32'h3b55cca3),
	.w5(32'hbb63e70e),
	.w6(32'hbb8c6bd6),
	.w7(32'h3b84fe48),
	.w8(32'hb95710e8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc1eb2),
	.w1(32'hbb98adef),
	.w2(32'hbbc40666),
	.w3(32'hbb7e4e4f),
	.w4(32'hbb4e35b3),
	.w5(32'hbaa08b34),
	.w6(32'hbb326c19),
	.w7(32'hbae62698),
	.w8(32'hbb28c457),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9939),
	.w1(32'h3a794d2c),
	.w2(32'hbb50c3d8),
	.w3(32'hbb7986ed),
	.w4(32'hbb58b331),
	.w5(32'hbb806c86),
	.w6(32'hbb559c7a),
	.w7(32'hbb60f9d6),
	.w8(32'hb9ef624a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a011b1d),
	.w1(32'h3bb384f0),
	.w2(32'hbb940c8c),
	.w3(32'hbb236734),
	.w4(32'h3b604849),
	.w5(32'hbbf2fee9),
	.w6(32'h3ada9e19),
	.w7(32'h38976aed),
	.w8(32'hbb7fc11e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc654a47),
	.w1(32'hba9a8e81),
	.w2(32'hba1349e4),
	.w3(32'hbc88cc9e),
	.w4(32'h3a929177),
	.w5(32'h3bf1b7d5),
	.w6(32'hbc937ae5),
	.w7(32'hbb27c2d9),
	.w8(32'h3a2600fa),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1119d7),
	.w1(32'hbb826534),
	.w2(32'h3b8fd687),
	.w3(32'hbb05a825),
	.w4(32'hbb496506),
	.w5(32'h3c1d184b),
	.w6(32'h3ae2dd34),
	.w7(32'h3c117531),
	.w8(32'h3c3d5e58),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4e616),
	.w1(32'h3a53409c),
	.w2(32'hb94ef3e7),
	.w3(32'h3c1661c6),
	.w4(32'h3b06a1ba),
	.w5(32'hb91ec357),
	.w6(32'h3bca6278),
	.w7(32'hbab04d79),
	.w8(32'hbb3ccf23),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39325952),
	.w1(32'h38d55a34),
	.w2(32'hbb0d822a),
	.w3(32'hbb2420b9),
	.w4(32'hbb399e74),
	.w5(32'hbb989212),
	.w6(32'hbb2e2ea5),
	.w7(32'h395bac4d),
	.w8(32'h393de78b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9939e1),
	.w1(32'hbc02aa70),
	.w2(32'hbbb71760),
	.w3(32'hbb26b4c9),
	.w4(32'hbae5eb56),
	.w5(32'hb948cf59),
	.w6(32'h3986940b),
	.w7(32'hbbf20934),
	.w8(32'hbba73c3c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977208c),
	.w1(32'h3bef6194),
	.w2(32'hbab03b6b),
	.w3(32'hbc0aedec),
	.w4(32'hb9460883),
	.w5(32'h3c726f62),
	.w6(32'hbb8ada84),
	.w7(32'hbc23f8ac),
	.w8(32'h3b6949ed),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ed54d),
	.w1(32'hbbd142dc),
	.w2(32'hbb886c4e),
	.w3(32'h3c05d235),
	.w4(32'h3addae52),
	.w5(32'h3b8d351d),
	.w6(32'h3b6c86e8),
	.w7(32'hbab5ab0a),
	.w8(32'hba185925),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba754ed),
	.w1(32'hba5732c8),
	.w2(32'hbbb15ec0),
	.w3(32'hbb397c20),
	.w4(32'hb9ab2914),
	.w5(32'h3b03fb60),
	.w6(32'hbbb6d28d),
	.w7(32'hbb846a41),
	.w8(32'h3bbf9cbf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cb053),
	.w1(32'h3bf5d36c),
	.w2(32'h3c3c88c1),
	.w3(32'hbc0dcc59),
	.w4(32'hbac20ee8),
	.w5(32'h3b6c8043),
	.w6(32'hbb8956fa),
	.w7(32'h3ace3b40),
	.w8(32'h3bb0e739),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8352c0),
	.w1(32'h3b08f85a),
	.w2(32'h3bb6f382),
	.w3(32'hba8c2713),
	.w4(32'hbb63fd27),
	.w5(32'hb8d3cb97),
	.w6(32'h3b6cfb01),
	.w7(32'hbb03ef70),
	.w8(32'hbb7d954c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a50a9),
	.w1(32'h3a021617),
	.w2(32'hbbb77edd),
	.w3(32'h3af92855),
	.w4(32'hbae11293),
	.w5(32'hbc16669e),
	.w6(32'hbb1f767e),
	.w7(32'hbc017732),
	.w8(32'hbbeb4b5a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe8df7),
	.w1(32'hbbff43cb),
	.w2(32'hbbc7ffca),
	.w3(32'hbb8d3d7f),
	.w4(32'hbc099f63),
	.w5(32'hbbe2553b),
	.w6(32'hbab0d127),
	.w7(32'hbbcb1675),
	.w8(32'hbb72bc05),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba065c4),
	.w1(32'h3b43ce69),
	.w2(32'h3b9b7a97),
	.w3(32'h3ada944d),
	.w4(32'h37260e38),
	.w5(32'h3b883752),
	.w6(32'h3a12fe29),
	.w7(32'h3a8bcaef),
	.w8(32'hbb3ffd33),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e66217),
	.w1(32'h3a91fd2f),
	.w2(32'h3c519317),
	.w3(32'hbb2541ae),
	.w4(32'hbbe83460),
	.w5(32'h3cd705cc),
	.w6(32'hbb950a5f),
	.w7(32'hbace9f32),
	.w8(32'h3c884af5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c827e),
	.w1(32'h3c7c01cf),
	.w2(32'h3c187a40),
	.w3(32'h3c853552),
	.w4(32'h3cf99782),
	.w5(32'h3d3522cb),
	.w6(32'h3bd01e70),
	.w7(32'h3b893d53),
	.w8(32'h3bbe53f3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdd33d),
	.w1(32'hbb69b1f7),
	.w2(32'hbb9dd939),
	.w3(32'h3bea46d0),
	.w4(32'h3a2a2449),
	.w5(32'h39bf9764),
	.w6(32'hbb524113),
	.w7(32'hbb0840ce),
	.w8(32'hbb724b4c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dcbc0),
	.w1(32'h38ed9eaf),
	.w2(32'h3a86406c),
	.w3(32'hbc1ff4ea),
	.w4(32'h3ac63bfe),
	.w5(32'h3b3980cf),
	.w6(32'hbc209d96),
	.w7(32'h394aff9b),
	.w8(32'h3a27d9ce),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b68fa3),
	.w1(32'h3a2e51ea),
	.w2(32'h3b122f94),
	.w3(32'h3a8c75fd),
	.w4(32'hbaed7858),
	.w5(32'h3c493e95),
	.w6(32'hbb11ea93),
	.w7(32'hba921307),
	.w8(32'h3bcaa072),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec822a),
	.w1(32'hb737be40),
	.w2(32'hbb9614c8),
	.w3(32'hbb10dbce),
	.w4(32'h3bac9771),
	.w5(32'h3b69e118),
	.w6(32'h3a40a0d9),
	.w7(32'hbb9111cf),
	.w8(32'h3b81c2f7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2b0c0),
	.w1(32'hba1ceceb),
	.w2(32'hba4cbc53),
	.w3(32'h3a4591a0),
	.w4(32'h3ab1b2c9),
	.w5(32'h3bc28051),
	.w6(32'hbb01d1ba),
	.w7(32'hb9a215e0),
	.w8(32'h3b3688f5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb190c22),
	.w1(32'h3b2a0689),
	.w2(32'h3a516980),
	.w3(32'h39b11f93),
	.w4(32'hba830e6f),
	.w5(32'hbb7e8e06),
	.w6(32'h3b1d6cce),
	.w7(32'hb9b2ce85),
	.w8(32'hbae92897),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de498),
	.w1(32'h3a9e639f),
	.w2(32'hbac43ba7),
	.w3(32'hba4ef13b),
	.w4(32'h3a8a588f),
	.w5(32'hbb06feba),
	.w6(32'h3aced105),
	.w7(32'h37fd5ccd),
	.w8(32'hbb553579),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ebec5),
	.w1(32'hbbaeff49),
	.w2(32'hbbb49edf),
	.w3(32'hbafc61b0),
	.w4(32'hbba0bd10),
	.w5(32'hbb925246),
	.w6(32'h39831177),
	.w7(32'h393e533c),
	.w8(32'hbb06237a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b542),
	.w1(32'h3be68a86),
	.w2(32'h3b7cc0d9),
	.w3(32'hbb0f5995),
	.w4(32'h3bb0e0ab),
	.w5(32'h3c5394a0),
	.w6(32'hbb0422ed),
	.w7(32'h3afcc5a8),
	.w8(32'h3c1e6a8e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e4f8),
	.w1(32'h3bf75a7e),
	.w2(32'h3bbdf049),
	.w3(32'hbaa6894e),
	.w4(32'h3ae3f111),
	.w5(32'h3b88212f),
	.w6(32'h3b61ae09),
	.w7(32'h3a5c46e8),
	.w8(32'h3b28f735),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5362c),
	.w1(32'hbac3049f),
	.w2(32'hba8bf1e7),
	.w3(32'hb9ec8c05),
	.w4(32'hbb7f30a1),
	.w5(32'hbb33b4d9),
	.w6(32'h39832fa5),
	.w7(32'hbaea472b),
	.w8(32'hbbec1ba4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe17fe7),
	.w1(32'hb9a35ea2),
	.w2(32'h3c0fa036),
	.w3(32'hbbf02298),
	.w4(32'h3be428f9),
	.w5(32'h3c96c83b),
	.w6(32'hbae8a2f5),
	.w7(32'h3b58f58b),
	.w8(32'h3ba061c5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7fe0),
	.w1(32'hbbe46324),
	.w2(32'hb937ba4f),
	.w3(32'h3c15c7ac),
	.w4(32'hbb5b6e01),
	.w5(32'hbb348d91),
	.w6(32'hbbaaae02),
	.w7(32'hbb715e79),
	.w8(32'hbbe88d33),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb887dcbb),
	.w1(32'hbbdfd7cb),
	.w2(32'hbb78f855),
	.w3(32'h3a6ca7c0),
	.w4(32'hbbf93fb9),
	.w5(32'hbb8b4897),
	.w6(32'h3baf7eab),
	.w7(32'hb9fe8e95),
	.w8(32'hba47fb63),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55be30),
	.w1(32'hbbf9c91c),
	.w2(32'hba6fdc00),
	.w3(32'hbb401b1a),
	.w4(32'hbb248113),
	.w5(32'hbb52b212),
	.w6(32'hbb24a345),
	.w7(32'hbb16b95e),
	.w8(32'hbaf87a3e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993b6d),
	.w1(32'h3c273368),
	.w2(32'h3bf36a4b),
	.w3(32'h3958598f),
	.w4(32'h3b5e6770),
	.w5(32'h3b0f0771),
	.w6(32'hbb88ba38),
	.w7(32'h3abd6396),
	.w8(32'h3b8a8b50),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95c6b1),
	.w1(32'hbb491bf1),
	.w2(32'hbb6eaf30),
	.w3(32'h3abe5c32),
	.w4(32'hb70cd38c),
	.w5(32'hbb9b36f8),
	.w6(32'h3b5c7827),
	.w7(32'hbad69759),
	.w8(32'hbbc0914e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d4137),
	.w1(32'hbb47d955),
	.w2(32'hbab704ac),
	.w3(32'hbb26dfdf),
	.w4(32'hbaac000d),
	.w5(32'h3b4dd224),
	.w6(32'hbafcde1d),
	.w7(32'hba35b0a0),
	.w8(32'h3b13086f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1fadd),
	.w1(32'h38a4fc9f),
	.w2(32'h3b00c45d),
	.w3(32'hbb9b90f1),
	.w4(32'hba4288b9),
	.w5(32'h3bf40342),
	.w6(32'hbb2e4f3a),
	.w7(32'hb95b7700),
	.w8(32'hba0d6a71),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bdf5d),
	.w1(32'hbbae7222),
	.w2(32'hba87a0b4),
	.w3(32'h3bbd7c22),
	.w4(32'hbae1ee6f),
	.w5(32'hbae9a0fd),
	.w6(32'hbac112cd),
	.w7(32'h3b8d626e),
	.w8(32'h3bb2c49c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba77208),
	.w1(32'h3b5c6d2b),
	.w2(32'hbb3023a4),
	.w3(32'hba5e2adc),
	.w4(32'h3a543421),
	.w5(32'hbb9d189a),
	.w6(32'hb957abfa),
	.w7(32'h3b10ede3),
	.w8(32'hba473d30),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaee73),
	.w1(32'h3b49876c),
	.w2(32'h3b107ef7),
	.w3(32'h3b8ef9c6),
	.w4(32'h3b371bf4),
	.w5(32'h3b92d462),
	.w6(32'h3b8fd2e1),
	.w7(32'h3b03b654),
	.w8(32'h3b73aafa),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b99cb),
	.w1(32'hbc001063),
	.w2(32'hbc10f05a),
	.w3(32'hbbe890a8),
	.w4(32'hbad2dc48),
	.w5(32'hb9b490c9),
	.w6(32'hba5988ab),
	.w7(32'hbb8955a1),
	.w8(32'hbafe3830),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81efbf),
	.w1(32'hbb643135),
	.w2(32'hbaa84ea4),
	.w3(32'hbb29d4c5),
	.w4(32'hbb9dae9c),
	.w5(32'hbb928a6f),
	.w6(32'hbbd2740b),
	.w7(32'hbb809d69),
	.w8(32'hbbb8e636),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb349463),
	.w1(32'hbb5ef5bd),
	.w2(32'hbab06617),
	.w3(32'hbb84a7e0),
	.w4(32'hbba9703e),
	.w5(32'h3b8a04f0),
	.w6(32'hbb39e5c0),
	.w7(32'hbb637123),
	.w8(32'hbac6e759),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2f62),
	.w1(32'hbb849004),
	.w2(32'hbaa792a7),
	.w3(32'hb8bbe320),
	.w4(32'hbb99ef18),
	.w5(32'hbb3ab6bf),
	.w6(32'h3962b127),
	.w7(32'hbaa552d5),
	.w8(32'hb91fc9d3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76048c),
	.w1(32'hbc8467f2),
	.w2(32'hbbf42cd5),
	.w3(32'hbb0e06b4),
	.w4(32'hbbb39071),
	.w5(32'hbc0b7175),
	.w6(32'hbc21648b),
	.w7(32'hbb92ce68),
	.w8(32'hbc2ce063),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44b062),
	.w1(32'h39950546),
	.w2(32'hba264e5b),
	.w3(32'h3a9a1e12),
	.w4(32'h39c27743),
	.w5(32'hbb2105b3),
	.w6(32'hba38a143),
	.w7(32'h3bb4725e),
	.w8(32'h3affdddb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6f302),
	.w1(32'h3ab4f0dd),
	.w2(32'h3a05f72c),
	.w3(32'h3b3e5daf),
	.w4(32'hb9a38973),
	.w5(32'h3be14b1d),
	.w6(32'h3c2526cc),
	.w7(32'h3a967862),
	.w8(32'h3b28e006),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule