module layer_8_featuremap_182(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7882b),
	.w1(32'hbaa97a33),
	.w2(32'hbc2a088b),
	.w3(32'h3b130e5f),
	.w4(32'hbb6d1fba),
	.w5(32'hbbea80ae),
	.w6(32'h3a8e1574),
	.w7(32'hbba9162c),
	.w8(32'hbc4e2ff5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9512e6),
	.w1(32'hbab42faf),
	.w2(32'hbb732894),
	.w3(32'h3bb5a75d),
	.w4(32'h3a20e0e3),
	.w5(32'hba765556),
	.w6(32'h3aa100f6),
	.w7(32'hbac6e583),
	.w8(32'hbb191a87),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8d23),
	.w1(32'h3c09bb92),
	.w2(32'h3c4f664e),
	.w3(32'hbbae0784),
	.w4(32'h3a42b866),
	.w5(32'hb9843120),
	.w6(32'h3b029f60),
	.w7(32'hbaf33270),
	.w8(32'h3b057ab9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b8af),
	.w1(32'h3a5806ba),
	.w2(32'h3ae1e505),
	.w3(32'hbc3dc6fe),
	.w4(32'hbb9c4732),
	.w5(32'hb9cea985),
	.w6(32'hbba40c50),
	.w7(32'hbb242682),
	.w8(32'hbc5daffb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84a8a6),
	.w1(32'hbb1edaa3),
	.w2(32'hbbb0a19f),
	.w3(32'hbc31358b),
	.w4(32'h35816385),
	.w5(32'hbb673ed4),
	.w6(32'hba4a83b3),
	.w7(32'hbb100518),
	.w8(32'hbae4ac7c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843ae9),
	.w1(32'hbba09451),
	.w2(32'hbbd3b157),
	.w3(32'hbb258918),
	.w4(32'hbb410836),
	.w5(32'hbb519afe),
	.w6(32'hbc3aa431),
	.w7(32'hbc48fd5a),
	.w8(32'hbc1e628b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99565c),
	.w1(32'h3aebd86e),
	.w2(32'h3b2fb3f7),
	.w3(32'h3ce4e118),
	.w4(32'hba8f9b73),
	.w5(32'hb90790e1),
	.w6(32'hbaee0da1),
	.w7(32'h3aa6ccac),
	.w8(32'h3a40402b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35252c),
	.w1(32'h3bc22407),
	.w2(32'h3b7226c1),
	.w3(32'h391e3213),
	.w4(32'hbb8afd79),
	.w5(32'hbcc79c51),
	.w6(32'h3b8786bd),
	.w7(32'h3c402be2),
	.w8(32'hbc96937c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb3cbb),
	.w1(32'hba78cbab),
	.w2(32'hbb7e13f3),
	.w3(32'h3c9259c2),
	.w4(32'hb94c61b8),
	.w5(32'h3a3d5025),
	.w6(32'h3aa28667),
	.w7(32'hbb1b9ec8),
	.w8(32'hbb52416e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d7fc9),
	.w1(32'hbba2bfe3),
	.w2(32'hbbb740fc),
	.w3(32'h3ab0272f),
	.w4(32'hbb8a7d98),
	.w5(32'hba0aac01),
	.w6(32'hbb9f335c),
	.w7(32'h3af0d907),
	.w8(32'h3b6ee690),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cbc57),
	.w1(32'hbad4397b),
	.w2(32'hbbc7b38e),
	.w3(32'hbc34a485),
	.w4(32'hbb3cc4f9),
	.w5(32'h3b25d4d6),
	.w6(32'h3a8c34e9),
	.w7(32'hbc14c2d4),
	.w8(32'hbc1f8a4a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb87843),
	.w1(32'hbb301cf5),
	.w2(32'h3b0447f4),
	.w3(32'h3b60bdb9),
	.w4(32'h3aba3a12),
	.w5(32'h3a342f15),
	.w6(32'hb82c6393),
	.w7(32'h3a00c689),
	.w8(32'hba3224f4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba023ee),
	.w1(32'h3b5ba8bb),
	.w2(32'h3bb0bb94),
	.w3(32'hb9fc9934),
	.w4(32'h3baad289),
	.w5(32'h3bc90244),
	.w6(32'hbba46b39),
	.w7(32'hbb156aca),
	.w8(32'h3abe5055),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d1c2),
	.w1(32'hbb406000),
	.w2(32'hbb5257d3),
	.w3(32'h3b127119),
	.w4(32'hbba2e4cb),
	.w5(32'hbc329f3e),
	.w6(32'hbb1e4b0d),
	.w7(32'h3aa62fc5),
	.w8(32'h3b8e88f9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c44d0),
	.w1(32'h39a57490),
	.w2(32'h3b938101),
	.w3(32'hbc83eaed),
	.w4(32'hb9fdacd3),
	.w5(32'h3b0e5692),
	.w6(32'h3a269b5a),
	.w7(32'h3afb0133),
	.w8(32'h3b2baad3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b7638),
	.w1(32'hbbbd6682),
	.w2(32'hbbf60299),
	.w3(32'hba520730),
	.w4(32'hbbdc9ab6),
	.w5(32'h3a7a8f91),
	.w6(32'h3bb18d7e),
	.w7(32'hbb8748c8),
	.w8(32'hbb73c1a3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43aa10),
	.w1(32'hba2a94d8),
	.w2(32'h3d11c32b),
	.w3(32'hbbad0c38),
	.w4(32'h3cd60f49),
	.w5(32'h3d17331f),
	.w6(32'hbc08b25a),
	.w7(32'h3a888298),
	.w8(32'h3cc59d30),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1dc2e5),
	.w1(32'h3be6da92),
	.w2(32'h3bd7a288),
	.w3(32'hbb07a63a),
	.w4(32'h3c4dbdd9),
	.w5(32'h3c4d0d69),
	.w6(32'h3b12670b),
	.w7(32'h3c087f25),
	.w8(32'h3b3f3b88),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc505387),
	.w1(32'hb7deba71),
	.w2(32'h3abf2116),
	.w3(32'hbc5a8a28),
	.w4(32'hbb73cfe1),
	.w5(32'h3b646349),
	.w6(32'h39a2c6fc),
	.w7(32'h3c08546f),
	.w8(32'h3b9f54d8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1446f),
	.w1(32'hb9f5f058),
	.w2(32'h3ae31f51),
	.w3(32'hbb5f9b5e),
	.w4(32'hbaefb188),
	.w5(32'hb9b8d9a3),
	.w6(32'hbb855882),
	.w7(32'hbb3b403c),
	.w8(32'hbaa7962a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d3562),
	.w1(32'h3b0c3179),
	.w2(32'hbbf2c344),
	.w3(32'hba4ce6e2),
	.w4(32'hbc20eade),
	.w5(32'hbbe3844d),
	.w6(32'h3c03037f),
	.w7(32'h3a376da0),
	.w8(32'h3bc36073),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be487),
	.w1(32'hbc3aa8cb),
	.w2(32'hba2ea876),
	.w3(32'hbc3a6877),
	.w4(32'hbc652a11),
	.w5(32'h3cb6f36e),
	.w6(32'hbc8cdef6),
	.w7(32'hbc7674dd),
	.w8(32'h3bb97125),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d377d4a),
	.w1(32'h3b48b940),
	.w2(32'h3ba687a9),
	.w3(32'h3d01837e),
	.w4(32'h3c2ec558),
	.w5(32'h3cda59ae),
	.w6(32'h3b1e5aa8),
	.w7(32'hbbcd1cfd),
	.w8(32'h3c3a9226),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea7ebb),
	.w1(32'hbc7f9214),
	.w2(32'hbbcb6ab2),
	.w3(32'hbbfc7808),
	.w4(32'hbc908df6),
	.w5(32'h3cc012b1),
	.w6(32'hbc252509),
	.w7(32'hbbdb2cf3),
	.w8(32'hbabc7f13),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d25b33b),
	.w1(32'hbb8cca65),
	.w2(32'hba3f2f50),
	.w3(32'h3d03aa69),
	.w4(32'h34711a97),
	.w5(32'h3bfbbd5a),
	.w6(32'hbb91adc7),
	.w7(32'hbb51440c),
	.w8(32'hbadefb8c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c912a),
	.w1(32'hbad05c7a),
	.w2(32'hbbf5c222),
	.w3(32'hbba3113c),
	.w4(32'h3a4d255b),
	.w5(32'h3b45d5ce),
	.w6(32'h3b184267),
	.w7(32'hbb9a064a),
	.w8(32'hb854adcf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16a718),
	.w1(32'h3c1692a2),
	.w2(32'h3b0c70d7),
	.w3(32'h3bc52c56),
	.w4(32'h3ba98f07),
	.w5(32'h3b1c085f),
	.w6(32'hbacdeb55),
	.w7(32'hbc27bc78),
	.w8(32'hbc916f51),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2575c0),
	.w1(32'hbaa52163),
	.w2(32'hbc2131d2),
	.w3(32'h3bc11e48),
	.w4(32'h3b21848c),
	.w5(32'hbbf8b2ad),
	.w6(32'hbb60d66c),
	.w7(32'hbc01b4b3),
	.w8(32'hbbc4ce9a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977a93),
	.w1(32'h3b8a28df),
	.w2(32'h3aebf7d8),
	.w3(32'hbad11c45),
	.w4(32'h39ea6c3b),
	.w5(32'h3b99b942),
	.w6(32'h3bce8ab4),
	.w7(32'h3b85338d),
	.w8(32'h3bbebaf2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be49477),
	.w1(32'hbbe2cc56),
	.w2(32'hbbebe905),
	.w3(32'h3bb574d8),
	.w4(32'h3bd2fc7f),
	.w5(32'h3c0516f9),
	.w6(32'h390538ff),
	.w7(32'hbb7dd717),
	.w8(32'hbb07f9a2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9969c5),
	.w1(32'h3a9e1f7c),
	.w2(32'h3afa5667),
	.w3(32'h3c5be0ca),
	.w4(32'hbb41d61f),
	.w5(32'h3a221a75),
	.w6(32'h384e3cf7),
	.w7(32'h3ba50438),
	.w8(32'hba3b98b7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2de829),
	.w1(32'h3b80abde),
	.w2(32'h3b392f38),
	.w3(32'hbba2e0e4),
	.w4(32'hbb5e1034),
	.w5(32'hbbd3594d),
	.w6(32'h3b177e0a),
	.w7(32'h3b059fa2),
	.w8(32'h3b6ecc64),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17e2e),
	.w1(32'h3b6c730b),
	.w2(32'hbb903ccb),
	.w3(32'hbc1e9816),
	.w4(32'hba86e519),
	.w5(32'h3b7e8b6a),
	.w6(32'hb8f91e92),
	.w7(32'hbafb8cb8),
	.w8(32'hbb9443fb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc975a0a),
	.w1(32'hbc83d24c),
	.w2(32'hbbff4b33),
	.w3(32'hbc24aeed),
	.w4(32'hbc14045c),
	.w5(32'h3a66661d),
	.w6(32'hbc89746a),
	.w7(32'hbc3971ed),
	.w8(32'hbb97bf3f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91fe0e),
	.w1(32'hbb211b53),
	.w2(32'h3a994bbf),
	.w3(32'h3c7370c2),
	.w4(32'h3b22805b),
	.w5(32'h3b5412a8),
	.w6(32'h3c08ddcb),
	.w7(32'h3bbfe8e9),
	.w8(32'h3b8f0a9c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab72cc3),
	.w1(32'h3c3c4ae0),
	.w2(32'h3c077f69),
	.w3(32'hbacf32c8),
	.w4(32'h3c3974a2),
	.w5(32'hbac3c5aa),
	.w6(32'hbadb6dda),
	.w7(32'h3be8fbb6),
	.w8(32'h3bfb26e3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb9ddc),
	.w1(32'hbb3e5103),
	.w2(32'h3912d2f8),
	.w3(32'hbc9d0b24),
	.w4(32'h3a859d98),
	.w5(32'h3ba05561),
	.w6(32'hbb041d94),
	.w7(32'hbb011ec9),
	.w8(32'hbb1a985f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b4ce),
	.w1(32'hbacfe466),
	.w2(32'h3b10f702),
	.w3(32'h3ba92224),
	.w4(32'hbaac7cf3),
	.w5(32'h3b0af2de),
	.w6(32'hba91666d),
	.w7(32'h398c7e2c),
	.w8(32'h3ad43fe8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b368e59),
	.w1(32'hbbd68c11),
	.w2(32'hbc354033),
	.w3(32'hbaa3a070),
	.w4(32'hbb9d4232),
	.w5(32'hbcbef25a),
	.w6(32'hbba2a3c5),
	.w7(32'hbc3724f8),
	.w8(32'h3ae1b336),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3828b),
	.w1(32'hbc737a13),
	.w2(32'hbc438d83),
	.w3(32'hbbb25e5f),
	.w4(32'hbc8a8360),
	.w5(32'h3c3eaa0e),
	.w6(32'hbc79689c),
	.w7(32'hbc5432f0),
	.w8(32'hbc2df0e4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77389f),
	.w1(32'h3a38d812),
	.w2(32'h39b651ec),
	.w3(32'h3cd57c54),
	.w4(32'h39c78336),
	.w5(32'hbaac1d0b),
	.w6(32'h3b870a6a),
	.w7(32'h3b92a4e4),
	.w8(32'h3b68ae68),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae721b2),
	.w1(32'hbb8b87b3),
	.w2(32'hbb60cdd6),
	.w3(32'hbb34bb51),
	.w4(32'hba3986e0),
	.w5(32'h3b65b3a4),
	.w6(32'hbad950dc),
	.w7(32'h3a3280fe),
	.w8(32'h39afe6f4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba974ae2),
	.w1(32'h3a187f93),
	.w2(32'hbc3fee7c),
	.w3(32'h3b2cd70f),
	.w4(32'hba8a0366),
	.w5(32'hbbd18bc8),
	.w6(32'hb9480cca),
	.w7(32'hbaa7f258),
	.w8(32'hb9b3102a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95a1c3),
	.w1(32'h3cac4b02),
	.w2(32'h3c8682f8),
	.w3(32'h3c0845f8),
	.w4(32'h3cbe29e5),
	.w5(32'h3b7f09a0),
	.w6(32'h3be8ec27),
	.w7(32'h3beeab39),
	.w8(32'hbb847c8f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79624e),
	.w1(32'hbcde091c),
	.w2(32'hbc4c5b0c),
	.w3(32'hbc609f56),
	.w4(32'hbc81f4d8),
	.w5(32'h3c02ec57),
	.w6(32'hbc9aaf48),
	.w7(32'hbbecdd6c),
	.w8(32'hbacd6d0f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873619),
	.w1(32'hbb804a2e),
	.w2(32'hbb24e6db),
	.w3(32'h3c176550),
	.w4(32'hbbc334e2),
	.w5(32'hbbdeba02),
	.w6(32'hbb494152),
	.w7(32'hbb95b89f),
	.w8(32'hbb3f133c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989a22),
	.w1(32'h38c2ba92),
	.w2(32'h375c8217),
	.w3(32'hbb697a94),
	.w4(32'h398d9c78),
	.w5(32'hbba62d98),
	.w6(32'h3b100a63),
	.w7(32'hbae71a66),
	.w8(32'h391586d9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0230d3),
	.w1(32'hbc9cc01f),
	.w2(32'hbc415d4c),
	.w3(32'hbc1f43e1),
	.w4(32'h3c272601),
	.w5(32'h3d098ce7),
	.w6(32'hbcb27db0),
	.w7(32'hbc13fa7a),
	.w8(32'hbcbdcae7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eacc3),
	.w1(32'hbc7e7919),
	.w2(32'hbc513898),
	.w3(32'h3c23b783),
	.w4(32'h3cabc2d2),
	.w5(32'h3cdf25cc),
	.w6(32'hbc6e59a2),
	.w7(32'hbc2556d5),
	.w8(32'hbc5f73e2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03704e),
	.w1(32'h3c2f9d30),
	.w2(32'hbb9fc110),
	.w3(32'h3c4508b5),
	.w4(32'h3b01b8df),
	.w5(32'hbc4cf6ea),
	.w6(32'hbbba93f6),
	.w7(32'hbbdef84e),
	.w8(32'hbc531e5f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b13d0),
	.w1(32'h3a944ba6),
	.w2(32'h3b9e50df),
	.w3(32'hbc7331b5),
	.w4(32'h3a1f5b60),
	.w5(32'hba9cf432),
	.w6(32'h3ab91d6c),
	.w7(32'h3b0bda44),
	.w8(32'h3a7f89e0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bcb1b),
	.w1(32'h3b4761b9),
	.w2(32'h3ad0b8af),
	.w3(32'hb9bd120d),
	.w4(32'h3a39fcb0),
	.w5(32'h3c0955d7),
	.w6(32'hbaff8d41),
	.w7(32'h3a5f60b3),
	.w8(32'h36e1f808),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aadfb),
	.w1(32'hbb367c53),
	.w2(32'hb92de202),
	.w3(32'h3c0b1a1e),
	.w4(32'h3a918e77),
	.w5(32'hb917b6ae),
	.w6(32'h3a77d186),
	.w7(32'hb9ad8861),
	.w8(32'h3adfd1bf),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251cec),
	.w1(32'h3b7893e2),
	.w2(32'hbba2423b),
	.w3(32'hbb14aa7b),
	.w4(32'hbb975559),
	.w5(32'hbbe1cd36),
	.w6(32'h3c972d98),
	.w7(32'h3c9e95d6),
	.w8(32'hbb81d793),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc659cd2),
	.w1(32'hbb853b00),
	.w2(32'hbbb88a0e),
	.w3(32'hbaba5de3),
	.w4(32'h3bd449a8),
	.w5(32'h3bd53566),
	.w6(32'hbc00d81b),
	.w7(32'h3ac4d925),
	.w8(32'hbba765ea),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66ab30),
	.w1(32'h3c0ea38a),
	.w2(32'h3c1cc988),
	.w3(32'hbc279c8c),
	.w4(32'h3bc4940d),
	.w5(32'h3c6b0b84),
	.w6(32'hb8e63470),
	.w7(32'hbb48e47f),
	.w8(32'h3bb563de),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc667e11),
	.w1(32'h3b2770fe),
	.w2(32'h3bcec7aa),
	.w3(32'h3abd8c05),
	.w4(32'h3b6eaabf),
	.w5(32'h3c33a15a),
	.w6(32'h3bcb3b5a),
	.w7(32'hbba824d7),
	.w8(32'h3bbde518),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bb716),
	.w1(32'hbad8de13),
	.w2(32'h3b8b8eaa),
	.w3(32'hbbf1126f),
	.w4(32'hbab7d4f3),
	.w5(32'h3bc0e0eb),
	.w6(32'h399b0267),
	.w7(32'h3bc88ecd),
	.w8(32'h3b1eb99b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dd737),
	.w1(32'h3afbd33f),
	.w2(32'h3b095dda),
	.w3(32'h3a418ad9),
	.w4(32'h3b3ec18e),
	.w5(32'h3b37dcf8),
	.w6(32'h3b31be15),
	.w7(32'h3aeba204),
	.w8(32'h3b1bf000),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1daee2),
	.w1(32'hbc5739fe),
	.w2(32'hbc234fa9),
	.w3(32'h3b477a79),
	.w4(32'hbc804c42),
	.w5(32'h3ced4a45),
	.w6(32'hbc3bfd31),
	.w7(32'hbc8fb341),
	.w8(32'h39f8569b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bdf38),
	.w1(32'h3ac0d1f5),
	.w2(32'h3b6f4bb3),
	.w3(32'h3d13d1ec),
	.w4(32'h3bac6bcb),
	.w5(32'h3a7f463f),
	.w6(32'h3b935546),
	.w7(32'hbb6847e7),
	.w8(32'hbc1b79ae),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4e3fa),
	.w1(32'hbb99767c),
	.w2(32'h3aed086a),
	.w3(32'hbb88b855),
	.w4(32'hbbf31557),
	.w5(32'hbb74b451),
	.w6(32'h3b9d2f89),
	.w7(32'h3ad38d32),
	.w8(32'h3ae918f9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987864),
	.w1(32'h3bb88996),
	.w2(32'h3bf43ab6),
	.w3(32'hbbde56bb),
	.w4(32'h3b9c7e48),
	.w5(32'h3b5b02f8),
	.w6(32'h3b8f4f76),
	.w7(32'h3bdb7bf1),
	.w8(32'h3b3e1793),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af56e2b),
	.w1(32'hbb6a2aff),
	.w2(32'hbba58922),
	.w3(32'h3ac0bf32),
	.w4(32'hbaf2b728),
	.w5(32'hbb9e170f),
	.w6(32'h3917f488),
	.w7(32'hbb2a1497),
	.w8(32'h38a062cb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf541e),
	.w1(32'hb992dc00),
	.w2(32'h3add488b),
	.w3(32'hbb5a48fa),
	.w4(32'h3a14c6bf),
	.w5(32'h3a8432cd),
	.w6(32'h3ad84a2d),
	.w7(32'h3b2480cd),
	.w8(32'h3b674266),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b35002),
	.w1(32'hbcd48102),
	.w2(32'hbc993679),
	.w3(32'h3b03ca0f),
	.w4(32'hbc1d622b),
	.w5(32'h3cde8d32),
	.w6(32'hbc85c3bc),
	.w7(32'hbc9be6fb),
	.w8(32'hbc20e84a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c401e),
	.w1(32'hbb9105eb),
	.w2(32'hbb536a8b),
	.w3(32'h3c998193),
	.w4(32'h3b941bfc),
	.w5(32'h3bffce76),
	.w6(32'h3c10b276),
	.w7(32'h3a511020),
	.w8(32'h3ba61393),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef3a03),
	.w1(32'h3a6e883a),
	.w2(32'h3b822bef),
	.w3(32'hbc5912c2),
	.w4(32'h3c46041b),
	.w5(32'hbbdb74a8),
	.w6(32'h3bd37b42),
	.w7(32'hbaa0708f),
	.w8(32'h3b63170a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a3083),
	.w1(32'hbcbf9f81),
	.w2(32'hbc70bf0b),
	.w3(32'hba9703eb),
	.w4(32'hbc86add2),
	.w5(32'h3a755777),
	.w6(32'hbc8db75b),
	.w7(32'hbc68693a),
	.w8(32'hb96195d4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe50bc2),
	.w1(32'hbb8dea78),
	.w2(32'hbc354e7c),
	.w3(32'hbbca8de6),
	.w4(32'hbb479504),
	.w5(32'h3cd2680b),
	.w6(32'hbbcf254c),
	.w7(32'hbc09ae95),
	.w8(32'hbc4e1995),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd167c3),
	.w1(32'hbae2148a),
	.w2(32'hbb15882a),
	.w3(32'h3c941c16),
	.w4(32'h3bad9ddf),
	.w5(32'h3b44263b),
	.w6(32'h3a368ea2),
	.w7(32'hba35fb62),
	.w8(32'hbc057b31),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3eee),
	.w1(32'h3c6aff04),
	.w2(32'h3c4ed720),
	.w3(32'hbba6314c),
	.w4(32'hbb2ccd78),
	.w5(32'hbc9bc7c6),
	.w6(32'h3c2fc051),
	.w7(32'h3c7edabc),
	.w8(32'h3c2d82b2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18c2a8),
	.w1(32'h3c6ee7f7),
	.w2(32'h3c930627),
	.w3(32'hbc80c0e5),
	.w4(32'h3b61a88e),
	.w5(32'hbc43d175),
	.w6(32'hbb632c4a),
	.w7(32'h3af8ba8f),
	.w8(32'h3c0839b6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2cf3),
	.w1(32'h3c6d5007),
	.w2(32'hbb2b6d31),
	.w3(32'hbcd05421),
	.w4(32'h3a3cf9be),
	.w5(32'hbbf3f703),
	.w6(32'h3baca386),
	.w7(32'h3adf6344),
	.w8(32'hbc435bcd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6380e3),
	.w1(32'h3b25ba7e),
	.w2(32'h3bca24a1),
	.w3(32'hbc149e1e),
	.w4(32'h3b6b5bb6),
	.w5(32'h3c081f61),
	.w6(32'hbaaa6368),
	.w7(32'h3b0a356b),
	.w8(32'hbb0bbd74),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8256c),
	.w1(32'h3b85a62a),
	.w2(32'h3a620d98),
	.w3(32'hbbd920ec),
	.w4(32'hbb5945e1),
	.w5(32'hb834a254),
	.w6(32'hb9177fda),
	.w7(32'hbbd34c19),
	.w8(32'hba80b889),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc405f3),
	.w1(32'hb83c17ed),
	.w2(32'hbbab085c),
	.w3(32'h3b9a75c8),
	.w4(32'h39b109a1),
	.w5(32'h3be58f91),
	.w6(32'h3c0f958d),
	.w7(32'hb94b5cd8),
	.w8(32'hbbb5ef74),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1025b3),
	.w1(32'hba056ca0),
	.w2(32'hbbc0cd12),
	.w3(32'h3c0021d1),
	.w4(32'hba9965cf),
	.w5(32'h3a06b463),
	.w6(32'h3ab58f1e),
	.w7(32'h37e3f3c0),
	.w8(32'hbb19fa3e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e1b3),
	.w1(32'hbbab36cc),
	.w2(32'h39d6bf72),
	.w3(32'h3bb9eaec),
	.w4(32'hbb3f24f2),
	.w5(32'hba89caf0),
	.w6(32'hbc1d2f0c),
	.w7(32'hba3422f7),
	.w8(32'h3984dfa6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68b1a4),
	.w1(32'h3c0a4d46),
	.w2(32'h3a2c1196),
	.w3(32'h37c62c4b),
	.w4(32'h3c9f474f),
	.w5(32'hbacb8405),
	.w6(32'hbb13ec49),
	.w7(32'hb9c2aeb2),
	.w8(32'hbc03552a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc414d89),
	.w1(32'h3c3f9d96),
	.w2(32'h3bf189cc),
	.w3(32'hba366810),
	.w4(32'hbbe7d774),
	.w5(32'hbc1faac2),
	.w6(32'hbba9b0da),
	.w7(32'h3bb65eed),
	.w8(32'h3b97ad53),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfac63),
	.w1(32'hbc903e24),
	.w2(32'hbc508dd1),
	.w3(32'hbc252670),
	.w4(32'hbc4180e6),
	.w5(32'hbbae6609),
	.w6(32'hbc28dd64),
	.w7(32'hbc00157a),
	.w8(32'hbc27be68),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80342),
	.w1(32'h3bdc378f),
	.w2(32'hbbd9438a),
	.w3(32'hbbaae095),
	.w4(32'h3b96c2a8),
	.w5(32'hbc37024a),
	.w6(32'h3c03ecb7),
	.w7(32'hbaef7387),
	.w8(32'hbadaac42),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f151e),
	.w1(32'h3b2f5d04),
	.w2(32'hbbd45582),
	.w3(32'h3aa9cf49),
	.w4(32'hbc0f48a3),
	.w5(32'hbbbcef69),
	.w6(32'h3b352c60),
	.w7(32'h3c461c5e),
	.w8(32'hbb41a12f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bd3bc),
	.w1(32'h3ab55fc0),
	.w2(32'h3c190bd2),
	.w3(32'h3c879afb),
	.w4(32'hbba5cb34),
	.w5(32'hbc8d47f8),
	.w6(32'hbc2dbc1c),
	.w7(32'h3bd19720),
	.w8(32'h3b9e247d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09ed6),
	.w1(32'hba8a7c46),
	.w2(32'hbb5a0bd0),
	.w3(32'hbcca37cf),
	.w4(32'hbbb7b9df),
	.w5(32'hbab1975f),
	.w6(32'hbb4d323f),
	.w7(32'hbbd46fac),
	.w8(32'hbc14dc41),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942523c),
	.w1(32'hbaac8606),
	.w2(32'hbaab2598),
	.w3(32'h3c48b885),
	.w4(32'h3b5048c6),
	.w5(32'h3bf3799b),
	.w6(32'hba4f78ae),
	.w7(32'h3ad30f66),
	.w8(32'hb841cb60),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a2064),
	.w1(32'h372f826d),
	.w2(32'h3995d1e0),
	.w3(32'h3bbc3f43),
	.w4(32'hbae42f5d),
	.w5(32'h39bcc9bc),
	.w6(32'hbac2e1bb),
	.w7(32'hbb453158),
	.w8(32'hbba7e42d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e0722),
	.w1(32'hbb78ccba),
	.w2(32'hbb6f0a14),
	.w3(32'h3bb31c95),
	.w4(32'h3b76148d),
	.w5(32'h3bc63847),
	.w6(32'hbb3df007),
	.w7(32'hba675b13),
	.w8(32'hbb4b3080),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcdb59),
	.w1(32'h3999a445),
	.w2(32'h3c1550ec),
	.w3(32'h3b32511c),
	.w4(32'h3bc5948f),
	.w5(32'h3be081ab),
	.w6(32'hbbeab8d7),
	.w7(32'h3b329785),
	.w8(32'h3ac2c529),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b032ac8),
	.w1(32'h3c9ae37b),
	.w2(32'h3c772710),
	.w3(32'hbb94a9e1),
	.w4(32'h3c11835a),
	.w5(32'hbc38a1c0),
	.w6(32'h3c45c889),
	.w7(32'h3be7c2df),
	.w8(32'h3c32c05b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0119),
	.w1(32'hbc318379),
	.w2(32'hbc8358b8),
	.w3(32'hbcdaf2d3),
	.w4(32'hbb63eb22),
	.w5(32'h39f85b84),
	.w6(32'hbbc9dd17),
	.w7(32'hbbd914d5),
	.w8(32'hbb874ba4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c175078),
	.w1(32'h3abac3df),
	.w2(32'hba4e7818),
	.w3(32'h3c3141a5),
	.w4(32'h3b1d4270),
	.w5(32'hb9a9f293),
	.w6(32'hbb49537f),
	.w7(32'hbb878974),
	.w8(32'hbb85d621),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2c27),
	.w1(32'hba9ae397),
	.w2(32'hbb136e44),
	.w3(32'hbb037060),
	.w4(32'h395cee21),
	.w5(32'hba8839d8),
	.w6(32'hb9991d0a),
	.w7(32'hbaace4ec),
	.w8(32'hbb60225f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49eb8b),
	.w1(32'h3b283960),
	.w2(32'hbc2bfee8),
	.w3(32'hba92ff13),
	.w4(32'hbab4a4c0),
	.w5(32'h3ae0cbf5),
	.w6(32'h39ad340a),
	.w7(32'hbb897519),
	.w8(32'hbb231fe2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd62bf),
	.w1(32'h3b5ce3eb),
	.w2(32'h3ad191b7),
	.w3(32'h3c33322f),
	.w4(32'h39d95753),
	.w5(32'h3a0dbfc2),
	.w6(32'h3aa69d4d),
	.w7(32'h3b66af3d),
	.w8(32'h3b83fc0a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b65f31),
	.w1(32'hbbe6db2c),
	.w2(32'hba5a7ba8),
	.w3(32'hbb83f30b),
	.w4(32'hb9ccbf89),
	.w5(32'h3c744d3a),
	.w6(32'hb9aa6014),
	.w7(32'hbc32b317),
	.w8(32'hb9923f3d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c844672),
	.w1(32'h3c7dafe4),
	.w2(32'h3b470cd2),
	.w3(32'h3c07efc7),
	.w4(32'h39eae311),
	.w5(32'hbcd9e642),
	.w6(32'h3c286b91),
	.w7(32'h3ba91482),
	.w8(32'hbb960ddb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10c2a8),
	.w1(32'h3c74b9b7),
	.w2(32'h3ba173d5),
	.w3(32'hbb5989dd),
	.w4(32'h3bcdfcdb),
	.w5(32'hbcd5a7f7),
	.w6(32'h3c918cd3),
	.w7(32'h3b27a648),
	.w8(32'h3888d435),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60305b),
	.w1(32'h3b809eef),
	.w2(32'hbb2d2f1f),
	.w3(32'hbc9a10e4),
	.w4(32'h3bf7e1db),
	.w5(32'hbbfc7a96),
	.w6(32'hbbcd217f),
	.w7(32'hbbf2ebe2),
	.w8(32'hbc85c602),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196351),
	.w1(32'hbb443dca),
	.w2(32'hbb99f7b7),
	.w3(32'hbbc5d583),
	.w4(32'hbb72f232),
	.w5(32'hbaa6173d),
	.w6(32'hbab438dc),
	.w7(32'hbbdbae05),
	.w8(32'hbb2c6a83),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb830c52),
	.w1(32'h3c13ea78),
	.w2(32'h3cd1c525),
	.w3(32'hba735a9c),
	.w4(32'hb8c95197),
	.w5(32'hbc5c4f58),
	.w6(32'h3c112900),
	.w7(32'h3c80cc51),
	.w8(32'h3c266b76),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c6149),
	.w1(32'hbc1367b3),
	.w2(32'hbb1dc162),
	.w3(32'hbc99dae0),
	.w4(32'hbbb83b68),
	.w5(32'hbc4860c2),
	.w6(32'h3a4c28d0),
	.w7(32'h3a5f0efe),
	.w8(32'hba4b6cb3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9253e8),
	.w1(32'hbc1ba323),
	.w2(32'h3c16f149),
	.w3(32'hba05292f),
	.w4(32'h3c8dc123),
	.w5(32'h3cef23f6),
	.w6(32'hbc3022ba),
	.w7(32'hbc1ef1aa),
	.w8(32'hbb2e217a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ea0f6),
	.w1(32'h3b354dbf),
	.w2(32'hbc098093),
	.w3(32'hbc615d9e),
	.w4(32'hbc045e46),
	.w5(32'hbc8bf8d4),
	.w6(32'h3c1553c9),
	.w7(32'h3b2603fe),
	.w8(32'h3c877762),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9478bb),
	.w1(32'hba9e9a99),
	.w2(32'hb984bc61),
	.w3(32'hbc6b7fe1),
	.w4(32'hba6cdffa),
	.w5(32'hbaf9e63c),
	.w6(32'hbbdbd278),
	.w7(32'hbb8dc189),
	.w8(32'h3a0addc0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9372e17),
	.w1(32'hbb7cc148),
	.w2(32'hbb92a003),
	.w3(32'hbb312ac5),
	.w4(32'hba83a8a9),
	.w5(32'h3b8b93ff),
	.w6(32'hbb0414bc),
	.w7(32'hbb558b0d),
	.w8(32'hbc10f5d5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba054625),
	.w1(32'hbb18aaa6),
	.w2(32'hbb53caf7),
	.w3(32'h3b77da6e),
	.w4(32'h3b031a48),
	.w5(32'h3b9fe14d),
	.w6(32'hbb5944e9),
	.w7(32'hb9c7f889),
	.w8(32'hbc198909),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02b372),
	.w1(32'h3b8a85fd),
	.w2(32'h3bf74cbf),
	.w3(32'h3affdea5),
	.w4(32'h3baeb367),
	.w5(32'hbb97b020),
	.w6(32'h3c79a949),
	.w7(32'h3c5d71bf),
	.w8(32'h3c0fb4e8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae89f1b),
	.w1(32'hba92a0f5),
	.w2(32'hba34c26d),
	.w3(32'hbafe4555),
	.w4(32'h3a73e547),
	.w5(32'h38ad6709),
	.w6(32'hba8ca994),
	.w7(32'hb915cfab),
	.w8(32'h39b8873d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17f4ce),
	.w1(32'hba2e7f67),
	.w2(32'h3bab9383),
	.w3(32'h3abf9c60),
	.w4(32'hbba60d35),
	.w5(32'hbc0150cc),
	.w6(32'h3ad2e729),
	.w7(32'h3b5700c4),
	.w8(32'h3aba7459),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36d4a4),
	.w1(32'hbbbe760b),
	.w2(32'hbb913176),
	.w3(32'hbc28fdd8),
	.w4(32'hbbd1905a),
	.w5(32'hbbb442df),
	.w6(32'hbb7eb534),
	.w7(32'hbb978fe1),
	.w8(32'hbbc1e63c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb979b00),
	.w1(32'hbba8ce82),
	.w2(32'h3aec6e29),
	.w3(32'hbb001f6b),
	.w4(32'hbbade520),
	.w5(32'h3c187569),
	.w6(32'hbb661836),
	.w7(32'hbb8bac1c),
	.w8(32'h3bd028e6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c180601),
	.w1(32'h3b990d7a),
	.w2(32'hbadbb5e0),
	.w3(32'h3b82f255),
	.w4(32'h3c55af2d),
	.w5(32'h3b1faceb),
	.w6(32'h3b7e4c98),
	.w7(32'h3bbba4c3),
	.w8(32'hbafe165a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90b151),
	.w1(32'hbb427134),
	.w2(32'hbb600288),
	.w3(32'hbbbe0ac1),
	.w4(32'h3b59eb08),
	.w5(32'h3b9c425d),
	.w6(32'hbab1cc3b),
	.w7(32'hbb2bd0f1),
	.w8(32'hbbfc2e25),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb324393),
	.w1(32'hbaed8ff8),
	.w2(32'hbadc0ca2),
	.w3(32'h3b4e8f5f),
	.w4(32'hba6b986f),
	.w5(32'hbaa923a1),
	.w6(32'hbb091747),
	.w7(32'hbb0ee4b3),
	.w8(32'hbadf50c4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb662c12),
	.w1(32'h3b834935),
	.w2(32'hbb926918),
	.w3(32'hb9c0c6ad),
	.w4(32'h3aee3183),
	.w5(32'h3aabb13e),
	.w6(32'h3c39c300),
	.w7(32'h3be53eb8),
	.w8(32'h3b76402a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa7a5),
	.w1(32'h3a8c0f3a),
	.w2(32'h3ba16524),
	.w3(32'h3c20024d),
	.w4(32'h3a850acb),
	.w5(32'h3b85cd08),
	.w6(32'h3bee5b72),
	.w7(32'hbaecb093),
	.w8(32'hbb67a4f1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b198391),
	.w1(32'hbbe02b07),
	.w2(32'hbc0fdd69),
	.w3(32'hba0e6dec),
	.w4(32'hbc185551),
	.w5(32'hbc4d65ad),
	.w6(32'hba88f30f),
	.w7(32'hbc39bc14),
	.w8(32'hba5b550b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27229c),
	.w1(32'hbb154275),
	.w2(32'h3ba2a2bf),
	.w3(32'hbba5acef),
	.w4(32'hbb77f36e),
	.w5(32'h3bc1ff0a),
	.w6(32'hbb6b9576),
	.w7(32'hbac9397b),
	.w8(32'h3a04f6b6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc701ad),
	.w1(32'hbc0f01aa),
	.w2(32'hbc4fd5f0),
	.w3(32'hbad558cc),
	.w4(32'hbafe055c),
	.w5(32'h3b5a9e7b),
	.w6(32'hbc1aff95),
	.w7(32'hbc059a79),
	.w8(32'hbba8bbc7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf447bc),
	.w1(32'hbac7aa28),
	.w2(32'h3ae40c95),
	.w3(32'h3b815fd1),
	.w4(32'hb9a8019b),
	.w5(32'hbbcccf20),
	.w6(32'hba989d8f),
	.w7(32'h3b7a2a72),
	.w8(32'hba05b0cc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe34779),
	.w1(32'hbb3dfa85),
	.w2(32'hbb91977d),
	.w3(32'hbb95662d),
	.w4(32'hbad8c804),
	.w5(32'hbb8f8758),
	.w6(32'h3ab61332),
	.w7(32'h359f3711),
	.w8(32'hbb2afa11),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfdf7c),
	.w1(32'hbc29565b),
	.w2(32'hba58055f),
	.w3(32'hbb976007),
	.w4(32'hbbe0eed3),
	.w5(32'h3bdf41d8),
	.w6(32'hb90a6515),
	.w7(32'hbb7a069a),
	.w8(32'h3912a4f6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c504293),
	.w1(32'hbc46b78c),
	.w2(32'hbc875d96),
	.w3(32'h3b9fee87),
	.w4(32'hbc94994f),
	.w5(32'hbc7a3a39),
	.w6(32'h3b1367c1),
	.w7(32'h3b39234a),
	.w8(32'h3c562b2b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16b89d),
	.w1(32'hbc937e00),
	.w2(32'hbc712525),
	.w3(32'h38f49497),
	.w4(32'h3c4082c9),
	.w5(32'h3d1a226c),
	.w6(32'hbca9a006),
	.w7(32'hbc5e290c),
	.w8(32'hbc52cf45),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024fb0),
	.w1(32'hbbb6822e),
	.w2(32'hbd0cddb1),
	.w3(32'h3cb7cfae),
	.w4(32'hbc1393c8),
	.w5(32'hbcde5133),
	.w6(32'h3c45c727),
	.w7(32'h3bc30706),
	.w8(32'h3bfa795a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc778e22),
	.w1(32'h3b3e583e),
	.w2(32'h3c8b585d),
	.w3(32'hbc80f784),
	.w4(32'h39c85c9a),
	.w5(32'h3c4d3878),
	.w6(32'h3b7f8749),
	.w7(32'h3b392f7e),
	.w8(32'h3b940e46),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule