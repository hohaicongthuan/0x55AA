module layer_10_featuremap_31(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa617d),
	.w1(32'h3b6ddab1),
	.w2(32'hbb5f9c03),
	.w3(32'hbb7bb5ec),
	.w4(32'hbbd02ced),
	.w5(32'hbc367238),
	.w6(32'hbb87b4f6),
	.w7(32'h3b08f6fb),
	.w8(32'hbaab62f6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38de9d),
	.w1(32'hba45a5e8),
	.w2(32'hbbc71d42),
	.w3(32'hbc497b70),
	.w4(32'hbad264c8),
	.w5(32'hbc420b93),
	.w6(32'hbc2a69f8),
	.w7(32'h3a99361b),
	.w8(32'hbbe158a3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ded64),
	.w1(32'h3bebdd4d),
	.w2(32'h3bff5200),
	.w3(32'hbb8b0e07),
	.w4(32'h3c983953),
	.w5(32'h3c307abd),
	.w6(32'h3b805bd0),
	.w7(32'h3c6ec367),
	.w8(32'h3bce9964),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba385829),
	.w1(32'h3ac062e8),
	.w2(32'hbb87426b),
	.w3(32'h3c3c036c),
	.w4(32'hba919703),
	.w5(32'hbc679159),
	.w6(32'h3c1c12be),
	.w7(32'h3b21200a),
	.w8(32'hbc387d36),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdecf83),
	.w1(32'hbbec94fd),
	.w2(32'hbb007bff),
	.w3(32'hbc6a5c35),
	.w4(32'hbb93d808),
	.w5(32'hba879d55),
	.w6(32'hb97d223c),
	.w7(32'h3c064308),
	.w8(32'hbc14cb36),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c321a),
	.w1(32'h3c305018),
	.w2(32'hbb7fd48c),
	.w3(32'hbb418d7c),
	.w4(32'h3c49ce84),
	.w5(32'hbb05a29f),
	.w6(32'h388077df),
	.w7(32'h3c63528e),
	.w8(32'h3aa642d7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc5b46),
	.w1(32'h3a0fe383),
	.w2(32'hbc1f845f),
	.w3(32'hbb9b1c2b),
	.w4(32'h3aa1050d),
	.w5(32'hbaa9aa1e),
	.w6(32'hba8f8112),
	.w7(32'h3b87d696),
	.w8(32'hb9a177f3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62cace),
	.w1(32'hba38fdd9),
	.w2(32'hbb59270f),
	.w3(32'hb9d1954f),
	.w4(32'h3ba0649d),
	.w5(32'hbb961b26),
	.w6(32'h3bef6580),
	.w7(32'h3b81f740),
	.w8(32'hbb02753f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85924b),
	.w1(32'hbb9819ba),
	.w2(32'h3a314520),
	.w3(32'hb904fd19),
	.w4(32'hba6757bf),
	.w5(32'hbb676fc0),
	.w6(32'hbb43035e),
	.w7(32'h3b0f134f),
	.w8(32'hba332391),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934e14),
	.w1(32'hbc0bd278),
	.w2(32'h3a077849),
	.w3(32'hbbd38dbc),
	.w4(32'hbc42c900),
	.w5(32'h38f41a74),
	.w6(32'hbb985ac6),
	.w7(32'hbc156278),
	.w8(32'h39ab44a8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c67165),
	.w1(32'hbae05b4f),
	.w2(32'h3b171577),
	.w3(32'hba4bb193),
	.w4(32'hba98df6a),
	.w5(32'h3b7fc13e),
	.w6(32'hba548215),
	.w7(32'hbb28c6d4),
	.w8(32'h3b1c0506),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac26795),
	.w1(32'hbb3ce374),
	.w2(32'hba69cd93),
	.w3(32'h3c1969d9),
	.w4(32'h3bb6fb05),
	.w5(32'hbb727ab2),
	.w6(32'h38089fec),
	.w7(32'h3b966a41),
	.w8(32'hbb778911),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac21d7),
	.w1(32'hbb8762b0),
	.w2(32'hbbbec5df),
	.w3(32'hbbdd009f),
	.w4(32'hbb9fb6bd),
	.w5(32'hbc246eed),
	.w6(32'hbbdd4aea),
	.w7(32'hbba2b4fc),
	.w8(32'hbbfd6115),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8099f1),
	.w1(32'hbb741e17),
	.w2(32'hbbb5900c),
	.w3(32'hbc28d764),
	.w4(32'h3b2ea5b6),
	.w5(32'hbc657dd6),
	.w6(32'h3b64ad01),
	.w7(32'h3b82ed5e),
	.w8(32'hbb996779),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c7dc6),
	.w1(32'hbc1cdf24),
	.w2(32'h3b9a770b),
	.w3(32'hbc4d34e9),
	.w4(32'h3b200192),
	.w5(32'h3bd378ca),
	.w6(32'hb92f473f),
	.w7(32'h3c39aa58),
	.w8(32'h3bc31bfe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44be06),
	.w1(32'h3b004141),
	.w2(32'h3ae11287),
	.w3(32'h3bc6f018),
	.w4(32'h3b6f0ac4),
	.w5(32'h3a902146),
	.w6(32'h3bd36fd7),
	.w7(32'h3b0452cb),
	.w8(32'h3acd7b45),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a523e38),
	.w1(32'hb986bd6c),
	.w2(32'hbb63c416),
	.w3(32'hb9c1f2fb),
	.w4(32'h39a6716b),
	.w5(32'hba859cc7),
	.w6(32'hb99e3dd0),
	.w7(32'hba011ad0),
	.w8(32'hbb8e4711),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03ea1f),
	.w1(32'hb8e3c6f3),
	.w2(32'hbbb390b3),
	.w3(32'hbaab1254),
	.w4(32'h3a178f74),
	.w5(32'hbb6ac930),
	.w6(32'hbbabb729),
	.w7(32'hbbaa044a),
	.w8(32'h3b00e5b9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47c24),
	.w1(32'hbaa2ce8a),
	.w2(32'hbc689438),
	.w3(32'hbaccd627),
	.w4(32'h3b9b5567),
	.w5(32'hbc75faaa),
	.w6(32'h3aadadeb),
	.w7(32'h3bcd4a8e),
	.w8(32'hbc111dfb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd445f4),
	.w1(32'hbbfe3cb3),
	.w2(32'hbafcadf8),
	.w3(32'hbc234bf0),
	.w4(32'h39a28b6c),
	.w5(32'h3a399292),
	.w6(32'hbc192891),
	.w7(32'hb9d06228),
	.w8(32'h3b06973b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88e739),
	.w1(32'hba5a8b71),
	.w2(32'hbbaef329),
	.w3(32'h3affa920),
	.w4(32'h39a3e5dc),
	.w5(32'h3b5cb40a),
	.w6(32'h3b2807b7),
	.w7(32'h3b802578),
	.w8(32'h3b0a6797),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54ea78),
	.w1(32'h3a826dbf),
	.w2(32'h3bae6ee4),
	.w3(32'h3c040ac8),
	.w4(32'h3b2804c5),
	.w5(32'h3b9ac5da),
	.w6(32'hba9947ca),
	.w7(32'hbbf8ab0b),
	.w8(32'h3c13ac51),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becb796),
	.w1(32'h3a877953),
	.w2(32'h3af7ca09),
	.w3(32'h3b9f1a4b),
	.w4(32'hbaf4270e),
	.w5(32'h3a879a43),
	.w6(32'h3badc5ab),
	.w7(32'hba2e8deb),
	.w8(32'h3a46ef68),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da875),
	.w1(32'hb9691976),
	.w2(32'hbb568c86),
	.w3(32'h3b23a37d),
	.w4(32'hba4ffdba),
	.w5(32'hbb87bc1c),
	.w6(32'h3a4dd7f4),
	.w7(32'hbb00a042),
	.w8(32'hba46abae),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81abb7),
	.w1(32'h3b0013f7),
	.w2(32'hbba0e017),
	.w3(32'hbaf78b35),
	.w4(32'h3c08fa3a),
	.w5(32'hbbacbbee),
	.w6(32'h3b25794c),
	.w7(32'h3ba7c493),
	.w8(32'hbbeb0915),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028194),
	.w1(32'h3b4a492b),
	.w2(32'hbb4aa976),
	.w3(32'hbbdce21d),
	.w4(32'hbb99097e),
	.w5(32'h3bef9aca),
	.w6(32'hbc5c510c),
	.w7(32'h3a8ad3a1),
	.w8(32'h3ba527d2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8adaf),
	.w1(32'h3be997b4),
	.w2(32'h3a6ce1b3),
	.w3(32'h3bd389c1),
	.w4(32'h3c046da8),
	.w5(32'hbab0bbb9),
	.w6(32'hba9c8cd8),
	.w7(32'h3b212200),
	.w8(32'h39c6fd8c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb90f9),
	.w1(32'h3a080465),
	.w2(32'hbbbfc796),
	.w3(32'h3a9eabc2),
	.w4(32'hba8357bd),
	.w5(32'h3c0c5a1f),
	.w6(32'h3b140aa5),
	.w7(32'hb8a84f4a),
	.w8(32'h3c6b3371),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa82a92),
	.w1(32'h3bc10127),
	.w2(32'h3c0333da),
	.w3(32'hb98b227d),
	.w4(32'h3bd04772),
	.w5(32'h3cba9cf5),
	.w6(32'h3b570364),
	.w7(32'h3bc1917e),
	.w8(32'hbb8cc4f5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a5e16),
	.w1(32'hbbb264fd),
	.w2(32'hbb148a80),
	.w3(32'hbb3f0ae8),
	.w4(32'hbbe64e64),
	.w5(32'hba8b34d8),
	.w6(32'h3c90902c),
	.w7(32'hbb9075f4),
	.w8(32'h3a80148c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41f01e),
	.w1(32'h3abfa393),
	.w2(32'hbc51d65d),
	.w3(32'h3b17f5ff),
	.w4(32'h3afa47a0),
	.w5(32'hbbe11215),
	.w6(32'hbb0a0b57),
	.w7(32'h3a8c9fc8),
	.w8(32'h3a9c2e80),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8937eec),
	.w1(32'h3a903cf3),
	.w2(32'hbc4e8125),
	.w3(32'hbb6df649),
	.w4(32'h3b0792af),
	.w5(32'h3c0b4611),
	.w6(32'hbc00bfec),
	.w7(32'hbbb3086a),
	.w8(32'hbb95c508),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47532e),
	.w1(32'hbc081166),
	.w2(32'hb6cef31d),
	.w3(32'hbc5d56b9),
	.w4(32'hbb058fd8),
	.w5(32'hbb3b35df),
	.w6(32'hbba859bc),
	.w7(32'hbc04ad0d),
	.w8(32'hbb0cb099),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc09f),
	.w1(32'hba849e95),
	.w2(32'hbacbdd36),
	.w3(32'hb93ddae6),
	.w4(32'hbac33251),
	.w5(32'h3b112124),
	.w6(32'hbae81436),
	.w7(32'hba04e2f1),
	.w8(32'h3b7a38dc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6940f3),
	.w1(32'h3b073afe),
	.w2(32'hbae10c8d),
	.w3(32'hbc175cab),
	.w4(32'h3b03aed5),
	.w5(32'hbb6a3491),
	.w6(32'hbb858516),
	.w7(32'h3c162fa9),
	.w8(32'hbb0a8664),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b0493),
	.w1(32'hbb7d972f),
	.w2(32'hbc118b75),
	.w3(32'hbb420add),
	.w4(32'hbb595565),
	.w5(32'hbb9ce78c),
	.w6(32'hba9c852c),
	.w7(32'hbaa57b8c),
	.w8(32'hbc4f832a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2565e8),
	.w1(32'hbb2be402),
	.w2(32'hbb90a54b),
	.w3(32'h3bc6be4a),
	.w4(32'hbc370f48),
	.w5(32'hbb96d24a),
	.w6(32'h3c24a47c),
	.w7(32'h3bcadc6d),
	.w8(32'hbb62d8d2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215aca),
	.w1(32'h3a1f9b5a),
	.w2(32'h3bb1e20b),
	.w3(32'h3b56b372),
	.w4(32'h3b973416),
	.w5(32'hbc4b9eac),
	.w6(32'hbad3bd3d),
	.w7(32'h3ba0e9a8),
	.w8(32'hbbf55a61),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed33b0),
	.w1(32'hbb8f7d0a),
	.w2(32'hbc635505),
	.w3(32'h3bc988be),
	.w4(32'hbbe657e0),
	.w5(32'h3cbacf50),
	.w6(32'hbb808a86),
	.w7(32'h3cbcb521),
	.w8(32'h3cdb482b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45fcf),
	.w1(32'h3bbaaead),
	.w2(32'hb9d82dd7),
	.w3(32'hbcd2c47d),
	.w4(32'h3c549e8f),
	.w5(32'hbbcc985a),
	.w6(32'hbbf23e12),
	.w7(32'hbc0b25e1),
	.w8(32'hbb9823fc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4b814),
	.w1(32'h36a339f7),
	.w2(32'hbb11f108),
	.w3(32'h3ad7074e),
	.w4(32'hb9e2befc),
	.w5(32'hbb8fc5ba),
	.w6(32'h3b8015cd),
	.w7(32'hbb40a451),
	.w8(32'hbaab89cc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e4aa),
	.w1(32'hbbc8c375),
	.w2(32'hbc031c3a),
	.w3(32'h39ce8148),
	.w4(32'h3b9b604c),
	.w5(32'hbc66280f),
	.w6(32'hbbb38c4b),
	.w7(32'h3c93f64f),
	.w8(32'hbc95749c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90555d),
	.w1(32'h3b181330),
	.w2(32'hba308d7d),
	.w3(32'hbcb3a8fc),
	.w4(32'hbc0dd296),
	.w5(32'h3a0eebfa),
	.w6(32'h3920c7b9),
	.w7(32'hbbac919b),
	.w8(32'h3b902140),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae036be),
	.w1(32'hbb71fdc7),
	.w2(32'h3c8004f1),
	.w3(32'h394d7f24),
	.w4(32'hbb36865c),
	.w5(32'h3c17c3ef),
	.w6(32'h3b487560),
	.w7(32'h3b57ed13),
	.w8(32'hbaa8b41b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bdfbc),
	.w1(32'h3c175616),
	.w2(32'hbcbbc733),
	.w3(32'hbc704fa7),
	.w4(32'hbb71605f),
	.w5(32'hbbc63e75),
	.w6(32'h3b643bd9),
	.w7(32'hbcb39e37),
	.w8(32'h3c39407f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf01ce4),
	.w1(32'hbc404e2f),
	.w2(32'h3c941443),
	.w3(32'h3b368661),
	.w4(32'h3bda2d0e),
	.w5(32'h3c5caec8),
	.w6(32'hbc4581e5),
	.w7(32'h3c6f28d8),
	.w8(32'hbbe95931),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc455830),
	.w1(32'hbb6895df),
	.w2(32'h3b9707fe),
	.w3(32'h3c1a5f86),
	.w4(32'hbcb59178),
	.w5(32'hbccdf747),
	.w6(32'h3cb5bbb0),
	.w7(32'hbce5ad5d),
	.w8(32'hbc94ab90),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c9793),
	.w1(32'hbc5dd068),
	.w2(32'hbac35f53),
	.w3(32'h3d0c6fb4),
	.w4(32'hbbcf92e1),
	.w5(32'h39a0284a),
	.w6(32'hbb651218),
	.w7(32'h3cea25a0),
	.w8(32'h3b2c0385),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f0954),
	.w1(32'hbb08a737),
	.w2(32'hbb0166ae),
	.w3(32'h37c6d222),
	.w4(32'h3ac5393b),
	.w5(32'h3afa6414),
	.w6(32'h3a224963),
	.w7(32'h3b6c8056),
	.w8(32'h39646727),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0c7b1),
	.w1(32'h3c2875be),
	.w2(32'h3b81bad0),
	.w3(32'h3b8d57fd),
	.w4(32'hbb67e5d0),
	.w5(32'h3bcac892),
	.w6(32'hbc06f84d),
	.w7(32'hbb98a892),
	.w8(32'h3bbb4e86),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44592d),
	.w1(32'h3bfa4286),
	.w2(32'hbc3b965d),
	.w3(32'hbb00fb3d),
	.w4(32'h3c1f0016),
	.w5(32'hbc631eee),
	.w6(32'hbbced114),
	.w7(32'h3c499956),
	.w8(32'hbb6c8518),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb731),
	.w1(32'hbc0af94d),
	.w2(32'h3c1d374c),
	.w3(32'hbc1ed0f1),
	.w4(32'hbbd48026),
	.w5(32'h3b4a84d9),
	.w6(32'h3b05fe85),
	.w7(32'hbbe1b548),
	.w8(32'h3bfc581e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0efbd0),
	.w1(32'hbb93a336),
	.w2(32'hba48503e),
	.w3(32'hbba8e102),
	.w4(32'h3c328d6d),
	.w5(32'hbb2e9421),
	.w6(32'hbb911e30),
	.w7(32'h3c8e9df9),
	.w8(32'hbac18e4b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c279475),
	.w1(32'hbba91a15),
	.w2(32'h3c064ef8),
	.w3(32'h3bd9111e),
	.w4(32'h3bce12ee),
	.w5(32'h3b90d647),
	.w6(32'hbb883118),
	.w7(32'hbb57dfeb),
	.w8(32'hbc46be8f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d68fc),
	.w1(32'h3a80c06b),
	.w2(32'h3afdf112),
	.w3(32'h3bd67880),
	.w4(32'hbc852c92),
	.w5(32'h3a985894),
	.w6(32'h3c652a37),
	.w7(32'hbb2dbef5),
	.w8(32'hbc0ec15c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a7d6e),
	.w1(32'h3b9032bc),
	.w2(32'h3a4347e0),
	.w3(32'hbb6c35f7),
	.w4(32'h3c055ca2),
	.w5(32'h3cf142a6),
	.w6(32'hbbfd6062),
	.w7(32'h3c11bbd1),
	.w8(32'h3c5ff479),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab159b),
	.w1(32'h3bd7e812),
	.w2(32'h3b18838a),
	.w3(32'hbcb038d4),
	.w4(32'h3c60fc2c),
	.w5(32'h3ac1665b),
	.w6(32'hbb10fe29),
	.w7(32'hbc3fe9fa),
	.w8(32'hb9984880),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b3f86),
	.w1(32'hbaa80c6f),
	.w2(32'h3ad5242e),
	.w3(32'hba044b5e),
	.w4(32'hbb996853),
	.w5(32'hba9b2024),
	.w6(32'hbb0f5a84),
	.w7(32'hbbe108a1),
	.w8(32'h3b26d069),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920ab3c),
	.w1(32'h3b968709),
	.w2(32'hbabce2cc),
	.w3(32'h3b193015),
	.w4(32'h3bcde454),
	.w5(32'hbb5507db),
	.w6(32'h3b2d9682),
	.w7(32'h3c233613),
	.w8(32'hba33f79d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d2c9c),
	.w1(32'hbb6c715b),
	.w2(32'hbc09e1e8),
	.w3(32'h3a528477),
	.w4(32'hbbab4ae9),
	.w5(32'hbc5f237a),
	.w6(32'h3a10fecb),
	.w7(32'hbb9cf10e),
	.w8(32'hbc0fe2ca),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c82f1),
	.w1(32'hbbd417e2),
	.w2(32'h3c975ab2),
	.w3(32'h3b821d4b),
	.w4(32'hbb48f8b7),
	.w5(32'h3c95704f),
	.w6(32'hbc0ca908),
	.w7(32'h3b6425e6),
	.w8(32'h3b6abe19),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd81049),
	.w1(32'h3c54d1b4),
	.w2(32'h3b9d8891),
	.w3(32'h3c3d9e1a),
	.w4(32'hba4a7000),
	.w5(32'hbb78d0c3),
	.w6(32'h3c0925e8),
	.w7(32'hbacf416d),
	.w8(32'hbc97b932),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca456d9),
	.w1(32'hbbf9975d),
	.w2(32'hbc3f8007),
	.w3(32'h3c536ddc),
	.w4(32'hbc660e27),
	.w5(32'hbc18a3b5),
	.w6(32'h3c12be7d),
	.w7(32'h38a7f706),
	.w8(32'hbb1c675b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c70b08),
	.w1(32'hbb943946),
	.w2(32'hbb71db0b),
	.w3(32'hbba9ebb7),
	.w4(32'hbb92eff0),
	.w5(32'h3b351b72),
	.w6(32'hbc2de6bf),
	.w7(32'h3a23370e),
	.w8(32'h3ba24201),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d657),
	.w1(32'hbba6a1ba),
	.w2(32'hb95604d8),
	.w3(32'h3c4a123d),
	.w4(32'h3c02c6b1),
	.w5(32'hbae17463),
	.w6(32'h3baab350),
	.w7(32'h3be9297a),
	.w8(32'h3a3004dd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801df4),
	.w1(32'h3c0846f1),
	.w2(32'hbb561657),
	.w3(32'hb9e6c1b2),
	.w4(32'h3c10ba8b),
	.w5(32'hbaf2c97c),
	.w6(32'h3a8e2cf8),
	.w7(32'h3b5bd63e),
	.w8(32'h3abf9ddc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0565d9),
	.w1(32'hbb80e8ac),
	.w2(32'hbc145005),
	.w3(32'hbb0380fb),
	.w4(32'hbbb7466d),
	.w5(32'hbc469d7b),
	.w6(32'hbb243938),
	.w7(32'hbb2a76a6),
	.w8(32'hbb9e2d47),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf930e),
	.w1(32'h3bc5d627),
	.w2(32'hbb58bc70),
	.w3(32'hbd003cc5),
	.w4(32'h3bf886f8),
	.w5(32'hba55928e),
	.w6(32'hbc85ea53),
	.w7(32'h3b9e9b60),
	.w8(32'hbc0826d0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a1ad3),
	.w1(32'hbc2182b2),
	.w2(32'hbb8f950f),
	.w3(32'hbbb6e9c4),
	.w4(32'hbb85aec0),
	.w5(32'hbb9fcfba),
	.w6(32'hbbbddbdd),
	.w7(32'h38e2ac17),
	.w8(32'hbb1e654e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad781e1),
	.w1(32'hbaefe592),
	.w2(32'h3bd177a4),
	.w3(32'hbbd89b9e),
	.w4(32'hbb824171),
	.w5(32'h3c69b701),
	.w6(32'hbbcf242b),
	.w7(32'hbb7e2b0d),
	.w8(32'h3b4a486a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00ae5),
	.w1(32'h3bcd5d31),
	.w2(32'h3b85e3bf),
	.w3(32'hbb4dbcc9),
	.w4(32'hbaf482c6),
	.w5(32'h3bf158f3),
	.w6(32'h3be11ca4),
	.w7(32'hbb766c27),
	.w8(32'hba513dd2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5652aa),
	.w1(32'h3c55d4e6),
	.w2(32'h3c614b1d),
	.w3(32'hbc77228d),
	.w4(32'h3bafee4e),
	.w5(32'hbc29218d),
	.w6(32'h3bb99226),
	.w7(32'hbc0222d0),
	.w8(32'hbcb50852),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79eaa9),
	.w1(32'h3a05b2eb),
	.w2(32'hbcac4515),
	.w3(32'hb83bb4a5),
	.w4(32'hbc860df7),
	.w5(32'hbc5f7800),
	.w6(32'h3c7a1db4),
	.w7(32'hbcdc5b01),
	.w8(32'h3c5e2c4d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81d169),
	.w1(32'h3b13bc1e),
	.w2(32'hbbe9eaaa),
	.w3(32'hbc982a26),
	.w4(32'h3ca86b7f),
	.w5(32'hbc07ed55),
	.w6(32'hbc9be6b7),
	.w7(32'h3bc5bb01),
	.w8(32'hbba85d0d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107ab3),
	.w1(32'hbb1c2853),
	.w2(32'h38fce19e),
	.w3(32'hbb7d0785),
	.w4(32'hb972a744),
	.w5(32'hbb4736f1),
	.w6(32'hbbceab55),
	.w7(32'hba0ab6e6),
	.w8(32'hbb62bca4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f79bf),
	.w1(32'hbbc822f2),
	.w2(32'hbb595d2b),
	.w3(32'hbc20805d),
	.w4(32'hbc033797),
	.w5(32'hbb7eb160),
	.w6(32'hbb8348b7),
	.w7(32'hbb1b5c43),
	.w8(32'h3b5b7750),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdf17b),
	.w1(32'hbabeee5b),
	.w2(32'hbc29350b),
	.w3(32'hbb9c1fe8),
	.w4(32'hbc72d75a),
	.w5(32'hbb44ddc5),
	.w6(32'h3b537dd9),
	.w7(32'hbbd0b97a),
	.w8(32'h3b8df15c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5268e),
	.w1(32'hbc743138),
	.w2(32'h3c210c03),
	.w3(32'hbb3511bc),
	.w4(32'hbc0988d3),
	.w5(32'h3b94d278),
	.w6(32'h3b0a4ec8),
	.w7(32'hbb87be71),
	.w8(32'hbc0337e7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc456bcf),
	.w1(32'h3b088dcc),
	.w2(32'h3ab8f8c8),
	.w3(32'h3c2793a3),
	.w4(32'hbc112ab0),
	.w5(32'hba8f759a),
	.w6(32'h3c3aa6c4),
	.w7(32'hbb29046b),
	.w8(32'h3a5342ca),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fad37),
	.w1(32'h3a08a769),
	.w2(32'hbab1f5fc),
	.w3(32'hbacaa346),
	.w4(32'hba6922b6),
	.w5(32'h36c3100d),
	.w6(32'h3b044176),
	.w7(32'hb8d0fd04),
	.w8(32'hbbf7d529),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcca86),
	.w1(32'h3ba45ccc),
	.w2(32'hbb175b72),
	.w3(32'hbaa97847),
	.w4(32'h3a422ea2),
	.w5(32'hbb483d2b),
	.w6(32'hbb4e77ea),
	.w7(32'h3a23a14c),
	.w8(32'hba6f4c5c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d0c45),
	.w1(32'hbacff99c),
	.w2(32'h3ba5bf56),
	.w3(32'h3a8a0210),
	.w4(32'hba98f435),
	.w5(32'hbc4e2c82),
	.w6(32'h38a4a6bb),
	.w7(32'hbac39d0d),
	.w8(32'hbc89e648),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a1c67),
	.w1(32'hbba989cc),
	.w2(32'h3c09e0ed),
	.w3(32'h3b2bb298),
	.w4(32'hbbd72867),
	.w5(32'hbbb3b371),
	.w6(32'h3b4fb465),
	.w7(32'hbc102d6d),
	.w8(32'hbc739f7a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dae41),
	.w1(32'hbc3f00f7),
	.w2(32'h3cf76afc),
	.w3(32'h3cecbd9c),
	.w4(32'hbc97d518),
	.w5(32'h3c3ad976),
	.w6(32'h3bfc8f1d),
	.w7(32'h3ba6052a),
	.w8(32'hbc0367cb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b610a),
	.w1(32'hbb34d67d),
	.w2(32'hbbdfea82),
	.w3(32'h3caefd60),
	.w4(32'hbc402fbb),
	.w5(32'hbaa3ae8f),
	.w6(32'h3cddc637),
	.w7(32'hbca53156),
	.w8(32'h3bc47503),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccb585),
	.w1(32'h3c0857ba),
	.w2(32'hbb15827f),
	.w3(32'hbc44772b),
	.w4(32'h38b7856c),
	.w5(32'hbb075c78),
	.w6(32'h3c07ca04),
	.w7(32'hbbf2551b),
	.w8(32'hbbc6f2b3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994cce),
	.w1(32'h3be356b0),
	.w2(32'h3a0bd907),
	.w3(32'hbb85b588),
	.w4(32'h3bb268bd),
	.w5(32'h397948ea),
	.w6(32'hbac408db),
	.w7(32'hbae5bc96),
	.w8(32'hbac6051e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8fa5a),
	.w1(32'h392c5408),
	.w2(32'h3ba195a8),
	.w3(32'hbad719cc),
	.w4(32'hba5eee2d),
	.w5(32'h3a0120e8),
	.w6(32'hbab768d6),
	.w7(32'h3ac31e1a),
	.w8(32'h3a31786a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1845de),
	.w1(32'h3b27a013),
	.w2(32'hbc124563),
	.w3(32'hbac30c9b),
	.w4(32'h3c2dbd7c),
	.w5(32'hbc02dc4d),
	.w6(32'h3b0458e6),
	.w7(32'h3c125a43),
	.w8(32'h3b42036f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54cdd9),
	.w1(32'hbc0a07b1),
	.w2(32'hbb05c305),
	.w3(32'hbbf98a2c),
	.w4(32'hbb3fb434),
	.w5(32'h3b487141),
	.w6(32'hbc10699a),
	.w7(32'hb7c50239),
	.w8(32'h3bcbfe5f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6b7b5),
	.w1(32'hba80f8e8),
	.w2(32'h3b42c743),
	.w3(32'h3ab8bfe5),
	.w4(32'hbb4b7dec),
	.w5(32'h3be55fc4),
	.w6(32'hbb72b70c),
	.w7(32'hbac50883),
	.w8(32'h3b501b5e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb71e1),
	.w1(32'hbb4d3f48),
	.w2(32'hba5744fb),
	.w3(32'h3c4e4393),
	.w4(32'h3b4ef0b9),
	.w5(32'h3a6d9ead),
	.w6(32'h3b462851),
	.w7(32'h3b466d84),
	.w8(32'h3a9b7b87),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bb589),
	.w1(32'hbb477276),
	.w2(32'hb7392c09),
	.w3(32'hba9c099a),
	.w4(32'hba3697fd),
	.w5(32'h3b907ac8),
	.w6(32'h3ae0b909),
	.w7(32'h3b1d7e7f),
	.w8(32'h3bab3c60),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8d5a3),
	.w1(32'h3ad27bc9),
	.w2(32'hbbbcc529),
	.w3(32'h3b5a5fe2),
	.w4(32'h3b04a558),
	.w5(32'hbb3e18da),
	.w6(32'h3afc4def),
	.w7(32'h3b196646),
	.w8(32'hbbbd8a7a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc259528),
	.w1(32'hbc2a7f32),
	.w2(32'h3a9fb540),
	.w3(32'hbc33dfd4),
	.w4(32'hbc75b72b),
	.w5(32'hbb83aff5),
	.w6(32'hbc012530),
	.w7(32'hbc425fcd),
	.w8(32'hbb12ea45),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb765e29),
	.w1(32'h3b90bc11),
	.w2(32'hbc0001ae),
	.w3(32'hbb858bf7),
	.w4(32'hbc3cda09),
	.w5(32'hbbe05769),
	.w6(32'hbc227b07),
	.w7(32'hbc96ea4e),
	.w8(32'hbb390e23),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bda79),
	.w1(32'hbaa6f075),
	.w2(32'h3ceb7e5f),
	.w3(32'hbc362872),
	.w4(32'hbc6d3952),
	.w5(32'h3c608736),
	.w6(32'hb98d28c1),
	.w7(32'hbc12b25e),
	.w8(32'hbcbcee15),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98edd7),
	.w1(32'hbbe7e9eb),
	.w2(32'hbb481329),
	.w3(32'h3cc646b7),
	.w4(32'hbc94f628),
	.w5(32'hbb74982f),
	.w6(32'h3cee6290),
	.w7(32'hbb45dad9),
	.w8(32'h3bcbf6cf),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd95a2),
	.w1(32'hbbcc23c5),
	.w2(32'hbb47ec10),
	.w3(32'hba7d833f),
	.w4(32'hbb8050d7),
	.w5(32'hbaee50fa),
	.w6(32'hbc01236f),
	.w7(32'hbaaa2d69),
	.w8(32'hba55c86b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1283f9),
	.w1(32'hbbb5ed0d),
	.w2(32'hbb323a66),
	.w3(32'h3addf994),
	.w4(32'h3b2fa38b),
	.w5(32'hbc8aeee5),
	.w6(32'hba66a615),
	.w7(32'h3b6b49a8),
	.w8(32'h3bde371f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf96f6e),
	.w1(32'hba8fb318),
	.w2(32'h3b846491),
	.w3(32'hbb9b5b17),
	.w4(32'h3bd5dcc6),
	.w5(32'h3af0c27a),
	.w6(32'hbc651b04),
	.w7(32'h3b1449e4),
	.w8(32'h3c84662c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59f539),
	.w1(32'h3b09e597),
	.w2(32'hbc2307d3),
	.w3(32'h3c48fb2c),
	.w4(32'h3bd3084f),
	.w5(32'hbc497304),
	.w6(32'hbaa19894),
	.w7(32'h3b5dafc0),
	.w8(32'hbb6a3a56),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fe9b6),
	.w1(32'hb9842cf9),
	.w2(32'hba9f915d),
	.w3(32'hbbd62e94),
	.w4(32'h3b698ea8),
	.w5(32'hbadaa401),
	.w6(32'hbc502a21),
	.w7(32'hbb0ab698),
	.w8(32'hbbcb3718),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5df3c9),
	.w1(32'hbab8fda3),
	.w2(32'hbbc5717f),
	.w3(32'h3a76afb4),
	.w4(32'h38196b33),
	.w5(32'hbbfd5604),
	.w6(32'hbb8c5e0c),
	.w7(32'hba7d1b85),
	.w8(32'hbbb3e965),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43d3e7),
	.w1(32'hbc042550),
	.w2(32'hbae6efb0),
	.w3(32'hbc868a6a),
	.w4(32'hbc4b195c),
	.w5(32'h3af2cf41),
	.w6(32'hbc14fe0b),
	.w7(32'hbc523726),
	.w8(32'hbb206ab7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc160fbb),
	.w1(32'h3ba2d8d3),
	.w2(32'h3b3b2488),
	.w3(32'hba640f91),
	.w4(32'h3baac9ce),
	.w5(32'h3c07ddab),
	.w6(32'h3b937225),
	.w7(32'hba43c5e2),
	.w8(32'h3a6dc4cb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9ac83),
	.w1(32'h3bbf4d7e),
	.w2(32'h3b0cd2e8),
	.w3(32'h39f6db8b),
	.w4(32'hbab03fcd),
	.w5(32'hbabf0002),
	.w6(32'h3c28f2ab),
	.w7(32'hbbbef339),
	.w8(32'hbc243a66),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1868e9),
	.w1(32'h3be26780),
	.w2(32'h3c9cdbe6),
	.w3(32'hbb6c9034),
	.w4(32'hbc01ebec),
	.w5(32'h3d0c3884),
	.w6(32'h3be5cc4c),
	.w7(32'hbbbd5d2b),
	.w8(32'hba91ec8e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf35a9b),
	.w1(32'h3bad66fe),
	.w2(32'hbc1b1cff),
	.w3(32'hbc9a930f),
	.w4(32'hbbc26d62),
	.w5(32'hbc2362ac),
	.w6(32'h3c837311),
	.w7(32'hbce488e1),
	.w8(32'hbb843b1f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157901),
	.w1(32'hba53db89),
	.w2(32'h3b974e23),
	.w3(32'hbbba6d0b),
	.w4(32'h3a8d2eb2),
	.w5(32'h3c1c3f89),
	.w6(32'hbc005286),
	.w7(32'h3b399c2e),
	.w8(32'hbc35ca32),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a892a),
	.w1(32'h3b3702a5),
	.w2(32'hbb6f5041),
	.w3(32'hbc2c7bfe),
	.w4(32'hbc4ab38d),
	.w5(32'h3bf8fd73),
	.w6(32'h3c0315f6),
	.w7(32'hbb710f6f),
	.w8(32'hb84ba585),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d69f1),
	.w1(32'h3bafdde1),
	.w2(32'h3aa88673),
	.w3(32'hbc5f1216),
	.w4(32'h3ab1105a),
	.w5(32'hbc11143e),
	.w6(32'h3b92a6db),
	.w7(32'hbbea62cd),
	.w8(32'hbb1fb078),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad937f1),
	.w1(32'h38e286cb),
	.w2(32'hb9aa6582),
	.w3(32'hbac3afdc),
	.w4(32'hbbfaffad),
	.w5(32'h3b0fb052),
	.w6(32'hbbc5778d),
	.w7(32'hbc074fde),
	.w8(32'hbbdf4269),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d02b0),
	.w1(32'h3b8cc7e3),
	.w2(32'h3bd88772),
	.w3(32'hbc1cf487),
	.w4(32'hbc639c1e),
	.w5(32'h3c11f489),
	.w6(32'hbbe616bc),
	.w7(32'hbc0beedd),
	.w8(32'h3bad0612),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6883),
	.w1(32'hbb5465a6),
	.w2(32'h3bc75836),
	.w3(32'hbb7a8264),
	.w4(32'hba95bc6a),
	.w5(32'h3b81c9b6),
	.w6(32'hbbff9ab5),
	.w7(32'hbbaff4c8),
	.w8(32'h3bcc4d6a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0606e2),
	.w1(32'h3a802eb7),
	.w2(32'hbb769e73),
	.w3(32'h3bc33d65),
	.w4(32'h3b5515aa),
	.w5(32'h3b027860),
	.w6(32'h3bb58f66),
	.w7(32'h3b53f094),
	.w8(32'h3a3d9230),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca234e),
	.w1(32'hba2780f8),
	.w2(32'h3b825e59),
	.w3(32'hba17c06d),
	.w4(32'h3b8e70ef),
	.w5(32'h39c0096d),
	.w6(32'h3ab7f85f),
	.w7(32'h39da922d),
	.w8(32'h3b672fb9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf664f7),
	.w1(32'hb9a48efb),
	.w2(32'hbc8b4b0b),
	.w3(32'h3b8d5e2a),
	.w4(32'h3addbb6e),
	.w5(32'hbc1f2e8d),
	.w6(32'h3b91d564),
	.w7(32'h3b95f898),
	.w8(32'h3be3eb96),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c100dd2),
	.w1(32'hbb2162b6),
	.w2(32'h3bfe7d20),
	.w3(32'hbb9c3a46),
	.w4(32'h3b098791),
	.w5(32'hbb62d8b0),
	.w6(32'hbc3c0581),
	.w7(32'h3b27b2b9),
	.w8(32'h3c803a9f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c931d8b),
	.w1(32'hb9f3ed9b),
	.w2(32'hbbcbc293),
	.w3(32'h3be8f4af),
	.w4(32'h3ae336cb),
	.w5(32'hbbf9879a),
	.w6(32'h3985dd96),
	.w7(32'h3c311d17),
	.w8(32'hbc8e4acf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdb510),
	.w1(32'hbc4c118a),
	.w2(32'hbba9401d),
	.w3(32'hbc59fb5f),
	.w4(32'hbc9d9b3f),
	.w5(32'hbba60859),
	.w6(32'hbb7dceb1),
	.w7(32'hbc0418de),
	.w8(32'hbb52db76),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba046229),
	.w1(32'hbb32c0ef),
	.w2(32'hbaff6eba),
	.w3(32'hba24ba8d),
	.w4(32'h38ac7544),
	.w5(32'hba9aa75a),
	.w6(32'hbbba8098),
	.w7(32'hbb0d5677),
	.w8(32'hbb71b652),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea1e27),
	.w1(32'hb973a911),
	.w2(32'h3c123337),
	.w3(32'hbaaa05c9),
	.w4(32'hbade49dc),
	.w5(32'hbcaaae80),
	.w6(32'hbb93f3a9),
	.w7(32'hbb2787e1),
	.w8(32'hbcad1606),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c433270),
	.w1(32'hbc833c5a),
	.w2(32'hbbe1ec80),
	.w3(32'h3cebf33e),
	.w4(32'hbc36c34e),
	.w5(32'hbb3058c1),
	.w6(32'hba3458ea),
	.w7(32'h3c33ac10),
	.w8(32'hbb1a2e35),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c45c),
	.w1(32'h3b615176),
	.w2(32'hbb9a15a1),
	.w3(32'h38f361aa),
	.w4(32'h3ab4eac7),
	.w5(32'hbc2ebcee),
	.w6(32'hbb18076a),
	.w7(32'hbb1cbe49),
	.w8(32'hbc41c247),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63d88e),
	.w1(32'hbafc16a8),
	.w2(32'h39d0e67d),
	.w3(32'hbcc3187f),
	.w4(32'hbc23e295),
	.w5(32'hbc76d55c),
	.w6(32'hbc9d4baa),
	.w7(32'hbb8c199d),
	.w8(32'hbc1c04bc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89c958),
	.w1(32'h3ba8f2b1),
	.w2(32'hbb6a1415),
	.w3(32'hbcdc210f),
	.w4(32'hbb1e25c6),
	.w5(32'hbc90796e),
	.w6(32'hbc445352),
	.w7(32'hbc32cbfc),
	.w8(32'hbc678691),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68dd95),
	.w1(32'h3b6fc938),
	.w2(32'hbc22289b),
	.w3(32'hbc4faa26),
	.w4(32'h3bd33bcb),
	.w5(32'h3cd658ff),
	.w6(32'hbbce3175),
	.w7(32'hba89bbc1),
	.w8(32'h3c9ae101),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc897dc5),
	.w1(32'h3c8a1eef),
	.w2(32'h3cb1dfd2),
	.w3(32'hbc745237),
	.w4(32'h3c6519cf),
	.w5(32'h3ca54ca5),
	.w6(32'hbb6c00f1),
	.w7(32'hba8f0c4b),
	.w8(32'hbc2f0564),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8be023),
	.w1(32'hb9fd6a7c),
	.w2(32'hbcdec77d),
	.w3(32'h3a718c81),
	.w4(32'hbc34345c),
	.w5(32'hbc4bcaee),
	.w6(32'h3cb7cec9),
	.w7(32'hbc34a711),
	.w8(32'h3ca2871d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09a7a6),
	.w1(32'hbc07bd93),
	.w2(32'hbbeb0a16),
	.w3(32'h3c67dcaf),
	.w4(32'h3c3cf6a3),
	.w5(32'hbb7f14aa),
	.w6(32'hbcc2cb89),
	.w7(32'h3c650c75),
	.w8(32'hbc41d182),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc574190),
	.w1(32'hb8a66ebc),
	.w2(32'hbc7689bf),
	.w3(32'hbc9448ec),
	.w4(32'hbc99a1d9),
	.w5(32'hbc204c26),
	.w6(32'hbc61f3c2),
	.w7(32'hbbb3727f),
	.w8(32'hbb587235),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04ffe5),
	.w1(32'hbc85cc58),
	.w2(32'h3c4da6ee),
	.w3(32'hbaa30382),
	.w4(32'hbc1da8f3),
	.w5(32'h3cb78bdc),
	.w6(32'hbc21552f),
	.w7(32'hbc22be0e),
	.w8(32'h3cc4bbcd),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c444202),
	.w1(32'h3b606b2e),
	.w2(32'hba8c109f),
	.w3(32'hbc3ff2d1),
	.w4(32'h3c2446bf),
	.w5(32'hb84882ff),
	.w6(32'hbb9c1abf),
	.w7(32'hbc070fd8),
	.w8(32'hb8be14b9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e0d01),
	.w1(32'h394d8a19),
	.w2(32'h3aafd56c),
	.w3(32'h3b4203ed),
	.w4(32'h3b2c0495),
	.w5(32'hbb5477fb),
	.w6(32'h3b3cbb3e),
	.w7(32'h3b4cd33f),
	.w8(32'h3b8001fb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe6359),
	.w1(32'h3ae5d605),
	.w2(32'h3b322d56),
	.w3(32'h3c1cbe99),
	.w4(32'h3b35ad70),
	.w5(32'hbaf4ed09),
	.w6(32'h3b874de0),
	.w7(32'h3b275a08),
	.w8(32'hbc14d113),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e5a42),
	.w1(32'h3c1cd690),
	.w2(32'h3b4aff12),
	.w3(32'h3b6ec2b2),
	.w4(32'hb9b1dfdc),
	.w5(32'h3b06a8b0),
	.w6(32'h3c12dc2a),
	.w7(32'hbbef3f7c),
	.w8(32'hba4ef584),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07e1f5),
	.w1(32'h3a835921),
	.w2(32'hbafb07a6),
	.w3(32'h3bbd67ba),
	.w4(32'h3927aa69),
	.w5(32'h383e3cfc),
	.w6(32'h3c0d1e76),
	.w7(32'h3b9973fb),
	.w8(32'hb99f1fa3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac269f1),
	.w1(32'hbb45fc65),
	.w2(32'hbc8cdd50),
	.w3(32'hba26d3d7),
	.w4(32'hbb21ba84),
	.w5(32'hbbbcb278),
	.w6(32'hba5c2849),
	.w7(32'hbb6a657e),
	.w8(32'hbc57cd6b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba842c68),
	.w1(32'h3a04ac3d),
	.w2(32'hbb2a8d38),
	.w3(32'hbc2ecc5e),
	.w4(32'h378b2bca),
	.w5(32'hbb12db7e),
	.w6(32'hbc610f95),
	.w7(32'hbbed8e64),
	.w8(32'hbb6db877),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac44132),
	.w1(32'h39fb76f7),
	.w2(32'h3bd9ad02),
	.w3(32'h3a9421d2),
	.w4(32'h3b35fdfd),
	.w5(32'h3bbd5b3c),
	.w6(32'hbad457cc),
	.w7(32'h398ec3ce),
	.w8(32'h3c380cda),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5303ad),
	.w1(32'h3b54cbff),
	.w2(32'hbb1fd0b9),
	.w3(32'hbad2af91),
	.w4(32'hbb4541f9),
	.w5(32'hbae4758d),
	.w6(32'h3bbe6250),
	.w7(32'hbaf1eebc),
	.w8(32'hbad01708),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25dce3),
	.w1(32'h3aa3a047),
	.w2(32'h3b9ccff8),
	.w3(32'hbb00ef67),
	.w4(32'h3be9276d),
	.w5(32'hbb0872ca),
	.w6(32'hbb25d022),
	.w7(32'h3b442cd1),
	.w8(32'hbaf2bc5e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b310c6c),
	.w1(32'h3a8c231f),
	.w2(32'hbb2cd634),
	.w3(32'hba8f4d7d),
	.w4(32'hbb1e69eb),
	.w5(32'h389a7d64),
	.w6(32'h3b601227),
	.w7(32'hbb04c709),
	.w8(32'hba5b411f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa1fb),
	.w1(32'hbb3a2163),
	.w2(32'hbbf4f14b),
	.w3(32'hba834096),
	.w4(32'hbb264e6d),
	.w5(32'hbbf072cf),
	.w6(32'hbb18e4ec),
	.w7(32'hbb6cc9d3),
	.w8(32'h3b447398),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48d08b),
	.w1(32'hb901a6a4),
	.w2(32'h3bc25154),
	.w3(32'hbc20df0b),
	.w4(32'h3b6aa4e3),
	.w5(32'h3b1512d1),
	.w6(32'hbbfc7efc),
	.w7(32'hbb052043),
	.w8(32'hbb3e305f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca4418),
	.w1(32'h3a6b5b3d),
	.w2(32'h3cf2e17a),
	.w3(32'h3bb8791e),
	.w4(32'hb90acc64),
	.w5(32'h3ab7469c),
	.w6(32'h3c07a3f2),
	.w7(32'hbb23b48a),
	.w8(32'hbcdd5eda),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc277ee),
	.w1(32'hbbadb958),
	.w2(32'h3b681f6c),
	.w3(32'h3c87b0b5),
	.w4(32'hbbfd47bd),
	.w5(32'h3a85b4d5),
	.w6(32'h3cbb4dea),
	.w7(32'h3c580f16),
	.w8(32'hbb27e69d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d7e2d),
	.w1(32'h3ae532c9),
	.w2(32'h3d0d06e4),
	.w3(32'h3b7153f2),
	.w4(32'h3bb189a7),
	.w5(32'h3cb7ee23),
	.w6(32'hba268d40),
	.w7(32'h3b94dec1),
	.w8(32'hbc67df9d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82b580),
	.w1(32'h3b5d4ed6),
	.w2(32'h3b6f6442),
	.w3(32'h3ce16863),
	.w4(32'hbc316823),
	.w5(32'h3beeec18),
	.w6(32'h3cf03383),
	.w7(32'h3a9a08f5),
	.w8(32'hbbb0aec8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f6bef),
	.w1(32'hbba73541),
	.w2(32'hba289b80),
	.w3(32'hbb16b0be),
	.w4(32'hbb82d3ab),
	.w5(32'hba5b36ea),
	.w6(32'h3be1db58),
	.w7(32'hbb54b5f9),
	.w8(32'hba880514),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420ea7),
	.w1(32'h3b23534e),
	.w2(32'h3c0db4ab),
	.w3(32'h3b6d290a),
	.w4(32'h3b84ba44),
	.w5(32'h3b710dfe),
	.w6(32'h3a2df65e),
	.w7(32'h3ba7c5a1),
	.w8(32'h3bd0597e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be58b4e),
	.w1(32'h3b0b886e),
	.w2(32'h3bd17a4b),
	.w3(32'h3c0ededa),
	.w4(32'h3b777ee0),
	.w5(32'hbcda92f4),
	.w6(32'h3b10ae22),
	.w7(32'h3aacd6cb),
	.w8(32'hbc680b27),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a211b),
	.w1(32'hbc57347d),
	.w2(32'hbb8e0335),
	.w3(32'h3bde00fe),
	.w4(32'hbc856b51),
	.w5(32'hbab61c67),
	.w6(32'hbc560f1b),
	.w7(32'h3c2a2383),
	.w8(32'h3ba88e15),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20538),
	.w1(32'hbc16c65e),
	.w2(32'h3a62688b),
	.w3(32'hbb3d6e67),
	.w4(32'hbc284cd3),
	.w5(32'h3c3acdcc),
	.w6(32'hbb04fcb5),
	.w7(32'hbc1d1519),
	.w8(32'h3b5a73d9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c772a85),
	.w1(32'h3b525862),
	.w2(32'hbbc41296),
	.w3(32'h3d329137),
	.w4(32'h3c8afa57),
	.w5(32'hbb9fa18b),
	.w6(32'h3cbb267d),
	.w7(32'h3bb5c07a),
	.w8(32'hbbe1c5cf),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d42b),
	.w1(32'hba6ce802),
	.w2(32'h3b8e8815),
	.w3(32'hbbc946fb),
	.w4(32'h3ba63da8),
	.w5(32'h3a91f27f),
	.w6(32'hbb5abe8f),
	.w7(32'h3bfb60d5),
	.w8(32'h3bbe97ee),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd28b4),
	.w1(32'h3b6fee1a),
	.w2(32'hbb8aebc7),
	.w3(32'h3c09443e),
	.w4(32'h3bbb1e01),
	.w5(32'hbb52731c),
	.w6(32'h3b48ebdc),
	.w7(32'h3c245299),
	.w8(32'hbb978bd6),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93e05d),
	.w1(32'hb9cbafb0),
	.w2(32'h3a396824),
	.w3(32'h3befb348),
	.w4(32'h3b9c79e8),
	.w5(32'h3ab00bba),
	.w6(32'h3b8bd41f),
	.w7(32'h3aa9086e),
	.w8(32'h3be02e5b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d9887),
	.w1(32'hbb82d065),
	.w2(32'h3b348991),
	.w3(32'h3bc92fb1),
	.w4(32'h3aa74399),
	.w5(32'h3ab353f4),
	.w6(32'h3af86159),
	.w7(32'hb994b284),
	.w8(32'hba82a1a4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd20b3),
	.w1(32'h3b32805e),
	.w2(32'h3cc2fbaf),
	.w3(32'h3c06e0be),
	.w4(32'h3bca5a80),
	.w5(32'h3c5e0ab9),
	.w6(32'hbbc7e285),
	.w7(32'hbb503f95),
	.w8(32'h3c17ff9c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca10f53),
	.w1(32'h3cb6c2f4),
	.w2(32'h3b1c4eb7),
	.w3(32'h3b93a3c9),
	.w4(32'h3c17e48e),
	.w5(32'hbb164c95),
	.w6(32'h3a9d72ae),
	.w7(32'h3be752a8),
	.w8(32'h3a1ec3ae),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31566c),
	.w1(32'hbbbf7cbe),
	.w2(32'h3bbdd0f5),
	.w3(32'hbc0a4aba),
	.w4(32'hbb2c015e),
	.w5(32'h3b342893),
	.w6(32'hba6f8f48),
	.w7(32'h3bbc5ec8),
	.w8(32'h3b31042a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c00d7),
	.w1(32'h3a6c5e13),
	.w2(32'hbb8e25da),
	.w3(32'hbbbc4e53),
	.w4(32'hbb035e20),
	.w5(32'hbb891d62),
	.w6(32'hbb8fde60),
	.w7(32'hba77976d),
	.w8(32'hbbc946fd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb591240),
	.w1(32'hbbb3e7ff),
	.w2(32'h3bfa4543),
	.w3(32'h3abc1e27),
	.w4(32'h3b49deae),
	.w5(32'hb998be32),
	.w6(32'hbaa59b86),
	.w7(32'hba3f671d),
	.w8(32'hba87c355),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc18c),
	.w1(32'h3b3b82d0),
	.w2(32'h3b790ce5),
	.w3(32'hbb81745e),
	.w4(32'hbafce9d3),
	.w5(32'h39140671),
	.w6(32'hbb602c45),
	.w7(32'hbab0dea6),
	.w8(32'hbb099236),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b138ce7),
	.w1(32'h3ab716c3),
	.w2(32'hbc0342db),
	.w3(32'h3bcbc703),
	.w4(32'h3c04a0c2),
	.w5(32'hbbb49ea0),
	.w6(32'h3b64a9a2),
	.w7(32'h3b80dca1),
	.w8(32'hbbd03968),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dd168),
	.w1(32'hbbba523d),
	.w2(32'h3b9984ae),
	.w3(32'hbbf165bb),
	.w4(32'hbbe693a4),
	.w5(32'h39d4bf90),
	.w6(32'hbad06cc5),
	.w7(32'hba461f9c),
	.w8(32'h3b493f4b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d550c),
	.w1(32'hb9a2243a),
	.w2(32'h3b38f43a),
	.w3(32'hbbbc3653),
	.w4(32'hbae0ee89),
	.w5(32'hbae96083),
	.w6(32'h37fb3504),
	.w7(32'h3b15d4e1),
	.w8(32'hbb244b32),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8583),
	.w1(32'h3b40cfa7),
	.w2(32'hbb6765ae),
	.w3(32'h3a26c0c0),
	.w4(32'hbb7ef2a7),
	.w5(32'hbbe58874),
	.w6(32'hba32797b),
	.w7(32'hb982bfb8),
	.w8(32'h3a4fc835),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c98bf),
	.w1(32'hba9fed30),
	.w2(32'h3bb887c4),
	.w3(32'hbaa5f082),
	.w4(32'hbb22c3fc),
	.w5(32'h3cbbdb02),
	.w6(32'hbab2ce6e),
	.w7(32'hbae4d5cc),
	.w8(32'h3c9ede46),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9695b1),
	.w1(32'h3c592b91),
	.w2(32'h3aba4ad1),
	.w3(32'h3d5391c0),
	.w4(32'h3d2d048c),
	.w5(32'h3b4359d2),
	.w6(32'h3d3d398d),
	.w7(32'h3d1a5363),
	.w8(32'h3aea29de),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1b51d),
	.w1(32'h3be59331),
	.w2(32'h3b87c9d5),
	.w3(32'h3bbea345),
	.w4(32'h3bf47a4f),
	.w5(32'h3bdad5e7),
	.w6(32'h3b5cfd37),
	.w7(32'h3ba6c788),
	.w8(32'h3bf8b0e9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d82aa),
	.w1(32'hbb3202dd),
	.w2(32'h3ab7dd9e),
	.w3(32'h3c276eb5),
	.w4(32'h3a34e834),
	.w5(32'h3b41d66a),
	.w6(32'h3b881c34),
	.w7(32'h3af05686),
	.w8(32'h3a627585),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088427),
	.w1(32'hb8201816),
	.w2(32'h3c018ae1),
	.w3(32'hbb36a9b8),
	.w4(32'hbaa560ad),
	.w5(32'h3bc8bde4),
	.w6(32'hbb934d89),
	.w7(32'hbaefebe8),
	.w8(32'h3b6f4e80),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4147e0),
	.w1(32'h3b880a12),
	.w2(32'h3bd29e4f),
	.w3(32'h3b337cd4),
	.w4(32'h3bc267a3),
	.w5(32'h3be3d2f3),
	.w6(32'h3aa4564c),
	.w7(32'h3b942510),
	.w8(32'h3c32e5c0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f3c8a),
	.w1(32'h3ba19385),
	.w2(32'hb9b6a664),
	.w3(32'hbb09abee),
	.w4(32'h3ae03eba),
	.w5(32'h3aeff738),
	.w6(32'h3b65e0d8),
	.w7(32'h3bf2bad3),
	.w8(32'h3aad5858),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2b131),
	.w1(32'hba867cf2),
	.w2(32'hbbb1dbb6),
	.w3(32'h3bc79135),
	.w4(32'h3b64b384),
	.w5(32'hbc053ef2),
	.w6(32'h3b005154),
	.w7(32'h3aff8674),
	.w8(32'hbb31dcf0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb2516),
	.w1(32'hbb8e9705),
	.w2(32'h38c9630f),
	.w3(32'hbb2d1290),
	.w4(32'hbb920545),
	.w5(32'h3b4aee30),
	.w6(32'hbad88cc5),
	.w7(32'hba46f01a),
	.w8(32'hba3bcb3f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d72a2),
	.w1(32'hbb109ff0),
	.w2(32'hbb9f91cd),
	.w3(32'hbb0dcbfa),
	.w4(32'hbb206447),
	.w5(32'h3b2215d8),
	.w6(32'h3a5dadaa),
	.w7(32'hbac595cb),
	.w8(32'hb83110e9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabab1b5),
	.w1(32'hbc1d5a9d),
	.w2(32'h3b558921),
	.w3(32'hbb6d63cf),
	.w4(32'h3aec4f71),
	.w5(32'h3b65c422),
	.w6(32'h3b08924d),
	.w7(32'hba24b4a5),
	.w8(32'h3aeea72c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc939ba),
	.w1(32'h39fe788e),
	.w2(32'h3ba406ba),
	.w3(32'hb956f8ef),
	.w4(32'hbac75048),
	.w5(32'h3adeeaae),
	.w6(32'h3a9bf63f),
	.w7(32'hbb3a3e83),
	.w8(32'h3bcea616),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c110c4f),
	.w1(32'h3c031741),
	.w2(32'hbaa665ca),
	.w3(32'h3c3beb80),
	.w4(32'h3c04e44c),
	.w5(32'hbaf8601f),
	.w6(32'h3c006121),
	.w7(32'h3be06335),
	.w8(32'h3aff2d27),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12b670),
	.w1(32'hbaf393d8),
	.w2(32'h3a73b3f1),
	.w3(32'h3b4a1fd1),
	.w4(32'h3b9a4445),
	.w5(32'hbabff429),
	.w6(32'h3bb3371b),
	.w7(32'h3c03b490),
	.w8(32'hbaecb9c6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c8a3),
	.w1(32'h3a0fa6a1),
	.w2(32'hbc85ba19),
	.w3(32'h3b5ce5df),
	.w4(32'h3ba9ea17),
	.w5(32'hbcaaf092),
	.w6(32'hbb57c71f),
	.w7(32'h3b3f7f13),
	.w8(32'hbc9c3aeb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8caae3),
	.w1(32'hbc371cfc),
	.w2(32'h3b105b8d),
	.w3(32'hbc95809e),
	.w4(32'hbbdf5862),
	.w5(32'h3b864e6f),
	.w6(32'hbc4c8a8b),
	.w7(32'hbb29d39f),
	.w8(32'h3c1db340),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35445e),
	.w1(32'h3bb2a9a6),
	.w2(32'hbc13b66a),
	.w3(32'h3c981d37),
	.w4(32'h3c8df07b),
	.w5(32'hbc7835fc),
	.w6(32'h3cc63e5b),
	.w7(32'h3cf16b47),
	.w8(32'hbc14f615),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a14e5),
	.w1(32'hbc5f5239),
	.w2(32'hbc148e8b),
	.w3(32'hbc9df8e0),
	.w4(32'hbc8f9d68),
	.w5(32'hbc5201b5),
	.w6(32'hbbb93745),
	.w7(32'hbbef7459),
	.w8(32'hbc2b1195),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc508864),
	.w1(32'hbc3329df),
	.w2(32'hba6af752),
	.w3(32'hbc53cbd1),
	.w4(32'hbc34d037),
	.w5(32'h3aa1ba28),
	.w6(32'hbc230009),
	.w7(32'hbbf3972f),
	.w8(32'h3bc70094),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcb2fd),
	.w1(32'h3a58348e),
	.w2(32'h3b4c90e1),
	.w3(32'h3c04b3cb),
	.w4(32'h3bd73588),
	.w5(32'h3b92f085),
	.w6(32'h3bedf55d),
	.w7(32'h3b02f98e),
	.w8(32'h3bf7e6f3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea80e8),
	.w1(32'h3c09bf81),
	.w2(32'hba6fc6fe),
	.w3(32'h3a26b6c4),
	.w4(32'h3befa050),
	.w5(32'h3c142121),
	.w6(32'h39ab6474),
	.w7(32'h3c0b3ee6),
	.w8(32'h3aa41e44),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e78fc),
	.w1(32'hbb202426),
	.w2(32'h3aeb7455),
	.w3(32'h3c639c18),
	.w4(32'h3c378393),
	.w5(32'h39ebeb4c),
	.w6(32'h3bb7b142),
	.w7(32'h3b9075d1),
	.w8(32'hbaca35f2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4084a),
	.w1(32'h3b1d0964),
	.w2(32'hbb17281d),
	.w3(32'hbaf1982b),
	.w4(32'h3a2db731),
	.w5(32'hba097348),
	.w6(32'hbb69d6cd),
	.w7(32'hba135fb0),
	.w8(32'hbbbc4e37),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab683df),
	.w1(32'h3b858e52),
	.w2(32'h3d07161c),
	.w3(32'h3a0b3cae),
	.w4(32'h3bb8c0b0),
	.w5(32'h3d52a1e4),
	.w6(32'hbb3cdf85),
	.w7(32'h3b1ad9de),
	.w8(32'h3d30e818),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5b2c34),
	.w1(32'h3d39acd0),
	.w2(32'hbaa3ef03),
	.w3(32'h3dc148ee),
	.w4(32'h3d9deff5),
	.w5(32'hb9685bf6),
	.w6(32'h3da48f9a),
	.w7(32'h3d83ea08),
	.w8(32'hb9999db9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8082ac),
	.w1(32'hba2ff8ea),
	.w2(32'h3be00730),
	.w3(32'h3a06448b),
	.w4(32'hbb71529c),
	.w5(32'h3baa6f42),
	.w6(32'h3be0bd37),
	.w7(32'h3b343aa1),
	.w8(32'h3b0b8138),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26295b),
	.w1(32'h3b827370),
	.w2(32'hbbae01a8),
	.w3(32'hb8ed16af),
	.w4(32'h3b97e296),
	.w5(32'hbaeb68d4),
	.w6(32'h3a5bf475),
	.w7(32'h3b97f461),
	.w8(32'hba64e780),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05ac3),
	.w1(32'hbbbae8cd),
	.w2(32'h3aace68c),
	.w3(32'h3ae3d639),
	.w4(32'hba91cba7),
	.w5(32'hbb174197),
	.w6(32'h3b3d281b),
	.w7(32'hbab0f2fc),
	.w8(32'hba8ea154),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacd5c6),
	.w1(32'hbc55d663),
	.w2(32'hba37076c),
	.w3(32'hbbf6e04a),
	.w4(32'hbc8d44c1),
	.w5(32'hb9336437),
	.w6(32'hbba26589),
	.w7(32'hbc9163bd),
	.w8(32'hbb4616c8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43f0de),
	.w1(32'hbaa62e0b),
	.w2(32'h3b046c60),
	.w3(32'hbc079e3c),
	.w4(32'hbb4e8d70),
	.w5(32'hb9bff53e),
	.w6(32'hbbbb6bf8),
	.w7(32'hbabdd935),
	.w8(32'h3aa3d4c6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e9705),
	.w1(32'hba00d5c7),
	.w2(32'hbbae2cec),
	.w3(32'hba3f9e6f),
	.w4(32'h3948d3bb),
	.w5(32'hbbda82f6),
	.w6(32'hb8b39ec1),
	.w7(32'h3b1cd2d8),
	.w8(32'hbb91117b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0aa46),
	.w1(32'hbb8328c7),
	.w2(32'h3aa83ad3),
	.w3(32'hbb5b4b09),
	.w4(32'hbbc274df),
	.w5(32'h3c02629e),
	.w6(32'hba142b30),
	.w7(32'hbbc4b552),
	.w8(32'h3be3f0a0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f91c4),
	.w1(32'hbb187379),
	.w2(32'h3b0b3504),
	.w3(32'h3c3afdb5),
	.w4(32'h3bd00af5),
	.w5(32'hbb4cf934),
	.w6(32'h3c4ad757),
	.w7(32'h3ba1225c),
	.w8(32'hbb5c7234),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f041f),
	.w1(32'hbb82cc34),
	.w2(32'hbab8f69a),
	.w3(32'hbc144761),
	.w4(32'hbc084f5a),
	.w5(32'h3b03e829),
	.w6(32'hbbe83618),
	.w7(32'hbc086e96),
	.w8(32'h3a943b6b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b640f08),
	.w1(32'hbbad0bda),
	.w2(32'hba78c6a9),
	.w3(32'h3adf1d66),
	.w4(32'h3b03e748),
	.w5(32'h3a5f9f57),
	.w6(32'h3b2042b5),
	.w7(32'h3b6b8caf),
	.w8(32'hbb20779c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b73cb),
	.w1(32'hbaac508a),
	.w2(32'h3b378b73),
	.w3(32'hbbf14da2),
	.w4(32'hbb158390),
	.w5(32'h3b80353d),
	.w6(32'hbb938091),
	.w7(32'h3a3d0a56),
	.w8(32'h3b74c615),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9a4dc),
	.w1(32'h3bc99a9e),
	.w2(32'h3bbe6728),
	.w3(32'hbbbccc32),
	.w4(32'h3b7f9cce),
	.w5(32'h3ba774d6),
	.w6(32'hbb73ec3f),
	.w7(32'h3b45e752),
	.w8(32'h3c27633a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf320f),
	.w1(32'h3c0d352f),
	.w2(32'h3b90197d),
	.w3(32'h3cf5a1c2),
	.w4(32'h3c754ca8),
	.w5(32'h3bad6908),
	.w6(32'h3c95b912),
	.w7(32'h3c52ee7b),
	.w8(32'h3b0e6521),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f77a71),
	.w1(32'hb9e41322),
	.w2(32'h3b47f958),
	.w3(32'hbaabc645),
	.w4(32'hb88ffacb),
	.w5(32'h3cd92a7e),
	.w6(32'h3a2e9e77),
	.w7(32'h3a0ddf82),
	.w8(32'h3c85fcd2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1206ed),
	.w1(32'h3ca2be23),
	.w2(32'h3ae29f9a),
	.w3(32'h3db7d26d),
	.w4(32'h3d82749d),
	.w5(32'h3b8d4384),
	.w6(32'h3d93b34e),
	.w7(32'h3d3340d5),
	.w8(32'hba88057a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b455fcc),
	.w1(32'h3c1c2b80),
	.w2(32'h3ad1895f),
	.w3(32'h3beeaece),
	.w4(32'h3c09b2f7),
	.w5(32'h3bd85b7c),
	.w6(32'h3bc54b87),
	.w7(32'h3befabfa),
	.w8(32'h3bd9b5fd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ae23),
	.w1(32'h3ab23aa2),
	.w2(32'hbba7444d),
	.w3(32'h3b9d4210),
	.w4(32'hba8026f4),
	.w5(32'hba573f5e),
	.w6(32'h3c2325be),
	.w7(32'hba03af9e),
	.w8(32'h3a946263),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6372dd),
	.w1(32'hbb0588ce),
	.w2(32'hbb152f34),
	.w3(32'hbb6329f9),
	.w4(32'h3a0f86a4),
	.w5(32'hbaa29ceb),
	.w6(32'hbbf89418),
	.w7(32'hbb714cfd),
	.w8(32'h3a87bb5d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd35920),
	.w1(32'h3b37bc4e),
	.w2(32'hb933ef36),
	.w3(32'hba8520fc),
	.w4(32'h3b2878a5),
	.w5(32'h3b10ed4a),
	.w6(32'h3b0b7fad),
	.w7(32'h3c0942ea),
	.w8(32'hba1bc98e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6b8d),
	.w1(32'h3ae07d1b),
	.w2(32'h3c2a31a2),
	.w3(32'h3c0aa615),
	.w4(32'h3bbfe421),
	.w5(32'h3c880556),
	.w6(32'h3c325249),
	.w7(32'h3c065982),
	.w8(32'h3c878ea9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ea51c),
	.w1(32'h3c609971),
	.w2(32'hbac72720),
	.w3(32'h3cb72aac),
	.w4(32'h3cb3e9e7),
	.w5(32'h3a0231f2),
	.w6(32'h3cc31436),
	.w7(32'h3caf8e90),
	.w8(32'h3b337db5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70ae72),
	.w1(32'h3b3dc83f),
	.w2(32'hba0d1dd4),
	.w3(32'hbb2e85e8),
	.w4(32'hbb2bb1d6),
	.w5(32'hbb22066f),
	.w6(32'h3ad3eefd),
	.w7(32'h3b916ef2),
	.w8(32'h3bb1401e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb653b8e),
	.w1(32'hbb57b540),
	.w2(32'hbb6d1c8d),
	.w3(32'hba9f8814),
	.w4(32'hba8922a6),
	.w5(32'hba220e82),
	.w6(32'h3b243ffa),
	.w7(32'hb89fc2ac),
	.w8(32'hbc1d323c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7c98),
	.w1(32'h3b25bb9c),
	.w2(32'hbc858449),
	.w3(32'h3c09399b),
	.w4(32'h3be6fdec),
	.w5(32'hbcc5593c),
	.w6(32'hbb22fc31),
	.w7(32'hbbb6ef96),
	.w8(32'hbcbb9e5b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc44122),
	.w1(32'hbc795fa9),
	.w2(32'h3b8335ad),
	.w3(32'hbcd62c97),
	.w4(32'hbc92f85f),
	.w5(32'h3ba09c7d),
	.w6(32'hbcce1dac),
	.w7(32'hbc6e0772),
	.w8(32'h3bb32769),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac53876),
	.w1(32'hbb295da3),
	.w2(32'h3b6db726),
	.w3(32'h3b5045de),
	.w4(32'h3a95cd96),
	.w5(32'h3c8fffcb),
	.w6(32'h3b2c20d1),
	.w7(32'h3a234b1e),
	.w8(32'h3c85e103),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e7547),
	.w1(32'h3c1390a5),
	.w2(32'h3be9ece7),
	.w3(32'h3d3c0531),
	.w4(32'h3d0b09bc),
	.w5(32'h3bad7f6c),
	.w6(32'h3d2be5b7),
	.w7(32'h3cf9ecb2),
	.w8(32'h3bc55a53),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acac1a1),
	.w1(32'h3a89b61c),
	.w2(32'h3a325add),
	.w3(32'hbb3e7a2c),
	.w4(32'h3a6b6a8d),
	.w5(32'h3c0930b9),
	.w6(32'h3af3c015),
	.w7(32'h3b41dc50),
	.w8(32'h3aef7f82),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c6c80b),
	.w1(32'h3b900b08),
	.w2(32'h3bc70f03),
	.w3(32'h3b866b1b),
	.w4(32'h3b625b09),
	.w5(32'h3b156876),
	.w6(32'h3bf7d73b),
	.w7(32'h3b785689),
	.w8(32'h3b513479),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d4b43),
	.w1(32'h3b668e14),
	.w2(32'hbbe33bb0),
	.w3(32'h3a91bc43),
	.w4(32'h3b276ea4),
	.w5(32'hbb80ae17),
	.w6(32'h3a918dbd),
	.w7(32'hba7d82f9),
	.w8(32'hbba61fec),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad721cc),
	.w1(32'h3a9a3be4),
	.w2(32'h3a88ae9b),
	.w3(32'hbb7f8b85),
	.w4(32'hbb594357),
	.w5(32'h3b7063b4),
	.w6(32'hbb01e812),
	.w7(32'hbb2711c4),
	.w8(32'h3b42d88a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a015),
	.w1(32'hbaf4ca91),
	.w2(32'h3b668962),
	.w3(32'h3c2ef1d3),
	.w4(32'h3b53f3a3),
	.w5(32'h3bb19ae8),
	.w6(32'h3bb42591),
	.w7(32'hbb9ed046),
	.w8(32'h3b953cde),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa4aa9),
	.w1(32'hbb9bdb7c),
	.w2(32'h3b0944be),
	.w3(32'h3c7906d9),
	.w4(32'hb98d3fbb),
	.w5(32'hbb92d503),
	.w6(32'h3c648dab),
	.w7(32'hbb10845a),
	.w8(32'h3a81fd37),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b466f67),
	.w1(32'h3ab90c5a),
	.w2(32'hb964aa95),
	.w3(32'hbbc12e1e),
	.w4(32'hbc04467b),
	.w5(32'hbbb5fa84),
	.w6(32'hba81e0b7),
	.w7(32'hbabdaca5),
	.w8(32'hb99c8173),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53ec7d),
	.w1(32'hbb5e9c49),
	.w2(32'h3b124cb2),
	.w3(32'hbc2641ad),
	.w4(32'hbb92bed1),
	.w5(32'h3b99850b),
	.w6(32'hbb2a5ba4),
	.w7(32'hbb2d8185),
	.w8(32'h3b44897e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c324a1e),
	.w1(32'h3b9fd924),
	.w2(32'h3a2215b9),
	.w3(32'h3c579961),
	.w4(32'h3b89b13d),
	.w5(32'h3bb259e0),
	.w6(32'h3c7da5ab),
	.w7(32'h3ba11ad3),
	.w8(32'h3aaf4f49),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada8ada),
	.w1(32'hbb9f6dc7),
	.w2(32'hbb44b429),
	.w3(32'h3b283c04),
	.w4(32'hbb877de1),
	.w5(32'hbb666b8c),
	.w6(32'h3ac3796e),
	.w7(32'hbc3d717c),
	.w8(32'hbb4fee8a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0cf9d),
	.w1(32'hbb6f69ac),
	.w2(32'h3bfe40b5),
	.w3(32'h3b33fd06),
	.w4(32'h39f6d994),
	.w5(32'h3be574f0),
	.w6(32'h3b188cd8),
	.w7(32'hb9a59e08),
	.w8(32'h3bb44c07),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6494d0),
	.w1(32'h3b57f802),
	.w2(32'h3b8684ae),
	.w3(32'h3b01baf5),
	.w4(32'h3b709dbe),
	.w5(32'h3ba75347),
	.w6(32'h3b9d852f),
	.w7(32'h3bdba9cd),
	.w8(32'h3b3afe61),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d58e4),
	.w1(32'h3b66ac17),
	.w2(32'h3ae667f5),
	.w3(32'hbabe93f9),
	.w4(32'h3bb9f655),
	.w5(32'h39cbbb0f),
	.w6(32'hb9984e01),
	.w7(32'h3b9c3021),
	.w8(32'h3b43e246),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ee54),
	.w1(32'hbbb62148),
	.w2(32'h3a1ba4bf),
	.w3(32'hb970aa0f),
	.w4(32'hbc0498a6),
	.w5(32'h3a867c0a),
	.w6(32'h3b9fa61d),
	.w7(32'hbb5e8ec4),
	.w8(32'h3aa4a068),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18fda5),
	.w1(32'h3b0f93df),
	.w2(32'h3b8ba3d4),
	.w3(32'hbac8ede3),
	.w4(32'h3b5e8058),
	.w5(32'hb9e8b989),
	.w6(32'hbb23ee7e),
	.w7(32'h3af148f6),
	.w8(32'h3b3b0151),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58d2f6),
	.w1(32'h3a8a9ca5),
	.w2(32'hbbb37c8d),
	.w3(32'hbab80ac8),
	.w4(32'h39b2f782),
	.w5(32'hbb9cb612),
	.w6(32'hbb8128d1),
	.w7(32'hbb8ed772),
	.w8(32'hbb9b3305),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb783bf5),
	.w1(32'h3b0fba74),
	.w2(32'hbb6489fc),
	.w3(32'hbad0d03c),
	.w4(32'hbb4ed295),
	.w5(32'h3a10f594),
	.w6(32'hbac55879),
	.w7(32'hbb6357be),
	.w8(32'h3996ef1f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb838901),
	.w1(32'hbb91e4b5),
	.w2(32'h3bcdaea5),
	.w3(32'hba7868db),
	.w4(32'hbb450159),
	.w5(32'h3b986543),
	.w6(32'h3b2f7804),
	.w7(32'hbbae9366),
	.w8(32'h3baca87e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c044a90),
	.w1(32'h3aa1be64),
	.w2(32'hba51b2b8),
	.w3(32'h3bdb52ad),
	.w4(32'h3b57c6b8),
	.w5(32'hbabe6e27),
	.w6(32'h3bb342e6),
	.w7(32'h3be0bbef),
	.w8(32'hbad92448),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc574e),
	.w1(32'h3b09eda6),
	.w2(32'h3ab4e24e),
	.w3(32'h3b334152),
	.w4(32'hbb52a35e),
	.w5(32'hbb8f759a),
	.w6(32'hba93f009),
	.w7(32'h3ac03b23),
	.w8(32'h3aba3c79),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f61de),
	.w1(32'hb9b88160),
	.w2(32'hbb9a38a5),
	.w3(32'h3b7c799a),
	.w4(32'hbaa37b5c),
	.w5(32'hbb795900),
	.w6(32'h3af3f161),
	.w7(32'h3c1bb68d),
	.w8(32'h39618d58),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0798d),
	.w1(32'hbc1ce00a),
	.w2(32'hbb8be413),
	.w3(32'hbbaebad4),
	.w4(32'hbc0e1db9),
	.w5(32'hbbe0773d),
	.w6(32'h3a9af256),
	.w7(32'hbaed4ade),
	.w8(32'hbc76b914),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8b3f5),
	.w1(32'hbbab4fdc),
	.w2(32'hbb78d636),
	.w3(32'hbbc2fe03),
	.w4(32'hbc00e435),
	.w5(32'h3a8144bd),
	.w6(32'hbc6b5e77),
	.w7(32'hbc752cb3),
	.w8(32'h3a2719fc),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed7c04),
	.w1(32'hbbb6d5d0),
	.w2(32'h3b107a86),
	.w3(32'h3b0df1c2),
	.w4(32'h3b504e16),
	.w5(32'hbb5a8722),
	.w6(32'h3b15d5ce),
	.w7(32'h3bb50491),
	.w8(32'h3bce98bd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc163),
	.w1(32'h39fb205c),
	.w2(32'hbab436a6),
	.w3(32'hbabf9f0b),
	.w4(32'h3ad76a5c),
	.w5(32'hb994e232),
	.w6(32'h3b7d94cc),
	.w7(32'h3b6f0635),
	.w8(32'h3b584268),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacdd79),
	.w1(32'hbb0031d1),
	.w2(32'h3baba4c0),
	.w3(32'hbad1aa15),
	.w4(32'h3b0642a9),
	.w5(32'hba4def51),
	.w6(32'h3b1546af),
	.w7(32'hb9153da1),
	.w8(32'h3b8b828a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fc710),
	.w1(32'h3be9d5ba),
	.w2(32'hbb942ae1),
	.w3(32'hbb60c219),
	.w4(32'hb719d01a),
	.w5(32'hbbbd7987),
	.w6(32'h3b85a702),
	.w7(32'h3c026677),
	.w8(32'hbbb6c075),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceb23e),
	.w1(32'hbbd92855),
	.w2(32'hba0acd35),
	.w3(32'hbc456457),
	.w4(32'hbc5a364a),
	.w5(32'hbba49708),
	.w6(32'hbc4f3bd5),
	.w7(32'hbc393c5a),
	.w8(32'hbb418448),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dd42b),
	.w1(32'hbbbf3de6),
	.w2(32'hbad15a7b),
	.w3(32'hbc2e19f6),
	.w4(32'hbc1358f2),
	.w5(32'h3c0fa86c),
	.w6(32'hbc1222df),
	.w7(32'hbc0fa116),
	.w8(32'h3ba07b30),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253cfd),
	.w1(32'hbb6a2f67),
	.w2(32'hbba10161),
	.w3(32'h3ba22185),
	.w4(32'h3b5023f1),
	.w5(32'hbb8a1c07),
	.w6(32'h3c22f004),
	.w7(32'h3bd9f8f4),
	.w8(32'h39b580c4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcb24b),
	.w1(32'h3b7d45d7),
	.w2(32'h3c064956),
	.w3(32'hbb775b31),
	.w4(32'h3b6d1e6c),
	.w5(32'h3bba6567),
	.w6(32'hb7ab773e),
	.w7(32'h3c0abe65),
	.w8(32'h3c2488cc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b538952),
	.w1(32'h3a47bc31),
	.w2(32'hbb398391),
	.w3(32'h3c060d29),
	.w4(32'h3be9ca1e),
	.w5(32'h3a9370be),
	.w6(32'h3c15a9d5),
	.w7(32'h3bf44c43),
	.w8(32'hba950c58),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74b39d),
	.w1(32'hbb97e7bb),
	.w2(32'h3b0c2f63),
	.w3(32'h39f2f6bc),
	.w4(32'hbb204f49),
	.w5(32'h3ab08d74),
	.w6(32'h3acfc808),
	.w7(32'h3aa08eb4),
	.w8(32'hbb0a881c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eccec),
	.w1(32'hbb8cdfd8),
	.w2(32'hbb58f40a),
	.w3(32'hbc28dfc6),
	.w4(32'h3aa1fe56),
	.w5(32'hbadef5d1),
	.w6(32'hbbd7df66),
	.w7(32'hbba7c7b7),
	.w8(32'h3afa704e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule