module layer_6_featuremap_9(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96cdfa),
	.w1(32'hbb55f963),
	.w2(32'h3bbd39c1),
	.w3(32'h397213b5),
	.w4(32'hbb77a46b),
	.w5(32'hbbd82162),
	.w6(32'h3accda08),
	.w7(32'h3c57ba7b),
	.w8(32'h3c09066c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a95c),
	.w1(32'hba88afe7),
	.w2(32'hba9e663c),
	.w3(32'hbb6235d4),
	.w4(32'hbab67aa7),
	.w5(32'hbab579a5),
	.w6(32'h3b242247),
	.w7(32'h3b39fa9b),
	.w8(32'h3b842611),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38bf34),
	.w1(32'hbc0640ee),
	.w2(32'h3af0dd97),
	.w3(32'hba3d9703),
	.w4(32'hbc4f7193),
	.w5(32'hbc246ba1),
	.w6(32'h3b85d4c6),
	.w7(32'hbaa62c4b),
	.w8(32'hbbbf0ce9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59fe21),
	.w1(32'h3abcb6fd),
	.w2(32'h3abbf6b8),
	.w3(32'h3b6eb911),
	.w4(32'h3bf8c01e),
	.w5(32'h3bc40227),
	.w6(32'hbae753ff),
	.w7(32'h3badd5b8),
	.w8(32'h3ac92a99),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaffc9b),
	.w1(32'hbc21ec39),
	.w2(32'hbbb20851),
	.w3(32'hbbda85a4),
	.w4(32'hbc1f1d41),
	.w5(32'hbba51a14),
	.w6(32'hbb01cd09),
	.w7(32'h3ae93f66),
	.w8(32'h3b907033),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b950c72),
	.w1(32'h39e94686),
	.w2(32'hba44ec61),
	.w3(32'h3b826532),
	.w4(32'h3b2558a7),
	.w5(32'h3ad8a6b4),
	.w6(32'h3b8c3c8c),
	.w7(32'h3aeaa3b3),
	.w8(32'h3a528e20),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a880884),
	.w1(32'h3b20e0b6),
	.w2(32'h3a9279fd),
	.w3(32'h3a8549c3),
	.w4(32'hbaf801f8),
	.w5(32'hbb1b57f8),
	.w6(32'hbb89f20f),
	.w7(32'hbb1d911b),
	.w8(32'hbaedbbde),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9043f2),
	.w1(32'h3b14e195),
	.w2(32'h3bfd5379),
	.w3(32'hbb1bef1e),
	.w4(32'h3bc6b782),
	.w5(32'h3be4a06f),
	.w6(32'h3b8edddb),
	.w7(32'h3c1b5cf7),
	.w8(32'h3b0989fd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c7e8),
	.w1(32'hbab700db),
	.w2(32'h3be8dd97),
	.w3(32'hba226e79),
	.w4(32'hbbb63d99),
	.w5(32'h3adaa1f7),
	.w6(32'h3bbdebd7),
	.w7(32'h3b2d8f49),
	.w8(32'hbacedbd8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc1184),
	.w1(32'h3aa905b0),
	.w2(32'hbad7607c),
	.w3(32'h3b99ad9e),
	.w4(32'hba4311f4),
	.w5(32'hbb322341),
	.w6(32'hbb32299f),
	.w7(32'hbac5f20f),
	.w8(32'hbb8680f2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88e1a8),
	.w1(32'hbca7bc65),
	.w2(32'hbc590511),
	.w3(32'hbc989ff5),
	.w4(32'hbcb5ee5c),
	.w5(32'hbc57e066),
	.w6(32'hbc502285),
	.w7(32'hbc7a9e8a),
	.w8(32'hbc250d97),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fb586),
	.w1(32'h3c233f24),
	.w2(32'h3b63593b),
	.w3(32'h3ae32700),
	.w4(32'h3c7268ff),
	.w5(32'h3afc8f8b),
	.w6(32'h3bc87cf2),
	.w7(32'h3bd3868c),
	.w8(32'h3be850d9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab81be6),
	.w1(32'hbba4a479),
	.w2(32'hbbad0810),
	.w3(32'hbbb2f256),
	.w4(32'hbb994dc9),
	.w5(32'hbade200d),
	.w6(32'hbb869841),
	.w7(32'hbbbe1ab2),
	.w8(32'hbb72eb8d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85a338),
	.w1(32'hbd03748a),
	.w2(32'hbcaf703f),
	.w3(32'hbc7fe3ad),
	.w4(32'hbd0ba148),
	.w5(32'hbcf1b855),
	.w6(32'hbc650c2d),
	.w7(32'hbc9b19d5),
	.w8(32'hbc90c9e4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fcae8),
	.w1(32'h3bcb5f45),
	.w2(32'h3b7d58ca),
	.w3(32'hbbcb914b),
	.w4(32'h3b1c87a7),
	.w5(32'hb9943874),
	.w6(32'h3bc1d423),
	.w7(32'h3bb78134),
	.w8(32'hba5cd072),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8f8a4),
	.w1(32'hbb09c1db),
	.w2(32'hbb2ed77e),
	.w3(32'hbc1595e4),
	.w4(32'hbb9f5849),
	.w5(32'hbb462cf2),
	.w6(32'h3ae2094f),
	.w7(32'hbb53fe26),
	.w8(32'hbb95d585),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc393312),
	.w1(32'hbc089878),
	.w2(32'h3b1a9f0f),
	.w3(32'hbc31022f),
	.w4(32'hbcc00a64),
	.w5(32'hbb416825),
	.w6(32'h3bc481b8),
	.w7(32'hbb68e6a5),
	.w8(32'hbaeecb08),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48469),
	.w1(32'h3b1e4526),
	.w2(32'h3bb82768),
	.w3(32'hbaa2bea0),
	.w4(32'h3b899bb0),
	.w5(32'h3bcd3f00),
	.w6(32'h3b2d7c92),
	.w7(32'h3bf2d4d5),
	.w8(32'h3c596522),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ee968),
	.w1(32'h3c3af50f),
	.w2(32'h3c66afbf),
	.w3(32'h3c94a1d9),
	.w4(32'h3c0d3d76),
	.w5(32'h3c59b0db),
	.w6(32'h3c09d6ba),
	.w7(32'h3c412332),
	.w8(32'h3c27fde5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0df6b8),
	.w1(32'hba359300),
	.w2(32'hbbc9549a),
	.w3(32'h3c210bab),
	.w4(32'h37b25f5f),
	.w5(32'hbb2adcf2),
	.w6(32'h3bb60847),
	.w7(32'hbb819a69),
	.w8(32'hbb8ebec6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d336),
	.w1(32'hbbdea4db),
	.w2(32'hbb9042c6),
	.w3(32'hbb91641d),
	.w4(32'hba83bc1f),
	.w5(32'hbb1c5c68),
	.w6(32'hbaeb7018),
	.w7(32'h3bdf5328),
	.w8(32'hbb0d91b3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9af5c4),
	.w1(32'hbc8397a8),
	.w2(32'hbad21a56),
	.w3(32'hbc2d368f),
	.w4(32'hbc8b991b),
	.w5(32'hbb94dbb5),
	.w6(32'h3b8b88cd),
	.w7(32'hb90560b8),
	.w8(32'hbb8e86d3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd2f2),
	.w1(32'h3b16ec82),
	.w2(32'h3b9ad557),
	.w3(32'h3c1f0f24),
	.w4(32'hba81db30),
	.w5(32'h3a041ce0),
	.w6(32'h3af16737),
	.w7(32'h3b833aac),
	.w8(32'h3b2774c3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd273014),
	.w1(32'hbd5d734d),
	.w2(32'hbc9d9dcc),
	.w3(32'hbd0fafee),
	.w4(32'hbd122187),
	.w5(32'hbcec9401),
	.w6(32'hbca2e8ab),
	.w7(32'hbc508cd0),
	.w8(32'hbce79d4e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf42e28),
	.w1(32'hbc849d32),
	.w2(32'hbbc02141),
	.w3(32'hbbd1ef05),
	.w4(32'hbc1bc637),
	.w5(32'hbb03ff10),
	.w6(32'h3b211010),
	.w7(32'h3c35476a),
	.w8(32'hba81341e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54d9b3),
	.w1(32'h3923813e),
	.w2(32'h392aa1c7),
	.w3(32'h3c0538ab),
	.w4(32'hb8ab0555),
	.w5(32'h3bdad46d),
	.w6(32'h388a5522),
	.w7(32'hbb0d0916),
	.w8(32'hbc018c76),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81d2b8),
	.w1(32'hbc34d6f1),
	.w2(32'hbbecfd93),
	.w3(32'hbbc8af0c),
	.w4(32'hbae77bc1),
	.w5(32'hbc75c545),
	.w6(32'hbb242ad2),
	.w7(32'h3b21ead4),
	.w8(32'hbb8b7850),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac23ec7),
	.w1(32'h3a773567),
	.w2(32'h3b284066),
	.w3(32'h3b08cf3b),
	.w4(32'hbb791bbb),
	.w5(32'hbb1d83df),
	.w6(32'hb934daf0),
	.w7(32'h3b45cfc9),
	.w8(32'h3a88a961),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb208542),
	.w1(32'h3ad45189),
	.w2(32'hbb5f6a1f),
	.w3(32'hbb9f5774),
	.w4(32'hbb110b84),
	.w5(32'hbb29222e),
	.w6(32'h3b4babff),
	.w7(32'hbb5d6f7a),
	.w8(32'hbb347559),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca019f),
	.w1(32'hbd2fc879),
	.w2(32'hbd1fe133),
	.w3(32'hbc78550c),
	.w4(32'h3c89945a),
	.w5(32'h3c61a881),
	.w6(32'hbca8e1bb),
	.w7(32'h3ce817a9),
	.w8(32'h3c7b386e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9773daa),
	.w1(32'hb926c639),
	.w2(32'hb88d7114),
	.w3(32'hba02ec7a),
	.w4(32'hb919ad1e),
	.w5(32'hb901a84c),
	.w6(32'hb7df1054),
	.w7(32'hb82572f2),
	.w8(32'hb8574d6b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4aebd),
	.w1(32'h3bf8d4f4),
	.w2(32'h3bf1ab39),
	.w3(32'h3bff23d7),
	.w4(32'h3c112d24),
	.w5(32'h3c11037a),
	.w6(32'h3bc25281),
	.w7(32'h3bf5e6ff),
	.w8(32'h3c073033),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8891448),
	.w1(32'hb90e8998),
	.w2(32'hb9339973),
	.w3(32'hb81c7612),
	.w4(32'hb90589de),
	.w5(32'hb9537dda),
	.w6(32'hb81e72a4),
	.w7(32'hb8c536bc),
	.w8(32'hb916460f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9503f6d),
	.w1(32'hb9919d95),
	.w2(32'hb946bec3),
	.w3(32'hb97ba5c9),
	.w4(32'hb8cf1779),
	.w5(32'hb7ea908a),
	.w6(32'hb93c1a15),
	.w7(32'hb846331a),
	.w8(32'h39082a2d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c00cd1),
	.w1(32'hb949d085),
	.w2(32'hb8a135cb),
	.w3(32'h390a245f),
	.w4(32'hb8bd8d23),
	.w5(32'hb879a998),
	.w6(32'hb83ebaf6),
	.w7(32'hb7c43e96),
	.w8(32'hb72f5ffa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b040a),
	.w1(32'hbba42f9a),
	.w2(32'hbc5a91a0),
	.w3(32'hba5276a3),
	.w4(32'hbb0e39c1),
	.w5(32'hbb1a1184),
	.w6(32'h3ab789fa),
	.w7(32'hbbb4af7c),
	.w8(32'hbbfe45fc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb304d64),
	.w1(32'hbb0cda51),
	.w2(32'hba37a915),
	.w3(32'hbb6aba75),
	.w4(32'hbb500680),
	.w5(32'hbaadb029),
	.w6(32'hbb4d80b5),
	.w7(32'hbb42310d),
	.w8(32'hbad30577),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61422c),
	.w1(32'hbbb28130),
	.w2(32'hbbc667df),
	.w3(32'hbbadc2c3),
	.w4(32'hbb283e4e),
	.w5(32'h3a2b3b8b),
	.w6(32'hba0f5ac2),
	.w7(32'hbaa42439),
	.w8(32'h392c3e2b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72abc1),
	.w1(32'h3b661bdc),
	.w2(32'h3b5494b8),
	.w3(32'h3b3ad50f),
	.w4(32'h3b14e93c),
	.w5(32'h3b012d81),
	.w6(32'h3b0f3aea),
	.w7(32'h3ac8e8f3),
	.w8(32'h3b00dcd3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac1c07),
	.w1(32'hbcb26771),
	.w2(32'h3c04360a),
	.w3(32'hbbd3009a),
	.w4(32'hbd1a1ffc),
	.w5(32'hbc6d2648),
	.w6(32'h3bbb4e43),
	.w7(32'hbc04361b),
	.w8(32'hbc4648af),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad35f1),
	.w1(32'h3c0c368b),
	.w2(32'h39a07c84),
	.w3(32'h3ab968e6),
	.w4(32'h3ae958ab),
	.w5(32'hbb5c16d9),
	.w6(32'h3b8bdfc0),
	.w7(32'h3b0dc5ed),
	.w8(32'hbbe829db),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5379bb),
	.w1(32'hbb867443),
	.w2(32'hbbe3c2e3),
	.w3(32'hbb43badc),
	.w4(32'hbade13cf),
	.w5(32'hbb01c091),
	.w6(32'h39b6ccb8),
	.w7(32'h3932f7b3),
	.w8(32'hba550a94),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb822b126),
	.w1(32'hb828a20a),
	.w2(32'hb6c40072),
	.w3(32'hb8598d7f),
	.w4(32'hb8659ee4),
	.w5(32'hb785ee86),
	.w6(32'hb80d265c),
	.w7(32'hb83f3c8f),
	.w8(32'hb7aba4df),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32675f),
	.w1(32'hbc372804),
	.w2(32'hbd154a90),
	.w3(32'hbb471a6a),
	.w4(32'h3c1a7ba8),
	.w5(32'h3bdaf62b),
	.w6(32'hbafe45c2),
	.w7(32'h3ba86dbf),
	.w8(32'hbabe2c07),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917ecb),
	.w1(32'hbc4d7c5c),
	.w2(32'h3b3bf220),
	.w3(32'h3c1a292b),
	.w4(32'hbc2188a3),
	.w5(32'hbbaae9e5),
	.w6(32'h397c832e),
	.w7(32'hbb633289),
	.w8(32'hbc108750),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b1920),
	.w1(32'h37f573ad),
	.w2(32'hb8f8cdf4),
	.w3(32'hb95c7489),
	.w4(32'hb91f79d3),
	.w5(32'hb93bcd2c),
	.w6(32'hb8823f23),
	.w7(32'hb91caad5),
	.w8(32'hb96a3fd8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb861901d),
	.w1(32'hb87a73cd),
	.w2(32'hb8f04c53),
	.w3(32'hb82d2b85),
	.w4(32'hb7c08b37),
	.w5(32'hb8075b4a),
	.w6(32'hb71e3806),
	.w7(32'h3682993e),
	.w8(32'hb7056d23),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bfb17),
	.w1(32'hbcad681d),
	.w2(32'hbc8b2e23),
	.w3(32'hbbc13e2e),
	.w4(32'hbb449ee1),
	.w5(32'hba126649),
	.w6(32'hba9d2970),
	.w7(32'h3b9d8474),
	.w8(32'h3c4af277),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ce7b0),
	.w1(32'hbab7d13c),
	.w2(32'hba4ec519),
	.w3(32'hbb3a8e54),
	.w4(32'hba19df68),
	.w5(32'h3a11e2f7),
	.w6(32'h3a50b151),
	.w7(32'h3b571817),
	.w8(32'h3bab0c5a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b4d2f),
	.w1(32'hbc650041),
	.w2(32'hbc10302b),
	.w3(32'hbb8dd116),
	.w4(32'hbc45b947),
	.w5(32'hbc126ca4),
	.w6(32'hbb3b5c39),
	.w7(32'hbba7b897),
	.w8(32'hbb6b0c5c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9b82),
	.w1(32'hb64aa413),
	.w2(32'h3a1de913),
	.w3(32'hbb22033a),
	.w4(32'hb94f9ac6),
	.w5(32'h3b69439e),
	.w6(32'hbb6e484d),
	.w7(32'hbb3ff6bf),
	.w8(32'hbaeee731),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99b1a),
	.w1(32'hbb41b3a9),
	.w2(32'hbc44a677),
	.w3(32'hbc1fe5fd),
	.w4(32'hbc10cb88),
	.w5(32'hbc349f62),
	.w6(32'hbc0243ae),
	.w7(32'hbc2b9790),
	.w8(32'hbc8899b3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccc463),
	.w1(32'hbcc2bd25),
	.w2(32'hbc803f0b),
	.w3(32'hbcc0ebd9),
	.w4(32'hbcf49327),
	.w5(32'hbcb211b8),
	.w6(32'hbc4d39ee),
	.w7(32'hbc5423b1),
	.w8(32'hbbee67c5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02da21),
	.w1(32'h3bad01d6),
	.w2(32'h3c038e1e),
	.w3(32'h3ba9bd78),
	.w4(32'h3bb656e3),
	.w5(32'h3c1b6888),
	.w6(32'h3bceb139),
	.w7(32'h3c1370cf),
	.w8(32'h3c9197f2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d160e),
	.w1(32'h3c198e2b),
	.w2(32'h3c20f3e6),
	.w3(32'h3c056686),
	.w4(32'h3bd82cce),
	.w5(32'h3bdf4e89),
	.w6(32'h3bff6505),
	.w7(32'h3ba2fcb1),
	.w8(32'h3bc8b8a4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e74e8),
	.w1(32'h3a281346),
	.w2(32'hbb6f3933),
	.w3(32'h38fc0276),
	.w4(32'h3b20e248),
	.w5(32'h3b805ffa),
	.w6(32'h3b3b210a),
	.w7(32'h3a7ecc1a),
	.w8(32'hbb5b1456),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b95b),
	.w1(32'hbba8e779),
	.w2(32'hbb561eac),
	.w3(32'hbbab3fcc),
	.w4(32'hbaf8a9f8),
	.w5(32'hba81c40f),
	.w6(32'hbb8642ae),
	.w7(32'hbaad11b2),
	.w8(32'hba0e18cd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b329ae3),
	.w1(32'h3afa87f1),
	.w2(32'h3b16b604),
	.w3(32'h3b466837),
	.w4(32'h3af36f54),
	.w5(32'h3b43e736),
	.w6(32'h3b67d93c),
	.w7(32'h3b469161),
	.w8(32'h3b4cddb9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33613e),
	.w1(32'h3ae8aecb),
	.w2(32'h3acaf199),
	.w3(32'h3b2dc87d),
	.w4(32'h3b11ca44),
	.w5(32'h3aefce3c),
	.w6(32'h3b0078e3),
	.w7(32'h3aa68f40),
	.w8(32'h3abf2f25),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a823c99),
	.w1(32'h3c2911fd),
	.w2(32'h3be90154),
	.w3(32'h3bed6bf8),
	.w4(32'hbb8df35e),
	.w5(32'hbc089709),
	.w6(32'h3c760aca),
	.w7(32'h3b853b82),
	.w8(32'hbc3dc018),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4560),
	.w1(32'h3a99e36a),
	.w2(32'h3b8e64db),
	.w3(32'h3ac35996),
	.w4(32'hb9e42af5),
	.w5(32'hba3976a5),
	.w6(32'hbb6c4c44),
	.w7(32'hbb8ba2bd),
	.w8(32'hbb761798),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb735be5),
	.w1(32'hbbd689bd),
	.w2(32'hbbf20541),
	.w3(32'h3a1fce14),
	.w4(32'hba33fbe5),
	.w5(32'h3b2206aa),
	.w6(32'h3b313efd),
	.w7(32'h3a543694),
	.w8(32'hba9df757),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac4142),
	.w1(32'hbbe12be9),
	.w2(32'hbcd2386e),
	.w3(32'h3cda5681),
	.w4(32'h3d0d09f2),
	.w5(32'h3ad0d660),
	.w6(32'h3c62ca11),
	.w7(32'h3c24b042),
	.w8(32'h3d369ab6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b717023),
	.w1(32'hbc3993d5),
	.w2(32'hbce57ca1),
	.w3(32'hbbee5bcd),
	.w4(32'hbc776514),
	.w5(32'h3bd717d5),
	.w6(32'hbc69f0c3),
	.w7(32'h3ae17309),
	.w8(32'h3c4b0914),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule