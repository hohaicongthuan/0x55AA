module layer_10_featuremap_125(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af700e5),
	.w1(32'h3cb4b49f),
	.w2(32'hbc61cea5),
	.w3(32'hba95ca6b),
	.w4(32'h3b2d4051),
	.w5(32'hbc8cde9e),
	.w6(32'h3c23674c),
	.w7(32'hbb252a3f),
	.w8(32'h3ba1fa52),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba957d),
	.w1(32'h3ba228c5),
	.w2(32'hbb1705af),
	.w3(32'hbc055aa7),
	.w4(32'h3b19938a),
	.w5(32'hbbae4827),
	.w6(32'h3b8eebd1),
	.w7(32'h3b034687),
	.w8(32'hbb1bbf66),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cee73),
	.w1(32'h3a97c27c),
	.w2(32'hbab57156),
	.w3(32'hbc1cc852),
	.w4(32'h3a3a81b9),
	.w5(32'hba7b6538),
	.w6(32'h3ab27b86),
	.w7(32'hbab64302),
	.w8(32'hb91fed97),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba962f85),
	.w1(32'h3a42b410),
	.w2(32'hbc1fb2ab),
	.w3(32'hbb0478eb),
	.w4(32'hbb1af861),
	.w5(32'hbbf4ebb0),
	.w6(32'h3bac0461),
	.w7(32'h3b3f48df),
	.w8(32'hbc0a9bee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84eb46),
	.w1(32'h3b6a3c43),
	.w2(32'h3b8c2392),
	.w3(32'hbb51a42e),
	.w4(32'h3bd46b61),
	.w5(32'h3bc621ce),
	.w6(32'h3b941983),
	.w7(32'h3c059dc8),
	.w8(32'h3bea91b1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9de326),
	.w1(32'h3ba1c701),
	.w2(32'h3c1fceaa),
	.w3(32'hbb946993),
	.w4(32'h3ae8f84b),
	.w5(32'h3a9844a6),
	.w6(32'h3bd37c51),
	.w7(32'h3c152d66),
	.w8(32'h3bf50226),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8885b),
	.w1(32'h3bbcf72c),
	.w2(32'h3b41d196),
	.w3(32'hbbd988fa),
	.w4(32'h3bd29790),
	.w5(32'hbb03ca54),
	.w6(32'h3b233482),
	.w7(32'h3baf1052),
	.w8(32'h3aa39c56),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7c1bd),
	.w1(32'hbb7d6ba9),
	.w2(32'hba453f92),
	.w3(32'hbbc74ffa),
	.w4(32'h3885d528),
	.w5(32'hb970d502),
	.w6(32'hbb8393ca),
	.w7(32'hbb2eef7b),
	.w8(32'h36b0efc5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36b0c9),
	.w1(32'h3aa5a09f),
	.w2(32'hbb8699c2),
	.w3(32'hb8cac1e4),
	.w4(32'hb9d92a3f),
	.w5(32'hbb958a9a),
	.w6(32'h3add260e),
	.w7(32'hbb38d4d7),
	.w8(32'hbb2b7631),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fa241),
	.w1(32'h3b89ad71),
	.w2(32'hbaea0426),
	.w3(32'hbabbbe02),
	.w4(32'h3a9d8d0e),
	.w5(32'h39ab726b),
	.w6(32'h3c0754dc),
	.w7(32'h3bbaae5e),
	.w8(32'h3b3d2b25),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e0f9d),
	.w1(32'hbbade8fb),
	.w2(32'hbbe4206c),
	.w3(32'hbaac9dce),
	.w4(32'hbb5d8a9b),
	.w5(32'h3b89175f),
	.w6(32'h3c108b32),
	.w7(32'h3b9aae3e),
	.w8(32'h3a955946),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9036),
	.w1(32'hbc820189),
	.w2(32'hbc6c8b25),
	.w3(32'hba09cdd8),
	.w4(32'hbc1da7fe),
	.w5(32'hbc5f3f0f),
	.w6(32'hbbd84dbe),
	.w7(32'hbbf95287),
	.w8(32'hbc0da308),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc732526),
	.w1(32'hbb0f7733),
	.w2(32'h39d2622f),
	.w3(32'hbc180c46),
	.w4(32'h3aea0a97),
	.w5(32'h3baac924),
	.w6(32'hbb815a56),
	.w7(32'hbb4b26b2),
	.w8(32'h395d85f0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b611),
	.w1(32'hbc3e0e2e),
	.w2(32'hbc2c39b4),
	.w3(32'h3a60fcd5),
	.w4(32'h3ac1026d),
	.w5(32'h3baf770a),
	.w6(32'hbc6a2e5c),
	.w7(32'hbc7275d4),
	.w8(32'hbad81dd0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a741836),
	.w1(32'hbc2b50de),
	.w2(32'hbc82d701),
	.w3(32'h3ba777c9),
	.w4(32'hbbb1dbcf),
	.w5(32'hbb4d2381),
	.w6(32'h3c1fe3f5),
	.w7(32'h3c4367e4),
	.w8(32'hbb8568fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc936c4d),
	.w1(32'h3ab1204b),
	.w2(32'hbb8891ba),
	.w3(32'hbb55783b),
	.w4(32'hbae4823d),
	.w5(32'hbbfe50d7),
	.w6(32'h3b633f36),
	.w7(32'hb99c4080),
	.w8(32'hbac74e20),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e3af),
	.w1(32'h3b49a3fd),
	.w2(32'h3baab8d3),
	.w3(32'hbb88045a),
	.w4(32'h3b97ecd1),
	.w5(32'hbab03781),
	.w6(32'h3b585d3f),
	.w7(32'h3b300bc7),
	.w8(32'h3b45b870),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc5926),
	.w1(32'h39174d1a),
	.w2(32'hbb42d9f4),
	.w3(32'hbab2ed51),
	.w4(32'hba8fc51b),
	.w5(32'hbbc53b24),
	.w6(32'h368f4f0a),
	.w7(32'h39b3de2d),
	.w8(32'hbab2934d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16be7a),
	.w1(32'h3b285784),
	.w2(32'h3b2031c3),
	.w3(32'hbbe65e73),
	.w4(32'h3b399037),
	.w5(32'h3b1b9c4b),
	.w6(32'h3a2c0b76),
	.w7(32'h3bb173f8),
	.w8(32'h3b14cda5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9858282),
	.w1(32'h3a15ce12),
	.w2(32'hbb7e79b5),
	.w3(32'h39710867),
	.w4(32'hba9a869c),
	.w5(32'hbb89eb29),
	.w6(32'h3b015ece),
	.w7(32'hbb141b48),
	.w8(32'hbad681ee),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb815885),
	.w1(32'hbbf221be),
	.w2(32'hbbe30c3b),
	.w3(32'hbb51620d),
	.w4(32'hb89f60cb),
	.w5(32'h3a267d5d),
	.w6(32'hbbb7912a),
	.w7(32'hbb889861),
	.w8(32'hba19f960),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1bec9),
	.w1(32'h3bc7e558),
	.w2(32'hbc39315c),
	.w3(32'h3b678596),
	.w4(32'hbae185a6),
	.w5(32'hbb6d4f65),
	.w6(32'hbbcbb185),
	.w7(32'hbca364da),
	.w8(32'hbc36279c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64fe22),
	.w1(32'h3b794ac1),
	.w2(32'hbb3fa715),
	.w3(32'hbc3a1b95),
	.w4(32'h3b0c7fed),
	.w5(32'hbb797f78),
	.w6(32'h3be75daa),
	.w7(32'h3b63635d),
	.w8(32'hb9c6defb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7e31),
	.w1(32'hbb1a4fcc),
	.w2(32'hbad7cca9),
	.w3(32'hbae5449e),
	.w4(32'h39c69860),
	.w5(32'hba64f0d4),
	.w6(32'hbb436bbc),
	.w7(32'hbb3d193e),
	.w8(32'hba56ebe3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb4e0f),
	.w1(32'h3b3fbb17),
	.w2(32'hbbdfa82d),
	.w3(32'hba8c2a2d),
	.w4(32'h3b0abc84),
	.w5(32'hbc2aaac9),
	.w6(32'h3c134be4),
	.w7(32'h3abd6604),
	.w8(32'hbb2664fb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc376c27),
	.w1(32'hbbfd2813),
	.w2(32'hba3128c9),
	.w3(32'hbbf2a616),
	.w4(32'hbb0f99cb),
	.w5(32'hbbd7c3ea),
	.w6(32'hbaf78d64),
	.w7(32'hba4b1219),
	.w8(32'hba24f5b7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a104895),
	.w1(32'h396c16fa),
	.w2(32'hbb6ceac3),
	.w3(32'hb723f965),
	.w4(32'hba5717f7),
	.w5(32'hbb79049a),
	.w6(32'h3afddda9),
	.w7(32'hb94a27b4),
	.w8(32'hba68181d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb452280),
	.w1(32'h3b95d269),
	.w2(32'hbb90fd18),
	.w3(32'hbb68d6d0),
	.w4(32'h399e8e30),
	.w5(32'hbbb4cd98),
	.w6(32'h3b9ffaec),
	.w7(32'h3ba94daa),
	.w8(32'h3b4a0507),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945832),
	.w1(32'h3b3704f2),
	.w2(32'hbb5d3978),
	.w3(32'hbab3be47),
	.w4(32'h3b9c0481),
	.w5(32'hbb4e1fd8),
	.w6(32'h3c6550ab),
	.w7(32'h3bf67e29),
	.w8(32'h3c0b6deb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb561aa6),
	.w1(32'h3b32c006),
	.w2(32'h3b322653),
	.w3(32'hbb12a58e),
	.w4(32'h3b4b7ec9),
	.w5(32'h3a1f1d8f),
	.w6(32'h3bbccdd3),
	.w7(32'h3b8f5fdf),
	.w8(32'h3b241518),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4735b),
	.w1(32'hbabbf9f6),
	.w2(32'hbb1da49b),
	.w3(32'hb842b30a),
	.w4(32'h3a71f658),
	.w5(32'h3a91e50f),
	.w6(32'hb9c86a8f),
	.w7(32'hba28e88f),
	.w8(32'h387a4b2a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ad449),
	.w1(32'hb8f9be90),
	.w2(32'h3abd53f0),
	.w3(32'h3a9cd12c),
	.w4(32'h3b00e761),
	.w5(32'h3b0c781e),
	.w6(32'h3a98144f),
	.w7(32'h3afb04c0),
	.w8(32'h3b2f7a8c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f3764),
	.w1(32'h3b6b7f69),
	.w2(32'hbb7bc7c5),
	.w3(32'h3a94b5d8),
	.w4(32'h3ab05652),
	.w5(32'h3af6d6b0),
	.w6(32'h3b122a86),
	.w7(32'hbc15c005),
	.w8(32'hbb15751e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab6fb4),
	.w1(32'hb7293c31),
	.w2(32'hba0aaef8),
	.w3(32'hbba02cc9),
	.w4(32'hb9009132),
	.w5(32'hbb99e0d9),
	.w6(32'h3bcabffe),
	.w7(32'hba8cfb27),
	.w8(32'hbbb7ef46),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ab3f8),
	.w1(32'h3c13a3ab),
	.w2(32'h3a287c8e),
	.w3(32'hbb8cc355),
	.w4(32'h3b02948d),
	.w5(32'hbb1eae0d),
	.w6(32'h3c2d349e),
	.w7(32'h3c24d3cd),
	.w8(32'h3bae197c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e7bc6),
	.w1(32'hbb7709ef),
	.w2(32'hbb9af2a1),
	.w3(32'hbbb0f8d7),
	.w4(32'hbb131798),
	.w5(32'hbba3728a),
	.w6(32'hba8d102e),
	.w7(32'hb8b01f52),
	.w8(32'hba0a8419),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e025d),
	.w1(32'h3be924f5),
	.w2(32'h3afc65a4),
	.w3(32'hbb914b69),
	.w4(32'h3ba63291),
	.w5(32'hbb8975b8),
	.w6(32'h3bfc3625),
	.w7(32'h3bec4b50),
	.w8(32'hbb73c5a6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56ad03),
	.w1(32'h3b117615),
	.w2(32'hbad2f4ed),
	.w3(32'hbc430aad),
	.w4(32'h3a3090e1),
	.w5(32'hbb90fa7f),
	.w6(32'h3acef9f5),
	.w7(32'h3b550548),
	.w8(32'hba81b5cf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b68ca),
	.w1(32'hbaaf3fac),
	.w2(32'hb9a2d729),
	.w3(32'hbbd859db),
	.w4(32'h39c18199),
	.w5(32'h39810925),
	.w6(32'hbad18256),
	.w7(32'hba229116),
	.w8(32'h39a34de7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fe498),
	.w1(32'h3b9a124c),
	.w2(32'h3a899f76),
	.w3(32'hb71a3069),
	.w4(32'h3b515994),
	.w5(32'hba3a60e9),
	.w6(32'h3b376cce),
	.w7(32'h3ba31eb6),
	.w8(32'hba9a00d5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd6673),
	.w1(32'h3bff8d9e),
	.w2(32'hb779f97a),
	.w3(32'hbba29f23),
	.w4(32'h3c03c44e),
	.w5(32'hba18cfa2),
	.w6(32'h3c2d9b58),
	.w7(32'h3bd2c3a9),
	.w8(32'h3ada774f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b083e),
	.w1(32'h3be50cb9),
	.w2(32'hba9e6588),
	.w3(32'hbb3091dd),
	.w4(32'h3abdba6f),
	.w5(32'hbb414b08),
	.w6(32'h3c042411),
	.w7(32'h3b4f3ff4),
	.w8(32'hbb167537),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba45c),
	.w1(32'h3b5b5296),
	.w2(32'h3b6c0c4f),
	.w3(32'hbb4d9d35),
	.w4(32'h3b981229),
	.w5(32'h3b9055f8),
	.w6(32'h391ea916),
	.w7(32'h3a81cd30),
	.w8(32'h3b4f2435),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d3a4e),
	.w1(32'h3bc162da),
	.w2(32'hbaacfa95),
	.w3(32'h3ab30124),
	.w4(32'h3b3e60b8),
	.w5(32'hbb9d874b),
	.w6(32'h3c421cf1),
	.w7(32'h3c025acf),
	.w8(32'h3bc5fa20),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d0552),
	.w1(32'hbb76edd0),
	.w2(32'hbc500751),
	.w3(32'hbb604a3b),
	.w4(32'hbb8e6cd7),
	.w5(32'hba138a72),
	.w6(32'hbb4d5414),
	.w7(32'hbc18c928),
	.w8(32'hbba0ead9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdfd37),
	.w1(32'h3b1d96ca),
	.w2(32'h3c1f49cb),
	.w3(32'hbb685d3c),
	.w4(32'h3b8b06c3),
	.w5(32'h3bbeabb3),
	.w6(32'hbb213599),
	.w7(32'h3ad90a51),
	.w8(32'h3bcc441f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43a3c),
	.w1(32'hbc285824),
	.w2(32'hbca0e72f),
	.w3(32'h3aae72f5),
	.w4(32'hbb4a3384),
	.w5(32'hbc6fb4e4),
	.w6(32'h3a7c0061),
	.w7(32'hbb39fa5a),
	.w8(32'hbbb17b22),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc811634),
	.w1(32'h3b862cf5),
	.w2(32'h3b0e331c),
	.w3(32'hbacc9a6c),
	.w4(32'h3b071339),
	.w5(32'hb9a776ab),
	.w6(32'h3c0c71c5),
	.w7(32'h3c1e2cb9),
	.w8(32'h3bb47d22),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0bbb),
	.w1(32'h3b21f47f),
	.w2(32'h3a46b8f2),
	.w3(32'hbb12c3bc),
	.w4(32'h3b216a92),
	.w5(32'hba1c718b),
	.w6(32'h3a3716a0),
	.w7(32'hb8efafcb),
	.w8(32'h3a92dbda),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2b9b6),
	.w1(32'hbb91f9c4),
	.w2(32'hbb265add),
	.w3(32'hbaed0ad7),
	.w4(32'h39a98337),
	.w5(32'h3a0834f4),
	.w6(32'hbb8e1970),
	.w7(32'hbba01933),
	.w8(32'hbb3efc42),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e698a7),
	.w1(32'hbbe38cdc),
	.w2(32'hbc0404ef),
	.w3(32'h3a68d35b),
	.w4(32'h3b10747f),
	.w5(32'hb94619cd),
	.w6(32'hbbce588b),
	.w7(32'hbbf8d969),
	.w8(32'hbb8c98f0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01d5db),
	.w1(32'hbbb2fc1b),
	.w2(32'hbc5023ad),
	.w3(32'h3b0e4ba0),
	.w4(32'hbc5d7689),
	.w5(32'hbce1070d),
	.w6(32'hbaae4ca9),
	.w7(32'hbc8b0ff2),
	.w8(32'hbc6d00a6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6fd6c),
	.w1(32'h3b9f1160),
	.w2(32'hbb14d1ba),
	.w3(32'hbccccae6),
	.w4(32'hba70a84b),
	.w5(32'hbc78f1bb),
	.w6(32'h3c226425),
	.w7(32'h3bdf678e),
	.w8(32'hba7035fd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f0f26),
	.w1(32'h3b6d3e39),
	.w2(32'h3c3c60b5),
	.w3(32'hbca5b513),
	.w4(32'h3c038b31),
	.w5(32'h3badd0ca),
	.w6(32'h3be953d3),
	.w7(32'h3c404ea6),
	.w8(32'h3b846507),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34f0ea),
	.w1(32'hbb34904b),
	.w2(32'hbbad9b0a),
	.w3(32'hbc3ce90a),
	.w4(32'hb9e8d80d),
	.w5(32'hbbb9ac9e),
	.w6(32'h3b63a824),
	.w7(32'h3a8dd835),
	.w8(32'hbb447e3e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0302d3),
	.w1(32'hba4e85ef),
	.w2(32'hbbfce55b),
	.w3(32'hbb91ba51),
	.w4(32'h3b1e7c31),
	.w5(32'hbbfb3823),
	.w6(32'h3bb982b3),
	.w7(32'h3886805c),
	.w8(32'hba2f80d2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaede2e),
	.w1(32'hbb801e5c),
	.w2(32'hbb4736b1),
	.w3(32'hbb7bb40b),
	.w4(32'h3b3278e6),
	.w5(32'h39a013a1),
	.w6(32'hbb628e83),
	.w7(32'hbba30b1e),
	.w8(32'h3b1ab94e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395e0b),
	.w1(32'hbb077ccd),
	.w2(32'h3bc6064e),
	.w3(32'h3a6a55cf),
	.w4(32'h3c06e2a7),
	.w5(32'h3c2df240),
	.w6(32'hbb0f3b6d),
	.w7(32'h3bbc47b2),
	.w8(32'h3c064604),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb930371),
	.w1(32'h3b804717),
	.w2(32'hbb8f30ee),
	.w3(32'h39101c4b),
	.w4(32'hba20202c),
	.w5(32'hbbeae038),
	.w6(32'h3b5d479b),
	.w7(32'h3888a896),
	.w8(32'hbb5b72fb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17950f),
	.w1(32'hba6828e9),
	.w2(32'hba9ab903),
	.w3(32'hbc10b923),
	.w4(32'h3a7da18c),
	.w5(32'h396872e2),
	.w6(32'hbb4023b3),
	.w7(32'hbb0d7369),
	.w8(32'hb985848d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e300a),
	.w1(32'h3b9475dd),
	.w2(32'h3b233a05),
	.w3(32'hba382a49),
	.w4(32'h3b3fe39c),
	.w5(32'hbb01d684),
	.w6(32'h3b9087d1),
	.w7(32'h3b988ec1),
	.w8(32'h3b0e6fda),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ed2c),
	.w1(32'hba316bb1),
	.w2(32'hbba6955a),
	.w3(32'hbb27a92d),
	.w4(32'h3ae7f069),
	.w5(32'h3b0c5644),
	.w6(32'hbaab8333),
	.w7(32'hbb60622e),
	.w8(32'hb90cedd0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb19c),
	.w1(32'h3c26a5a4),
	.w2(32'hbb81d897),
	.w3(32'h3b0ace99),
	.w4(32'hba647bc0),
	.w5(32'hbb741623),
	.w6(32'h3be4212f),
	.w7(32'hbb3a6561),
	.w8(32'hbba5a082),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc45541),
	.w1(32'h3baa1318),
	.w2(32'h382ed054),
	.w3(32'hba65c665),
	.w4(32'h3b198669),
	.w5(32'hbb27e0ec),
	.w6(32'h3c16fac8),
	.w7(32'h3bdf13e2),
	.w8(32'h3ba00273),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb088562),
	.w1(32'hbacffd8e),
	.w2(32'h3a8fb0ce),
	.w3(32'hbb1a2e32),
	.w4(32'hba98c4e7),
	.w5(32'h39c077c1),
	.w6(32'h39dc08cf),
	.w7(32'hb9f2bc4f),
	.w8(32'hba19e126),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe554c),
	.w1(32'hba9f81cd),
	.w2(32'h3c9f21cc),
	.w3(32'hba62c147),
	.w4(32'h3bd805ad),
	.w5(32'h3c2957ef),
	.w6(32'hbc287e83),
	.w7(32'hba3cdce1),
	.w8(32'h3c000cb3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be84674),
	.w1(32'h3c10d87c),
	.w2(32'h3b838244),
	.w3(32'hbb93dfca),
	.w4(32'h3c016ef4),
	.w5(32'h3b5da24c),
	.w6(32'h3c07bee7),
	.w7(32'h3bf3001a),
	.w8(32'h3b7ef13f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3838334d),
	.w1(32'h3be7e665),
	.w2(32'hbb22ea28),
	.w3(32'hba8b64a7),
	.w4(32'h3c20f918),
	.w5(32'hbb1c11bc),
	.w6(32'h3c16f90c),
	.w7(32'h3bf6ef36),
	.w8(32'h3af8aeb7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0eed3),
	.w1(32'h390c8be0),
	.w2(32'hbb0c1fe8),
	.w3(32'hbb5c83f7),
	.w4(32'h3a4c0a2d),
	.w5(32'hbbc48d50),
	.w6(32'h3b2fa7bd),
	.w7(32'h3abf1872),
	.w8(32'hba67dbc0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6d368),
	.w1(32'hba471ae2),
	.w2(32'h3c0500e8),
	.w3(32'hbba47a2f),
	.w4(32'h3c46a491),
	.w5(32'h3c439fcb),
	.w6(32'hbb9df362),
	.w7(32'h3af51d0b),
	.w8(32'h3bbcaa1c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a73e9),
	.w1(32'h3b87457f),
	.w2(32'hbb4e7e9b),
	.w3(32'h3c2d2019),
	.w4(32'h3a5ffabc),
	.w5(32'hbbb1b102),
	.w6(32'h3b665f94),
	.w7(32'h3af3c649),
	.w8(32'hbb1c4f50),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e034e),
	.w1(32'hbab0a8f6),
	.w2(32'h3abd293c),
	.w3(32'hbbf9766d),
	.w4(32'h3b0eef65),
	.w5(32'h39e1a369),
	.w6(32'hbaa0d5f0),
	.w7(32'hb9a5721e),
	.w8(32'h3b138fbc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2174e8),
	.w1(32'hba57c305),
	.w2(32'hba44b583),
	.w3(32'hbaa67c54),
	.w4(32'h39f8a59d),
	.w5(32'hba10c2a2),
	.w6(32'hbabcb880),
	.w7(32'hba85083b),
	.w8(32'h39eb7d13),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922e90f),
	.w1(32'hbb177464),
	.w2(32'hbaeb32aa),
	.w3(32'hba522119),
	.w4(32'hb8c31e26),
	.w5(32'h394db3b2),
	.w6(32'hb91ef32e),
	.w7(32'h3a1ba914),
	.w8(32'h39ff2712),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7f9d4),
	.w1(32'h3b21cdb5),
	.w2(32'hbbc45c21),
	.w3(32'hb9a2cab6),
	.w4(32'hba51e543),
	.w5(32'hbc26df51),
	.w6(32'h3b85191a),
	.w7(32'hba838886),
	.w8(32'hbb9e1962),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38c69b),
	.w1(32'hbbd8e24c),
	.w2(32'hbac0bd3a),
	.w3(32'hbc1d5f1f),
	.w4(32'hbb296ec7),
	.w5(32'hbc3f9f4d),
	.w6(32'h3b04c329),
	.w7(32'hbbfd5209),
	.w8(32'hbc0c4df5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0744),
	.w1(32'hbb6dc759),
	.w2(32'h3a225104),
	.w3(32'hbb2dd9e9),
	.w4(32'h3a899327),
	.w5(32'h3b907cfb),
	.w6(32'hbb31ef29),
	.w7(32'hbb2557f4),
	.w8(32'h3b5dfafd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87315d),
	.w1(32'h3a1f7c17),
	.w2(32'hbb339dcb),
	.w3(32'h3b890701),
	.w4(32'hbab3e229),
	.w5(32'hbb82f087),
	.w6(32'h39aac50b),
	.w7(32'hbaff184e),
	.w8(32'hbb30fcdd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ebf9),
	.w1(32'hbb8a0fd5),
	.w2(32'hbb27285e),
	.w3(32'hbafc1377),
	.w4(32'hbb1b6c07),
	.w5(32'hbbd2e374),
	.w6(32'h3b1f7bb2),
	.w7(32'hbb922125),
	.w8(32'hbb1b989c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb6366),
	.w1(32'hbb03d9f2),
	.w2(32'hbb4f7411),
	.w3(32'hbb06d21a),
	.w4(32'h3acd5d1b),
	.w5(32'h3b43cc2f),
	.w6(32'hba5d581e),
	.w7(32'hbb05f6b4),
	.w8(32'h3a0871d1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0380d3),
	.w1(32'h3c2bacd8),
	.w2(32'h39f4933a),
	.w3(32'h3ae53f61),
	.w4(32'h3c2b71f0),
	.w5(32'hbb040658),
	.w6(32'h3c55671a),
	.w7(32'h3c2c4b90),
	.w8(32'h3b879ef2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba185f4),
	.w1(32'h3bd8ce6b),
	.w2(32'h3a8e7c95),
	.w3(32'hbba7ae15),
	.w4(32'h3b913912),
	.w5(32'hbaebc094),
	.w6(32'h3be7f98a),
	.w7(32'h3b7f580a),
	.w8(32'hbaecff2c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870833),
	.w1(32'h3beedfe6),
	.w2(32'hbb1d00b5),
	.w3(32'hbb703492),
	.w4(32'h3b7b5299),
	.w5(32'hbbc9539b),
	.w6(32'h3c3f6087),
	.w7(32'h3bc0fbc0),
	.w8(32'h3afa1f0c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7ad9),
	.w1(32'h3b6b089d),
	.w2(32'hbb177d2b),
	.w3(32'hbbb52865),
	.w4(32'hbaf84c7b),
	.w5(32'hbc0188a9),
	.w6(32'h3b79520c),
	.w7(32'h3b0e19c5),
	.w8(32'hbab56387),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6bdb1),
	.w1(32'h3be1a419),
	.w2(32'h3c03a79e),
	.w3(32'hbbfc4a90),
	.w4(32'h38f0e70c),
	.w5(32'h3ba60ba9),
	.w6(32'h3bd31848),
	.w7(32'h3c52cd63),
	.w8(32'h397aec67),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8ec1),
	.w1(32'h3aaa68d9),
	.w2(32'hbae948b5),
	.w3(32'hba65fe5f),
	.w4(32'h3a990900),
	.w5(32'hbb9186ad),
	.w6(32'h3a827f37),
	.w7(32'hba835e38),
	.w8(32'hb99d2518),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71f85e),
	.w1(32'hbbc9bcb0),
	.w2(32'hbba6f0dd),
	.w3(32'hbb8d9014),
	.w4(32'hb9dad290),
	.w5(32'hbb0d0dc8),
	.w6(32'hbbcfbeaf),
	.w7(32'hbbf4948a),
	.w8(32'hbb6aa887),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba890ec9),
	.w1(32'hbb16bf8a),
	.w2(32'hbb06f211),
	.w3(32'hb95a4dc3),
	.w4(32'h3a17fd13),
	.w5(32'h3aab1502),
	.w6(32'hbaaf4b00),
	.w7(32'hba6df939),
	.w8(32'hb8385793),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92e5dc),
	.w1(32'h3b6df641),
	.w2(32'hbb3900e9),
	.w3(32'h3a94e063),
	.w4(32'h3b4a6ee0),
	.w5(32'hbbc22f28),
	.w6(32'h3bdd7b2f),
	.w7(32'h3b8cffbc),
	.w8(32'hb96bcfd0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0677a),
	.w1(32'hbb2a22b5),
	.w2(32'hbb3c26eb),
	.w3(32'hbbc07921),
	.w4(32'h39421c16),
	.w5(32'h3a06b309),
	.w6(32'hba46b0c3),
	.w7(32'hbaac59ce),
	.w8(32'h3ace48a8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398560cf),
	.w1(32'hbafc9a9f),
	.w2(32'hbab90df3),
	.w3(32'h3b7c2f8d),
	.w4(32'h3b06432b),
	.w5(32'h3b1052cd),
	.w6(32'hb9e79eb0),
	.w7(32'h39ebe1c2),
	.w8(32'h3a9acad0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993cede),
	.w1(32'h3927b4a2),
	.w2(32'hbb7cc3c2),
	.w3(32'h3ab6322a),
	.w4(32'hba797cc5),
	.w5(32'hbb5d8990),
	.w6(32'h3afe13df),
	.w7(32'h3a8a887f),
	.w8(32'hba0cbec7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf73c96),
	.w1(32'h3be91e6d),
	.w2(32'hbabcae83),
	.w3(32'hbba5d33f),
	.w4(32'h3759db31),
	.w5(32'hbc06b7c2),
	.w6(32'h3c19b96d),
	.w7(32'h3ba0af27),
	.w8(32'hbb046513),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc255dec),
	.w1(32'h3be0c6e6),
	.w2(32'hbbb48af1),
	.w3(32'hbc49d42a),
	.w4(32'h3bebc24f),
	.w5(32'hbbced859),
	.w6(32'h3c547955),
	.w7(32'h3bdbf55f),
	.w8(32'h3b7e7b9c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbabf50),
	.w1(32'h3b819a3e),
	.w2(32'hb9c0d37e),
	.w3(32'hbba5e9be),
	.w4(32'h3a01533e),
	.w5(32'hb9b0316d),
	.w6(32'h3b2cb954),
	.w7(32'h3aac79b0),
	.w8(32'h3a9347d3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f252d),
	.w1(32'h3bbc2399),
	.w2(32'h3cabc490),
	.w3(32'hba567363),
	.w4(32'h3af2ec2c),
	.w5(32'h3b4d0023),
	.w6(32'hbb1880a3),
	.w7(32'h3beafe32),
	.w8(32'h3bfc967e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c892b),
	.w1(32'h3b7b1920),
	.w2(32'h3a45c16f),
	.w3(32'hbc47ea71),
	.w4(32'h3aaff799),
	.w5(32'hbaf16945),
	.w6(32'h3b197171),
	.w7(32'h3ace38c2),
	.w8(32'hbc01a07b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee593f),
	.w1(32'h3b90a234),
	.w2(32'hbb2810d3),
	.w3(32'hbb188aed),
	.w4(32'h3b104cb8),
	.w5(32'hbaf7e519),
	.w6(32'h3bb0638a),
	.w7(32'hb95b3b6c),
	.w8(32'hbab3c920),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd010b0),
	.w1(32'h3c081e7c),
	.w2(32'h3badfb6d),
	.w3(32'hbb8be425),
	.w4(32'h3bc669a7),
	.w5(32'h3a94a73c),
	.w6(32'h3bc42b1b),
	.w7(32'h3bdd73df),
	.w8(32'hbaba3317),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bccbf),
	.w1(32'h3bb82808),
	.w2(32'hbb83219f),
	.w3(32'hbbae37ad),
	.w4(32'h3a76af97),
	.w5(32'hbc3a5d9f),
	.w6(32'h3c08bdba),
	.w7(32'h3bdefe84),
	.w8(32'hba9df62d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65134e),
	.w1(32'hbc5ce71f),
	.w2(32'hbc36f98a),
	.w3(32'hbc7521a0),
	.w4(32'hbb83e00d),
	.w5(32'hbba63a38),
	.w6(32'hbb87b633),
	.w7(32'hbc0a22c7),
	.w8(32'hbbf32664),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc829125),
	.w1(32'h3c5902c6),
	.w2(32'h3d1540c0),
	.w3(32'hbc72f627),
	.w4(32'h3b291c74),
	.w5(32'h3c324b69),
	.w6(32'h3851174b),
	.w7(32'h3ab7f63c),
	.w8(32'h3b49d4bc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8016ef),
	.w1(32'hbbae5e2e),
	.w2(32'h3a8ba477),
	.w3(32'hbc67a3ab),
	.w4(32'h3b06ae28),
	.w5(32'h3be5fbe3),
	.w6(32'hbb90384d),
	.w7(32'hbb7b4bc5),
	.w8(32'h3babc512),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2e7c3),
	.w1(32'hbb2269d4),
	.w2(32'h3a6b8213),
	.w3(32'h3bde0612),
	.w4(32'h3a004b81),
	.w5(32'h3a855c85),
	.w6(32'h3a7db970),
	.w7(32'h3af7fe47),
	.w8(32'h3ae5e2fb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b79ae),
	.w1(32'hbb29264c),
	.w2(32'h39d5be85),
	.w3(32'hba8a9f78),
	.w4(32'h3a25cbf9),
	.w5(32'h3b44ceb0),
	.w6(32'hbadda0c7),
	.w7(32'hbae53424),
	.w8(32'h3b221d20),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395317),
	.w1(32'hb9db615c),
	.w2(32'hbb6766a3),
	.w3(32'h3b33c21c),
	.w4(32'hb9f7f530),
	.w5(32'hbb29e691),
	.w6(32'hb96b7768),
	.w7(32'hbb22b386),
	.w8(32'hbafbe810),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d219b),
	.w1(32'h3afae68b),
	.w2(32'hbb812ed6),
	.w3(32'hbaea9b03),
	.w4(32'hba0af4f1),
	.w5(32'hbacbb745),
	.w6(32'h3b6082e9),
	.w7(32'h3a5cf225),
	.w8(32'hbb1a1fee),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d9b94),
	.w1(32'hbb9da127),
	.w2(32'hbbb66dc7),
	.w3(32'hbb146108),
	.w4(32'h3a0c3a16),
	.w5(32'h3a3d735f),
	.w6(32'hbaf7c1f5),
	.w7(32'hbb016a84),
	.w8(32'hba72d177),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc7a68),
	.w1(32'hbb37578f),
	.w2(32'h3a278236),
	.w3(32'h3b05ca23),
	.w4(32'h3aa24465),
	.w5(32'h3b77c83a),
	.w6(32'hbb290a04),
	.w7(32'hbb0ffa17),
	.w8(32'h3b2e1d89),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c89b),
	.w1(32'hbbffdd48),
	.w2(32'hbbaa6501),
	.w3(32'h3b596a09),
	.w4(32'hbb751926),
	.w5(32'hbac4f288),
	.w6(32'hbc1013fd),
	.w7(32'hbc323f21),
	.w8(32'hbb833041),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2b1c),
	.w1(32'hbb30574c),
	.w2(32'hbc18d27a),
	.w3(32'hbb57c94f),
	.w4(32'hbbae638d),
	.w5(32'hbc2a2b4c),
	.w6(32'hba0efb80),
	.w7(32'hbb870f00),
	.w8(32'hbb4a0ac7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8e4ac),
	.w1(32'hbb50b17c),
	.w2(32'hbc964eba),
	.w3(32'hbb9342d3),
	.w4(32'hbbb7e473),
	.w5(32'hbc6582e5),
	.w6(32'hbc07b0e0),
	.w7(32'hbcb2ade2),
	.w8(32'hbc014478),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc602f3a),
	.w1(32'hbb074042),
	.w2(32'hbbe07a34),
	.w3(32'hbc00dd06),
	.w4(32'hbba01757),
	.w5(32'hbc1f276b),
	.w6(32'h3b4a27a4),
	.w7(32'h3a87da4d),
	.w8(32'hbb40d32e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21a7a5),
	.w1(32'h3a2b5176),
	.w2(32'hbb5c2e7b),
	.w3(32'hbbd64bbe),
	.w4(32'hbadc5d64),
	.w5(32'h3aeb299e),
	.w6(32'h3aecfee9),
	.w7(32'hbb3281ee),
	.w8(32'hbaeeeb57),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dfdf3),
	.w1(32'h39bfab38),
	.w2(32'hbb989fb0),
	.w3(32'h3b6c535a),
	.w4(32'h3ba1e826),
	.w5(32'h39faf745),
	.w6(32'hbb02c63e),
	.w7(32'hbbbfcb7a),
	.w8(32'h3a50b17f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ef787),
	.w1(32'hbb7bb03f),
	.w2(32'h3a71d057),
	.w3(32'h36db96f7),
	.w4(32'h3ab674d4),
	.w5(32'h3baa0924),
	.w6(32'hbb3f0efe),
	.w7(32'hbb3193c7),
	.w8(32'h3b83886b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1dd31),
	.w1(32'h39a0e5d2),
	.w2(32'h3b35d0a6),
	.w3(32'h3ba0ee99),
	.w4(32'h3aa95453),
	.w5(32'h3b004c39),
	.w6(32'hb9fca4ca),
	.w7(32'h39d98cd5),
	.w8(32'h3b338a1f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a0611),
	.w1(32'h3a6d51e6),
	.w2(32'h3b62722e),
	.w3(32'h3a126c22),
	.w4(32'h3a90a880),
	.w5(32'h3b3b4e2f),
	.w6(32'h3a3fcebb),
	.w7(32'h3ad80866),
	.w8(32'h3b64afaa),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b283eb6),
	.w1(32'h3b802249),
	.w2(32'hbadb8a34),
	.w3(32'hb9a3a218),
	.w4(32'h3bcdbe9a),
	.w5(32'h3bb67be3),
	.w6(32'hbb851dbc),
	.w7(32'hbc0131f1),
	.w8(32'h3a995c4e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dd204),
	.w1(32'hbb7945a2),
	.w2(32'h3ac5553e),
	.w3(32'hba414766),
	.w4(32'h3a4fcebe),
	.w5(32'hba2d6318),
	.w6(32'hbbc959d0),
	.w7(32'h3b08ef34),
	.w8(32'h38e355c4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7f77c),
	.w1(32'h3b9d994d),
	.w2(32'h3a6f1d85),
	.w3(32'hbb691ffe),
	.w4(32'h3abd19b6),
	.w5(32'hb99717e4),
	.w6(32'h3c051c9a),
	.w7(32'h3c15fecc),
	.w8(32'h3b690c0a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb55b3),
	.w1(32'h3c04f721),
	.w2(32'hbaf6414d),
	.w3(32'hbc0f3cb5),
	.w4(32'h3a154a96),
	.w5(32'hbbb2310c),
	.w6(32'h3bab9144),
	.w7(32'h3b03e245),
	.w8(32'hba424d02),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fc2a4),
	.w1(32'hbaff2418),
	.w2(32'hba5f98fd),
	.w3(32'hbc024026),
	.w4(32'h39cbbf14),
	.w5(32'h39303b5c),
	.w6(32'hbb4a71d6),
	.w7(32'hbb3b5bf8),
	.w8(32'hba6114ce),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a874f61),
	.w1(32'h3c8c7fb0),
	.w2(32'h3c8a253c),
	.w3(32'hba061039),
	.w4(32'h3b941c02),
	.w5(32'h3b0f81af),
	.w6(32'h3bbe4c50),
	.w7(32'h3ba0cf03),
	.w8(32'h3c4832c0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7d1e4),
	.w1(32'h3c0d2221),
	.w2(32'h3c55a541),
	.w3(32'h3bc1cca2),
	.w4(32'h3a8aa0ac),
	.w5(32'hbbc5d611),
	.w6(32'h3c61ac8d),
	.w7(32'h3c5eae42),
	.w8(32'h3b51b937),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ceeb),
	.w1(32'hbb8d2f44),
	.w2(32'hbb50804b),
	.w3(32'hbca19818),
	.w4(32'hb9a2ffa9),
	.w5(32'h3b01195b),
	.w6(32'hbb2355b4),
	.w7(32'hba16895e),
	.w8(32'hba83fa75),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07786c),
	.w1(32'hb8b351b9),
	.w2(32'hb8e00876),
	.w3(32'h393f0106),
	.w4(32'hb8529436),
	.w5(32'hb8a01aad),
	.w6(32'hb8860aeb),
	.w7(32'hb89497b6),
	.w8(32'hb8ddf7f9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86097a6),
	.w1(32'hb87fa173),
	.w2(32'hb8c2666f),
	.w3(32'hb7b8ac59),
	.w4(32'hb79441ed),
	.w5(32'hb82e7afb),
	.w6(32'hb81b26d6),
	.w7(32'hb80d94b1),
	.w8(32'hb871563e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c11127),
	.w1(32'hba01e842),
	.w2(32'hb9f0e3bd),
	.w3(32'hb98718dd),
	.w4(32'hb9d066be),
	.w5(32'hb9e2d507),
	.w6(32'hb9a0bd69),
	.w7(32'hb9dfd8fa),
	.w8(32'hb9ec9620),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3576a235),
	.w1(32'h34bad35a),
	.w2(32'h352ee31a),
	.w3(32'hb5e50f6e),
	.w4(32'hb5a0b78d),
	.w5(32'hb4e06528),
	.w6(32'h35c5eb46),
	.w7(32'hb648c3a6),
	.w8(32'hb5b1dc23),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836f494),
	.w1(32'h3517486c),
	.w2(32'hb787747d),
	.w3(32'h35095802),
	.w4(32'h37de9de6),
	.w5(32'h378a60f8),
	.w6(32'h370a22c6),
	.w7(32'h38177efe),
	.w8(32'h369d3307),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71afe5d),
	.w1(32'h342e137e),
	.w2(32'hb689a5e4),
	.w3(32'hb5f254eb),
	.w4(32'h36d80ea8),
	.w5(32'h33ab5b0b),
	.w6(32'hb6e5badd),
	.w7(32'h367d9ca7),
	.w8(32'hb57fdfaa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee956d),
	.w1(32'hb8ec4d23),
	.w2(32'hb9131c4f),
	.w3(32'hb8c7190c),
	.w4(32'hb8c8024d),
	.w5(32'hb8fe320b),
	.w6(32'hb8afd72c),
	.w7(32'hb8837c5e),
	.w8(32'hb8c94519),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9162af7),
	.w1(32'hb95c522f),
	.w2(32'hb9323732),
	.w3(32'hb8b8c3f8),
	.w4(32'hb924982a),
	.w5(32'hb95882b5),
	.w6(32'hb8d5ea0f),
	.w7(32'hb92b168f),
	.w8(32'hb91b3572),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94eab51),
	.w1(32'hb94418ba),
	.w2(32'hb96bf731),
	.w3(32'hb91b14ef),
	.w4(32'hb8f25cad),
	.w5(32'hb93750ab),
	.w6(32'hb92bb579),
	.w7(32'hb920208f),
	.w8(32'hb95a53e7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92859ab),
	.w1(32'hb916ffc0),
	.w2(32'hb92108dd),
	.w3(32'hb8cf98f2),
	.w4(32'hb8ad6ff9),
	.w5(32'hb9030582),
	.w6(32'hb8ab70ed),
	.w7(32'hb88aad01),
	.w8(32'hb8f7da08),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c0ceb),
	.w1(32'hb96028c6),
	.w2(32'hb94c4dd9),
	.w3(32'hb9292fd1),
	.w4(32'hb931825b),
	.w5(32'hb93da754),
	.w6(32'hb93b0644),
	.w7(32'hb96143a6),
	.w8(32'hb9628f0e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5b19f),
	.w1(32'hb90a67aa),
	.w2(32'hb9259ac5),
	.w3(32'hb88e625c),
	.w4(32'hb8b669a0),
	.w5(32'hb907bf4d),
	.w6(32'hb8a9ede1),
	.w7(32'hb8b572de),
	.w8(32'hb91f789c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf9eb4),
	.w1(32'hb81d6f14),
	.w2(32'hb8112cf1),
	.w3(32'hb884324e),
	.w4(32'hb723bc31),
	.w5(32'hb747587c),
	.w6(32'hb891efe3),
	.w7(32'hb7fc1941),
	.w8(32'hb82e8672),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96269e3),
	.w1(32'hb9769a1c),
	.w2(32'hb986ede8),
	.w3(32'hb93ffcb4),
	.w4(32'hb9354245),
	.w5(32'hb960bbe2),
	.w6(32'hb949f669),
	.w7(32'hb946e696),
	.w8(32'hb984ae7e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d2a93),
	.w1(32'hb86c4b40),
	.w2(32'hb89d7ace),
	.w3(32'hb81adef0),
	.w4(32'hb817e8ba),
	.w5(32'hb87bf0bc),
	.w6(32'hb8380133),
	.w7(32'hb83e580a),
	.w8(32'hb89455b8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ed13f),
	.w1(32'hb93042aa),
	.w2(32'hb9394d8d),
	.w3(32'hb91b8095),
	.w4(32'hb8cc8156),
	.w5(32'hb913b3c5),
	.w6(32'hb91f5462),
	.w7(32'hb9094b4a),
	.w8(32'hb93606ce),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8933058),
	.w1(32'hb88e8482),
	.w2(32'hb8a324d6),
	.w3(32'hb85629dc),
	.w4(32'hb87ca1f6),
	.w5(32'hb868b43e),
	.w6(32'hb86893e9),
	.w7(32'hb8776a11),
	.w8(32'hb86e3831),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36db58b9),
	.w1(32'h369cd50d),
	.w2(32'h3674fd5d),
	.w3(32'h365029da),
	.w4(32'h363aca7e),
	.w5(32'h359082ba),
	.w6(32'h368b8ee7),
	.w7(32'h36c488d9),
	.w8(32'hb4072724),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36279073),
	.w1(32'h36971133),
	.w2(32'h361f2934),
	.w3(32'h357001a1),
	.w4(32'h36aa97be),
	.w5(32'h362117f9),
	.w6(32'h368087a5),
	.w7(32'h36e3a4f9),
	.w8(32'h35c5adeb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7067989),
	.w1(32'h3610f545),
	.w2(32'h3628e587),
	.w3(32'hb6802d1c),
	.w4(32'hb5657337),
	.w5(32'h3507c7b8),
	.w6(32'hb6655bfe),
	.w7(32'hb66a91be),
	.w8(32'hb2796f4c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdea3f),
	.w1(32'hb8206536),
	.w2(32'hb89b8aff),
	.w3(32'hb8a52f8c),
	.w4(32'hb78bdfc4),
	.w5(32'hb8345718),
	.w6(32'hb8b0841a),
	.w7(32'hb8468c2c),
	.w8(32'hb867add2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918f92a),
	.w1(32'hb92474a6),
	.w2(32'hb947d5e6),
	.w3(32'hb8f232d7),
	.w4(32'hb8d84855),
	.w5(32'hb92b320c),
	.w6(32'hb90110d3),
	.w7(32'hb916f7c1),
	.w8(32'hb93a1203),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e67ea4),
	.w1(32'hb5bbf4f6),
	.w2(32'hb5b74b71),
	.w3(32'hb52d2147),
	.w4(32'hb6b80e83),
	.w5(32'hb6f96b5a),
	.w6(32'h35a83c9c),
	.w7(32'hb5aaac91),
	.w8(32'hb680b6ce),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9746272),
	.w1(32'hb98012de),
	.w2(32'hb990ee7b),
	.w3(32'hb93cfedf),
	.w4(32'hb92e3fde),
	.w5(32'hb95aee33),
	.w6(32'hb94fac45),
	.w7(32'hb952dee2),
	.w8(32'hb98366b2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995e266),
	.w1(32'hb9b8bb77),
	.w2(32'hb9d9caa0),
	.w3(32'hb98f27bb),
	.w4(32'hb9a4054f),
	.w5(32'hb9c3586d),
	.w6(32'hb9b324d8),
	.w7(32'hb9d454a7),
	.w8(32'hb9f55041),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9232f85),
	.w1(32'hb947b69a),
	.w2(32'hb985326b),
	.w3(32'hb9099636),
	.w4(32'hb91269e5),
	.w5(32'hb96a4c39),
	.w6(32'hb90d6b7d),
	.w7(32'hb9299004),
	.w8(32'hb9847e9b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9a3a6),
	.w1(32'hb799e9b9),
	.w2(32'hb81eef57),
	.w3(32'hb82af08a),
	.w4(32'h3829c61e),
	.w5(32'hb64ff356),
	.w6(32'hb8211cea),
	.w7(32'h3797ebb5),
	.w8(32'hb731c599),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b3671),
	.w1(32'hb8c41a5d),
	.w2(32'hb62c042e),
	.w3(32'hb8ac73dd),
	.w4(32'hb887cab1),
	.w5(32'hb7d0ca86),
	.w6(32'hb9192b1e),
	.w7(32'hb9108cf7),
	.w8(32'hb90f3587),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6d163),
	.w1(32'hb8732adf),
	.w2(32'hb75e9c06),
	.w3(32'hb8d224fd),
	.w4(32'hb93bcb93),
	.w5(32'hb8ef0042),
	.w6(32'hb844d96b),
	.w7(32'hb95b7fb4),
	.w8(32'hb8ae764d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cfc80c),
	.w1(32'hb818d645),
	.w2(32'hb7851c78),
	.w3(32'hb6a21bfa),
	.w4(32'h373adb51),
	.w5(32'hb8192583),
	.w6(32'h38afb05b),
	.w7(32'h385b6c74),
	.w8(32'hb8b6337e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722d2f9),
	.w1(32'h38660be3),
	.w2(32'h37af0e0c),
	.w3(32'h3803ce4c),
	.w4(32'h389fb3f2),
	.w5(32'h3846c5cf),
	.w6(32'h378aceaf),
	.w7(32'h381e7435),
	.w8(32'h3770e51c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38232e82),
	.w1(32'h38c3c792),
	.w2(32'h3795dd9e),
	.w3(32'h38b9699a),
	.w4(32'h3919e3d8),
	.w5(32'h38a5694e),
	.w6(32'h38aae975),
	.w7(32'h390f8eb2),
	.w8(32'h388d1de1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5643389),
	.w1(32'h36e2fe1b),
	.w2(32'hb71bf0af),
	.w3(32'h368799e1),
	.w4(32'h36d8d5e3),
	.w5(32'hb7174ae2),
	.w6(32'h369726b6),
	.w7(32'h3692151f),
	.w8(32'hb6f610e3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34c6845b),
	.w1(32'h35eec71c),
	.w2(32'h3620ebca),
	.w3(32'h354fce25),
	.w4(32'h35851804),
	.w5(32'h35c787ca),
	.w6(32'h36201e32),
	.w7(32'h349ea774),
	.w8(32'h360ea8be),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9142f23),
	.w1(32'hb912dbc3),
	.w2(32'hb92d045c),
	.w3(32'hb8b27794),
	.w4(32'hb8afcb7f),
	.w5(32'hb9030203),
	.w6(32'hb8ee9d73),
	.w7(32'hb8ee3e4f),
	.w8(32'hb91b66b0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb673cf16),
	.w1(32'h368f820b),
	.w2(32'hb66bd309),
	.w3(32'hb43acdb4),
	.w4(32'h35e52cc4),
	.w5(32'hb6ab4a51),
	.w6(32'h376399cc),
	.w7(32'h3712a926),
	.w8(32'h345df348),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d86082),
	.w1(32'hb8d0d7f3),
	.w2(32'hb8d42cf6),
	.w3(32'hb89c6f17),
	.w4(32'hb8a4e76b),
	.w5(32'hb8c27ed5),
	.w6(32'hb8b48fa1),
	.w7(32'hb8a61163),
	.w8(32'hb8db3032),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a3c68f),
	.w1(32'h38610ee7),
	.w2(32'hb7e24e81),
	.w3(32'h37fc597f),
	.w4(32'h38a0b3c8),
	.w5(32'h38203a60),
	.w6(32'h37ec4116),
	.w7(32'h388224b4),
	.w8(32'h36fddd84),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a810a),
	.w1(32'h39020c9b),
	.w2(32'hb6e454ba),
	.w3(32'h38d4abb9),
	.w4(32'h392979b6),
	.w5(32'h3802f607),
	.w6(32'h38338f7e),
	.w7(32'h38cdbda3),
	.w8(32'hb7f67413),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853b852),
	.w1(32'hb83d5009),
	.w2(32'hb726a783),
	.w3(32'hb86d0b08),
	.w4(32'hb82f397c),
	.w5(32'hb75bb3dc),
	.w6(32'hb889b64e),
	.w7(32'hb84bad62),
	.w8(32'hb8036ef3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d888c2),
	.w1(32'hb7f16ebc),
	.w2(32'hb8303383),
	.w3(32'h37cb507a),
	.w4(32'hb76b9eb9),
	.w5(32'hb7f87989),
	.w6(32'h36d4a5e2),
	.w7(32'hb7c2a442),
	.w8(32'hb874cb5e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904d0cc),
	.w1(32'hb9343e4d),
	.w2(32'hb9645f57),
	.w3(32'hb854f12b),
	.w4(32'hb8e064f3),
	.w5(32'hb960fb5f),
	.w6(32'hb86ee36d),
	.w7(32'hb8835776),
	.w8(32'hb94e1b81),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b53072),
	.w1(32'hb9a70735),
	.w2(32'hb9b25469),
	.w3(32'hb99e33f3),
	.w4(32'hb98b0452),
	.w5(32'hb9a7fc07),
	.w6(32'hb9d09147),
	.w7(32'hb9cc539f),
	.w8(32'hb9e304b3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d3765),
	.w1(32'h376fb142),
	.w2(32'hb7985b66),
	.w3(32'h3876aa28),
	.w4(32'h38e12d47),
	.w5(32'h383a441b),
	.w6(32'h39018bdf),
	.w7(32'h39116ade),
	.w8(32'h37ee3cf7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991ceed),
	.w1(32'hb992781e),
	.w2(32'hb9da415a),
	.w3(32'hb93f30a3),
	.w4(32'hb9367e33),
	.w5(32'hb9bcdfaa),
	.w6(32'hb96f0b9f),
	.w7(32'hb94a2fc8),
	.w8(32'hb9c7a141),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb857cfa1),
	.w1(32'hb83ad7b9),
	.w2(32'hb8687163),
	.w3(32'hb8108e92),
	.w4(32'hb79be49b),
	.w5(32'hb825af01),
	.w6(32'hb8077002),
	.w7(32'hb8007eb7),
	.w8(32'hb85ab940),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946bd01),
	.w1(32'hb8e9d0c6),
	.w2(32'hb9425966),
	.w3(32'hb8ae38b0),
	.w4(32'h370064df),
	.w5(32'hb879bee2),
	.w6(32'hb8b57409),
	.w7(32'hb7fd16d7),
	.w8(32'hb89c2c09),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9937a1b),
	.w1(32'hb9589723),
	.w2(32'hb9abf71c),
	.w3(32'hb91d3a11),
	.w4(32'hb88ad410),
	.w5(32'hb96e9858),
	.w6(32'hb9341294),
	.w7(32'hb8ef0a66),
	.w8(32'hb972c1c1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990119d),
	.w1(32'hb993e4f2),
	.w2(32'hb9d0e05c),
	.w3(32'hb968d3c5),
	.w4(32'hb9843105),
	.w5(32'hb9bd780e),
	.w6(32'hb988022e),
	.w7(32'hb98e821d),
	.w8(32'hb9d2ff0b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883bcc5),
	.w1(32'h3509ef32),
	.w2(32'h37de4e70),
	.w3(32'hb8a5cb07),
	.w4(32'hb5237aa7),
	.w5(32'h37becc6a),
	.w6(32'hb83d7380),
	.w7(32'h382cc42c),
	.w8(32'h384930c7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f4ac8b),
	.w1(32'hb91317e9),
	.w2(32'hb90e3b01),
	.w3(32'hb8e658cd),
	.w4(32'hb915d966),
	.w5(32'hb9134842),
	.w6(32'hb8ea2d74),
	.w7(32'hb93091fd),
	.w8(32'hb9409674),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36caee63),
	.w1(32'h3692f0c9),
	.w2(32'h36e83edf),
	.w3(32'h35f73d7d),
	.w4(32'h34a8e996),
	.w5(32'h362be79c),
	.w6(32'h3615e38c),
	.w7(32'hb5bb80a8),
	.w8(32'h35a3f91d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d5e5aa),
	.w1(32'hb6411bac),
	.w2(32'hb7ff5edf),
	.w3(32'hb7ae0661),
	.w4(32'h36c2a0dd),
	.w5(32'hb78ca283),
	.w6(32'hb7ad9557),
	.w7(32'h371608f5),
	.w8(32'hb780d612),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da70a0),
	.w1(32'hb7533a3d),
	.w2(32'hb7df07e9),
	.w3(32'hb7873cf5),
	.w4(32'hb7168527),
	.w5(32'hb7c89240),
	.w6(32'hb78d4a12),
	.w7(32'hb739542c),
	.w8(32'hb79506f8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c27086),
	.w1(32'hb8782d5c),
	.w2(32'hb8b1c85d),
	.w3(32'hb85f8b2e),
	.w4(32'hb7135400),
	.w5(32'hb8368d6d),
	.w6(32'hb86f270e),
	.w7(32'hb766f531),
	.w8(32'hb84a7c2a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb519a1e0),
	.w1(32'hb4f2ec79),
	.w2(32'h35fd759c),
	.w3(32'hb5f89669),
	.w4(32'hb678f421),
	.w5(32'hb5c60ab2),
	.w6(32'hb5529674),
	.w7(32'hb5c72736),
	.w8(32'h352a8081),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cd28ce),
	.w1(32'hb6c8047b),
	.w2(32'hb5bab248),
	.w3(32'hb4bd6278),
	.w4(32'hb69cf71c),
	.w5(32'hb689a106),
	.w6(32'hb588697e),
	.w7(32'h353a5e65),
	.w8(32'hb651138c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67aaebf),
	.w1(32'h36b4db7e),
	.w2(32'h36a5612e),
	.w3(32'hb5785348),
	.w4(32'h3692f0bb),
	.w5(32'h368e7746),
	.w6(32'h35d9cec5),
	.w7(32'h35f74cc6),
	.w8(32'h36cfbee4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3e095),
	.w1(32'hb86bf618),
	.w2(32'hb91a9f32),
	.w3(32'hb87a5f88),
	.w4(32'h364332cb),
	.w5(32'hb8ab649c),
	.w6(32'hb8426933),
	.w7(32'hb68f5b9e),
	.w8(32'hb8da909c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d669e6),
	.w1(32'hb6b2fc4e),
	.w2(32'hb6f76b7c),
	.w3(32'h357ef44f),
	.w4(32'hb74b780b),
	.w5(32'hb72346ee),
	.w6(32'h357c781c),
	.w7(32'hb799aed9),
	.w8(32'hb7f1fefe),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bf0df0),
	.w1(32'hb6b4b891),
	.w2(32'hb6e1e1c7),
	.w3(32'hb70164e4),
	.w4(32'h36b63b74),
	.w5(32'hb494620d),
	.w6(32'hb685c381),
	.w7(32'h34a21d94),
	.w8(32'hb65750e1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f71a37),
	.w1(32'hb9de9733),
	.w2(32'hb9b19ace),
	.w3(32'hb9c89a60),
	.w4(32'hb9b65d43),
	.w5(32'hb9999555),
	.w6(32'hb9a72994),
	.w7(32'hb99bc46f),
	.w8(32'hb9965bcd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dc78b),
	.w1(32'hb93bd3e3),
	.w2(32'hb9391233),
	.w3(32'hb975a2de),
	.w4(32'hb902b30c),
	.w5(32'hb9262ff2),
	.w6(32'hb960bc93),
	.w7(32'hb89dacaf),
	.w8(32'hb9044f07),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7adaff0),
	.w1(32'hb7a97648),
	.w2(32'h34dd0060),
	.w3(32'hb74afde1),
	.w4(32'hb769e230),
	.w5(32'h35aaa134),
	.w6(32'hb6d3c4b0),
	.w7(32'hb76f1af4),
	.w8(32'hb6e0bfd0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34599196),
	.w1(32'h35820bbc),
	.w2(32'h34f6c10a),
	.w3(32'h366b3645),
	.w4(32'h353a05c2),
	.w5(32'h34048334),
	.w6(32'h3616f2e0),
	.w7(32'hb580d3fe),
	.w8(32'hb58ba047),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71cf894),
	.w1(32'hb610f03a),
	.w2(32'hb808cb38),
	.w3(32'h37ca42a0),
	.w4(32'h38074ab7),
	.w5(32'hb7d64596),
	.w6(32'h37ec1770),
	.w7(32'h37b0c6da),
	.w8(32'hb7a92741),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3739155a),
	.w1(32'h3713e699),
	.w2(32'h36d0f1d3),
	.w3(32'h3725b1a0),
	.w4(32'h371bcf5d),
	.w5(32'h36bcea7b),
	.w6(32'h363e1f41),
	.w7(32'h36250715),
	.w8(32'h34ca9dd0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0aadd),
	.w1(32'hb885b96b),
	.w2(32'hb8e962b8),
	.w3(32'hb8935b3c),
	.w4(32'hb807ed3b),
	.w5(32'hb89c632f),
	.w6(32'hb8771801),
	.w7(32'hb8196256),
	.w8(32'hb8bd73e6),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971348a),
	.w1(32'hb93656d0),
	.w2(32'hb979cfbe),
	.w3(32'hb95cb050),
	.w4(32'hb5b7a63b),
	.w5(32'hb8563a44),
	.w6(32'hb9406b35),
	.w7(32'hb912b982),
	.w8(32'hb92b4533),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9894f2c),
	.w1(32'hb9a0323a),
	.w2(32'hb995107c),
	.w3(32'hb9706f05),
	.w4(32'hb983cea5),
	.w5(32'hb9973394),
	.w6(32'hb95f5b80),
	.w7(32'hb9864ce5),
	.w8(32'hb992f80d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b1b4f),
	.w1(32'hb88e465b),
	.w2(32'hb8b756a7),
	.w3(32'hb8cc1d45),
	.w4(32'hb823eb2a),
	.w5(32'hb814419b),
	.w6(32'hb90c39d1),
	.w7(32'hb8d8cf82),
	.w8(32'hb8f66d08),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e6326),
	.w1(32'hb999e3c0),
	.w2(32'hb9aa367f),
	.w3(32'hb975fffc),
	.w4(32'hb9449f6d),
	.w5(32'hb96cdefc),
	.w6(32'hb988f197),
	.w7(32'hb9302d4f),
	.w8(32'hb97e6d72),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8962f62),
	.w1(32'hb88ce831),
	.w2(32'hb8855396),
	.w3(32'hb82573b6),
	.w4(32'hb812f59f),
	.w5(32'hb81f2aa1),
	.w6(32'hb7f05ce3),
	.w7(32'hb7e87829),
	.w8(32'hb82d07bc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cf3ed0),
	.w1(32'h36a284a1),
	.w2(32'h3736dc1f),
	.w3(32'h3626bbd7),
	.w4(32'h34c60cac),
	.w5(32'h36e12518),
	.w6(32'h36551486),
	.w7(32'h3549881c),
	.w8(32'h36c99962),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374074d7),
	.w1(32'h3687aae3),
	.w2(32'h37930bc8),
	.w3(32'hb62dc80f),
	.w4(32'hb704f332),
	.w5(32'h37391d1f),
	.w6(32'hb55c7b24),
	.w7(32'hb69a26da),
	.w8(32'h371b4e44),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a94a26),
	.w1(32'h3776360a),
	.w2(32'h37c781cd),
	.w3(32'h3716ce94),
	.w4(32'h3642c286),
	.w5(32'h375d66d1),
	.w6(32'h37400bd1),
	.w7(32'h3667def8),
	.w8(32'h377173e7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914567c),
	.w1(32'hb9019044),
	.w2(32'hb94acf85),
	.w3(32'hb8b50c4d),
	.w4(32'hb88adf36),
	.w5(32'hb91bf570),
	.w6(32'hb8d6c55f),
	.w7(32'hb8bcd3bc),
	.w8(32'hb926b8c3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8d933),
	.w1(32'h369fa5eb),
	.w2(32'hb8e1be7b),
	.w3(32'h36cf9bf1),
	.w4(32'h391397df),
	.w5(32'h3717cd8f),
	.w6(32'h36ada0bf),
	.w7(32'h390762b6),
	.w8(32'h3706a9d5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98679d4),
	.w1(32'hb9513616),
	.w2(32'hb9a34410),
	.w3(32'hb90414ad),
	.w4(32'hb8892d9a),
	.w5(32'hb9502c9f),
	.w6(32'hb8fee124),
	.w7(32'hb89f8bff),
	.w8(32'hb9649013),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3799094d),
	.w1(32'h37c5e796),
	.w2(32'h3730316d),
	.w3(32'h37b2e80c),
	.w4(32'h37ddaf74),
	.w5(32'h3791aeb2),
	.w6(32'h37ac6902),
	.w7(32'h37d817a4),
	.w8(32'h3742c33f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9510e10),
	.w1(32'hb94cc4ce),
	.w2(32'hb96689e1),
	.w3(32'hb9139abb),
	.w4(32'hb905d0bf),
	.w5(32'hb9438cc0),
	.w6(32'hb904066e),
	.w7(32'hb907d5bd),
	.w8(32'hb955c345),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968bd3d),
	.w1(32'hb9840f56),
	.w2(32'hb965371b),
	.w3(32'hb940851c),
	.w4(32'hb96dce62),
	.w5(32'hb95063fe),
	.w6(32'hb94c5e9e),
	.w7(32'hb95c52de),
	.w8(32'hb9658d08),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ba7ab),
	.w1(32'hb918acf9),
	.w2(32'hb92fd2c6),
	.w3(32'hb95d9552),
	.w4(32'hb8e1ccaf),
	.w5(32'hb8d33783),
	.w6(32'hb944058e),
	.w7(32'hb8e0c6dc),
	.w8(32'hb8f9cc81),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37638c68),
	.w1(32'h360d8538),
	.w2(32'hb80331fd),
	.w3(32'h377e2e7d),
	.w4(32'h3703e97e),
	.w5(32'hb7a6f601),
	.w6(32'h37deb885),
	.w7(32'h37aaf254),
	.w8(32'hb6b368d4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365bb355),
	.w1(32'h35c81e5f),
	.w2(32'h36050178),
	.w3(32'h362fb45d),
	.w4(32'h3552948f),
	.w5(32'h35a0c2ef),
	.w6(32'h35854afa),
	.w7(32'h354a33ea),
	.w8(32'h36105e8c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968be5f),
	.w1(32'hb8a3e8b3),
	.w2(32'hb9698b44),
	.w3(32'hb8dc2288),
	.w4(32'h38737937),
	.w5(32'hb8a8f6ea),
	.w6(32'hb8f6bbe8),
	.w7(32'h38382a40),
	.w8(32'hb8dc7a77),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f87ffb),
	.w1(32'hb9f22989),
	.w2(32'hba15c098),
	.w3(32'hb9a456ed),
	.w4(32'hb99144c6),
	.w5(32'hb9d7bc1f),
	.w6(32'hb9b2b70e),
	.w7(32'hb99f3c91),
	.w8(32'hb9ff28a0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cc87e),
	.w1(32'hb92e4794),
	.w2(32'hb985d36b),
	.w3(32'hb9264010),
	.w4(32'hb8910701),
	.w5(32'hb93a6b3a),
	.w6(32'hb9171bfe),
	.w7(32'hb8b89043),
	.w8(32'hb950b8a2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37521749),
	.w1(32'h35c76947),
	.w2(32'h378bc671),
	.w3(32'h35e6b475),
	.w4(32'hb6fdbb26),
	.w5(32'hb6dab87c),
	.w6(32'h376ec575),
	.w7(32'hb6fd4553),
	.w8(32'h370164d6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36964846),
	.w1(32'h3510368a),
	.w2(32'h37104fde),
	.w3(32'hb5de5034),
	.w4(32'hb681f183),
	.w5(32'h361682de),
	.w6(32'hb6914cf1),
	.w7(32'hb6640a0c),
	.w8(32'h365d075f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77384cd),
	.w1(32'h35d3b831),
	.w2(32'h3595cdc3),
	.w3(32'hb766060a),
	.w4(32'hb6e334c3),
	.w5(32'h36bc294d),
	.w6(32'hb6e7935e),
	.w7(32'hb60611dc),
	.w8(32'h36cc0a35),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797165f),
	.w1(32'h36191cf2),
	.w2(32'hb7868c36),
	.w3(32'h37e1b12b),
	.w4(32'h37e97a6a),
	.w5(32'h379ea1c0),
	.w6(32'h37b4cb6a),
	.w7(32'h37d1275b),
	.w8(32'h36d134d7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2160e),
	.w1(32'hb8d1850a),
	.w2(32'hb906fbfe),
	.w3(32'hb8b7630d),
	.w4(32'hb87eea96),
	.w5(32'hb886a94e),
	.w6(32'hb9068cd5),
	.w7(32'hb89b1c9c),
	.w8(32'hb8acbb81),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362a9869),
	.w1(32'hb717a0d9),
	.w2(32'hb716e40f),
	.w3(32'h37419147),
	.w4(32'hb77c17fc),
	.w5(32'hb72497b7),
	.w6(32'h35fdaa9f),
	.w7(32'hb7fbc0b8),
	.w8(32'hb7a693a8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884eb93),
	.w1(32'hb695f0b2),
	.w2(32'hb889de2a),
	.w3(32'h361d219f),
	.w4(32'h387ad017),
	.w5(32'hb70f66fb),
	.w6(32'h3659f420),
	.w7(32'h38810356),
	.w8(32'hb710d22e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900f2bb),
	.w1(32'hb85059d3),
	.w2(32'hb8dc5228),
	.w3(32'hb88a2ed5),
	.w4(32'hb506e07b),
	.w5(32'hb8897929),
	.w6(32'hb8892c9d),
	.w7(32'hb7a14412),
	.w8(32'hb8a8d072),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360ee0e1),
	.w1(32'h36810dc3),
	.w2(32'h3684fa95),
	.w3(32'h338c4477),
	.w4(32'h364e74dc),
	.w5(32'h36707378),
	.w6(32'h36470456),
	.w7(32'h3633fcc3),
	.w8(32'h363e2e22),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3671d6d8),
	.w1(32'h3670f73b),
	.w2(32'h36b5111c),
	.w3(32'h35c54fd7),
	.w4(32'h3619c72e),
	.w5(32'h36543a28),
	.w6(32'h363beab2),
	.w7(32'h35f45657),
	.w8(32'h3671614e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3672fbfd),
	.w1(32'h35ab4e78),
	.w2(32'hb65a78eb),
	.w3(32'h36a043b5),
	.w4(32'h3626763e),
	.w5(32'h34bd32f1),
	.w6(32'h372d4d7f),
	.w7(32'h35e4212f),
	.w8(32'h355c2835),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35db9b9d),
	.w1(32'h36677445),
	.w2(32'h36cd82c9),
	.w3(32'hb59cea29),
	.w4(32'hb5759c57),
	.w5(32'h3683177c),
	.w6(32'hb59477d7),
	.w7(32'hb6187031),
	.w8(32'h35d1137f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72761c6),
	.w1(32'hb6d25924),
	.w2(32'hb7c1ddfe),
	.w3(32'h35ec22e6),
	.w4(32'h369b2ed5),
	.w5(32'hb7225b8a),
	.w6(32'h370d9f9a),
	.w7(32'h36e150d7),
	.w8(32'hb71c9d24),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cb19c),
	.w1(32'hb985060d),
	.w2(32'hb9a06c31),
	.w3(32'hb92539c2),
	.w4(32'hb92e7846),
	.w5(32'hb9708fc7),
	.w6(32'hb9644b3f),
	.w7(32'hb957adc8),
	.w8(32'hb99a71e6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a8885),
	.w1(32'hb94d80ab),
	.w2(32'hb9599fe4),
	.w3(32'hb9188d44),
	.w4(32'hb90e9498),
	.w5(32'hb9248a6f),
	.w6(32'hb90a8971),
	.w7(32'hb8ff39ff),
	.w8(32'hb9391044),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366e1ce0),
	.w1(32'hb5183bff),
	.w2(32'h368a75f0),
	.w3(32'h355a539e),
	.w4(32'hb5ca7d55),
	.w5(32'h35c7f7c6),
	.w6(32'h35054f08),
	.w7(32'h359f9415),
	.w8(32'h3693dfac),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ec1b5),
	.w1(32'hb90d5202),
	.w2(32'hb9731fd0),
	.w3(32'hb8d324b9),
	.w4(32'hb8c2d79e),
	.w5(32'hb929342a),
	.w6(32'hb8d06d8c),
	.w7(32'hb901b88e),
	.w8(32'hb944a79e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf8443),
	.w1(32'hb8c40a11),
	.w2(32'hb8d01117),
	.w3(32'hb89e8c7c),
	.w4(32'hb84ce377),
	.w5(32'hb89a4c8a),
	.w6(32'hb8a25c4a),
	.w7(32'hb8700ba2),
	.w8(32'hb89cf6e2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8762877),
	.w1(32'hb8ac359c),
	.w2(32'hb8f04691),
	.w3(32'hb880d54c),
	.w4(32'hb8ee3f4a),
	.w5(32'hb915e2f0),
	.w6(32'hb869afbd),
	.w7(32'hb8bd1a62),
	.w8(32'hb8f06592),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899c6a1),
	.w1(32'hb88c3903),
	.w2(32'hb8c1787b),
	.w3(32'hb8306a68),
	.w4(32'hb821408a),
	.w5(32'hb8793c70),
	.w6(32'hb83d3710),
	.w7(32'hb81aa827),
	.w8(32'hb8710399),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370ded39),
	.w1(32'h37b62eaa),
	.w2(32'h37249f01),
	.w3(32'h37fbff4c),
	.w4(32'h383c8443),
	.w5(32'h37b04aa8),
	.w6(32'h379ec324),
	.w7(32'h378f43f9),
	.w8(32'h367060bd),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb702bbbd),
	.w1(32'h3757904c),
	.w2(32'hb687b807),
	.w3(32'hb7f7850b),
	.w4(32'hb6b04285),
	.w5(32'hb78403f2),
	.w6(32'hb8274a14),
	.w7(32'hb7a91b7e),
	.w8(32'hb7bf6176),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3619b2c6),
	.w1(32'h35c572cf),
	.w2(32'h3602074c),
	.w3(32'h34f21725),
	.w4(32'hb5d525a8),
	.w5(32'h355e75f4),
	.w6(32'h3577a7a3),
	.w7(32'hb6e93e82),
	.w8(32'hb5efd341),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37437806),
	.w1(32'h37a52fe9),
	.w2(32'h372a642b),
	.w3(32'h372a6062),
	.w4(32'h378ab99a),
	.w5(32'h36ff5ac5),
	.w6(32'h36b1bf5c),
	.w7(32'h37201bb6),
	.w8(32'hb632af81),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df6eb4),
	.w1(32'hb78788c3),
	.w2(32'hb71d717f),
	.w3(32'hb876255c),
	.w4(32'h388d7b8d),
	.w5(32'h383f1f68),
	.w6(32'hb903ab39),
	.w7(32'h376c04a3),
	.w8(32'h371683c7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4a5ec),
	.w1(32'hb9c6101c),
	.w2(32'hb9c832c0),
	.w3(32'hb9a18326),
	.w4(32'hb99d3e99),
	.w5(32'hb9b23eb8),
	.w6(32'hb99b5288),
	.w7(32'hb99ccc02),
	.w8(32'hb9c92247),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966e97a),
	.w1(32'hb98897a6),
	.w2(32'hb9876ba0),
	.w3(32'hb95c0f5c),
	.w4(32'hb97312c8),
	.w5(32'hb981bb88),
	.w6(32'hb95ffccb),
	.w7(32'hb97db1af),
	.w8(32'hb98cef68),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967ca5f),
	.w1(32'hb99e56f2),
	.w2(32'hb99a993e),
	.w3(32'hb9609ca9),
	.w4(32'hb987e148),
	.w5(32'hb9886deb),
	.w6(32'hb9505a01),
	.w7(32'hb985f548),
	.w8(32'hb9921103),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5963397),
	.w1(32'h36ee4826),
	.w2(32'hb68a0feb),
	.w3(32'h36930ab2),
	.w4(32'h3745740b),
	.w5(32'hb547ff8c),
	.w6(32'h36a78c86),
	.w7(32'h372855b5),
	.w8(32'hb5f7d3f7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3617dfb3),
	.w1(32'h3507e2f9),
	.w2(32'h35900307),
	.w3(32'h350f8e8a),
	.w4(32'hb4272bdc),
	.w5(32'h363522f6),
	.w6(32'h35c6b7d0),
	.w7(32'h34d9e978),
	.w8(32'h35d31fdb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b3e728),
	.w1(32'hb42563dc),
	.w2(32'h339ef73a),
	.w3(32'h36b6fdd7),
	.w4(32'hb71393ca),
	.w5(32'hb6ac5b3a),
	.w6(32'h361e3b37),
	.w7(32'hb6104203),
	.w8(32'h3488322a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3626ab2c),
	.w1(32'h36a07444),
	.w2(32'h3681f693),
	.w3(32'h35920248),
	.w4(32'h35e9e537),
	.w5(32'h362b7f67),
	.w6(32'h36b94d36),
	.w7(32'h36a3a6cd),
	.w8(32'h3646465d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd9c8f),
	.w1(32'hb515d133),
	.w2(32'hb8421e4f),
	.w3(32'hb8c482bb),
	.w4(32'h387016ac),
	.w5(32'hb7305f09),
	.w6(32'hb8cb52bb),
	.w7(32'h38034540),
	.w8(32'hb74b01cb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368cb8a2),
	.w1(32'h3722b8b7),
	.w2(32'hb77e1af8),
	.w3(32'hb643638f),
	.w4(32'hb7f60add),
	.w5(32'hb83186bd),
	.w6(32'h37a39b27),
	.w7(32'h356a979d),
	.w8(32'hb8044b5c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c579d7),
	.w1(32'h3825a45d),
	.w2(32'h3752bac5),
	.w3(32'h3828b74f),
	.w4(32'h384f7de3),
	.w5(32'h37c915b9),
	.w6(32'h3858d914),
	.w7(32'h3839a6ed),
	.w8(32'h37698f93),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3742fdb7),
	.w1(32'h37895035),
	.w2(32'h3753e5d5),
	.w3(32'h37ae381e),
	.w4(32'h37ba8c4a),
	.w5(32'h37906adb),
	.w6(32'h386fa7db),
	.w7(32'h3871e42e),
	.w8(32'h381682b6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7867bdf),
	.w1(32'hb7a4b99e),
	.w2(32'hb7cb2969),
	.w3(32'h3719bacc),
	.w4(32'hb729b202),
	.w5(32'hb7e53b68),
	.w6(32'h37b34b24),
	.w7(32'h33248778),
	.w8(32'hb791b7fc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78f5767),
	.w1(32'hb71fe504),
	.w2(32'hb6b5476c),
	.w3(32'hb76c512e),
	.w4(32'hb74848d9),
	.w5(32'hb6dcb0e0),
	.w6(32'hb7a52e9b),
	.w7(32'hb77afdb0),
	.w8(32'hb6fa2e85),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34c69d0a),
	.w1(32'h35942798),
	.w2(32'hb56acf29),
	.w3(32'h33615491),
	.w4(32'hb235409b),
	.w5(32'hb5f453a6),
	.w6(32'h361e3f8d),
	.w7(32'hb5ac30d0),
	.w8(32'hb5e5333c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9343c80),
	.w1(32'hb94fa067),
	.w2(32'hb9346ac5),
	.w3(32'hb92410eb),
	.w4(32'hb920722e),
	.w5(32'hb9308dad),
	.w6(32'hb8f751f0),
	.w7(32'hb90a80c7),
	.w8(32'hb9243d1b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70eeaa3),
	.w1(32'hb7248e10),
	.w2(32'hb7d54321),
	.w3(32'hb78f1cb7),
	.w4(32'hb7237914),
	.w5(32'hb802e8c4),
	.w6(32'hb77ec5e7),
	.w7(32'hb7baaa18),
	.w8(32'hb80c2695),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca6428),
	.w1(32'hb9239996),
	.w2(32'hb8a8570d),
	.w3(32'hb97c62e1),
	.w4(32'hb922d2fc),
	.w5(32'hb8adb7f0),
	.w6(32'hb9a40de6),
	.w7(32'hb931cbd7),
	.w8(32'hb8eb4cc2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule