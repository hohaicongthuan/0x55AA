module layer_8_featuremap_194(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c749a58),
	.w1(32'h3acdb9d6),
	.w2(32'h3a858959),
	.w3(32'hbc12098e),
	.w4(32'h3b7e7492),
	.w5(32'hbb167062),
	.w6(32'h3bba318b),
	.w7(32'h3c25ea7d),
	.w8(32'hbafcf9f7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc261cc1),
	.w1(32'hbc6d0a2b),
	.w2(32'h3b343b81),
	.w3(32'hbbb76f6f),
	.w4(32'h3d4f8427),
	.w5(32'h3e0cd5e4),
	.w6(32'hbd80d60d),
	.w7(32'hbddc1bd6),
	.w8(32'hbda59946),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba7d62),
	.w1(32'hbc334e9f),
	.w2(32'hbba12086),
	.w3(32'h3d872580),
	.w4(32'hbc69a7fd),
	.w5(32'hbc23795e),
	.w6(32'hbacffeb1),
	.w7(32'hbbbce4c8),
	.w8(32'hba4917b4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb661da),
	.w1(32'hbc1f4dae),
	.w2(32'hbb5f1aeb),
	.w3(32'hbb85937d),
	.w4(32'hbba5c0d4),
	.w5(32'hbc09dbdb),
	.w6(32'hbb36e16a),
	.w7(32'hbaf5780e),
	.w8(32'hbb0108e3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5998ba),
	.w1(32'hbc52c45c),
	.w2(32'h3b9e070a),
	.w3(32'h3bb76962),
	.w4(32'h3d4a4940),
	.w5(32'h3e122c78),
	.w6(32'hbd6e6bea),
	.w7(32'hbddc37b2),
	.w8(32'hbda2c8ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8115bf),
	.w1(32'hbb631271),
	.w2(32'hbb489ae3),
	.w3(32'h3d8e47cd),
	.w4(32'hbb3b961e),
	.w5(32'h398fec89),
	.w6(32'h3a228f75),
	.w7(32'hbaf1825f),
	.w8(32'h3b840814),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfce819),
	.w1(32'hbab73eac),
	.w2(32'hbbbfc87b),
	.w3(32'h3be2c298),
	.w4(32'hbcf9d7be),
	.w5(32'hbd972307),
	.w6(32'h3d03f1b8),
	.w7(32'h3d6b2c21),
	.w8(32'h3d294748),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5f5ec),
	.w1(32'hbc0beba0),
	.w2(32'hbb2252d5),
	.w3(32'hbd42718f),
	.w4(32'h3903f32c),
	.w5(32'h3971ae05),
	.w6(32'h3b99e1bf),
	.w7(32'h3bc8a9fa),
	.w8(32'hba1a578c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f717),
	.w1(32'hbcc432c4),
	.w2(32'hbbf26ce1),
	.w3(32'hbbf0a026),
	.w4(32'h3cc69286),
	.w5(32'h3dd5b299),
	.w6(32'hbd0bb1b0),
	.w7(32'hbd8f8c7a),
	.w8(32'hbd462611),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd08bc0d),
	.w1(32'hbbf8b5ac),
	.w2(32'hbc0c6a12),
	.w3(32'h3d0bd132),
	.w4(32'hbc830401),
	.w5(32'h3b195689),
	.w6(32'hbc58d02d),
	.w7(32'hbc39d34c),
	.w8(32'hbc0b2191),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd1612),
	.w1(32'hbb88a333),
	.w2(32'hbbc5f618),
	.w3(32'h3c40ffb8),
	.w4(32'h3b0a9a61),
	.w5(32'hb990ed84),
	.w6(32'h3c9c831d),
	.w7(32'h3cac7c12),
	.w8(32'h3c48e7f4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d0678),
	.w1(32'h39d5a7fa),
	.w2(32'h3b44ea6c),
	.w3(32'h3b33508d),
	.w4(32'h3c83403e),
	.w5(32'h3c5be9d3),
	.w6(32'hba5511ac),
	.w7(32'hbc0bbb5f),
	.w8(32'hbba35ac7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf601e),
	.w1(32'hbc835c1e),
	.w2(32'hbc8c27ae),
	.w3(32'h3c060ba8),
	.w4(32'hbad82956),
	.w5(32'h3b7e569f),
	.w6(32'hbc9b45ad),
	.w7(32'hbca614c3),
	.w8(32'hbc1f0b0e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bba5c),
	.w1(32'h3a90181a),
	.w2(32'h3b052e5d),
	.w3(32'hbb88674a),
	.w4(32'h3a815f67),
	.w5(32'hbae8d9f1),
	.w6(32'h3c2c4c2f),
	.w7(32'h3bf65572),
	.w8(32'h3c02c869),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc65aa),
	.w1(32'h3b78bf3c),
	.w2(32'hbc49aeb3),
	.w3(32'hbb9e941e),
	.w4(32'hbd5e6fb6),
	.w5(32'hbe0345b2),
	.w6(32'h3d82dba0),
	.w7(32'h3dd8c0e0),
	.w8(32'h3da26ce0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f56e6),
	.w1(32'h3b02a4f7),
	.w2(32'h3baa7007),
	.w3(32'hbd860a8d),
	.w4(32'h3af5120f),
	.w5(32'h39beb8ca),
	.w6(32'h3b3e9b33),
	.w7(32'h3a52860e),
	.w8(32'h3c1703c2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb4124),
	.w1(32'hbb038485),
	.w2(32'hbaeb0db2),
	.w3(32'hbb72f7ec),
	.w4(32'hbb2ace37),
	.w5(32'hbb90de59),
	.w6(32'hbbd758c3),
	.w7(32'hbbbadb67),
	.w8(32'hbaf36294),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb660b08),
	.w1(32'h3b46418b),
	.w2(32'h388c6df3),
	.w3(32'hbc02ae5c),
	.w4(32'h3b89d101),
	.w5(32'h3bb29771),
	.w6(32'h3b71717d),
	.w7(32'h3a40795a),
	.w8(32'h3a760f4d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b924d8d),
	.w1(32'h3b641431),
	.w2(32'hb8ac8ec9),
	.w3(32'h3b8bb09b),
	.w4(32'h3c067239),
	.w5(32'h3c3b01fd),
	.w6(32'h3c958f46),
	.w7(32'h3c88c6ca),
	.w8(32'h3bbaf00e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5be1),
	.w1(32'h3aa36f9d),
	.w2(32'hbc0663aa),
	.w3(32'h3c1af812),
	.w4(32'hbd765639),
	.w5(32'hbe18bb6a),
	.w6(32'h3daefc3c),
	.w7(32'h3e08ab9d),
	.w8(32'h3dd9d55f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cb54b),
	.w1(32'h3b9a7237),
	.w2(32'h3ba91eb4),
	.w3(32'hbda7b99b),
	.w4(32'h3b90050d),
	.w5(32'h3b5abe73),
	.w6(32'h3c12e671),
	.w7(32'h3ba50970),
	.w8(32'h3bd90628),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f1132),
	.w1(32'hbbe89ab6),
	.w2(32'hbc122e93),
	.w3(32'hbb836d65),
	.w4(32'hbc344631),
	.w5(32'hbbd0e79a),
	.w6(32'hbc27a4ec),
	.w7(32'hbbf853db),
	.w8(32'h3a9f6a94),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b810f),
	.w1(32'hbaef2d1c),
	.w2(32'hba931200),
	.w3(32'h3c021324),
	.w4(32'h3bbd69ed),
	.w5(32'hba9b77df),
	.w6(32'h3c8e957c),
	.w7(32'h3c5e8148),
	.w8(32'h3bc3293f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942fd8a),
	.w1(32'hbbd9f5c9),
	.w2(32'hba7428dc),
	.w3(32'h3b7a1a77),
	.w4(32'h3a894c9d),
	.w5(32'hbb1d94b7),
	.w6(32'h3c07da6a),
	.w7(32'h3ab7db08),
	.w8(32'h3b483494),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91039a),
	.w1(32'hbc685e9d),
	.w2(32'hbce8071a),
	.w3(32'hbaaaae98),
	.w4(32'h3b0871c4),
	.w5(32'hbb4ca429),
	.w6(32'hbbb1fb7b),
	.w7(32'h3a4e397e),
	.w8(32'h3bafc986),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab73ed3),
	.w1(32'h3aac8379),
	.w2(32'hbc93aa4d),
	.w3(32'h3c7cc9fa),
	.w4(32'h3b8d2402),
	.w5(32'h3bc09a05),
	.w6(32'h3b7410ee),
	.w7(32'h3b0a73c6),
	.w8(32'h3bb946c2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d71e3),
	.w1(32'hbbcc648b),
	.w2(32'hbb0a29a4),
	.w3(32'hbbcf2a9b),
	.w4(32'hbb83a80c),
	.w5(32'hba93756e),
	.w6(32'hba8e339b),
	.w7(32'hbc1fd28f),
	.w8(32'hba9909df),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6fa1e),
	.w1(32'h3c25c977),
	.w2(32'hbbf5cf89),
	.w3(32'h3cc06d1d),
	.w4(32'h3cad4b37),
	.w5(32'h3b888462),
	.w6(32'h3d0209f5),
	.w7(32'h3cf0e7d4),
	.w8(32'h3c2c0f85),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567c59),
	.w1(32'hbad8546b),
	.w2(32'hbb38b2ba),
	.w3(32'hbb32dae7),
	.w4(32'h3ae5f188),
	.w5(32'h3c2e9e46),
	.w6(32'h3cb77a37),
	.w7(32'h3c3e0a8e),
	.w8(32'h3be7cb8d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3382bc),
	.w1(32'hbc2f04b8),
	.w2(32'hbbbe1aec),
	.w3(32'hbb242961),
	.w4(32'h3c4559ad),
	.w5(32'h3cbd6f31),
	.w6(32'hbabe4082),
	.w7(32'h3b4c126a),
	.w8(32'hbb83bf02),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc501064),
	.w1(32'hbc8f54f1),
	.w2(32'hbcf9d395),
	.w3(32'h3c6de8fd),
	.w4(32'hbc8481a3),
	.w5(32'hbc324065),
	.w6(32'hbb773e16),
	.w7(32'hbc1e1d50),
	.w8(32'hbb35a4a5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc946326),
	.w1(32'hbb4fcce0),
	.w2(32'hbb562586),
	.w3(32'hbbc9fac4),
	.w4(32'hbbd3162c),
	.w5(32'hbb8aefb0),
	.w6(32'h3c7e5e51),
	.w7(32'h3cc03d7d),
	.w8(32'h3caaf95e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba610da),
	.w1(32'hbb9cded3),
	.w2(32'hbbcc03a2),
	.w3(32'hbc02c14d),
	.w4(32'hbb016aeb),
	.w5(32'h3acebe38),
	.w6(32'hbabd7313),
	.w7(32'hbb2c4ee1),
	.w8(32'hba8a4a12),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f6261),
	.w1(32'hbba75e17),
	.w2(32'h3ae03ef7),
	.w3(32'h3bc3f12f),
	.w4(32'hbbccf7d8),
	.w5(32'h3b35d5c4),
	.w6(32'hbbba7b1d),
	.w7(32'hbb4369db),
	.w8(32'h3b03dc25),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdddb58),
	.w1(32'hbc2665d8),
	.w2(32'hbc79b9c4),
	.w3(32'h3bd5db64),
	.w4(32'h3beec14d),
	.w5(32'h3c4da87c),
	.w6(32'h3b3c46dd),
	.w7(32'h3bda7156),
	.w8(32'hb8d75773),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca47e63),
	.w1(32'hbb74dcc4),
	.w2(32'hbb9c24b4),
	.w3(32'h3c61db82),
	.w4(32'h3a81eda2),
	.w5(32'hbb3763ff),
	.w6(32'h3bef6334),
	.w7(32'h3bfd8b13),
	.w8(32'h3b49802a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ffad),
	.w1(32'hbbc0538c),
	.w2(32'hbc1d3643),
	.w3(32'hbbe4a8d2),
	.w4(32'h3b6d0a2f),
	.w5(32'hbb2660f0),
	.w6(32'hbb7ad474),
	.w7(32'hbba8e2b1),
	.w8(32'h3b5d715e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc676730),
	.w1(32'hbbc74284),
	.w2(32'h39e19cc9),
	.w3(32'hbc039078),
	.w4(32'hbba535c3),
	.w5(32'h3c4f5161),
	.w6(32'h3b6a12ae),
	.w7(32'h3b54759d),
	.w8(32'h3b52a56b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4842f),
	.w1(32'hbb5dfb5f),
	.w2(32'h3b463cb9),
	.w3(32'h3be016d2),
	.w4(32'hb9f79069),
	.w5(32'h3bdb4457),
	.w6(32'h3b87b35d),
	.w7(32'h3c6535fb),
	.w8(32'h3c03ec0a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef9e29),
	.w1(32'h3ab01780),
	.w2(32'hb8ad4670),
	.w3(32'hbbac768b),
	.w4(32'h3b258d07),
	.w5(32'hbb126883),
	.w6(32'hbb11ba8b),
	.w7(32'hbb6b9225),
	.w8(32'hba97dfee),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab65052),
	.w1(32'h3be928e3),
	.w2(32'h3b83cf53),
	.w3(32'h3b5448ce),
	.w4(32'h3bfc7a90),
	.w5(32'h3b9c718f),
	.w6(32'h3c059e5a),
	.w7(32'hb9b52332),
	.w8(32'h3c0944f3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6c0d),
	.w1(32'hbc0dd8e0),
	.w2(32'hbb325704),
	.w3(32'h3b87c4d3),
	.w4(32'hba32f639),
	.w5(32'h3bd5cb8f),
	.w6(32'hbb185fe9),
	.w7(32'hbb9e9087),
	.w8(32'h3c1468c0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339765),
	.w1(32'hbbc672ab),
	.w2(32'hbbcc9243),
	.w3(32'h3b38ff3d),
	.w4(32'hbb02ba8e),
	.w5(32'h3b560375),
	.w6(32'hbb90a209),
	.w7(32'hbb9625d3),
	.w8(32'hbb142a98),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9429),
	.w1(32'hbafec788),
	.w2(32'h3b7c2702),
	.w3(32'h3b7d81d2),
	.w4(32'h3b26a3d4),
	.w5(32'h3c276d77),
	.w6(32'h3b9420c2),
	.w7(32'h3bfa4465),
	.w8(32'h3bdaf938),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48d6c5),
	.w1(32'hbacaf3de),
	.w2(32'h3970adbb),
	.w3(32'h3be31a35),
	.w4(32'h3abab69c),
	.w5(32'h3c4e2f3c),
	.w6(32'h3c473128),
	.w7(32'h3c9ac514),
	.w8(32'h3c567dd0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23e024),
	.w1(32'hbaad60f2),
	.w2(32'hbc9f34b3),
	.w3(32'h3c0f59eb),
	.w4(32'hbd2b79d9),
	.w5(32'hbddc6f88),
	.w6(32'h3d0cad32),
	.w7(32'h3d8171c5),
	.w8(32'h3d4c6c30),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f7bd1),
	.w1(32'h390661e5),
	.w2(32'h3b9a892b),
	.w3(32'hbd769186),
	.w4(32'h3b21312a),
	.w5(32'h3ba23e34),
	.w6(32'h39367435),
	.w7(32'h3be8683c),
	.w8(32'h3c054a23),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b470282),
	.w1(32'h3bb426e5),
	.w2(32'h3bae2167),
	.w3(32'h3c1ee543),
	.w4(32'h3bc22d62),
	.w5(32'h3b8514e8),
	.w6(32'h3c6415e0),
	.w7(32'h3c5cfb31),
	.w8(32'h3c9d553c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f126a),
	.w1(32'hb8b49973),
	.w2(32'hbb53d910),
	.w3(32'hbbc465ed),
	.w4(32'hbb82c2c9),
	.w5(32'hbb1588d4),
	.w6(32'hbb17b2be),
	.w7(32'h3b97b0cb),
	.w8(32'h3b70c965),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72b6a0),
	.w1(32'hb795ba9b),
	.w2(32'hbaf1b5d1),
	.w3(32'hbb523d4d),
	.w4(32'h3c6e417a),
	.w5(32'h3a491859),
	.w6(32'h3bdffc30),
	.w7(32'h3b76fc05),
	.w8(32'h3aa83435),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc912bf2),
	.w1(32'hbb882d9c),
	.w2(32'hbc6fad6c),
	.w3(32'hbc932946),
	.w4(32'hbaafccb7),
	.w5(32'hbbbec91a),
	.w6(32'hbc1a53f7),
	.w7(32'hbc5010f1),
	.w8(32'h3b4879b4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ddf19),
	.w1(32'h3be64aac),
	.w2(32'hba19e5cc),
	.w3(32'h3c4662b2),
	.w4(32'h3a8ec666),
	.w5(32'h3b5f0469),
	.w6(32'h3ccabe7f),
	.w7(32'h3c0c2f90),
	.w8(32'h3c6407f5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a18d0),
	.w1(32'hbbfca0d3),
	.w2(32'hbb9ff81d),
	.w3(32'h3c93343d),
	.w4(32'h3cd8f304),
	.w5(32'h3d97fe59),
	.w6(32'hbc2cf185),
	.w7(32'hbd2a999b),
	.w8(32'hbcf0a261),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfc8d8),
	.w1(32'hbb79299a),
	.w2(32'h3b4a53cd),
	.w3(32'h3ce80a52),
	.w4(32'hb9ea1ac6),
	.w5(32'h3bcb3000),
	.w6(32'h3c1e20dc),
	.w7(32'h3b58c973),
	.w8(32'h3a93bfad),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d947a),
	.w1(32'h3b93aa28),
	.w2(32'h3a475ff6),
	.w3(32'h3b5a292f),
	.w4(32'hbb5c7a38),
	.w5(32'h3c3b9f71),
	.w6(32'h3bbfc499),
	.w7(32'h3b7dcf6b),
	.w8(32'h3b6c2076),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdfc86),
	.w1(32'h39a70fdb),
	.w2(32'hbba4c59d),
	.w3(32'h3aa39a48),
	.w4(32'hbaf49548),
	.w5(32'hba6b53c6),
	.w6(32'h3c665dac),
	.w7(32'h3b892af3),
	.w8(32'hbb3efc48),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e9ba0),
	.w1(32'hbc69d96e),
	.w2(32'hb9f70483),
	.w3(32'hbba28712),
	.w4(32'hbac0919f),
	.w5(32'hb98eb0eb),
	.w6(32'hbb897569),
	.w7(32'hbb043021),
	.w8(32'hbb7a86a8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158a16),
	.w1(32'hbaff99c5),
	.w2(32'hbbcd5e1d),
	.w3(32'h3aec3c70),
	.w4(32'hbb172eef),
	.w5(32'hbba47305),
	.w6(32'h37838cd6),
	.w7(32'hbbe91ff7),
	.w8(32'hbc1668e5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22336),
	.w1(32'hbb8fa507),
	.w2(32'hbb0be478),
	.w3(32'hbbd493f9),
	.w4(32'hb732fc42),
	.w5(32'hbb93de4c),
	.w6(32'h39cedecf),
	.w7(32'hba8cd69d),
	.w8(32'h3acb3493),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cebb5d),
	.w1(32'hba918d29),
	.w2(32'hbb94db94),
	.w3(32'hbb42b16f),
	.w4(32'h3a284457),
	.w5(32'hbb8f5e87),
	.w6(32'h3994f84f),
	.w7(32'h3bc96160),
	.w8(32'hba8b839e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb669a4a),
	.w1(32'hbb8950f5),
	.w2(32'hbbfcd372),
	.w3(32'hb9c84561),
	.w4(32'hbb08029e),
	.w5(32'hbb452d5f),
	.w6(32'h3ba41517),
	.w7(32'h3b1a8996),
	.w8(32'h3bf74f63),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a5460),
	.w1(32'hbd1e8d7f),
	.w2(32'hbd5f9077),
	.w3(32'hba977394),
	.w4(32'hbc427f35),
	.w5(32'hbce98953),
	.w6(32'hbb6d046a),
	.w7(32'hbb48c895),
	.w8(32'hbb8ca871),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd30dde8),
	.w1(32'hb942676a),
	.w2(32'h3c6c9d3c),
	.w3(32'hbc947e3d),
	.w4(32'h3b2de8a8),
	.w5(32'hba164367),
	.w6(32'h3cf4f037),
	.w7(32'h3d416033),
	.w8(32'h3d1db476),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babe5dd),
	.w1(32'h3994e95d),
	.w2(32'hb97a5559),
	.w3(32'hbbddc6b2),
	.w4(32'h39d9997c),
	.w5(32'h3b5f2c2d),
	.w6(32'hbb6925db),
	.w7(32'hbc27bd9f),
	.w8(32'hbbe2289d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7896c0),
	.w1(32'hbacd56e4),
	.w2(32'hbbfd9064),
	.w3(32'h3c03c318),
	.w4(32'hbb443b59),
	.w5(32'hbca7ad5a),
	.w6(32'h3c09f437),
	.w7(32'h3c4b7e15),
	.w8(32'h3c0fc4ad),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc9ef),
	.w1(32'hb9f95733),
	.w2(32'hbabc3f68),
	.w3(32'hbc40ac93),
	.w4(32'hbb55d0b3),
	.w5(32'hbc4653a7),
	.w6(32'h3b00b301),
	.w7(32'h3b227a0c),
	.w8(32'h3a2e5e84),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92184e),
	.w1(32'hb895a2ee),
	.w2(32'h3bbdf765),
	.w3(32'hbbe27713),
	.w4(32'hba6e901a),
	.w5(32'h3b803e50),
	.w6(32'hba7f93ee),
	.w7(32'hbad48474),
	.w8(32'h3b8a032e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91cf08),
	.w1(32'h3bb38180),
	.w2(32'h3ad8ac01),
	.w3(32'h3b738288),
	.w4(32'h3c1a5c7a),
	.w5(32'h3a7b574f),
	.w6(32'h3c254321),
	.w7(32'h3b930411),
	.w8(32'hb8e2f391),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4007ce),
	.w1(32'hbbbbaf77),
	.w2(32'h3ba8ea1f),
	.w3(32'hba58ae5b),
	.w4(32'h3923fc32),
	.w5(32'h3b83f230),
	.w6(32'h3b8e5315),
	.w7(32'h3b99749e),
	.w8(32'h3bde6cba),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77e0cf),
	.w1(32'h3b712c11),
	.w2(32'hbb7e3df7),
	.w3(32'h3bb89b2b),
	.w4(32'h3b2fca9e),
	.w5(32'h3a8322b5),
	.w6(32'h3c9b5c91),
	.w7(32'h3c40f9da),
	.w8(32'h3b8ea9bc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d465f),
	.w1(32'h3b7d1d1d),
	.w2(32'h3c110066),
	.w3(32'hbbaccca2),
	.w4(32'hbc644607),
	.w5(32'h3b02378e),
	.w6(32'h3cc2e19c),
	.w7(32'h3cbc04f4),
	.w8(32'h3b9e2bd4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09dffe),
	.w1(32'hbb872e23),
	.w2(32'hbaaa5aa4),
	.w3(32'h3c3be8db),
	.w4(32'hbb89f6ca),
	.w5(32'hbb95ab6e),
	.w6(32'h3c028ad2),
	.w7(32'h3bf10a3c),
	.w8(32'h3aec879a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc083959),
	.w1(32'hbb501e57),
	.w2(32'hbb0307df),
	.w3(32'hbc182302),
	.w4(32'hbaa25b52),
	.w5(32'hbabe7e2a),
	.w6(32'h397a73d1),
	.w7(32'h3b11dde3),
	.w8(32'h39f14f72),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb40bc),
	.w1(32'h3ad6d585),
	.w2(32'h3b01922b),
	.w3(32'hbc8ecf88),
	.w4(32'h3ac5495d),
	.w5(32'h3b25901a),
	.w6(32'h3b82a1a8),
	.w7(32'h3c08f844),
	.w8(32'hbba3566e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea8c8),
	.w1(32'hbc2ea634),
	.w2(32'hbcfa2b8b),
	.w3(32'h3bc7f3dd),
	.w4(32'hbc6773a4),
	.w5(32'hbc4fddc0),
	.w6(32'h3b11980f),
	.w7(32'hbc392f06),
	.w8(32'hbbe8afe9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7009a9),
	.w1(32'h3b44813b),
	.w2(32'hbb8d58f3),
	.w3(32'h3c1cb0f3),
	.w4(32'h39ffb9ed),
	.w5(32'hbafb28ef),
	.w6(32'h3c06d4d6),
	.w7(32'h3c14a8fd),
	.w8(32'h3a84a84a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36b63),
	.w1(32'h3b84dc14),
	.w2(32'hbc08104c),
	.w3(32'hbb805a14),
	.w4(32'hba3c6bbd),
	.w5(32'h3b07027d),
	.w6(32'h39f7dcc5),
	.w7(32'hbbb95c8c),
	.w8(32'hbc2b50fc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61bdc7),
	.w1(32'h3b3a0fb1),
	.w2(32'h39e32b0d),
	.w3(32'h3bac0506),
	.w4(32'h3c5978dd),
	.w5(32'h3c1f417c),
	.w6(32'h3b8b28f5),
	.w7(32'h3bcecf32),
	.w8(32'h3c076d5a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac810b9),
	.w1(32'h3bf737c5),
	.w2(32'h3b94b986),
	.w3(32'hbb88cad2),
	.w4(32'h3b93d6f3),
	.w5(32'h3c5661d2),
	.w6(32'h3c31e5c6),
	.w7(32'h3bebb6cd),
	.w8(32'h3c0757e8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6af6a),
	.w1(32'hb9f7af9d),
	.w2(32'hbb904feb),
	.w3(32'h3c1b00af),
	.w4(32'h3a9cdcfb),
	.w5(32'hbc02cdf2),
	.w6(32'h3b055aea),
	.w7(32'h3bd18c0d),
	.w8(32'h3bf74504),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f268),
	.w1(32'hbc09cd97),
	.w2(32'hbc5ce661),
	.w3(32'hbaa6fb6c),
	.w4(32'hba25a17c),
	.w5(32'hbbcf212c),
	.w6(32'h3b20b7b4),
	.w7(32'hbba5099f),
	.w8(32'hba928260),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14b483),
	.w1(32'h39b8421d),
	.w2(32'h3b5b5dca),
	.w3(32'hbbe3b796),
	.w4(32'hbb92cd4e),
	.w5(32'h39275709),
	.w6(32'h3c2d12aa),
	.w7(32'h3c653e94),
	.w8(32'h3c2080b5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8a164),
	.w1(32'hbbdf7f91),
	.w2(32'hb7d59e46),
	.w3(32'h3c0636e4),
	.w4(32'hbab9ade5),
	.w5(32'h3be5e594),
	.w6(32'h3c8978e1),
	.w7(32'h3c7583f4),
	.w8(32'h3bfda762),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c622),
	.w1(32'h3c08949d),
	.w2(32'hbb8895ba),
	.w3(32'h3bf8dd36),
	.w4(32'h3ba7b28a),
	.w5(32'h39ef2f61),
	.w6(32'h3c068004),
	.w7(32'h3bd40598),
	.w8(32'hbaf69af9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c136039),
	.w1(32'hb9c7d8d8),
	.w2(32'hbba8940e),
	.w3(32'h3c255e88),
	.w4(32'h3bfdaf01),
	.w5(32'h3bdfba8d),
	.w6(32'h3c7e4ddb),
	.w7(32'h3c9f39fb),
	.w8(32'h3c533583),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c9812),
	.w1(32'h3c5fcb89),
	.w2(32'h3b57f1e5),
	.w3(32'h3bd55e70),
	.w4(32'h3c5c7705),
	.w5(32'h3c22aed7),
	.w6(32'h3cc146c6),
	.w7(32'h3c2a7a18),
	.w8(32'h3c613038),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d699),
	.w1(32'h3c5ae622),
	.w2(32'h3c9e6469),
	.w3(32'hb982f5ce),
	.w4(32'h3b5b187a),
	.w5(32'h3bf2b443),
	.w6(32'h3c0b1a2e),
	.w7(32'h3c0ae13a),
	.w8(32'h3c20b483),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a1a4b),
	.w1(32'h3b5d3d77),
	.w2(32'h3bbc24d0),
	.w3(32'h3c11a0a6),
	.w4(32'h3c699147),
	.w5(32'h3caa5478),
	.w6(32'h3bd64d92),
	.w7(32'h3c29721b),
	.w8(32'h3c82d5fd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001964),
	.w1(32'hb9f788f1),
	.w2(32'hbabe06a7),
	.w3(32'h3c92ada2),
	.w4(32'h3c2c7363),
	.w5(32'h3c573f89),
	.w6(32'h3bede5c4),
	.w7(32'h3c0a9014),
	.w8(32'h3bb75424),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffae6a),
	.w1(32'h3af22521),
	.w2(32'h3af0348a),
	.w3(32'h3c9ab114),
	.w4(32'hbbdd3e6e),
	.w5(32'h3bca3468),
	.w6(32'h3a6ea66a),
	.w7(32'h3ba84303),
	.w8(32'h3bfde41d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0b0b),
	.w1(32'h3996a638),
	.w2(32'hbaaad02a),
	.w3(32'h3ac4cdc4),
	.w4(32'hb94727b7),
	.w5(32'hbb7a89d5),
	.w6(32'h3b3e9deb),
	.w7(32'h3c0122c2),
	.w8(32'h3b510c80),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27aeb3),
	.w1(32'hbb42d649),
	.w2(32'h3b260236),
	.w3(32'hbbdd8fb4),
	.w4(32'h3a18e351),
	.w5(32'h3a845293),
	.w6(32'hbae6277d),
	.w7(32'h3b04b794),
	.w8(32'h3b49e054),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9a865),
	.w1(32'h3c0003aa),
	.w2(32'h3c077695),
	.w3(32'hbb69e775),
	.w4(32'h3c9ec0b9),
	.w5(32'h3d152697),
	.w6(32'hbc2e6d9a),
	.w7(32'hbcbf1298),
	.w8(32'hbc96b88b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7a3b2),
	.w1(32'hbb88468f),
	.w2(32'h3c02fbd5),
	.w3(32'h3ccab969),
	.w4(32'h3cf0a2a0),
	.w5(32'h3d8ef21d),
	.w6(32'hbcb3ef2b),
	.w7(32'hbd1ead21),
	.w8(32'hbce1cdf5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f49ca),
	.w1(32'h3bb2d41f),
	.w2(32'h3a1e8fff),
	.w3(32'h3d230596),
	.w4(32'h3b5ad0bd),
	.w5(32'h3bab79ee),
	.w6(32'h3b3837ef),
	.w7(32'h3ab153b0),
	.w8(32'hbb03f98d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07eadd),
	.w1(32'h3c9791a2),
	.w2(32'h3c3b47b9),
	.w3(32'h3b12e3e0),
	.w4(32'h3c3fe99e),
	.w5(32'h3bef9886),
	.w6(32'h3c7bd2f2),
	.w7(32'h3be85fe2),
	.w8(32'h3b41417b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6a2bd),
	.w1(32'h3baedde9),
	.w2(32'h3c399239),
	.w3(32'h3bf4f9c9),
	.w4(32'h3c601eb9),
	.w5(32'h3c93b4dc),
	.w6(32'h3ca71ec4),
	.w7(32'h3cb2b56c),
	.w8(32'h3cba6492),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2114),
	.w1(32'h3b0a9f82),
	.w2(32'hbb33d506),
	.w3(32'hba0e21c4),
	.w4(32'hbb8a24d8),
	.w5(32'h3b23d854),
	.w6(32'h3c201df6),
	.w7(32'h3c38f5ee),
	.w8(32'h3c428171),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfe93b),
	.w1(32'hba051512),
	.w2(32'h3b7a6901),
	.w3(32'hba5177c7),
	.w4(32'hba7f9aea),
	.w5(32'h3b809cde),
	.w6(32'h3bbefe75),
	.w7(32'h3c005eca),
	.w8(32'h3be38f0d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb521ebe),
	.w1(32'hbb32709c),
	.w2(32'hba73abfc),
	.w3(32'h3b82c964),
	.w4(32'hbb991ac9),
	.w5(32'hba3bd1a8),
	.w6(32'h3b251d4d),
	.w7(32'hbbe6bf5b),
	.w8(32'hba4f641d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f8ef),
	.w1(32'h3bbff412),
	.w2(32'hbb8a111a),
	.w3(32'h3b603240),
	.w4(32'h3be37233),
	.w5(32'h3b5472e2),
	.w6(32'h3b80f585),
	.w7(32'h3a856464),
	.w8(32'h3a84c468),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90f77),
	.w1(32'hba84c20a),
	.w2(32'hbbcd0cc6),
	.w3(32'hbafda0b5),
	.w4(32'hbae84538),
	.w5(32'h3b671427),
	.w6(32'hb9a245f7),
	.w7(32'hba1abedd),
	.w8(32'hba97ad47),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050980),
	.w1(32'h3b0f8a2c),
	.w2(32'h3b210706),
	.w3(32'h3bd5688a),
	.w4(32'hba861899),
	.w5(32'h3b6dcfed),
	.w6(32'h3bb48e93),
	.w7(32'h3bc1d1e1),
	.w8(32'h3bf30af7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a4697),
	.w1(32'hbbd43fd5),
	.w2(32'h3bb66dcb),
	.w3(32'hbc02580c),
	.w4(32'hbb4e5bf9),
	.w5(32'hba43c5ec),
	.w6(32'hbab7c420),
	.w7(32'hbb3e3af1),
	.w8(32'h3bbbb098),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f47f8),
	.w1(32'hb8fc5198),
	.w2(32'hbb8de207),
	.w3(32'hbb5bc20f),
	.w4(32'h39c2a2ad),
	.w5(32'hbb647bd7),
	.w6(32'h3c0180bf),
	.w7(32'hbb64b5de),
	.w8(32'hbc000b88),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901646),
	.w1(32'h3be7e792),
	.w2(32'hbc91de89),
	.w3(32'h3ad9b7ad),
	.w4(32'hbcbed818),
	.w5(32'hbdbdf050),
	.w6(32'h3d57c1aa),
	.w7(32'h3d9ba614),
	.w8(32'h3d6bf546),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4f1a5),
	.w1(32'h3be3e8eb),
	.w2(32'h3ac47f72),
	.w3(32'hbd19b918),
	.w4(32'h3b89afc1),
	.w5(32'h3bbd366f),
	.w6(32'h3c1deb73),
	.w7(32'h3bae34cd),
	.w8(32'h3c4497d2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c141d52),
	.w1(32'hbc9c501e),
	.w2(32'hbccda1e4),
	.w3(32'h3bca6920),
	.w4(32'hbb5159f7),
	.w5(32'hbb9497da),
	.w6(32'hbb3a663b),
	.w7(32'h3a28527e),
	.w8(32'h3c280f4f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35804b),
	.w1(32'hbacaf73c),
	.w2(32'hbb60052d),
	.w3(32'hbba39a1e),
	.w4(32'h3b6c1d14),
	.w5(32'hbb1e6d5a),
	.w6(32'h3aa3e155),
	.w7(32'h3b4c2c73),
	.w8(32'hb98106e0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269568),
	.w1(32'hbb39ff34),
	.w2(32'h3c3ee1cf),
	.w3(32'hbbe164f8),
	.w4(32'h3d007f16),
	.w5(32'h3db03c0e),
	.w6(32'hbcdc6cd7),
	.w7(32'hbd4f80ab),
	.w8(32'hbd1dccc2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39059720),
	.w1(32'hbace962b),
	.w2(32'h3c12fe07),
	.w3(32'h3d437cee),
	.w4(32'h3a08a54d),
	.w5(32'h3a9a3c5d),
	.w6(32'h3c1ef715),
	.w7(32'h3bd6054f),
	.w8(32'h3b32d55c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92dccb7),
	.w1(32'hbc300838),
	.w2(32'hbc93de98),
	.w3(32'h3adcc41b),
	.w4(32'hbc34761b),
	.w5(32'hbd08ea0c),
	.w6(32'h3bc722bd),
	.w7(32'h3c041f57),
	.w8(32'h3bd591d3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5c7c1),
	.w1(32'hbc2b4fef),
	.w2(32'hbc239f39),
	.w3(32'hbcc102f5),
	.w4(32'hbc0c3ba9),
	.w5(32'hbbd4c35c),
	.w6(32'hbc284e00),
	.w7(32'hbb97f5b7),
	.w8(32'hbba58686),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd1a72),
	.w1(32'hbc0d44eb),
	.w2(32'hbc747c94),
	.w3(32'hbb86aecf),
	.w4(32'hbae55cc1),
	.w5(32'hba97db7b),
	.w6(32'hbaaa5d94),
	.w7(32'hbc8a7083),
	.w8(32'hbc0ba40d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc358ea7),
	.w1(32'hbb377ab7),
	.w2(32'hbbed519d),
	.w3(32'hbb99860c),
	.w4(32'h3a422569),
	.w5(32'h3b3f8431),
	.w6(32'h3bc21f4a),
	.w7(32'h3b93bfcd),
	.w8(32'h3c171b10),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55c510),
	.w1(32'hba8e9489),
	.w2(32'h3bfd8b5b),
	.w3(32'h3b9752fd),
	.w4(32'h3ca34e72),
	.w5(32'h3d64891c),
	.w6(32'hbc678c53),
	.w7(32'hbcfe974d),
	.w8(32'hbcc77406),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e2f08),
	.w1(32'h3b4b7550),
	.w2(32'hbbf39082),
	.w3(32'h3d0371fa),
	.w4(32'hbb962834),
	.w5(32'hbc039a3f),
	.w6(32'h3c1e85a9),
	.w7(32'h3c1ad9b6),
	.w8(32'h3bd37919),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109644),
	.w1(32'hbac230f8),
	.w2(32'hbb9f6972),
	.w3(32'hbbfa2d0d),
	.w4(32'hbb9a2ec1),
	.w5(32'hbb95fc94),
	.w6(32'hbb7b20d0),
	.w7(32'hba794816),
	.w8(32'hbb4485df),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7d5b),
	.w1(32'hbbc3c7a9),
	.w2(32'hbc7564c1),
	.w3(32'hbb754fa6),
	.w4(32'hbbcb4dcc),
	.w5(32'hbb6ee793),
	.w6(32'hbc3eaac8),
	.w7(32'hbba7ff4e),
	.w8(32'hba4ae6b9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0634f5),
	.w1(32'h3b453c08),
	.w2(32'hbb65ee35),
	.w3(32'hbc19b29a),
	.w4(32'hbad9ba5d),
	.w5(32'hbb25ebc5),
	.w6(32'h3c364ae3),
	.w7(32'h3c19568c),
	.w8(32'h3b86404e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba78d64),
	.w1(32'hbb9de613),
	.w2(32'h3a7def82),
	.w3(32'hbb1cb3e5),
	.w4(32'h3a40b5df),
	.w5(32'h3ae88ebc),
	.w6(32'hbb1dc96c),
	.w7(32'hb9b1fe48),
	.w8(32'h3bf5334c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f1754),
	.w1(32'hb990f6ab),
	.w2(32'h3be0f208),
	.w3(32'h3bf1f490),
	.w4(32'hbb07dd51),
	.w5(32'h3bb8c3be),
	.w6(32'h3b9a7277),
	.w7(32'h3b265c55),
	.w8(32'h3bd4a41e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb77cfb),
	.w1(32'hbc5d28e6),
	.w2(32'h38e228b3),
	.w3(32'h3acf23d1),
	.w4(32'h3ce7cd81),
	.w5(32'h3da61fde),
	.w6(32'hbd10ccae),
	.w7(32'hbd8367f6),
	.w8(32'hbd3e6741),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69b330),
	.w1(32'hbb90e2a2),
	.w2(32'hbbd0c3c9),
	.w3(32'h3d219fea),
	.w4(32'hbbfd76fa),
	.w5(32'hbb0455d6),
	.w6(32'hbadcf810),
	.w7(32'hbb2aaac9),
	.w8(32'hbbb6cd60),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78df0),
	.w1(32'hbaa70bd1),
	.w2(32'h3b08561c),
	.w3(32'hbbd0fab9),
	.w4(32'hbba0e22f),
	.w5(32'hbc749390),
	.w6(32'hbc08aefe),
	.w7(32'h3b9d78b0),
	.w8(32'hba07e057),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f62d),
	.w1(32'hbae3387a),
	.w2(32'h3b61720b),
	.w3(32'hbbefef88),
	.w4(32'h3b9cebec),
	.w5(32'hb95377c8),
	.w6(32'h3998250a),
	.w7(32'h3c19e73c),
	.w8(32'h3b84ca47),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58da9f),
	.w1(32'hbac5a436),
	.w2(32'h3abccfdd),
	.w3(32'hbc4f8bc0),
	.w4(32'hbafc2d21),
	.w5(32'h3a21995f),
	.w6(32'hbb006819),
	.w7(32'h393c9682),
	.w8(32'hbace4560),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb856f934),
	.w1(32'h3b2d76a4),
	.w2(32'hbbf983cd),
	.w3(32'h39ea3a60),
	.w4(32'h3a005dec),
	.w5(32'hb9a2ac96),
	.w6(32'h3be23099),
	.w7(32'hbc046973),
	.w8(32'hb9ff8080),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule