module layer_8_featuremap_89(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ac996),
	.w1(32'h3a33fe00),
	.w2(32'h3aec4380),
	.w3(32'h3b239484),
	.w4(32'hbc40bc0e),
	.w5(32'hbb643d60),
	.w6(32'hbaa5d034),
	.w7(32'hba287c54),
	.w8(32'hbc297ae0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02f082),
	.w1(32'h3a3dffe2),
	.w2(32'h3d529a58),
	.w3(32'hba93329d),
	.w4(32'h3bce85f2),
	.w5(32'hbad9bd1a),
	.w6(32'h3b744e1e),
	.w7(32'hb98dc3c1),
	.w8(32'h3aee22f1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37c6a0),
	.w1(32'hbc0c68c1),
	.w2(32'hba303032),
	.w3(32'hbb13d7a4),
	.w4(32'hba9a181d),
	.w5(32'hbbb6d306),
	.w6(32'h39124980),
	.w7(32'hbc407b08),
	.w8(32'hbc1f9f41),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be069ad),
	.w1(32'hbb9903cf),
	.w2(32'hbb750c68),
	.w3(32'hbc128452),
	.w4(32'hbc955b9a),
	.w5(32'h3bb13592),
	.w6(32'hbc196fcd),
	.w7(32'hbbfed658),
	.w8(32'hbb66fd22),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b5b6f),
	.w1(32'hbbb6bc5b),
	.w2(32'h3bc47ba9),
	.w3(32'hbad27bfe),
	.w4(32'h3b2dd6b2),
	.w5(32'hba6ca896),
	.w6(32'hbbef6552),
	.w7(32'h3786541b),
	.w8(32'hbbc7bef5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6d7e9),
	.w1(32'h3c2c43fe),
	.w2(32'hbc620349),
	.w3(32'hbc482699),
	.w4(32'h3ccd937c),
	.w5(32'hbb15de38),
	.w6(32'hbc066e78),
	.w7(32'hbb270dbc),
	.w8(32'hbc444c2b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ababacc),
	.w1(32'h3bd7b60d),
	.w2(32'hba620a52),
	.w3(32'h3b80e736),
	.w4(32'hbb43b820),
	.w5(32'h3c42eaa2),
	.w6(32'hbb7ae774),
	.w7(32'hba3aa252),
	.w8(32'h3c1fa7fb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a02a8),
	.w1(32'hbb38f1f9),
	.w2(32'h3b61a4de),
	.w3(32'h3bc11776),
	.w4(32'hbb4834ad),
	.w5(32'hb95e733f),
	.w6(32'hbbbc536c),
	.w7(32'hbbb99d15),
	.w8(32'hbbd7789c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a1caf),
	.w1(32'h3b55948b),
	.w2(32'hbc546876),
	.w3(32'h3b6eba54),
	.w4(32'h3bb1479f),
	.w5(32'hbb5403ec),
	.w6(32'h3b842da5),
	.w7(32'hbae59838),
	.w8(32'h3c0593ac),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc86f8a),
	.w1(32'hbc542998),
	.w2(32'hbbcc4f35),
	.w3(32'h399e2fea),
	.w4(32'hbb9e2d18),
	.w5(32'hbb7bd30f),
	.w6(32'hbc6264d0),
	.w7(32'h3bd2e527),
	.w8(32'h3ba321cc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b905d5c),
	.w1(32'h3c1a955b),
	.w2(32'h3b2112eb),
	.w3(32'hbcb109d2),
	.w4(32'hbc73cb4e),
	.w5(32'h3acf596f),
	.w6(32'hbbf10e24),
	.w7(32'hbc2dfafc),
	.w8(32'hbb06373d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176000),
	.w1(32'hbd48c893),
	.w2(32'hbc050a4c),
	.w3(32'hbbacc4de),
	.w4(32'hbbb58369),
	.w5(32'hb9fec042),
	.w6(32'h3ba47f6f),
	.w7(32'h3bd16c73),
	.w8(32'hbb455c4c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e71b),
	.w1(32'hbae9b966),
	.w2(32'hbca552ad),
	.w3(32'h3aa4e594),
	.w4(32'h3b949783),
	.w5(32'h3ab375f8),
	.w6(32'hbb4e4370),
	.w7(32'hbabcd1d4),
	.w8(32'hbc2763e6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb711889),
	.w1(32'hb78f8ec6),
	.w2(32'h3c00fd2e),
	.w3(32'hbaff383b),
	.w4(32'hbc340b90),
	.w5(32'hbb10e8cd),
	.w6(32'h3bb1b30a),
	.w7(32'hbb48c993),
	.w8(32'hbb7f2bdd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55c252),
	.w1(32'h3bd507ba),
	.w2(32'h3a0788b3),
	.w3(32'hbb292d55),
	.w4(32'hbca7486b),
	.w5(32'hbbe98121),
	.w6(32'hbbdb4e7e),
	.w7(32'h3cf675aa),
	.w8(32'h3be0d503),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038bd4),
	.w1(32'hbca844d9),
	.w2(32'h3b79707b),
	.w3(32'hbc6858a6),
	.w4(32'hbbd96108),
	.w5(32'h3b03ab77),
	.w6(32'hbb546298),
	.w7(32'hbc9a83ef),
	.w8(32'hbc2d11f7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94f04a),
	.w1(32'h3cd5d9f7),
	.w2(32'h3c01d845),
	.w3(32'h3ba6125c),
	.w4(32'hbbc85166),
	.w5(32'hbb30e74c),
	.w6(32'hbc0fe133),
	.w7(32'hbc5641c5),
	.w8(32'hbd0f4183),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45349b),
	.w1(32'h3bbd4d71),
	.w2(32'hb98fb419),
	.w3(32'h39718d91),
	.w4(32'hbc3be3c4),
	.w5(32'hbb320174),
	.w6(32'h3b353b34),
	.w7(32'h3d00fea9),
	.w8(32'hbbe1b53e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7623b0),
	.w1(32'h3c655b09),
	.w2(32'h3ce90252),
	.w3(32'hbd598a85),
	.w4(32'hbd08c5ad),
	.w5(32'h3d1aa5a9),
	.w6(32'h3c0f12d9),
	.w7(32'hbc1fc223),
	.w8(32'hbb57e56b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7612e2),
	.w1(32'hbce1a1f8),
	.w2(32'hbc8f47e7),
	.w3(32'h3b6fe19c),
	.w4(32'hb9e26679),
	.w5(32'hbbffefd6),
	.w6(32'h3bbcb822),
	.w7(32'h3c8645dd),
	.w8(32'hbbabffa5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b7b78),
	.w1(32'h3c5dda03),
	.w2(32'hbc41020a),
	.w3(32'hbc05c1ba),
	.w4(32'hbad2d2e3),
	.w5(32'hbd3b190e),
	.w6(32'h3d551bad),
	.w7(32'hbbc40555),
	.w8(32'hbba45950),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73ab88),
	.w1(32'h3cb8339f),
	.w2(32'h3c9fda63),
	.w3(32'h3bde4b70),
	.w4(32'h3d0bfafa),
	.w5(32'h3d419d55),
	.w6(32'h3c4e3e4a),
	.w7(32'h3bca063e),
	.w8(32'h3b1634fd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4a5b8),
	.w1(32'hbc394804),
	.w2(32'hbbbfada4),
	.w3(32'h3b34936d),
	.w4(32'hbcbd02ff),
	.w5(32'h3bef79ab),
	.w6(32'hba192658),
	.w7(32'hbd0da92a),
	.w8(32'hba830d7e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfe2e9),
	.w1(32'h3c069a2c),
	.w2(32'hbb628193),
	.w3(32'hbc926f30),
	.w4(32'hbc2be831),
	.w5(32'h3d440396),
	.w6(32'hbbb98fbb),
	.w7(32'hbc8db547),
	.w8(32'hbd1dfa8c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf24d0),
	.w1(32'h3bbf56ae),
	.w2(32'h3c60b4c5),
	.w3(32'hbc709b46),
	.w4(32'hbd2ee7bd),
	.w5(32'hbb23ed85),
	.w6(32'hbb9633dc),
	.w7(32'h3bfb6e6e),
	.w8(32'hbaa3a880),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f3c64),
	.w1(32'h3ada6f16),
	.w2(32'h3b18f55c),
	.w3(32'hbaa94eaf),
	.w4(32'hbc38890a),
	.w5(32'hbac8351f),
	.w6(32'h3c4c49ec),
	.w7(32'hba67a97e),
	.w8(32'h3a012f8b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3d441),
	.w1(32'hbb93bc2f),
	.w2(32'h3c4b78b9),
	.w3(32'h3c982d56),
	.w4(32'h3c859fdd),
	.w5(32'hbca6bd2e),
	.w6(32'hbb69b095),
	.w7(32'hbc230a50),
	.w8(32'hbbd25da5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9cabe),
	.w1(32'h3d24dd42),
	.w2(32'hbd1436c1),
	.w3(32'hba948d70),
	.w4(32'hbe370d80),
	.w5(32'hbd3ebfdb),
	.w6(32'h3cf97662),
	.w7(32'h3d158ae7),
	.w8(32'hbdda974b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3b8c63),
	.w1(32'h3b7b9195),
	.w2(32'hbaa4ec75),
	.w3(32'hbd14eaa7),
	.w4(32'hbc101c21),
	.w5(32'hbcb6c545),
	.w6(32'hbc4704c9),
	.w7(32'hbd387489),
	.w8(32'hbd76ead6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd45f2b),
	.w1(32'hbdcd820e),
	.w2(32'hbbf8fe56),
	.w3(32'h3c8508e2),
	.w4(32'hbd10335d),
	.w5(32'h3bb9b2e2),
	.w6(32'hbcb1fdfa),
	.w7(32'h3ccc59d9),
	.w8(32'hbd089431),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd371d0f),
	.w1(32'h3ca37545),
	.w2(32'hbc20b96a),
	.w3(32'h3d46868b),
	.w4(32'h3bf4adb8),
	.w5(32'h3c303c48),
	.w6(32'h3cba664d),
	.w7(32'h3b1478de),
	.w8(32'hbb2a03e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabbacf),
	.w1(32'hbbc9e5ee),
	.w2(32'hbd24644e),
	.w3(32'hbd459fa3),
	.w4(32'h3c1ee38b),
	.w5(32'h3ca77109),
	.w6(32'hbbeb59bd),
	.w7(32'h3ca0f232),
	.w8(32'h3b85f31f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc5177),
	.w1(32'hbd3f3cbd),
	.w2(32'h3c6bca7e),
	.w3(32'hbc201908),
	.w4(32'hbcb7afed),
	.w5(32'hbcb8400d),
	.w6(32'hbb50ad45),
	.w7(32'hbc9ba9a6),
	.w8(32'hbcc3f639),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd60b51),
	.w1(32'hbc707a8c),
	.w2(32'h3ce6d60c),
	.w3(32'hbc864a8a),
	.w4(32'hbce7975e),
	.w5(32'h3ccff2d2),
	.w6(32'hbbc736b5),
	.w7(32'hbb950fb7),
	.w8(32'h3bbb7145),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b533c61),
	.w1(32'hbc9c6851),
	.w2(32'h3c9e4497),
	.w3(32'h3b07b289),
	.w4(32'hbbbcb276),
	.w5(32'h3cdb9eb1),
	.w6(32'h3ce8601e),
	.w7(32'h3d569028),
	.w8(32'h3c876b99),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5767c5),
	.w1(32'h3bff1ce0),
	.w2(32'hbd280745),
	.w3(32'hbca2414b),
	.w4(32'hbb5c4b80),
	.w5(32'h3c82c5c1),
	.w6(32'hbd502f92),
	.w7(32'hbca6e917),
	.w8(32'hbab9082b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdd571ec),
	.w1(32'hbbe626b9),
	.w2(32'h3ca9ed19),
	.w3(32'hbc8dbad0),
	.w4(32'h3d015280),
	.w5(32'h3c13756b),
	.w6(32'hbcec9e98),
	.w7(32'h3ce1c4d9),
	.w8(32'h3cd47760),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1bf62),
	.w1(32'h3dc9f367),
	.w2(32'hbc5f292a),
	.w3(32'h3bec205a),
	.w4(32'h3c1b18f9),
	.w5(32'hbd8af904),
	.w6(32'hbacaed1a),
	.w7(32'hbc817845),
	.w8(32'h3d98d9fe),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53109),
	.w1(32'hbc0005c8),
	.w2(32'h3c33995f),
	.w3(32'h3d21553b),
	.w4(32'hbd6e81c4),
	.w5(32'h3c545b3c),
	.w6(32'h3b80d75a),
	.w7(32'h3af06565),
	.w8(32'h3bbc9dcb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a890),
	.w1(32'h3c03ba4b),
	.w2(32'h3c5d8b2b),
	.w3(32'h3b3187a2),
	.w4(32'h3c713636),
	.w5(32'hbce0296e),
	.w6(32'h3b00005d),
	.w7(32'h3b0623d5),
	.w8(32'h3b0532c9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc925643),
	.w1(32'hbcac7584),
	.w2(32'h3ba66568),
	.w3(32'hbd6d6833),
	.w4(32'hbc582de1),
	.w5(32'hbcc7a30a),
	.w6(32'hbcaa169e),
	.w7(32'hbacc52ad),
	.w8(32'hbc2070a4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b3bfc),
	.w1(32'hbc42b224),
	.w2(32'hbc15a92e),
	.w3(32'h3c5399e3),
	.w4(32'h3ccbc8b6),
	.w5(32'hbacd3a89),
	.w6(32'hbb688224),
	.w7(32'h3a37077b),
	.w8(32'hbb60a662),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd47301),
	.w1(32'hbcac22f8),
	.w2(32'h3a3c1321),
	.w3(32'h3c59b6f7),
	.w4(32'hbc17de0b),
	.w5(32'hbc32d7f7),
	.w6(32'h3ba5b3bd),
	.w7(32'hbb5fa940),
	.w8(32'hbcc2734c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03503f),
	.w1(32'hbc519865),
	.w2(32'hbcb6a60b),
	.w3(32'h3c845f2c),
	.w4(32'hbd068e1f),
	.w5(32'h3c84094c),
	.w6(32'hbc3e724a),
	.w7(32'hbc6560e6),
	.w8(32'h3c6d60ec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbfe917),
	.w1(32'h3cb4dfa9),
	.w2(32'h3d1e2335),
	.w3(32'hbcdfe759),
	.w4(32'hbc699461),
	.w5(32'h3c69f263),
	.w6(32'hbbac7ef8),
	.w7(32'h3b9b5a27),
	.w8(32'h3a4f60b6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd087999),
	.w1(32'hbcc45147),
	.w2(32'hbc3eec6b),
	.w3(32'h3ba4ae28),
	.w4(32'hbc16dbdf),
	.w5(32'h3c3c9132),
	.w6(32'hbbd4ebda),
	.w7(32'hba2a244b),
	.w8(32'hbd130f36),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ab99b),
	.w1(32'hbca901ad),
	.w2(32'hba17956c),
	.w3(32'hbaefd688),
	.w4(32'hbd46638f),
	.w5(32'h3a653446),
	.w6(32'hbce29061),
	.w7(32'h3b948f9e),
	.w8(32'hbb254cce),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c390c5f),
	.w1(32'hbcbac57a),
	.w2(32'hbcc922fa),
	.w3(32'h3bb998a2),
	.w4(32'hbb887042),
	.w5(32'hbb804a81),
	.w6(32'hbbcd0a7e),
	.w7(32'hbb9a1a47),
	.w8(32'hbb385937),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e56ac),
	.w1(32'hbc16313d),
	.w2(32'hbbc5db66),
	.w3(32'hbc067259),
	.w4(32'hbc342ce7),
	.w5(32'hbd0b22fb),
	.w6(32'hb9bbdcac),
	.w7(32'hbcd5e156),
	.w8(32'hbc80c941),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3969d),
	.w1(32'hbbab8235),
	.w2(32'hb926dec4),
	.w3(32'hbd34b4af),
	.w4(32'hbcd7be41),
	.w5(32'h3cb16928),
	.w6(32'hbbe4b230),
	.w7(32'hbad6e43f),
	.w8(32'hbc9deb82),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e8f0d),
	.w1(32'h3ab73c3f),
	.w2(32'h3b504811),
	.w3(32'h3d3d4e08),
	.w4(32'h3d2bc474),
	.w5(32'hbbac4b24),
	.w6(32'hbbb96456),
	.w7(32'hbc493c03),
	.w8(32'h3b2a46d9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d8994),
	.w1(32'h3aea6fa2),
	.w2(32'hbca40c42),
	.w3(32'hbd7e69bb),
	.w4(32'hbd18f814),
	.w5(32'hbcd2aa4c),
	.w6(32'h3cebbabe),
	.w7(32'hbcc1fa09),
	.w8(32'hbd17c8ef),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfdbc96),
	.w1(32'h3c40fb46),
	.w2(32'hbc27e144),
	.w3(32'hbc25af49),
	.w4(32'h3d8ad6ed),
	.w5(32'h3c2317e2),
	.w6(32'h3cb85346),
	.w7(32'hbcca8c78),
	.w8(32'h3ca254b0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc208c1),
	.w1(32'h3d7a254f),
	.w2(32'hbbbbe97d),
	.w3(32'h3cf70e69),
	.w4(32'h3bb46055),
	.w5(32'hbb2160e5),
	.w6(32'h3b88b4a6),
	.w7(32'h3c6b917d),
	.w8(32'h3c220bb3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc203329),
	.w1(32'hbc31dd44),
	.w2(32'h3c0f6cf2),
	.w3(32'h3b34faa5),
	.w4(32'hbba28d09),
	.w5(32'h3c2fe9fc),
	.w6(32'h3c8d7e7e),
	.w7(32'hbc850206),
	.w8(32'h3c9ae1b9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0831c2),
	.w1(32'h3bce69b5),
	.w2(32'hbc8a5897),
	.w3(32'hbadca919),
	.w4(32'hbca8bd5a),
	.w5(32'hbce93b00),
	.w6(32'hbc8998ff),
	.w7(32'hbaadc0e5),
	.w8(32'hbd36b9d1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73dd78),
	.w1(32'hbd364284),
	.w2(32'h3b621e1f),
	.w3(32'hbc109f38),
	.w4(32'h3d2a7cf3),
	.w5(32'hbaeb76f6),
	.w6(32'h3b052edf),
	.w7(32'hbc67e579),
	.w8(32'hbb6af69d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94f583),
	.w1(32'hbca0f1d3),
	.w2(32'hbd13ffb4),
	.w3(32'hbd0d1a8b),
	.w4(32'hbc0fbbc5),
	.w5(32'hbd6f28cb),
	.w6(32'h3d431ac9),
	.w7(32'hbca4306d),
	.w8(32'hbd53de90),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bb869),
	.w1(32'h3c8fe252),
	.w2(32'hbc000c46),
	.w3(32'hbce54fd5),
	.w4(32'hbc6fb132),
	.w5(32'hbbea8870),
	.w6(32'h3ca0c445),
	.w7(32'h3c3bf0ef),
	.w8(32'h3c15eb05),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceda4c2),
	.w1(32'hbb075ffd),
	.w2(32'hbd19202d),
	.w3(32'hbbd34806),
	.w4(32'hb96deef8),
	.w5(32'hbc0f9a62),
	.w6(32'hbcf23e5a),
	.w7(32'hbd74364d),
	.w8(32'h3a4abbd0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf31589),
	.w1(32'h3b9614ea),
	.w2(32'hbc99fe29),
	.w3(32'h3c1d760f),
	.w4(32'hbcc6ccdd),
	.w5(32'h3ce6140a),
	.w6(32'h3c8e81e3),
	.w7(32'hbcd10fe3),
	.w8(32'hbc837405),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b3854),
	.w1(32'hbd1c90c6),
	.w2(32'hbbd44fd0),
	.w3(32'h3aed3d35),
	.w4(32'h3d64598c),
	.w5(32'h3bbde4cc),
	.w6(32'h3d108aa9),
	.w7(32'hbbb1d023),
	.w8(32'hbd54030d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9acc10),
	.w1(32'hbbc3efa5),
	.w2(32'hbd27e285),
	.w3(32'hbc5f167a),
	.w4(32'hbc953782),
	.w5(32'hbc529ec8),
	.w6(32'hbbc1f2a8),
	.w7(32'hbd2e285d),
	.w8(32'h3ccb45c1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a3fdb),
	.w1(32'hbcf8e8b3),
	.w2(32'h3c935119),
	.w3(32'h3b82c760),
	.w4(32'hbc567068),
	.w5(32'h3d209a10),
	.w6(32'hbd2aee9c),
	.w7(32'hbbae2ed0),
	.w8(32'h3cdea6a1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdc508),
	.w1(32'h3b85bd81),
	.w2(32'hbbf321ff),
	.w3(32'h3d66c282),
	.w4(32'hbc619183),
	.w5(32'hbc548ac2),
	.w6(32'hbc9fc193),
	.w7(32'hbbc47d18),
	.w8(32'hbc4281c4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddb2a1),
	.w1(32'hbcf052aa),
	.w2(32'hbc6d7008),
	.w3(32'hbc927aaf),
	.w4(32'h3bc60bb2),
	.w5(32'hb926c28d),
	.w6(32'hbd21cdfc),
	.w7(32'h3b5c7aac),
	.w8(32'h3c10796d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc353e1),
	.w1(32'h3bfc5197),
	.w2(32'hbc95ad14),
	.w3(32'hbd2ab249),
	.w4(32'h3ceaf9ef),
	.w5(32'hbbe77298),
	.w6(32'hbd39c16b),
	.w7(32'hbd76b06a),
	.w8(32'h3c54edff),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb129e8b),
	.w1(32'h3b0c58e0),
	.w2(32'hba314fea),
	.w3(32'hbd287b03),
	.w4(32'hbc42ccd3),
	.w5(32'h3c707664),
	.w6(32'h3d036d4e),
	.w7(32'h3bcb1f2d),
	.w8(32'hbd104313),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ca049),
	.w1(32'h3c96a4c1),
	.w2(32'h3cf6c585),
	.w3(32'h3b3db3a3),
	.w4(32'h3c2dcb2d),
	.w5(32'hbc4cf9d7),
	.w6(32'hbba297ee),
	.w7(32'hbc830c48),
	.w8(32'hba5bcf11),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c083a),
	.w1(32'h3aefffb0),
	.w2(32'hbc4ffd1e),
	.w3(32'hbd2fbeeb),
	.w4(32'hbc63b46a),
	.w5(32'h3cdda1f5),
	.w6(32'hbd27cf0c),
	.w7(32'hbcc60863),
	.w8(32'h3c1162cc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be25a4b),
	.w1(32'hbb482bb9),
	.w2(32'hbbff21f1),
	.w3(32'hba25e904),
	.w4(32'hbc4f203f),
	.w5(32'hbb9df687),
	.w6(32'h3bb2bc68),
	.w7(32'hbd8192e0),
	.w8(32'hbd7efca0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842c2c),
	.w1(32'h3c0b4f57),
	.w2(32'hb911daac),
	.w3(32'h3cb68c21),
	.w4(32'h3b830548),
	.w5(32'hbc37563a),
	.w6(32'hbcbabbb1),
	.w7(32'h3d417c73),
	.w8(32'h3c657dd4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d082bbe),
	.w1(32'hbc49f362),
	.w2(32'h3c9aafb1),
	.w3(32'h3cd966f0),
	.w4(32'hbc09c851),
	.w5(32'hbbb3e10c),
	.w6(32'h3c1b6624),
	.w7(32'hbae2f757),
	.w8(32'hbbd47bb7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90aad4),
	.w1(32'hbd2b6ace),
	.w2(32'h3c22c25f),
	.w3(32'hbcd027b6),
	.w4(32'h3c8be3ff),
	.w5(32'h3c21f672),
	.w6(32'h3c63db94),
	.w7(32'hb93d7674),
	.w8(32'h3bbb7556),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff6499),
	.w1(32'hbc6b831e),
	.w2(32'h3d16b4ec),
	.w3(32'h3be00837),
	.w4(32'h3a31e86f),
	.w5(32'h39762d6d),
	.w6(32'hbcea2511),
	.w7(32'hbcb6cd1c),
	.w8(32'h3d852791),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45ecbd),
	.w1(32'hbc1d1e75),
	.w2(32'h39a4fde1),
	.w3(32'hbb92fe0b),
	.w4(32'hbd362d03),
	.w5(32'hbcc53b8c),
	.w6(32'hbbe4e446),
	.w7(32'h3c782da0),
	.w8(32'h3c62728b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560c76),
	.w1(32'h3d093af7),
	.w2(32'h3bc01926),
	.w3(32'hbc05d5a4),
	.w4(32'hbc5b405d),
	.w5(32'h3c8fbccf),
	.w6(32'h3d403c2d),
	.w7(32'hbb98f404),
	.w8(32'h3d198a95),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe167df),
	.w1(32'h3c48f78e),
	.w2(32'hbba59163),
	.w3(32'h3b041301),
	.w4(32'h3c506dab),
	.w5(32'hbb9feeb2),
	.w6(32'hbc9a7890),
	.w7(32'h3d2ec25d),
	.w8(32'hbb92acf4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53e8e7),
	.w1(32'hbb7e34c4),
	.w2(32'h3c5e88f3),
	.w3(32'h38169a25),
	.w4(32'hbc3f0539),
	.w5(32'h3c3566fb),
	.w6(32'hbbe2b71c),
	.w7(32'h3c4a5cb3),
	.w8(32'hba9f6a30),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ba6b1),
	.w1(32'h39e63754),
	.w2(32'h3c4a85e4),
	.w3(32'hb9e41f33),
	.w4(32'hbd01ece5),
	.w5(32'hbc927470),
	.w6(32'hbc7cdd23),
	.w7(32'h3b319541),
	.w8(32'h3c601085),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd020eb0),
	.w1(32'hbb5ca152),
	.w2(32'hb8eb0cfd),
	.w3(32'hbba81705),
	.w4(32'hbb837259),
	.w5(32'hbc033e43),
	.w6(32'hbb41a68a),
	.w7(32'h3cb2b0e9),
	.w8(32'h3c268aca),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9737a0),
	.w1(32'h3c6587c5),
	.w2(32'h3c45b77e),
	.w3(32'hbc54bff0),
	.w4(32'hbc74521a),
	.w5(32'h3bd9fa34),
	.w6(32'hbc799535),
	.w7(32'hb90bcd7c),
	.w8(32'h3c65ed05),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbaeed5),
	.w1(32'hbc113c4f),
	.w2(32'hbb2a90b4),
	.w3(32'hbc5bbbf9),
	.w4(32'hbbb70e4b),
	.w5(32'h3d41c95b),
	.w6(32'hbbcaa83b),
	.w7(32'h3c8463d9),
	.w8(32'h3c2aa787),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd200861),
	.w1(32'h3afc0b1c),
	.w2(32'hbcaf7cb9),
	.w3(32'hbc23c25d),
	.w4(32'h3c872a58),
	.w5(32'hbd179085),
	.w6(32'h3a9c2bdb),
	.w7(32'hbc1a0750),
	.w8(32'hbc5edb41),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d16ac9a),
	.w1(32'h3c1bec3e),
	.w2(32'hbd451255),
	.w3(32'hbaba09d8),
	.w4(32'hbaec9a77),
	.w5(32'h3d070e2e),
	.w6(32'h3c3a8903),
	.w7(32'h3b25cdf5),
	.w8(32'h3b8959a1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f60ed),
	.w1(32'h3c194086),
	.w2(32'h3d2ac2cf),
	.w3(32'hb8966e6d),
	.w4(32'h3b141b27),
	.w5(32'h3ca684ba),
	.w6(32'h3d71e747),
	.w7(32'hbbe85ba3),
	.w8(32'hbd06a151),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77b956),
	.w1(32'h3d847e8a),
	.w2(32'hbb627b15),
	.w3(32'h3d7d686e),
	.w4(32'h3ca2ff2b),
	.w5(32'hbb9ce85a),
	.w6(32'h3d13661d),
	.w7(32'h3bebb26f),
	.w8(32'hbc7964e8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99fab5),
	.w1(32'h3ce839d5),
	.w2(32'h3cd4a253),
	.w3(32'hbb63e928),
	.w4(32'hbb2455a1),
	.w5(32'hbc568b78),
	.w6(32'hbb0c04c9),
	.w7(32'hbcc8cbe6),
	.w8(32'hbb4ab1f6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d62cf62),
	.w1(32'hbb838fd2),
	.w2(32'hbca05edf),
	.w3(32'h3ccd5559),
	.w4(32'h3c86c03c),
	.w5(32'hbc6b25bb),
	.w6(32'hbd32b3d4),
	.w7(32'h3d8ba34e),
	.w8(32'h3d7eb783),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d83a3f7),
	.w1(32'hbc53860a),
	.w2(32'hbc98f4ea),
	.w3(32'h3d50099b),
	.w4(32'h3c638797),
	.w5(32'h3c1bbfc5),
	.w6(32'h3b353239),
	.w7(32'hb930ead4),
	.w8(32'h3d299ea1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5c435),
	.w1(32'h3d80024a),
	.w2(32'hbd6d973a),
	.w3(32'hbc955f3a),
	.w4(32'h3d019df3),
	.w5(32'hbcc60030),
	.w6(32'h3b9129fa),
	.w7(32'hbd2c8d9c),
	.w8(32'hbc8be4a6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd4af4),
	.w1(32'h3d83e69b),
	.w2(32'h3d37c66f),
	.w3(32'hbbd43c32),
	.w4(32'h3d29bec5),
	.w5(32'h3c941610),
	.w6(32'hbb8f7dc3),
	.w7(32'hbcb04d2e),
	.w8(32'h3c886af7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9010d3),
	.w1(32'h3c2ddf51),
	.w2(32'h3c4013cf),
	.w3(32'h3d863a5e),
	.w4(32'h3cc48d8b),
	.w5(32'h3d5575c0),
	.w6(32'h3cc81ca0),
	.w7(32'h3d14d256),
	.w8(32'h3c90193a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e4a8d),
	.w1(32'hbc964c91),
	.w2(32'h3d59bd3e),
	.w3(32'h3cc8edd0),
	.w4(32'hbb48c053),
	.w5(32'h3cf2167a),
	.w6(32'hba3abda5),
	.w7(32'hbb2bc5a9),
	.w8(32'h3bb0c8c0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc640),
	.w1(32'hbc4d6e61),
	.w2(32'h3d2c12ed),
	.w3(32'h3ccdddfe),
	.w4(32'h3d8087e1),
	.w5(32'h3ca4d1ce),
	.w6(32'h3ce5e879),
	.w7(32'h3d648634),
	.w8(32'hbc2ee9d0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd35cb19),
	.w1(32'hbcce5f87),
	.w2(32'h3c8856df),
	.w3(32'h3d0fcf8d),
	.w4(32'h3af9309a),
	.w5(32'hbd316ac1),
	.w6(32'h3c893c1b),
	.w7(32'h3d1d8dd0),
	.w8(32'h3c8b429d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2437c1),
	.w1(32'hbb19dd38),
	.w2(32'hbcd37e41),
	.w3(32'hbc2bbd99),
	.w4(32'h3aba5e29),
	.w5(32'hbd0bc6de),
	.w6(32'hbd3fb9a9),
	.w7(32'hbb051185),
	.w8(32'h3b703fb7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8f335),
	.w1(32'hbcbd4fff),
	.w2(32'h3d68f6e6),
	.w3(32'h3d31e0a7),
	.w4(32'hbd0bef81),
	.w5(32'h37b45e74),
	.w6(32'h3d1554cb),
	.w7(32'h3c4ec489),
	.w8(32'h3c6dc240),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9252d),
	.w1(32'hbd2e7c08),
	.w2(32'h3b6017dd),
	.w3(32'h3bf0867d),
	.w4(32'h3b2f9caf),
	.w5(32'h3b49ebc9),
	.w6(32'hbc7aa963),
	.w7(32'h3aff3743),
	.w8(32'h3c0131e6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdea0bc1),
	.w1(32'hbd389c22),
	.w2(32'h3ad1c4f1),
	.w3(32'h3d1efaf5),
	.w4(32'hbd411e2c),
	.w5(32'h3c2c5bbc),
	.w6(32'hbc6376a0),
	.w7(32'hbb87f7e2),
	.w8(32'h3c7c7475),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93c202),
	.w1(32'h3c893720),
	.w2(32'hbc2aa480),
	.w3(32'h3c196232),
	.w4(32'hbc7a6d3b),
	.w5(32'hbc7bcbc6),
	.w6(32'hbaa21031),
	.w7(32'h3c931cbe),
	.w8(32'h3cce1cbf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bfdc4),
	.w1(32'hbc7bdf33),
	.w2(32'hbcafa86d),
	.w3(32'hbbc918a1),
	.w4(32'h3d084fdc),
	.w5(32'hbc07903d),
	.w6(32'h3cfba9ec),
	.w7(32'hbc9ff098),
	.w8(32'h3c1bfe34),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014a17),
	.w1(32'h3c8c4b37),
	.w2(32'h3c9bccdf),
	.w3(32'hbbf25446),
	.w4(32'hbbace803),
	.w5(32'hbc9c215b),
	.w6(32'h3d0d6f12),
	.w7(32'h3b5abf05),
	.w8(32'hbbfd8b37),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4bbaa),
	.w1(32'hbcdb45d2),
	.w2(32'h3ca861aa),
	.w3(32'hbba5f914),
	.w4(32'hbc33ed8c),
	.w5(32'h3bc196ae),
	.w6(32'hbbf2ac4d),
	.w7(32'hbb61cf9d),
	.w8(32'h3c03e949),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd37126),
	.w1(32'hbc2d70cf),
	.w2(32'h3dbfdac0),
	.w3(32'hbd1a5508),
	.w4(32'hbbe91c1e),
	.w5(32'h3b0504d0),
	.w6(32'hbb49d9bd),
	.w7(32'h3c9cd6a5),
	.w8(32'h3c179f9a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca0765),
	.w1(32'hbca69802),
	.w2(32'hbc248781),
	.w3(32'hbc1b4063),
	.w4(32'hbcdf7d0a),
	.w5(32'h3c4fa0f8),
	.w6(32'h3bd41e85),
	.w7(32'hbd6d703e),
	.w8(32'hbd514ecc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2286d2),
	.w1(32'h3cffdcc3),
	.w2(32'hbd34a18e),
	.w3(32'hbc7dc54d),
	.w4(32'h3c0ba205),
	.w5(32'hbd22e0d9),
	.w6(32'hbbc8c654),
	.w7(32'h3bd47be5),
	.w8(32'hbcc6a936),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40ced4),
	.w1(32'hbe0d28ac),
	.w2(32'hbcc3f142),
	.w3(32'h395a209e),
	.w4(32'h3cba35e5),
	.w5(32'h39a4dfd1),
	.w6(32'hbc6b4bd1),
	.w7(32'h3c5a81cb),
	.w8(32'hbd39664c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd13a4a0),
	.w1(32'hbad84f76),
	.w2(32'h3ca00055),
	.w3(32'hbc6fc8bd),
	.w4(32'h3d21bf18),
	.w5(32'h3d20284f),
	.w6(32'hbc107bd2),
	.w7(32'h3a1758bf),
	.w8(32'h3cd10423),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d179eb0),
	.w1(32'hbc742316),
	.w2(32'hbb21fbb8),
	.w3(32'hbd324c44),
	.w4(32'hbb210239),
	.w5(32'hbcf5deec),
	.w6(32'hbbc03b71),
	.w7(32'hbc914382),
	.w8(32'hbbd4bb50),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeeadf),
	.w1(32'h3bd064c5),
	.w2(32'hbc7363ca),
	.w3(32'hba22f453),
	.w4(32'h3bb04af9),
	.w5(32'h3b7bb918),
	.w6(32'hbac13f98),
	.w7(32'hbd70166f),
	.w8(32'h3b189472),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad60907),
	.w1(32'hbd735fb7),
	.w2(32'h3be545e8),
	.w3(32'hbd8be742),
	.w4(32'hbd03a2cc),
	.w5(32'hbc388d17),
	.w6(32'h3c90a1fc),
	.w7(32'hbab001da),
	.w8(32'hb81ba22c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac33c7),
	.w1(32'h3b261025),
	.w2(32'hba8b73e3),
	.w3(32'hbd4ed24a),
	.w4(32'h3c7ddc16),
	.w5(32'hbcc9b8ab),
	.w6(32'h3bb17829),
	.w7(32'h3bbfd13d),
	.w8(32'h3b518c65),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d96ee),
	.w1(32'h3c2a548f),
	.w2(32'hbbf19b11),
	.w3(32'h3c16aa5f),
	.w4(32'h3bbb5895),
	.w5(32'hbbc86d5c),
	.w6(32'hbb98563a),
	.w7(32'h3c898ba8),
	.w8(32'hbd389e74),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d4f82),
	.w1(32'hbab8d872),
	.w2(32'hbca2ab03),
	.w3(32'hbcd59436),
	.w4(32'hbb96075e),
	.w5(32'hbc6b6ffd),
	.w6(32'hbd08e5f0),
	.w7(32'hbc8c80e5),
	.w8(32'hbcf6362a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf46d05),
	.w1(32'hbd9c8271),
	.w2(32'h3d0f26e0),
	.w3(32'hbbeac932),
	.w4(32'h3b4828eb),
	.w5(32'hbb399931),
	.w6(32'hbc923e3f),
	.w7(32'hbc433cda),
	.w8(32'h3b6d98fd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becfb25),
	.w1(32'hbc81ce94),
	.w2(32'h3c982e8d),
	.w3(32'h3c3ea80f),
	.w4(32'hbd25af04),
	.w5(32'h3d215460),
	.w6(32'hbcc0241f),
	.w7(32'h3ba3b7a8),
	.w8(32'hbda2c90b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd023b8f),
	.w1(32'hbc9f2855),
	.w2(32'hbcaecffb),
	.w3(32'h3ce6973c),
	.w4(32'hbc046445),
	.w5(32'h391b8fee),
	.w6(32'hbb844d8b),
	.w7(32'hbc28925c),
	.w8(32'hbc4067f7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c865992),
	.w1(32'h3b261737),
	.w2(32'hbb03a88e),
	.w3(32'hbc41e6a1),
	.w4(32'hbb0ac201),
	.w5(32'h3b0d1140),
	.w6(32'hbd0fcd85),
	.w7(32'hbd87a51a),
	.w8(32'hbc35bf88),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78d7ee),
	.w1(32'h3a796fa6),
	.w2(32'hbc77c753),
	.w3(32'h3d13bb6a),
	.w4(32'hb9ca3c3f),
	.w5(32'h3bfaa336),
	.w6(32'hbc2c5c9b),
	.w7(32'hbbea38e3),
	.w8(32'hb9e17dac),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d33145d),
	.w1(32'hbd792620),
	.w2(32'hbdb746ca),
	.w3(32'h3cd6b2d1),
	.w4(32'h3b227aa1),
	.w5(32'hbdc1dabb),
	.w6(32'h3ca68fb7),
	.w7(32'hbd7d2b7d),
	.w8(32'hbb008005),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1454f6),
	.w1(32'hbd805de5),
	.w2(32'hbc344e09),
	.w3(32'h3be2d312),
	.w4(32'hbcb7ed59),
	.w5(32'hbc27db28),
	.w6(32'h3c9f2eca),
	.w7(32'hbc196dfc),
	.w8(32'h3b20ccc6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31f8c7),
	.w1(32'h3b85c7dd),
	.w2(32'hbd9f98ec),
	.w3(32'hbc1e8216),
	.w4(32'h3befbcad),
	.w5(32'hbd2aa5a7),
	.w6(32'h3c9d1f49),
	.w7(32'hbc11cc75),
	.w8(32'hbcdb2151),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd21120c),
	.w1(32'hbc23ff34),
	.w2(32'hbc32fdb8),
	.w3(32'hbcec7cee),
	.w4(32'h3d5b3c0b),
	.w5(32'hbc477631),
	.w6(32'hba261b57),
	.w7(32'h3c0ccbb2),
	.w8(32'h3c04a7a2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd219898),
	.w1(32'h3b8907ab),
	.w2(32'hbc6d98ba),
	.w3(32'hbd7b4889),
	.w4(32'h3c2e4351),
	.w5(32'hbc36731c),
	.w6(32'h3c83efd0),
	.w7(32'h3c6dc6cf),
	.w8(32'h3bf69ef2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e81df),
	.w1(32'hbbeab3e9),
	.w2(32'hbcc8fa86),
	.w3(32'h3ca03788),
	.w4(32'h3b834c84),
	.w5(32'h3c060a1c),
	.w6(32'hbb1a0586),
	.w7(32'h3c17ea9f),
	.w8(32'hbc48cd7f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c2d26),
	.w1(32'hbc8ec8df),
	.w2(32'h3c069afc),
	.w3(32'hbbec7d09),
	.w4(32'hbd133a45),
	.w5(32'hbb2ca04e),
	.w6(32'h3c195e3c),
	.w7(32'hbc01f565),
	.w8(32'h3bc91189),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5236a8),
	.w1(32'hbc547b70),
	.w2(32'hbd34eef8),
	.w3(32'hbb940aee),
	.w4(32'h3c3b988a),
	.w5(32'hbbde2294),
	.w6(32'hbd5de884),
	.w7(32'hbcb6556a),
	.w8(32'hbcfd1f6b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule