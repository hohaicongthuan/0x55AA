module layer_10_featuremap_424(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3141c),
	.w1(32'hbb978a6b),
	.w2(32'h3abc40ac),
	.w3(32'hbbafcf18),
	.w4(32'hbbe1f426),
	.w5(32'h3ae2d6db),
	.w6(32'h3bb946c6),
	.w7(32'hbbf35fb2),
	.w8(32'h3b2e3c8d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d20b4),
	.w1(32'hb9cd0b0f),
	.w2(32'hba2e7f67),
	.w3(32'hbb8333b6),
	.w4(32'hba64dc53),
	.w5(32'hbb1e12d5),
	.w6(32'hbb2e8b3a),
	.w7(32'hbb098fe4),
	.w8(32'hbb84631b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba183184),
	.w1(32'h3a9f4f9c),
	.w2(32'h39585f9e),
	.w3(32'hbae79d16),
	.w4(32'hba558d4d),
	.w5(32'hbb090c91),
	.w6(32'hbad2504b),
	.w7(32'hbc080914),
	.w8(32'hbb990824),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40b910),
	.w1(32'h3b9873a6),
	.w2(32'h3c2092da),
	.w3(32'h39f012a8),
	.w4(32'h3a35f632),
	.w5(32'h3cc4d7cf),
	.w6(32'hbb177e9a),
	.w7(32'h3b81b361),
	.w8(32'h3c4f59c6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73952e),
	.w1(32'hba852f4a),
	.w2(32'hbb311b9c),
	.w3(32'h3c422718),
	.w4(32'hbb1b9b98),
	.w5(32'hbbe2d509),
	.w6(32'h39608458),
	.w7(32'hbacdea95),
	.w8(32'hbbfc1de1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbf899),
	.w1(32'h3ac96995),
	.w2(32'h3af0a6b6),
	.w3(32'hbbc68eb3),
	.w4(32'h3bc5fec3),
	.w5(32'h3b32c21b),
	.w6(32'hbc232e03),
	.w7(32'h3aa5b090),
	.w8(32'hbb95caa2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08a94f),
	.w1(32'hbba46c70),
	.w2(32'hbb93a76f),
	.w3(32'hbaceb10b),
	.w4(32'hbbce4d9b),
	.w5(32'hbbf04f71),
	.w6(32'hbb832304),
	.w7(32'hbba8e612),
	.w8(32'h3b2a4fb5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffa795),
	.w1(32'hbbfe84a3),
	.w2(32'hba2c38c6),
	.w3(32'hbb103453),
	.w4(32'hbba992cf),
	.w5(32'h3c5dfa2a),
	.w6(32'h3b136332),
	.w7(32'hbb34670f),
	.w8(32'h3bfded58),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25feb6),
	.w1(32'h38d8920a),
	.w2(32'h39d2c710),
	.w3(32'h3b99a71e),
	.w4(32'h3ba122db),
	.w5(32'h3a277a5a),
	.w6(32'hbbabe082),
	.w7(32'h3b61f8ae),
	.w8(32'hbb0bb20e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c088796),
	.w1(32'h39bd12d9),
	.w2(32'hbae560dd),
	.w3(32'h3ab176e0),
	.w4(32'h389d307e),
	.w5(32'hb9e0d9e3),
	.w6(32'h3b8e6313),
	.w7(32'h3ac3abd4),
	.w8(32'h3a1b0511),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96371e5),
	.w1(32'hbab1cf04),
	.w2(32'hbb5dc670),
	.w3(32'hbb992f0b),
	.w4(32'h3af54338),
	.w5(32'h3a7e35c5),
	.w6(32'hb9ac38a4),
	.w7(32'hbab6b798),
	.w8(32'h3aeaf752),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08c808),
	.w1(32'h3b9337dd),
	.w2(32'hbc04e39b),
	.w3(32'h3a910e42),
	.w4(32'h3bac288c),
	.w5(32'hbc24c0a5),
	.w6(32'h3ae02e5f),
	.w7(32'hbaef59bc),
	.w8(32'hbc7c95b7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfba36),
	.w1(32'h3c213857),
	.w2(32'h3ba4fd04),
	.w3(32'h3b6e9b7b),
	.w4(32'h3b8136ab),
	.w5(32'h3bc1fca0),
	.w6(32'hb7eefec8),
	.w7(32'h3a1f0e96),
	.w8(32'h396682c9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944f272),
	.w1(32'hbabb36c4),
	.w2(32'h3b88b594),
	.w3(32'hbb8ee65a),
	.w4(32'h3b708747),
	.w5(32'h3b0f3968),
	.w6(32'hba125caa),
	.w7(32'h3b0c0ff5),
	.w8(32'h3ae08439),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2c010),
	.w1(32'hbaf4bc4c),
	.w2(32'hbac8b8f0),
	.w3(32'hb9bf38cf),
	.w4(32'h3b095bb0),
	.w5(32'hbb2998e6),
	.w6(32'h3b155355),
	.w7(32'h3ad8bc3d),
	.w8(32'hbacd3c84),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7716),
	.w1(32'hbb07d282),
	.w2(32'h3a6ef60c),
	.w3(32'hbb4230c6),
	.w4(32'h3b3c76bb),
	.w5(32'h3a76ed8c),
	.w6(32'hbb54cff0),
	.w7(32'hb8b3eb5a),
	.w8(32'h3a466951),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6689e1),
	.w1(32'h3a41f20c),
	.w2(32'hbb9182cc),
	.w3(32'h3a113eb1),
	.w4(32'h3b8352a5),
	.w5(32'hbb498c1d),
	.w6(32'hbb0bc30c),
	.w7(32'h3b1976a1),
	.w8(32'hba944804),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaada755),
	.w1(32'hbb674c90),
	.w2(32'h3bd5e321),
	.w3(32'hba39c397),
	.w4(32'hba8c9a83),
	.w5(32'h3c61af04),
	.w6(32'h39d57db9),
	.w7(32'hbc0b864b),
	.w8(32'h3c4ccd82),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432f43),
	.w1(32'hbb2799ec),
	.w2(32'hbbcc3e2f),
	.w3(32'h3b54dedd),
	.w4(32'hbbeff416),
	.w5(32'hbbcf894d),
	.w6(32'h38b83faf),
	.w7(32'hbbabf766),
	.w8(32'hbc2d105a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d5d9d),
	.w1(32'h3b515aa7),
	.w2(32'hbc34b129),
	.w3(32'hbb6c3cfe),
	.w4(32'h3bd3ccc3),
	.w5(32'hbbd48d18),
	.w6(32'hbb24e32f),
	.w7(32'hbaa81ca8),
	.w8(32'h3c371936),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525bf3),
	.w1(32'hbaba5784),
	.w2(32'hbb21dd44),
	.w3(32'h3aef2421),
	.w4(32'hbb86c279),
	.w5(32'hbb4b4958),
	.w6(32'hbb6c98bc),
	.w7(32'hbb50742f),
	.w8(32'hbc27a6a2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa906eb),
	.w1(32'hbb320da7),
	.w2(32'h3bc5f178),
	.w3(32'hb99c3ce1),
	.w4(32'hbb9688e3),
	.w5(32'h3a4023f7),
	.w6(32'h3872fb4a),
	.w7(32'hbb441944),
	.w8(32'h3b56a079),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79aefc),
	.w1(32'h3a71a7ad),
	.w2(32'hbc79f61a),
	.w3(32'hbbf8f66a),
	.w4(32'hb8ae330d),
	.w5(32'hbc81e2ef),
	.w6(32'hbb58dcf2),
	.w7(32'h3b596719),
	.w8(32'hbc7a61be),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95ebe0),
	.w1(32'hba987c19),
	.w2(32'h3b8be11f),
	.w3(32'hbc35951a),
	.w4(32'hbb9366cb),
	.w5(32'hbb26b43d),
	.w6(32'hbb4b1b03),
	.w7(32'hbbea3893),
	.w8(32'hbb4ea113),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e43d),
	.w1(32'h3c21dde9),
	.w2(32'h3b7a8b26),
	.w3(32'hbb8bc8ec),
	.w4(32'h3bad8ecf),
	.w5(32'h3c8d1897),
	.w6(32'hbb5f9269),
	.w7(32'h3bb7687f),
	.w8(32'h3b95d580),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61764f),
	.w1(32'hbbc592af),
	.w2(32'hbbd2d548),
	.w3(32'hbbb30294),
	.w4(32'hbc0ca5d8),
	.w5(32'hbbf1695d),
	.w6(32'hbbaad91f),
	.w7(32'hbb9b7757),
	.w8(32'hbbcbacb1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c26f8),
	.w1(32'h3b8a5444),
	.w2(32'hb9b283a7),
	.w3(32'hbbb12963),
	.w4(32'h3bba1080),
	.w5(32'h3a421046),
	.w6(32'hbbf79352),
	.w7(32'h3bf02d23),
	.w8(32'hbb3577f7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb599b23),
	.w1(32'h3a8588f7),
	.w2(32'h3b9dedc8),
	.w3(32'h3aafd549),
	.w4(32'hba907f6f),
	.w5(32'h3bec2eb0),
	.w6(32'h3b8b013f),
	.w7(32'hba4f0c6b),
	.w8(32'h3b3ef6ef),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85dab28),
	.w1(32'h3c15c904),
	.w2(32'hbc5e730d),
	.w3(32'h39ad3ab1),
	.w4(32'h3b3adcaf),
	.w5(32'hbc8199cb),
	.w6(32'h3af47f68),
	.w7(32'h3b27c1d2),
	.w8(32'hbbd4b6d3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8606fc),
	.w1(32'h3afba219),
	.w2(32'hbc23725a),
	.w3(32'hbb56e6f2),
	.w4(32'h3b1dd6c9),
	.w5(32'hbc395eb0),
	.w6(32'h3c86f92a),
	.w7(32'hbba161f2),
	.w8(32'hbc7f16c8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2199),
	.w1(32'hbbc07026),
	.w2(32'hbc09ad6a),
	.w3(32'hba5ab0f5),
	.w4(32'h3a52b8eb),
	.w5(32'hbbe21e22),
	.w6(32'hbb91e07b),
	.w7(32'hbbbd138a),
	.w8(32'hbb2c3a0a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d67e8),
	.w1(32'h3baf9ead),
	.w2(32'hba85e57d),
	.w3(32'hbb8e278f),
	.w4(32'h3c02e463),
	.w5(32'h37e981f4),
	.w6(32'hbb1ec141),
	.w7(32'h3bc13f11),
	.w8(32'h3b523b0e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d4e39),
	.w1(32'h3b3c712c),
	.w2(32'h3c092118),
	.w3(32'h3b01cf7a),
	.w4(32'h3b842f06),
	.w5(32'hbb498594),
	.w6(32'h3ba0064f),
	.w7(32'hbaef31f6),
	.w8(32'hba05f6a2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5adc21),
	.w1(32'hbb111e3f),
	.w2(32'hbbb540ab),
	.w3(32'hbb453ed8),
	.w4(32'hbb45cbad),
	.w5(32'hbbb733f1),
	.w6(32'h3b89eef8),
	.w7(32'hbbb2112d),
	.w8(32'hbb016b3c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0235),
	.w1(32'hbb8323ca),
	.w2(32'h3a590eb5),
	.w3(32'hbc0b6898),
	.w4(32'hbb855b6c),
	.w5(32'h3c92f77c),
	.w6(32'hbaa3cf2a),
	.w7(32'hbc1c9715),
	.w8(32'h3ba385c3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc6d21),
	.w1(32'h3b85be44),
	.w2(32'hbafb6883),
	.w3(32'h3ba1f909),
	.w4(32'hba07dd0b),
	.w5(32'hba721b5b),
	.w6(32'hb76858ac),
	.w7(32'hbb20ba2b),
	.w8(32'hba9f0ac8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947297),
	.w1(32'hbc08d064),
	.w2(32'h3b8b77e1),
	.w3(32'hba717d7f),
	.w4(32'hbc10103f),
	.w5(32'h3b2a8e6c),
	.w6(32'hbb558991),
	.w7(32'hbba0937c),
	.w8(32'h3b3894a1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e0ba2),
	.w1(32'h3b7817d9),
	.w2(32'h37f4d907),
	.w3(32'h3b895b27),
	.w4(32'h3bab4875),
	.w5(32'h3b28a0a6),
	.w6(32'h3b3ccfbb),
	.w7(32'h3b485ec6),
	.w8(32'h3b92542e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b367914),
	.w1(32'hbbc5b168),
	.w2(32'h3b664dfc),
	.w3(32'h3bbcb716),
	.w4(32'hba1cf7e7),
	.w5(32'h3c34ccde),
	.w6(32'h3b657028),
	.w7(32'h3b775b6c),
	.w8(32'h3b18267e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a3ef2),
	.w1(32'hbb37d19a),
	.w2(32'hb8a7b584),
	.w3(32'h39867074),
	.w4(32'hbb484235),
	.w5(32'h3c38de53),
	.w6(32'hbbcb012a),
	.w7(32'hb9b7644c),
	.w8(32'h3af2ee15),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b955fcd),
	.w1(32'h391abbf1),
	.w2(32'h3b1495fb),
	.w3(32'h3a111106),
	.w4(32'h3b1a8cd4),
	.w5(32'h3a26a38d),
	.w6(32'h3a81fb93),
	.w7(32'hb93780e0),
	.w8(32'hbac2b178),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b568d36),
	.w1(32'hbb54f875),
	.w2(32'hba956578),
	.w3(32'h3bab31c2),
	.w4(32'hbb145ed4),
	.w5(32'h3ad87eea),
	.w6(32'h3b53fe53),
	.w7(32'hbb1cc742),
	.w8(32'hbbac8dfc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901124e),
	.w1(32'hbab5d0ee),
	.w2(32'h3b1d2a61),
	.w3(32'hba718b3a),
	.w4(32'hbbafdc80),
	.w5(32'h3c20aa35),
	.w6(32'hbb594527),
	.w7(32'hbbb70bda),
	.w8(32'hbb696be5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3411c0),
	.w1(32'hbbc2e112),
	.w2(32'h3cc36a01),
	.w3(32'h3b6cf9e3),
	.w4(32'hbb842d28),
	.w5(32'h3d39b73c),
	.w6(32'h3b49d5e2),
	.w7(32'h3a217662),
	.w8(32'h3d2595ca),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c738e1b),
	.w1(32'h3b393f21),
	.w2(32'hbba25b39),
	.w3(32'h3c62e43d),
	.w4(32'h3b000e75),
	.w5(32'hbb8b5b87),
	.w6(32'h3be1ad62),
	.w7(32'h3a995c2f),
	.w8(32'hbb7940a7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75f6ad),
	.w1(32'hbb76bd13),
	.w2(32'hbaa89f01),
	.w3(32'h3b9cccae),
	.w4(32'h37e78bde),
	.w5(32'h39b333e5),
	.w6(32'h3bd74996),
	.w7(32'hbada368f),
	.w8(32'hbb86ff12),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b0de2),
	.w1(32'hbb987028),
	.w2(32'hbc0060f1),
	.w3(32'h3afb743c),
	.w4(32'hba1659c4),
	.w5(32'hbc9588e0),
	.w6(32'hbab87914),
	.w7(32'hbad86402),
	.w8(32'hbc4dc042),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50d9b4),
	.w1(32'h3bb573f2),
	.w2(32'h3b6c50d4),
	.w3(32'hbbdd55d8),
	.w4(32'h3b86599a),
	.w5(32'h3b6dc01c),
	.w6(32'hbb416876),
	.w7(32'h3b11b818),
	.w8(32'h3aa4b623),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf631c),
	.w1(32'h3b84dc04),
	.w2(32'h3b9f5e65),
	.w3(32'hbb98afb3),
	.w4(32'h3bacd692),
	.w5(32'h3b2d5993),
	.w6(32'hbb3cdd89),
	.w7(32'h3bcf401c),
	.w8(32'h3b4f3d53),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a186),
	.w1(32'hbc2ff84a),
	.w2(32'hbc078809),
	.w3(32'h3b1ab697),
	.w4(32'hbb67523f),
	.w5(32'hbc68a44a),
	.w6(32'h3b915b66),
	.w7(32'hbbb3d5ab),
	.w8(32'hbc51108d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae43a79),
	.w1(32'h3b99847d),
	.w2(32'hbbf4917b),
	.w3(32'h3af6704d),
	.w4(32'h3b15d946),
	.w5(32'hbc26b6eb),
	.w6(32'h3a9f9485),
	.w7(32'h3b8698fa),
	.w8(32'hbc349963),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dbbbb),
	.w1(32'h3b850ddf),
	.w2(32'h3b0adbb2),
	.w3(32'hbbcda452),
	.w4(32'h3c096582),
	.w5(32'h3a10dbb1),
	.w6(32'hbbaa3ed8),
	.w7(32'h3b9d52dc),
	.w8(32'h3af4df77),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb151b6c),
	.w1(32'hbb7d8db6),
	.w2(32'hbb09a140),
	.w3(32'h3ad21cda),
	.w4(32'hb90634d6),
	.w5(32'h3ba94c4b),
	.w6(32'hba4553f2),
	.w7(32'hba8dd0a2),
	.w8(32'hbb3c7a54),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4af9),
	.w1(32'hbadf39fa),
	.w2(32'h3b83d0c8),
	.w3(32'hbaad7eb3),
	.w4(32'hb985b7c3),
	.w5(32'h3c0f8364),
	.w6(32'hbaf3e4ec),
	.w7(32'hbbb8213f),
	.w8(32'hb9a3bd49),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77b3a),
	.w1(32'h393c1f33),
	.w2(32'hbb517f1f),
	.w3(32'hbb444f8f),
	.w4(32'hbaf9ce42),
	.w5(32'hb8d69931),
	.w6(32'hbb3013ba),
	.w7(32'hbaf664cb),
	.w8(32'hbb79e811),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc009c),
	.w1(32'h3b4ef354),
	.w2(32'h3c27d79e),
	.w3(32'h3b0cf026),
	.w4(32'hbb4adedc),
	.w5(32'h3b70baab),
	.w6(32'hbaff1566),
	.w7(32'hbb8d7e72),
	.w8(32'h3a1f8787),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fcfe6),
	.w1(32'hbad3c76a),
	.w2(32'hbbb2db49),
	.w3(32'hba80f196),
	.w4(32'hba64307c),
	.w5(32'hbbb372f8),
	.w6(32'h3b3ea7e4),
	.w7(32'hbaf2e6c8),
	.w8(32'hbc05cb62),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9b8e),
	.w1(32'hba0f12e3),
	.w2(32'hba486513),
	.w3(32'hbc155970),
	.w4(32'hbb4eb699),
	.w5(32'hbbc1a209),
	.w6(32'hbbee6cc3),
	.w7(32'hb720f32a),
	.w8(32'hbc134433),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52f422),
	.w1(32'hbbcdabdc),
	.w2(32'h3a36a476),
	.w3(32'h3ba8f91f),
	.w4(32'hbc4c4422),
	.w5(32'hbaab72e4),
	.w6(32'h3ac91afa),
	.w7(32'hbbb0ff18),
	.w8(32'hbb12fb7d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147162),
	.w1(32'hbb1b480a),
	.w2(32'hbc3bd336),
	.w3(32'hbbac96ab),
	.w4(32'hb9dbbd7a),
	.w5(32'hbc4363d7),
	.w6(32'h39339778),
	.w7(32'h3b890dae),
	.w8(32'hbc670687),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba648171),
	.w1(32'hbb83a08a),
	.w2(32'hbb95d340),
	.w3(32'hbc6b9db6),
	.w4(32'h3aadf44e),
	.w5(32'hbc0eaa19),
	.w6(32'hbc93ef06),
	.w7(32'h3a4ea3f0),
	.w8(32'hbb6f067f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e2308),
	.w1(32'h399d130e),
	.w2(32'h3adca960),
	.w3(32'hbbaa1959),
	.w4(32'hbaa6ce81),
	.w5(32'h3b3864ee),
	.w6(32'hbab44730),
	.w7(32'hbae7e495),
	.w8(32'h3b3a8560),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9abbad),
	.w1(32'hba9401a6),
	.w2(32'h3c1048a1),
	.w3(32'h3b10fb22),
	.w4(32'hbc0ef9a8),
	.w5(32'h3c8648a9),
	.w6(32'h3b9f48d6),
	.w7(32'hbbdab67f),
	.w8(32'h3c16909f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb973ec),
	.w1(32'hbb0a0c1f),
	.w2(32'hbbece9b0),
	.w3(32'h3b951fd9),
	.w4(32'hba4be8e4),
	.w5(32'hbc2f1ed8),
	.w6(32'h3b230f75),
	.w7(32'hbb93639b),
	.w8(32'hbc52f641),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5420b),
	.w1(32'hbb89c6f6),
	.w2(32'h3a4893e9),
	.w3(32'hbb8072f1),
	.w4(32'hbb539982),
	.w5(32'h3b5ee880),
	.w6(32'hbbddc8f8),
	.w7(32'hbb8b3f53),
	.w8(32'h3b8d22a3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d3699),
	.w1(32'hbc10130a),
	.w2(32'h3afcad6b),
	.w3(32'hbb6045d2),
	.w4(32'hbc1c4c54),
	.w5(32'h3c07f331),
	.w6(32'hbba05fcc),
	.w7(32'hbb520785),
	.w8(32'h3b5064d4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b5e62),
	.w1(32'hbb53c20c),
	.w2(32'hbbdaa939),
	.w3(32'h3c09b92f),
	.w4(32'hbba4ad6c),
	.w5(32'hbbac78f9),
	.w6(32'h3ba8fb10),
	.w7(32'hbb96f06b),
	.w8(32'hbb212f62),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688463),
	.w1(32'hbb4ce25c),
	.w2(32'hbc149140),
	.w3(32'hbb93474f),
	.w4(32'hbc16739f),
	.w5(32'hbc184840),
	.w6(32'hbaae703a),
	.w7(32'hbc62de5a),
	.w8(32'hbbf37723),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a0ed1),
	.w1(32'h3ba90875),
	.w2(32'h3b6e9836),
	.w3(32'hbb722bae),
	.w4(32'h3a95887b),
	.w5(32'h3b0156a3),
	.w6(32'hbb82ac19),
	.w7(32'h3a214093),
	.w8(32'h3bb2164a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cb36f),
	.w1(32'h3b375fc6),
	.w2(32'h3bd710ec),
	.w3(32'hb9fab914),
	.w4(32'h3a835a98),
	.w5(32'hbaf53101),
	.w6(32'h3bfff440),
	.w7(32'hbb21a067),
	.w8(32'hbb214a97),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32cf8e),
	.w1(32'hbb6a96a3),
	.w2(32'h3bf44fc6),
	.w3(32'h3c075e51),
	.w4(32'h3b74e2f6),
	.w5(32'h3bc7ae56),
	.w6(32'h3b8dba7d),
	.w7(32'hbb5676c6),
	.w8(32'hbc24d528),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baae895),
	.w1(32'h3b6ec264),
	.w2(32'h395c0206),
	.w3(32'hbb2e8d93),
	.w4(32'h3be6349c),
	.w5(32'h3cbb58dc),
	.w6(32'hbb8875bc),
	.w7(32'hba7289c4),
	.w8(32'h3b0174aa),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12400),
	.w1(32'h3c1bfc8f),
	.w2(32'h3b48c2ab),
	.w3(32'h3aa45037),
	.w4(32'h3b5c31a5),
	.w5(32'hbbf529aa),
	.w6(32'h3b81bce8),
	.w7(32'h3b2440f4),
	.w8(32'h3a1d82db),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be677e4),
	.w1(32'h3abea039),
	.w2(32'hbb888ac9),
	.w3(32'h3bba6323),
	.w4(32'hbc28b4b3),
	.w5(32'hbcc7dc1b),
	.w6(32'h394630d3),
	.w7(32'h3aa6e510),
	.w8(32'h3ce70a75),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3bfe),
	.w1(32'hba0e0d18),
	.w2(32'hbbed314a),
	.w3(32'h3aad5994),
	.w4(32'h3b088b62),
	.w5(32'h3c05e4fd),
	.w6(32'h3ca3aaee),
	.w7(32'h3bec23b3),
	.w8(32'h3bdc5b17),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb461a7c),
	.w1(32'hbb298c43),
	.w2(32'h3ad1c73e),
	.w3(32'h3a8ff697),
	.w4(32'hbc49e35d),
	.w5(32'hbc5b2096),
	.w6(32'h3ac20a82),
	.w7(32'h3b0f0cba),
	.w8(32'h3d2ee500),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88ab40),
	.w1(32'h3afe7e00),
	.w2(32'hbae36f60),
	.w3(32'hbb6dd90e),
	.w4(32'hbb88b304),
	.w5(32'hba6c7438),
	.w6(32'h3c9405e4),
	.w7(32'hb9152a74),
	.w8(32'hbb924b6f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb682bd8),
	.w1(32'h3b699b54),
	.w2(32'h3ba1f816),
	.w3(32'hbba8a627),
	.w4(32'h3b90d29e),
	.w5(32'hbbd96d59),
	.w6(32'hbbf23f2e),
	.w7(32'hbb1fc704),
	.w8(32'h3b8475bb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ffb1),
	.w1(32'hbbe455b6),
	.w2(32'hbb0af6db),
	.w3(32'hbc7fcf01),
	.w4(32'hbc18ea78),
	.w5(32'h3ba521ae),
	.w6(32'hbbac712d),
	.w7(32'hbc16e394),
	.w8(32'hbc2a53fa),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01ac43),
	.w1(32'h3b4af4bb),
	.w2(32'hbb0714f9),
	.w3(32'h3c5354b1),
	.w4(32'hbaafe0c5),
	.w5(32'hba03b8e5),
	.w6(32'hbb43ffd5),
	.w7(32'hbab01a04),
	.w8(32'h3baaa225),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8946fb),
	.w1(32'h3c8f94e7),
	.w2(32'h3c2c047e),
	.w3(32'h3a8a601a),
	.w4(32'h3c8754fa),
	.w5(32'h3b9c5b5b),
	.w6(32'h38be7ec4),
	.w7(32'h3c3af87a),
	.w8(32'hbbe40110),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c354f54),
	.w1(32'hbaaaaef4),
	.w2(32'hbb0020fd),
	.w3(32'h3bd10797),
	.w4(32'h3b970d6c),
	.w5(32'h39d16a54),
	.w6(32'h3a5f8242),
	.w7(32'h3b32f7a5),
	.w8(32'h3a2479b1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70826e),
	.w1(32'h3aa8e2e8),
	.w2(32'h3ca0880c),
	.w3(32'hbbafbb40),
	.w4(32'h3c113112),
	.w5(32'h3d2045ba),
	.w6(32'h3b4c0cb9),
	.w7(32'hbc3bb1ae),
	.w8(32'hbc98cf19),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff725),
	.w1(32'hb9ab0380),
	.w2(32'hbb2fb06a),
	.w3(32'hbc20421d),
	.w4(32'hbaa0d62a),
	.w5(32'hba862a16),
	.w6(32'hbca20529),
	.w7(32'hba62cb5e),
	.w8(32'hbb00c6d4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6c763),
	.w1(32'h3b212411),
	.w2(32'hbbcdca73),
	.w3(32'hbc217750),
	.w4(32'h3b1d73e4),
	.w5(32'h3bf59a01),
	.w6(32'h3bbdb9b2),
	.w7(32'h388fd943),
	.w8(32'hbba313d0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc361),
	.w1(32'h3bddde5d),
	.w2(32'h3ba517e1),
	.w3(32'h3c0459e3),
	.w4(32'h3b265993),
	.w5(32'h3b05b909),
	.w6(32'hba3aff14),
	.w7(32'h3b01e269),
	.w8(32'h3bab1122),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe1005),
	.w1(32'h3b0c8ef2),
	.w2(32'hbb64180e),
	.w3(32'h3b4158cb),
	.w4(32'h3a8e759f),
	.w5(32'h3b93bd84),
	.w6(32'h3bb18d04),
	.w7(32'hba89e22f),
	.w8(32'h3a5290da),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfffd20),
	.w1(32'hbbcb68a9),
	.w2(32'hbb90b275),
	.w3(32'h3b86732f),
	.w4(32'hbb705858),
	.w5(32'h3c6aafcc),
	.w6(32'hbbf44542),
	.w7(32'hbbafb9f7),
	.w8(32'h3b833998),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b7978),
	.w1(32'hbbed6825),
	.w2(32'hbc4eefb5),
	.w3(32'h3b2c4de7),
	.w4(32'hbc20107a),
	.w5(32'h3b13df09),
	.w6(32'hbb670790),
	.w7(32'hbc11099a),
	.w8(32'hbc64fdbe),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c9b2),
	.w1(32'hbbdddf92),
	.w2(32'h3b178322),
	.w3(32'hbbcb8f49),
	.w4(32'hbc2ca44c),
	.w5(32'hbc0504cc),
	.w6(32'hbc1c4300),
	.w7(32'hbb7a3362),
	.w8(32'h3ba87838),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc0931),
	.w1(32'hbb4287ec),
	.w2(32'hbaf7ea14),
	.w3(32'hbbdebfb7),
	.w4(32'h3bdc9ee4),
	.w5(32'hbb813eb8),
	.w6(32'hba960277),
	.w7(32'hbb970392),
	.w8(32'hbc46efe1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242070),
	.w1(32'hbbe9838d),
	.w2(32'hbc429f01),
	.w3(32'hbbe7db74),
	.w4(32'hba0b08f9),
	.w5(32'hbbf909b5),
	.w6(32'hbb0c80cb),
	.w7(32'h3981c717),
	.w8(32'h3b0e8bc9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc3db7),
	.w1(32'hbb54b496),
	.w2(32'hbb805b55),
	.w3(32'hbc0b380e),
	.w4(32'hb972e0a2),
	.w5(32'h3c764357),
	.w6(32'hbbaf6e5f),
	.w7(32'hbbf11a42),
	.w8(32'hbc2ac5fc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3da18a),
	.w1(32'hbc541bb0),
	.w2(32'hbcd4fb13),
	.w3(32'h3ba3ddb7),
	.w4(32'hbb4f44b9),
	.w5(32'hbc66e717),
	.w6(32'hbb22d96d),
	.w7(32'h3bd11cd3),
	.w8(32'h3d0857fc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99fb63),
	.w1(32'h3b2f14c3),
	.w2(32'hbbbe4317),
	.w3(32'hbc7b4ade),
	.w4(32'h3b4d4323),
	.w5(32'hbb125fee),
	.w6(32'h3bc7f9d4),
	.w7(32'h3b3817b8),
	.w8(32'h3b878c61),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58e809),
	.w1(32'h3c1e85b2),
	.w2(32'hbb0e4911),
	.w3(32'hbb3ea55b),
	.w4(32'h37cdab9a),
	.w5(32'hbc7d739c),
	.w6(32'h3ad14ee3),
	.w7(32'h3c1870fd),
	.w8(32'hbbebb78e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f35fa),
	.w1(32'h3b2ebfe0),
	.w2(32'hbab6ead1),
	.w3(32'h3ac17535),
	.w4(32'hbba15738),
	.w5(32'hbc888ccd),
	.w6(32'hbbca9aec),
	.w7(32'hbafec5c2),
	.w8(32'hbae554e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb22b7e),
	.w1(32'hbbd77c68),
	.w2(32'h3ad01b20),
	.w3(32'h3bafdb4a),
	.w4(32'h3a18e8c4),
	.w5(32'hbb22c5be),
	.w6(32'h3b3a8423),
	.w7(32'hbb97f927),
	.w8(32'h3b99f655),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5368f4),
	.w1(32'h3ab468ea),
	.w2(32'h3b7afa2e),
	.w3(32'hbaac5fb6),
	.w4(32'hbb260967),
	.w5(32'hbc030474),
	.w6(32'hbb1c5c03),
	.w7(32'h3b3d0eae),
	.w8(32'h3c1ad34f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92d4f7),
	.w1(32'h3b63e4d0),
	.w2(32'h3b4839e3),
	.w3(32'hba7d0eb8),
	.w4(32'hbbdbcb27),
	.w5(32'hbc306bb9),
	.w6(32'h3b9df366),
	.w7(32'hbb766777),
	.w8(32'h3bfc2305),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba20b0a),
	.w1(32'hbb9721ff),
	.w2(32'hbb12c9c4),
	.w3(32'hba9bb8b1),
	.w4(32'hbb93af21),
	.w5(32'hbc357cff),
	.w6(32'h3b8158c6),
	.w7(32'hb96d201c),
	.w8(32'h3cb02d43),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfcf7f),
	.w1(32'hba23fe90),
	.w2(32'hbbec18f2),
	.w3(32'h3b82c6bf),
	.w4(32'hbb7941b6),
	.w5(32'hbb91a050),
	.w6(32'h3c49e047),
	.w7(32'h3b7732a1),
	.w8(32'hbc04064d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57ddf8),
	.w1(32'hbc574f61),
	.w2(32'h3b2d7b65),
	.w3(32'hbb8ce59e),
	.w4(32'hbb6df466),
	.w5(32'h3d645395),
	.w6(32'hbbe8936d),
	.w7(32'hbc1ff6c3),
	.w8(32'hbc52bae9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990678b),
	.w1(32'h3beea93e),
	.w2(32'hbc4fefaf),
	.w3(32'hbc1ee51e),
	.w4(32'h3b7d4bb9),
	.w5(32'h3badcb81),
	.w6(32'hbb7504da),
	.w7(32'h3c849151),
	.w8(32'hbc86d381),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcedd1db),
	.w1(32'h3a6fe69e),
	.w2(32'h3ba0f3ce),
	.w3(32'h3ccc84cf),
	.w4(32'hba15ad28),
	.w5(32'h3c650c4c),
	.w6(32'hbca36ae3),
	.w7(32'hbb30112c),
	.w8(32'hbbe32066),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f207bb),
	.w1(32'h3a9bb85c),
	.w2(32'hbbe4db8c),
	.w3(32'hbaaf61c5),
	.w4(32'hbbedf440),
	.w5(32'hbbce018d),
	.w6(32'h3b05f673),
	.w7(32'h3ba0f4aa),
	.w8(32'h3c3222e3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8817),
	.w1(32'h3bb1ebd9),
	.w2(32'h3c82e71c),
	.w3(32'h3ba88b57),
	.w4(32'h3bd88529),
	.w5(32'hba5a2fd1),
	.w6(32'h3b3a9ec8),
	.w7(32'hbbe18593),
	.w8(32'hbac54f6e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbca39b),
	.w1(32'hbbb0d373),
	.w2(32'h3a99817a),
	.w3(32'hbb20deea),
	.w4(32'h3b95d1f3),
	.w5(32'h3ba95934),
	.w6(32'h3b8bc0b2),
	.w7(32'h3b46dd77),
	.w8(32'hba40df8f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb366ba3),
	.w1(32'h3ab60bde),
	.w2(32'h3b034f30),
	.w3(32'hb9e55856),
	.w4(32'hbb1f2f53),
	.w5(32'h3a997e5d),
	.w6(32'hbab87dc6),
	.w7(32'h3b741b4a),
	.w8(32'h3bbc5679),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c1569),
	.w1(32'hbb587445),
	.w2(32'hbba715d0),
	.w3(32'hbb98f32e),
	.w4(32'hbb7a1221),
	.w5(32'hbc00cbff),
	.w6(32'h3bf5c35c),
	.w7(32'hbc105ccd),
	.w8(32'h3a641203),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc155133),
	.w1(32'hbbbd58ee),
	.w2(32'h3c20f1f9),
	.w3(32'hbc85be43),
	.w4(32'hbb795b1a),
	.w5(32'hbb9e0f70),
	.w6(32'hbbab50ab),
	.w7(32'hbb19dcc5),
	.w8(32'hbac52262),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db26d),
	.w1(32'h3bfad6ff),
	.w2(32'h3ba5e856),
	.w3(32'hbad8ac5b),
	.w4(32'h3accc982),
	.w5(32'hbbfd5bfc),
	.w6(32'h3a8bdc5b),
	.w7(32'h3b968fc3),
	.w8(32'hbb34297d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ec67e),
	.w1(32'h3aad3b86),
	.w2(32'h3b6a3557),
	.w3(32'h3a1e2acf),
	.w4(32'h3c0b17e8),
	.w5(32'h3c1186a3),
	.w6(32'h3ab8a7d7),
	.w7(32'hb9e32c0b),
	.w8(32'hbb3da31e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdae91c),
	.w1(32'h3c3a454b),
	.w2(32'h3c9f11fd),
	.w3(32'hbc3333ea),
	.w4(32'h3b43c9bb),
	.w5(32'hbcf67fce),
	.w6(32'hbc463b4a),
	.w7(32'h3acee6c2),
	.w8(32'h3c9dad57),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fbcfa2),
	.w1(32'h3b86ea82),
	.w2(32'hbb4d25a6),
	.w3(32'h3c330f86),
	.w4(32'h3b807ba8),
	.w5(32'hbc327d87),
	.w6(32'h3c45fc2b),
	.w7(32'h396c54bd),
	.w8(32'h3a51c863),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96f88c),
	.w1(32'h3b532902),
	.w2(32'hbab31248),
	.w3(32'h3a7ed987),
	.w4(32'hbb40baf5),
	.w5(32'hbb7e014f),
	.w6(32'h3b4ffd86),
	.w7(32'hbb4cf8bd),
	.w8(32'hbb675c3a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a258),
	.w1(32'hbacfe0c5),
	.w2(32'hba38f5c0),
	.w3(32'hbc1253dd),
	.w4(32'h3a9b222b),
	.w5(32'hbc24c48d),
	.w6(32'hbc35848a),
	.w7(32'h3bdf4c52),
	.w8(32'h3bfa407e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d743a),
	.w1(32'hbc893eb1),
	.w2(32'hbcac062e),
	.w3(32'hbc24da71),
	.w4(32'hbbb4b3fd),
	.w5(32'hbb8cdd2a),
	.w6(32'hbb75374d),
	.w7(32'h3b59ebad),
	.w8(32'h3cf1958a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97a67d),
	.w1(32'hbbaf600b),
	.w2(32'hbb87dd29),
	.w3(32'hbabc2a7d),
	.w4(32'hbc4543fd),
	.w5(32'hbc1a84af),
	.w6(32'h3c89aa38),
	.w7(32'hbbcd9dea),
	.w8(32'h3b57c0ca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f232e),
	.w1(32'hbc42996f),
	.w2(32'h3b527e82),
	.w3(32'hbc6fb0b8),
	.w4(32'h3c814513),
	.w5(32'h3cd0c0f2),
	.w6(32'h3b17b9f1),
	.w7(32'hbbf3ff99),
	.w8(32'h3c1f5251),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47a638),
	.w1(32'h3afb3cc8),
	.w2(32'hbb324e16),
	.w3(32'hbc37c837),
	.w4(32'h3b98d4a5),
	.w5(32'h3bb8ff37),
	.w6(32'hb9e5d671),
	.w7(32'hbac97c73),
	.w8(32'hbc222565),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae7b7),
	.w1(32'hbb53a2a6),
	.w2(32'h3a769286),
	.w3(32'hbb903e74),
	.w4(32'hba987a2c),
	.w5(32'hbbac0561),
	.w6(32'hbba66196),
	.w7(32'hbbd470a7),
	.w8(32'hbbf8bfa0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39149164),
	.w1(32'hbbe5617e),
	.w2(32'h3a41fa5d),
	.w3(32'hbbd1f068),
	.w4(32'h3b5815cd),
	.w5(32'h3cd04688),
	.w6(32'h3ac36d65),
	.w7(32'hbc3eb16c),
	.w8(32'hbbf2cdbf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8df286),
	.w1(32'h3a8524c1),
	.w2(32'h3aac888c),
	.w3(32'hbb3b082c),
	.w4(32'hbb3ee06e),
	.w5(32'h3bcae3ca),
	.w6(32'hbb00b685),
	.w7(32'hbb7b2b40),
	.w8(32'h39c13fc5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a246e),
	.w1(32'hbbaf6d25),
	.w2(32'h3aad656f),
	.w3(32'hbbbb7d84),
	.w4(32'hbc5ebb2a),
	.w5(32'h3b003836),
	.w6(32'hbc0c8935),
	.w7(32'hba8a81d9),
	.w8(32'h3c8eb2c2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5f8bc),
	.w1(32'h3b3b5800),
	.w2(32'h3b4dac81),
	.w3(32'hbbf9dfe9),
	.w4(32'hbac3dd0e),
	.w5(32'hbbe78fdc),
	.w6(32'h3bdc381d),
	.w7(32'hbb626943),
	.w8(32'hba09ec2a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ec26),
	.w1(32'hbaabad44),
	.w2(32'hbb6b29e9),
	.w3(32'hbb9291df),
	.w4(32'hbaa02792),
	.w5(32'hbc8df1f1),
	.w6(32'hba43d29c),
	.w7(32'hbbb67173),
	.w8(32'hbbcabf24),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44054e),
	.w1(32'hbbe06dce),
	.w2(32'hbc2c3bcb),
	.w3(32'hbb74d213),
	.w4(32'hbc564297),
	.w5(32'hbc29aafe),
	.w6(32'hbc405c07),
	.w7(32'hbbe43906),
	.w8(32'h393e7de1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0f261),
	.w1(32'h3a993e3b),
	.w2(32'hb98f39a2),
	.w3(32'hbbd6db4d),
	.w4(32'h3ade1f33),
	.w5(32'hbad855db),
	.w6(32'h3bc5626f),
	.w7(32'h3b9056b3),
	.w8(32'h3c049219),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4cd2e),
	.w1(32'h3bb9edf6),
	.w2(32'h3b8b003a),
	.w3(32'hb9c5e04d),
	.w4(32'h39a14812),
	.w5(32'h3b14a352),
	.w6(32'h3be87a44),
	.w7(32'h3b9c812e),
	.w8(32'h3c016b23),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5f03f),
	.w1(32'hbc68cdaf),
	.w2(32'h3c4b3f51),
	.w3(32'h3b19f996),
	.w4(32'hbc34e3db),
	.w5(32'hbc36bab0),
	.w6(32'hbb63abfe),
	.w7(32'hbc147667),
	.w8(32'h3d3a652c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccda79a),
	.w1(32'hba66a129),
	.w2(32'hbb994fce),
	.w3(32'h3bd4850d),
	.w4(32'hbc109c34),
	.w5(32'hbc38abf5),
	.w6(32'h3c1fcd1d),
	.w7(32'h3b0e7b61),
	.w8(32'h3b02d4f4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966f19),
	.w1(32'h3a80dd52),
	.w2(32'hbbb2069b),
	.w3(32'h3c48996c),
	.w4(32'hbb455a76),
	.w5(32'h3b5182b9),
	.w6(32'h3c003cf7),
	.w7(32'hbacda317),
	.w8(32'hbb4b229f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1b25),
	.w1(32'h39d90363),
	.w2(32'hbc5309a6),
	.w3(32'h3affd90e),
	.w4(32'h3ba7ca3f),
	.w5(32'hbb3994ff),
	.w6(32'hbaf5805f),
	.w7(32'hbad5bfb1),
	.w8(32'hbbb83b5a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa2bf2),
	.w1(32'h3ba2a38e),
	.w2(32'h398c156e),
	.w3(32'hbb81d2d0),
	.w4(32'hbab04ffb),
	.w5(32'hbc4f3a16),
	.w6(32'hbc1106b1),
	.w7(32'h3b6724f7),
	.w8(32'h3c7670ee),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eb23b),
	.w1(32'hbc9abe62),
	.w2(32'hbcd66afd),
	.w3(32'hbbcd1883),
	.w4(32'hbae8edce),
	.w5(32'hbc9c1854),
	.w6(32'h3bbb7568),
	.w7(32'h3ca4010b),
	.w8(32'h3d456d8a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61d743),
	.w1(32'h3cc7cddf),
	.w2(32'h3b0f3297),
	.w3(32'hbc9b252f),
	.w4(32'h3c00eeda),
	.w5(32'h3b25ce78),
	.w6(32'h3c7ecfab),
	.w7(32'h3ca4e142),
	.w8(32'h3cc0a710),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bcddf),
	.w1(32'h3a820bf2),
	.w2(32'h3aacb981),
	.w3(32'h3d5bf370),
	.w4(32'h3b1eb041),
	.w5(32'h3b1d88b9),
	.w6(32'h3cab9bc4),
	.w7(32'h3bc7d59e),
	.w8(32'hbb88cd0b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7729ff),
	.w1(32'h3b831b3a),
	.w2(32'h3ba9c9c3),
	.w3(32'hbac1bed9),
	.w4(32'hbb8d7405),
	.w5(32'hba5dc231),
	.w6(32'hba39200d),
	.w7(32'h39dcb010),
	.w8(32'h3b51d381),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba195c21),
	.w1(32'h3bddf873),
	.w2(32'hbb83ab16),
	.w3(32'h3b7cdc4b),
	.w4(32'h39f46e77),
	.w5(32'h3ba8b969),
	.w6(32'h3c15456e),
	.w7(32'h3b1f2afd),
	.w8(32'h39e50d19),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9c2ef),
	.w1(32'hba830072),
	.w2(32'h3b0ac7e0),
	.w3(32'h3b83ae18),
	.w4(32'h3b1ecb57),
	.w5(32'hba8c162a),
	.w6(32'h3b44c8f6),
	.w7(32'h3a16e82e),
	.w8(32'hbbc8fe4e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3547e9),
	.w1(32'h3c12b170),
	.w2(32'h3b983e1f),
	.w3(32'hbc531d54),
	.w4(32'h3c1b1368),
	.w5(32'h3d514866),
	.w6(32'hbc1e0217),
	.w7(32'h3bb0079d),
	.w8(32'hbc8e7e57),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace05b8),
	.w1(32'hbc438eea),
	.w2(32'hbb5824d7),
	.w3(32'h3cd90fdc),
	.w4(32'hba9c0e65),
	.w5(32'hbad3077d),
	.w6(32'hbc5b8100),
	.w7(32'hbb227870),
	.w8(32'h3c91f572),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48f432),
	.w1(32'hba3d4b57),
	.w2(32'h3bb80848),
	.w3(32'hbbc4aae8),
	.w4(32'h3bc3aac1),
	.w5(32'h3a40387a),
	.w6(32'h3c1eb787),
	.w7(32'hbb19a48b),
	.w8(32'h3c272975),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c375530),
	.w1(32'h3b26a32b),
	.w2(32'h3bcc051d),
	.w3(32'hbb68334d),
	.w4(32'h3bd21dc8),
	.w5(32'h3bfddcf1),
	.w6(32'h3bb62977),
	.w7(32'h3a8a65dd),
	.w8(32'hb90fce92),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc11ade),
	.w1(32'hba256982),
	.w2(32'h3bcb0c86),
	.w3(32'h3bec379d),
	.w4(32'h3ac62f98),
	.w5(32'h3b5828ab),
	.w6(32'h3c244e17),
	.w7(32'h3b9b5cda),
	.w8(32'h3bd5c3b0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c3332),
	.w1(32'h3b428433),
	.w2(32'h3b5c1215),
	.w3(32'h3b384b88),
	.w4(32'hbc1d94bd),
	.w5(32'hbc68a782),
	.w6(32'h396d4ae4),
	.w7(32'hb7a066d2),
	.w8(32'hbb549b38),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba675224),
	.w1(32'hba761f71),
	.w2(32'h3bf59a04),
	.w3(32'h3bfef343),
	.w4(32'h3a3e958e),
	.w5(32'h3b7185c7),
	.w6(32'hba821a34),
	.w7(32'hbbc25516),
	.w8(32'hbbe8c501),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed33d),
	.w1(32'h3be79656),
	.w2(32'h3b44b0d6),
	.w3(32'hbba81f99),
	.w4(32'h3b04331d),
	.w5(32'hbbcb2a6e),
	.w6(32'hbae24373),
	.w7(32'h3b73d5d3),
	.w8(32'hbc0c6b19),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42959d),
	.w1(32'h3b2e59fb),
	.w2(32'h3b62f05a),
	.w3(32'h3a2dffb8),
	.w4(32'h3b86a4b1),
	.w5(32'hbbabef87),
	.w6(32'hbbf35e8f),
	.w7(32'h3a3c78c8),
	.w8(32'hbb5f1e02),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d91d7),
	.w1(32'h3a8c0171),
	.w2(32'h3a662715),
	.w3(32'hbb32c4f5),
	.w4(32'hbb9efe0d),
	.w5(32'hbb88e67e),
	.w6(32'hb9c40866),
	.w7(32'h3be1549a),
	.w8(32'h3b4e8c2d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d7e3c),
	.w1(32'h3c925df4),
	.w2(32'h3c49040f),
	.w3(32'hbb395e38),
	.w4(32'h3c9ae1d3),
	.w5(32'h3bdb48be),
	.w6(32'hbbd022d3),
	.w7(32'hba205845),
	.w8(32'hbb85b336),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec40d1),
	.w1(32'h3ad58fe8),
	.w2(32'h3bd5767a),
	.w3(32'h3c400348),
	.w4(32'hba2c356b),
	.w5(32'h3aacfa62),
	.w6(32'hbb6654e3),
	.w7(32'hbb635d38),
	.w8(32'hbb35907e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ad2b6),
	.w1(32'h3c1de5e0),
	.w2(32'h3bbbe719),
	.w3(32'h3c37b893),
	.w4(32'hb986c8b3),
	.w5(32'hbc964c58),
	.w6(32'h3aa63c18),
	.w7(32'h3b4ce287),
	.w8(32'hbbbe0cb5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981f80),
	.w1(32'h3b995fd0),
	.w2(32'h3bc5ebf7),
	.w3(32'hbb81e543),
	.w4(32'h3bdf20b5),
	.w5(32'hba20f310),
	.w6(32'h3b1d3e17),
	.w7(32'hba294b1d),
	.w8(32'hbaf82362),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38f2fb),
	.w1(32'h3b881814),
	.w2(32'hbad293c3),
	.w3(32'hbbee76c3),
	.w4(32'h3b1563b1),
	.w5(32'hbc2484f2),
	.w6(32'h3a449480),
	.w7(32'h3b0a128b),
	.w8(32'hbb58298a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbad9e8),
	.w1(32'hbb098866),
	.w2(32'hbbd5ba7b),
	.w3(32'hbb8ce748),
	.w4(32'hbb15ae1c),
	.w5(32'hbbbfb87c),
	.w6(32'h392c2e1a),
	.w7(32'h3c16dfd0),
	.w8(32'h3bd42cb0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ab52),
	.w1(32'hbc1a3b50),
	.w2(32'hbba7d2d3),
	.w3(32'hbbcb0154),
	.w4(32'hbb63c60a),
	.w5(32'h3c0d022e),
	.w6(32'h3b6d69f6),
	.w7(32'hbbf20737),
	.w8(32'hbbc1aaa9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb397f1),
	.w1(32'hbb6f24ca),
	.w2(32'hbc63cbb4),
	.w3(32'h39d7c237),
	.w4(32'hbae04e03),
	.w5(32'hbaba7e70),
	.w6(32'h3a731fba),
	.w7(32'h38edb579),
	.w8(32'hbb090ff0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37191),
	.w1(32'hbc14a0ad),
	.w2(32'h39e80d54),
	.w3(32'hbbfd9543),
	.w4(32'h3cc3395e),
	.w5(32'h3ba8b45d),
	.w6(32'hbaa72c0d),
	.w7(32'h3c8ec695),
	.w8(32'h3cb650c4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c964371),
	.w1(32'h3b7e9cc9),
	.w2(32'hbb579c62),
	.w3(32'hbb6b428c),
	.w4(32'hbb175b21),
	.w5(32'hbb493922),
	.w6(32'h3c2b8d58),
	.w7(32'h3a72a2be),
	.w8(32'hbb8537a9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba175d98),
	.w1(32'h3b41f334),
	.w2(32'h3ae9be81),
	.w3(32'h3b5b00e7),
	.w4(32'hbabfd2c2),
	.w5(32'hbc284acb),
	.w6(32'h3984da44),
	.w7(32'h3922391d),
	.w8(32'h3ae561db),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cdd0d),
	.w1(32'h3cabab24),
	.w2(32'h3d37dac9),
	.w3(32'h38da0a2c),
	.w4(32'h3c8baa1f),
	.w5(32'h3d4fcced),
	.w6(32'h3a6cd900),
	.w7(32'hbcaf2444),
	.w8(32'hbd513c50),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb99784),
	.w1(32'h3b3e1c0a),
	.w2(32'hbb043da0),
	.w3(32'h3be7ce2a),
	.w4(32'h3adfa0fb),
	.w5(32'hbbfa4b88),
	.w6(32'hbd3a2fff),
	.w7(32'h3b872c75),
	.w8(32'h3b446602),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33614a),
	.w1(32'hbb463265),
	.w2(32'hbc16a0a8),
	.w3(32'h3aebbe7e),
	.w4(32'hbbdb0eb3),
	.w5(32'hbbf633e9),
	.w6(32'hbafedea3),
	.w7(32'h3b464793),
	.w8(32'h3bd38914),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b555a00),
	.w1(32'h39f24737),
	.w2(32'hbb90d1ca),
	.w3(32'hbb3807b2),
	.w4(32'h3b9e246e),
	.w5(32'hbb0b9355),
	.w6(32'h3c471ea8),
	.w7(32'h3c169c09),
	.w8(32'h3c01c494),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118b74),
	.w1(32'h3c692051),
	.w2(32'h3bbe38f4),
	.w3(32'hbbefdd2f),
	.w4(32'hbb007951),
	.w5(32'hbc6e1233),
	.w6(32'h3bdda7c7),
	.w7(32'h3a1ab67c),
	.w8(32'hbbdf8443),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb923c2b),
	.w1(32'h3b44936d),
	.w2(32'hbb2969e5),
	.w3(32'hbba19c78),
	.w4(32'hbbe526cf),
	.w5(32'hbc0ba253),
	.w6(32'hbc42f07a),
	.w7(32'hbb5e7d2e),
	.w8(32'hbc079e8e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f558e),
	.w1(32'hbd167924),
	.w2(32'hbd31aa5f),
	.w3(32'h3b7f46e3),
	.w4(32'hbc748627),
	.w5(32'h3db0e167),
	.w6(32'hbb07ada2),
	.w7(32'hbc9ef782),
	.w8(32'hbbf8aa9f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca4437),
	.w1(32'hbc1924c7),
	.w2(32'hbbeaeeb4),
	.w3(32'hbaac2108),
	.w4(32'hba23108e),
	.w5(32'h3cc10a87),
	.w6(32'hbc20a026),
	.w7(32'hbc030f8f),
	.w8(32'h3c0a74a9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2f39b),
	.w1(32'hbbe43f03),
	.w2(32'hba0ebb9b),
	.w3(32'h3ba96c28),
	.w4(32'hba96eb07),
	.w5(32'hbb1d4adb),
	.w6(32'h3c35e2ef),
	.w7(32'hbbdefdf9),
	.w8(32'hbb96d1cf),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb799f6),
	.w1(32'h3bb4b45e),
	.w2(32'hbbb146cd),
	.w3(32'h3a82cf09),
	.w4(32'h3b61bf9b),
	.w5(32'hbaab3494),
	.w6(32'h3bb2ebe8),
	.w7(32'h3babe9b3),
	.w8(32'hbbca49f3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25819d),
	.w1(32'h3abb6ab9),
	.w2(32'h3ac342e3),
	.w3(32'h3b64cd2a),
	.w4(32'h3b846fad),
	.w5(32'h3a277b69),
	.w6(32'hb9cf2ab1),
	.w7(32'h3bc6e782),
	.w8(32'h3b88642f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39604243),
	.w1(32'hbb411ea3),
	.w2(32'h3b30b0ac),
	.w3(32'hbb50c8a6),
	.w4(32'h3a474654),
	.w5(32'hbbe95456),
	.w6(32'hbb50468a),
	.w7(32'hbb8348ae),
	.w8(32'hbaa06206),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27a24),
	.w1(32'hb9368804),
	.w2(32'h3bc6e8a3),
	.w3(32'h3b69e8c3),
	.w4(32'h3989766c),
	.w5(32'h3bc177aa),
	.w6(32'h3b838316),
	.w7(32'hbc266d9a),
	.w8(32'hbbe48ebb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd5372),
	.w1(32'hbb1be791),
	.w2(32'hbb2ca9fb),
	.w3(32'hba9ca20c),
	.w4(32'hbbf7ff8c),
	.w5(32'hbc60e661),
	.w6(32'hbc05690f),
	.w7(32'hbb5162ca),
	.w8(32'hbbbad49b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cc1c),
	.w1(32'hbb2b54bc),
	.w2(32'hbc17632b),
	.w3(32'hbba1dcc6),
	.w4(32'hbc255afe),
	.w5(32'hba4f7a6d),
	.w6(32'hbadd5e37),
	.w7(32'hbb8c283b),
	.w8(32'hbc7192c6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc2fa9),
	.w1(32'hbc925c88),
	.w2(32'hbb20dc41),
	.w3(32'h3c865545),
	.w4(32'h3bdd2d3f),
	.w5(32'h3cb5e294),
	.w6(32'hbc15900b),
	.w7(32'hbc219625),
	.w8(32'h3ad7a539),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc39aa),
	.w1(32'h3a9bfed0),
	.w2(32'hbb610f83),
	.w3(32'hbc9365b5),
	.w4(32'h3b66411e),
	.w5(32'hbbffacfb),
	.w6(32'hbc76939f),
	.w7(32'hbb6874b1),
	.w8(32'hbbc675ed),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd2fda),
	.w1(32'h3bf0ed60),
	.w2(32'h3a18109c),
	.w3(32'h3bfc2769),
	.w4(32'h3bc2aee1),
	.w5(32'hbb9b0817),
	.w6(32'hba185841),
	.w7(32'h3c5b740b),
	.w8(32'h3b99e146),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54a0de),
	.w1(32'h3a4e8c84),
	.w2(32'hbbbabe9e),
	.w3(32'h3ad04bb5),
	.w4(32'h3bbf9513),
	.w5(32'h3ba14059),
	.w6(32'h3a99ba66),
	.w7(32'h3b0648d4),
	.w8(32'hbb6d0366),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15f749),
	.w1(32'h3c25e06b),
	.w2(32'h3c12b965),
	.w3(32'h3b4c233d),
	.w4(32'h3bb3116b),
	.w5(32'h3bfb0c62),
	.w6(32'hbbdf89cb),
	.w7(32'hbbad67ff),
	.w8(32'hbcaa8142),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c348927),
	.w1(32'hbb9d30de),
	.w2(32'hbc0da0e9),
	.w3(32'h3c859c56),
	.w4(32'hbbe09b67),
	.w5(32'hbbefe403),
	.w6(32'hbc53b958),
	.w7(32'hbb69e83a),
	.w8(32'h3a859fc4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfa3dd),
	.w1(32'h3c2f7000),
	.w2(32'h3b93f1fc),
	.w3(32'hbbd24fe5),
	.w4(32'hbbfdafa8),
	.w5(32'hbb8768c5),
	.w6(32'hbb0f2654),
	.w7(32'h3bcc2c12),
	.w8(32'hbc1e2f2c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08390c),
	.w1(32'h3a6035f4),
	.w2(32'hb9b0417f),
	.w3(32'h3ca05c9d),
	.w4(32'h3a2ac1ec),
	.w5(32'hbb9d5b23),
	.w6(32'hbbb3db90),
	.w7(32'hbb3c32d2),
	.w8(32'h3880e826),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d0e9),
	.w1(32'h3bc13b97),
	.w2(32'h38c23030),
	.w3(32'hbbcc333a),
	.w4(32'hba0e5dd6),
	.w5(32'hbba194e4),
	.w6(32'hbb0e1391),
	.w7(32'hbac10164),
	.w8(32'hbae09c2e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7247ad),
	.w1(32'hbb1c5093),
	.w2(32'hbb9c11e9),
	.w3(32'h3ba514fc),
	.w4(32'h3b1382ab),
	.w5(32'h39c2bca1),
	.w6(32'h3a970e5b),
	.w7(32'hbb111f7d),
	.w8(32'h3b536dfc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6565e),
	.w1(32'h3bc203a0),
	.w2(32'h3b94077c),
	.w3(32'hbab6edbd),
	.w4(32'h3b34a31d),
	.w5(32'hbc41a1be),
	.w6(32'h3b843bbf),
	.w7(32'h3b0f73e1),
	.w8(32'h3bb425ac),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec132),
	.w1(32'h3b9b45c5),
	.w2(32'h3baa079d),
	.w3(32'hba9f6a0d),
	.w4(32'h3c205241),
	.w5(32'hbb109758),
	.w6(32'hbb9bcace),
	.w7(32'h3c8985ea),
	.w8(32'h3ba8d4d2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e55fb),
	.w1(32'hbb6cf95f),
	.w2(32'hbb93d8c4),
	.w3(32'hba3740b8),
	.w4(32'h3c380995),
	.w5(32'h3af14878),
	.w6(32'h3a982ca9),
	.w7(32'h3c30a407),
	.w8(32'h3c074d54),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8596d),
	.w1(32'hbbed6df2),
	.w2(32'h3b962bf7),
	.w3(32'hbc25dc00),
	.w4(32'h3b4a8f3c),
	.w5(32'h3c8be4f7),
	.w6(32'h3adea33e),
	.w7(32'hbc2385e9),
	.w8(32'h3a22f20c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05db32),
	.w1(32'h3b9288b2),
	.w2(32'hbae0f016),
	.w3(32'hbbe82ac3),
	.w4(32'hbb9d89e3),
	.w5(32'hbb495a90),
	.w6(32'hbb77b1fd),
	.w7(32'h3aae5dc6),
	.w8(32'h3ae664e8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cf67e),
	.w1(32'h3c3015ad),
	.w2(32'h3bd95085),
	.w3(32'hbb89d2b3),
	.w4(32'h3c34b6ac),
	.w5(32'h3c29cc50),
	.w6(32'hbb9378d4),
	.w7(32'h3bf45f7f),
	.w8(32'hbb44be39),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be895dd),
	.w1(32'h3c0ae7da),
	.w2(32'hbb977792),
	.w3(32'h3c175e8c),
	.w4(32'h3b1704c9),
	.w5(32'hbbfe8d98),
	.w6(32'hbad091e8),
	.w7(32'h3b8c3456),
	.w8(32'hbbd0f45c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7e1b9),
	.w1(32'h3b4857df),
	.w2(32'hbb77a04c),
	.w3(32'h3bc5a88e),
	.w4(32'hbbb584a6),
	.w5(32'hbc95937e),
	.w6(32'h38cd696f),
	.w7(32'h3b564fa6),
	.w8(32'h3b4c24cc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb7888),
	.w1(32'hbbdd7a83),
	.w2(32'h3c75efe9),
	.w3(32'hbbe07400),
	.w4(32'h3b05fa84),
	.w5(32'hbc6ffa14),
	.w6(32'hbb6be0bc),
	.w7(32'h3a47ad1a),
	.w8(32'h3a934200),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba540bf),
	.w1(32'hb91e8fb2),
	.w2(32'hbbb2227b),
	.w3(32'hbc9fb267),
	.w4(32'hbba695d5),
	.w5(32'hbc165f63),
	.w6(32'hbb8bcc79),
	.w7(32'hbaebf549),
	.w8(32'h3b5c1656),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5858a7),
	.w1(32'hbae3ebc7),
	.w2(32'hbad17402),
	.w3(32'h3b85b29e),
	.w4(32'hbaa4a44b),
	.w5(32'hbaa3174a),
	.w6(32'h3c423427),
	.w7(32'hbac574e2),
	.w8(32'hbae33ebf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace3ee5),
	.w1(32'hb79bfee5),
	.w2(32'h39eb3fd2),
	.w3(32'hbad0e45f),
	.w4(32'h3910a066),
	.w5(32'hb764e9b8),
	.w6(32'hbac8ede6),
	.w7(32'h3863c986),
	.w8(32'h39902601),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eaf8a8),
	.w1(32'h3804fed9),
	.w2(32'hb8f4726a),
	.w3(32'h3959c738),
	.w4(32'h38e292de),
	.w5(32'hba65a6cb),
	.w6(32'hb9578d8d),
	.w7(32'hb9bea15a),
	.w8(32'hba4aea74),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa0605),
	.w1(32'hba2257fd),
	.w2(32'hba0507a9),
	.w3(32'hb9d7dc90),
	.w4(32'hba19d2c9),
	.w5(32'hba9495ac),
	.w6(32'hba352335),
	.w7(32'hba0b6ec8),
	.w8(32'hba65f381),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc86dd),
	.w1(32'h3933b541),
	.w2(32'h397e8aa3),
	.w3(32'hba3ff384),
	.w4(32'h39642dd8),
	.w5(32'h3a02c1c1),
	.w6(32'hba5effad),
	.w7(32'h39c01dc1),
	.w8(32'h3a09da11),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dff030),
	.w1(32'h399d953e),
	.w2(32'hb8023b22),
	.w3(32'h39de0749),
	.w4(32'hba671698),
	.w5(32'hb93bb4b3),
	.w6(32'h39b13a2e),
	.w7(32'hba0f435a),
	.w8(32'hb9d27c73),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795b2e6),
	.w1(32'hba62b029),
	.w2(32'hba25db90),
	.w3(32'hb70a9bf0),
	.w4(32'hba147510),
	.w5(32'hba0d57c3),
	.w6(32'hb98d70e6),
	.w7(32'h391cedbe),
	.w8(32'h3a0271c0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba062dcc),
	.w1(32'hba97c1ce),
	.w2(32'hbae779c8),
	.w3(32'hb996316b),
	.w4(32'hbac5c701),
	.w5(32'hbad3c99f),
	.w6(32'h3989dd80),
	.w7(32'hbb0765e5),
	.w8(32'hbb0effd4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefe8fe),
	.w1(32'hba0879c3),
	.w2(32'hb9c9fbf4),
	.w3(32'hbb0b0809),
	.w4(32'hb941b22c),
	.w5(32'hbab64109),
	.w6(32'hbad937e0),
	.w7(32'h38e3e447),
	.w8(32'h36778097),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b918c1),
	.w1(32'h3aab4e5f),
	.w2(32'h3a8f5980),
	.w3(32'h38fbbe04),
	.w4(32'h3a68b59b),
	.w5(32'h39d487bb),
	.w6(32'hb8c643d8),
	.w7(32'h3a85b655),
	.w8(32'h3a0fb22f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84536c),
	.w1(32'hba017276),
	.w2(32'hb981c269),
	.w3(32'h3a2cb203),
	.w4(32'hb9b0342f),
	.w5(32'h39e56bc2),
	.w6(32'h3a5366c5),
	.w7(32'hba4791b9),
	.w8(32'hba074265),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03de38),
	.w1(32'h3aa9a401),
	.w2(32'h3a9226a2),
	.w3(32'hb9ececc2),
	.w4(32'h3aa62aec),
	.w5(32'h3aac1425),
	.w6(32'hba5e438e),
	.w7(32'h3aadd023),
	.w8(32'h3a7cc90e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27b0e6),
	.w1(32'h3979cb6c),
	.w2(32'hb863409e),
	.w3(32'h39d07cb4),
	.w4(32'h393fbee0),
	.w5(32'h38313a01),
	.w6(32'h39c188ef),
	.w7(32'h38d8e0c4),
	.w8(32'hb85e889e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3c9bf),
	.w1(32'h3a91ebcd),
	.w2(32'h3a56b545),
	.w3(32'hb9a7ddfb),
	.w4(32'h3a2fcb61),
	.w5(32'h3a49eb9b),
	.w6(32'hb99ec2f9),
	.w7(32'h39acc194),
	.w8(32'h39258b2c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e8cd9),
	.w1(32'hba13574d),
	.w2(32'hba262f00),
	.w3(32'h3a4404ce),
	.w4(32'hba112618),
	.w5(32'hbaba1537),
	.w6(32'h398ae744),
	.w7(32'hba7c22e8),
	.w8(32'hba53bcaf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cfb97),
	.w1(32'h3635ab5b),
	.w2(32'h38f9e0a0),
	.w3(32'hba902b8b),
	.w4(32'h385e1cb6),
	.w5(32'hba465bfe),
	.w6(32'hba763520),
	.w7(32'h39be7415),
	.w8(32'h39cddaf4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e943c2),
	.w1(32'hba3bf75d),
	.w2(32'hb99d18ed),
	.w3(32'hb8d17c9f),
	.w4(32'hba11b031),
	.w5(32'hbaa2b81c),
	.w6(32'hb9a97208),
	.w7(32'hb94ffe34),
	.w8(32'hb9da2156),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd7873),
	.w1(32'hb9eb8118),
	.w2(32'hb8f374e8),
	.w3(32'h39a19fa8),
	.w4(32'hb93956b5),
	.w5(32'hba4f55fa),
	.w6(32'h397caa3a),
	.w7(32'hba0ef1ca),
	.w8(32'hb9d362d5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dd464),
	.w1(32'hb9ed18c9),
	.w2(32'hb9b62e59),
	.w3(32'h39efabd8),
	.w4(32'h38e70e02),
	.w5(32'hba5ab5ff),
	.w6(32'h39d7ff88),
	.w7(32'hb99a2d5d),
	.w8(32'h397ec69a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a117e38),
	.w1(32'h3800743a),
	.w2(32'hb9a2f14a),
	.w3(32'h3a8f3702),
	.w4(32'hb80576bc),
	.w5(32'hb9403cbc),
	.w6(32'h3a9efdcc),
	.w7(32'hba27b759),
	.w8(32'hba23b7d0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9713912),
	.w1(32'hb91f85ea),
	.w2(32'hb92c0a48),
	.w3(32'hb9a5ecd4),
	.w4(32'hba77f003),
	.w5(32'hba31eb54),
	.w6(32'h39efc708),
	.w7(32'hba56def2),
	.w8(32'hba7a7563),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b8348),
	.w1(32'h394b6053),
	.w2(32'hb94da801),
	.w3(32'hb8e1031b),
	.w4(32'hb8287384),
	.w5(32'hb9cbc1c6),
	.w6(32'hb9c571de),
	.w7(32'hb98ccaae),
	.w8(32'h3961b37b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a154349),
	.w1(32'h3900e87e),
	.w2(32'hb925b7cc),
	.w3(32'h3a1c1545),
	.w4(32'hb8c7a3de),
	.w5(32'hba512add),
	.w6(32'h3a38e4d3),
	.w7(32'h391e8936),
	.w8(32'h39be7fa9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949876),
	.w1(32'h3a5b3a8d),
	.w2(32'h39dfe02e),
	.w3(32'hba1810fe),
	.w4(32'h3a241462),
	.w5(32'h38ed4b52),
	.w6(32'hb9718f44),
	.w7(32'h3a87d154),
	.w8(32'h38d229d9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eab48c),
	.w1(32'h397ad173),
	.w2(32'hb845a91d),
	.w3(32'h3a0c5c36),
	.w4(32'h3a0a82ac),
	.w5(32'hb8bca6af),
	.w6(32'hb90c6a88),
	.w7(32'h3a8966f0),
	.w8(32'h39fa9f6b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928c185),
	.w1(32'hba03a2e2),
	.w2(32'hb9f73834),
	.w3(32'hb8a9e60f),
	.w4(32'hba539ac7),
	.w5(32'hba872265),
	.w6(32'h39a91c96),
	.w7(32'hba5f5481),
	.w8(32'hba7a840f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6bbd4),
	.w1(32'h39f58ec8),
	.w2(32'h3a4165c2),
	.w3(32'hba308cb2),
	.w4(32'h3a935218),
	.w5(32'h3a788474),
	.w6(32'hba7dd1b0),
	.w7(32'h3a0c2f76),
	.w8(32'h3a529348),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01e9e3),
	.w1(32'h39b54cc4),
	.w2(32'h3a62c88b),
	.w3(32'h3a963d3d),
	.w4(32'h3a51c00d),
	.w5(32'h3a429e68),
	.w6(32'h3a4010fc),
	.w7(32'h39df5b75),
	.w8(32'h3a1e56c9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391321a6),
	.w1(32'hb89230d6),
	.w2(32'hba16f0c4),
	.w3(32'h3a20212c),
	.w4(32'hba05d5a8),
	.w5(32'hba4c5aac),
	.w6(32'h39df7995),
	.w7(32'hb8aafc86),
	.w8(32'hb984a569),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f556c4),
	.w1(32'hbadefdcd),
	.w2(32'hbaf1d54d),
	.w3(32'h38d00be8),
	.w4(32'hbb08de72),
	.w5(32'hbb2069b6),
	.w6(32'hb969e8d7),
	.w7(32'hbb00ebbe),
	.w8(32'hbb01aab3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07a5de),
	.w1(32'hba059bc2),
	.w2(32'hb9bfb073),
	.w3(32'hbb28e75d),
	.w4(32'hba382b7b),
	.w5(32'hba4af8b7),
	.w6(32'hbb12d6eb),
	.w7(32'hb889f823),
	.w8(32'hb855264b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7c3c6),
	.w1(32'hb940da27),
	.w2(32'h39a5c615),
	.w3(32'hb9b4b13b),
	.w4(32'h383fe3f8),
	.w5(32'hb85e3e5a),
	.w6(32'hb9a25aec),
	.w7(32'hb89599ec),
	.w8(32'hb9b7c441),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb795632c),
	.w1(32'hba03ddce),
	.w2(32'hb9c246c9),
	.w3(32'hb92dc310),
	.w4(32'hb9407bd5),
	.w5(32'hba642695),
	.w6(32'hb92a4450),
	.w7(32'hb9022501),
	.w8(32'hba0e349e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9a8e2),
	.w1(32'hba872bb7),
	.w2(32'hb9a6d95d),
	.w3(32'hb8d1a8a5),
	.w4(32'hba19bfb1),
	.w5(32'hb985638a),
	.w6(32'hb959e196),
	.w7(32'hba2e6de4),
	.w8(32'hb98014b8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f99a0b),
	.w1(32'hba6425bc),
	.w2(32'hb9413563),
	.w3(32'hb753684e),
	.w4(32'hba37fb0a),
	.w5(32'hba5adb8f),
	.w6(32'hba0f5b1b),
	.w7(32'hba399340),
	.w8(32'hba533dba),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1191f1),
	.w1(32'h39ec1a8f),
	.w2(32'h3a16b409),
	.w3(32'hba28ae03),
	.w4(32'h3915eee2),
	.w5(32'hb98a893e),
	.w6(32'hba909f1f),
	.w7(32'hb8f6be16),
	.w8(32'h37fb8bfa),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0420b),
	.w1(32'hb6f597b9),
	.w2(32'h388e4077),
	.w3(32'h39be0979),
	.w4(32'hb7fc40f4),
	.w5(32'hba08dd96),
	.w6(32'hb91f3456),
	.w7(32'h3703b065),
	.w8(32'hb9c97059),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39960e27),
	.w1(32'hb9b31c35),
	.w2(32'hb9e3929c),
	.w3(32'hb9bf4ae9),
	.w4(32'hba128582),
	.w5(32'hb988ede8),
	.w6(32'hb92538d7),
	.w7(32'hb981c404),
	.w8(32'hb8e61875),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad862e),
	.w1(32'h38408d27),
	.w2(32'hb93e90c9),
	.w3(32'hb995844c),
	.w4(32'h39705c7f),
	.w5(32'hb997c224),
	.w6(32'hb90be07d),
	.w7(32'hb8ee7370),
	.w8(32'hb881904f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876e127),
	.w1(32'h39909f93),
	.w2(32'h3a31e5f5),
	.w3(32'hb7a80b20),
	.w4(32'h391f021b),
	.w5(32'hb9cd452e),
	.w6(32'hb89f104e),
	.w7(32'h37aca04f),
	.w8(32'h39820ec7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38490226),
	.w1(32'hb9bfed6c),
	.w2(32'hb9fc0115),
	.w3(32'hb87b997c),
	.w4(32'hb9ee84ed),
	.w5(32'hbac9d799),
	.w6(32'hb937de2b),
	.w7(32'hba1dd282),
	.w8(32'hba1f1892),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880b492),
	.w1(32'hba24cddc),
	.w2(32'hba4cd2cd),
	.w3(32'hb82a1b62),
	.w4(32'hba085066),
	.w5(32'hb9d43d55),
	.w6(32'hba25194a),
	.w7(32'hba1ab4a9),
	.w8(32'hba03e342),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa10447),
	.w1(32'hba81801a),
	.w2(32'hba670e70),
	.w3(32'hba6bfb55),
	.w4(32'hba6716a4),
	.w5(32'hba8a5894),
	.w6(32'hba6e1adf),
	.w7(32'hba28d2de),
	.w8(32'hba36795d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2d86),
	.w1(32'hb97a1b03),
	.w2(32'h38fd409c),
	.w3(32'hba203e54),
	.w4(32'h387f5ba2),
	.w5(32'h3a2cde9f),
	.w6(32'hba4696bf),
	.w7(32'h3882c60d),
	.w8(32'h3a01145b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb78d7),
	.w1(32'hb97c148b),
	.w2(32'hb927f9ea),
	.w3(32'h3a0639eb),
	.w4(32'hb8b4599b),
	.w5(32'h3a377f13),
	.w6(32'h39ec702a),
	.w7(32'hb9b976f0),
	.w8(32'hb91862ac),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa366f5),
	.w1(32'h393e691c),
	.w2(32'hb8ea5134),
	.w3(32'hb9855641),
	.w4(32'h38d6c5ef),
	.w5(32'h3914a43b),
	.w6(32'h37ccdb96),
	.w7(32'h39de2ced),
	.w8(32'hba137dee),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff5dfe),
	.w1(32'hb9f38b11),
	.w2(32'hba3fe20a),
	.w3(32'hba3fcee0),
	.w4(32'hb9b77f38),
	.w5(32'hba376d46),
	.w6(32'hba7c558b),
	.w7(32'hb9ce7d9e),
	.w8(32'hba55ac9b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2688b5),
	.w1(32'h39bc3e2e),
	.w2(32'h38fe0689),
	.w3(32'hba03c250),
	.w4(32'h3a382ffb),
	.w5(32'hb99e6c64),
	.w6(32'hba20887b),
	.w7(32'h3a8a1203),
	.w8(32'h39a59f70),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a77a9),
	.w1(32'h39f3814a),
	.w2(32'hb9dc19f8),
	.w3(32'hb97b0241),
	.w4(32'h39bb3247),
	.w5(32'h3925ea93),
	.w6(32'h395dda0e),
	.w7(32'h3a0d5dd4),
	.w8(32'hb87d004d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9986bde),
	.w1(32'hb91eb2bf),
	.w2(32'h37e90de5),
	.w3(32'hb98df409),
	.w4(32'h3a40841c),
	.w5(32'h39b5231e),
	.w6(32'hb9e39f12),
	.w7(32'h39eb468b),
	.w8(32'h3a467e91),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934f4a3),
	.w1(32'h3a0e9346),
	.w2(32'h3a16d6fa),
	.w3(32'h3a6c5a8d),
	.w4(32'h3a4338c3),
	.w5(32'h38bd62f1),
	.w6(32'h3a4124a9),
	.w7(32'h39f67f1c),
	.w8(32'h39696371),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49291c),
	.w1(32'h396bb014),
	.w2(32'hba29861b),
	.w3(32'h398d7816),
	.w4(32'hb9e636c6),
	.w5(32'hba2454aa),
	.w6(32'h39073557),
	.w7(32'hb9fbd2c0),
	.w8(32'hba65c0f4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f544ee),
	.w1(32'h3990cd9e),
	.w2(32'h3a2154c2),
	.w3(32'hba3919fc),
	.w4(32'h3a0f2dba),
	.w5(32'h39c5c5ba),
	.w6(32'hb98666c3),
	.w7(32'h39064075),
	.w8(32'h37286f0a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac5c4f),
	.w1(32'hb8a7b2ef),
	.w2(32'hb8411d01),
	.w3(32'hb9046346),
	.w4(32'h387f300e),
	.w5(32'hb8844383),
	.w6(32'h390af2a9),
	.w7(32'hba01116d),
	.w8(32'hb82b474e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f3317),
	.w1(32'h3900e3da),
	.w2(32'h3a02888d),
	.w3(32'h39e04c50),
	.w4(32'h39f7a272),
	.w5(32'h399cf7ce),
	.w6(32'h391785d9),
	.w7(32'h3a451ec8),
	.w8(32'h3a7bc922),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f6de0),
	.w1(32'hba1f3e51),
	.w2(32'hba1f7c0f),
	.w3(32'h3a8cc198),
	.w4(32'hb9c383ca),
	.w5(32'hbadc152d),
	.w6(32'h3a728039),
	.w7(32'hb986bd25),
	.w8(32'hb7e79b5e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79cf2c),
	.w1(32'hb91fbd80),
	.w2(32'hba031fda),
	.w3(32'hba345284),
	.w4(32'hb93cd593),
	.w5(32'h394ea8cf),
	.w6(32'hba1e5162),
	.w7(32'hb9b85402),
	.w8(32'hb8a7ee25),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1631db),
	.w1(32'h3a089aa3),
	.w2(32'h39a39fe5),
	.w3(32'hb8f4bab3),
	.w4(32'h3999f40e),
	.w5(32'h3a11f6b0),
	.w6(32'hba40bf5a),
	.w7(32'h39b41b7b),
	.w8(32'h3a5e63b5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d64c9e),
	.w1(32'h397a92ac),
	.w2(32'h3a01b305),
	.w3(32'h39978d05),
	.w4(32'h39de94d7),
	.w5(32'h39ae9b3d),
	.w6(32'h3a0ef26a),
	.w7(32'hb841d485),
	.w8(32'h39bc3b2e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule