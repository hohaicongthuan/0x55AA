module layer_8_featuremap_228(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9e4f),
	.w1(32'h3baf1733),
	.w2(32'h3c02853e),
	.w3(32'hb9dbf270),
	.w4(32'hbb0dd6c7),
	.w5(32'h3a7901e3),
	.w6(32'hbb068cde),
	.w7(32'h39d31d64),
	.w8(32'hbab5f88f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc2e6b),
	.w1(32'h3b67ff62),
	.w2(32'h3b2069dc),
	.w3(32'hba4431a5),
	.w4(32'hbb880902),
	.w5(32'hbbaf436f),
	.w6(32'h3bbf9f2d),
	.w7(32'h3b995ae6),
	.w8(32'h3a8de7ee),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c760a),
	.w1(32'hba6b6080),
	.w2(32'hba594d76),
	.w3(32'hbac46a27),
	.w4(32'h3aeb8c08),
	.w5(32'hbb58fade),
	.w6(32'h3b7e4e9b),
	.w7(32'hbbd2d7bc),
	.w8(32'hbafc71eb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226b65),
	.w1(32'h3b146043),
	.w2(32'h3bb46a0d),
	.w3(32'hbb4f1bf9),
	.w4(32'hbbb1ce81),
	.w5(32'hbb4820a5),
	.w6(32'hb7df1098),
	.w7(32'h3b8033f8),
	.w8(32'h39d5fa3c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba84723),
	.w1(32'h3b5fb9a4),
	.w2(32'h3b37ce22),
	.w3(32'hbc2dcaaa),
	.w4(32'hbb7db814),
	.w5(32'hbb24831a),
	.w6(32'h3a27d184),
	.w7(32'hbaa70154),
	.w8(32'hbb359336),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d49fe),
	.w1(32'hbaba5d5f),
	.w2(32'hbac477fd),
	.w3(32'h3a7a3818),
	.w4(32'hbaa71739),
	.w5(32'hbb34ca25),
	.w6(32'h3aa97f8e),
	.w7(32'h3bb8da18),
	.w8(32'h3b69c3f8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9dc87),
	.w1(32'hb915244b),
	.w2(32'h39783358),
	.w3(32'hbb8cb517),
	.w4(32'hb989da15),
	.w5(32'h38a9f153),
	.w6(32'hba4f8e4c),
	.w7(32'h389a8968),
	.w8(32'hbac0c3b7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add32a0),
	.w1(32'h3b5594eb),
	.w2(32'h39bc1ded),
	.w3(32'h3b7807f4),
	.w4(32'h3a5f496e),
	.w5(32'hbb7ef4b2),
	.w6(32'h3b953020),
	.w7(32'h3b8b9737),
	.w8(32'hbb2b4970),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a49fd0),
	.w1(32'h3b7e7820),
	.w2(32'hbad7c05d),
	.w3(32'h3ae81e18),
	.w4(32'hbb4697c1),
	.w5(32'hbc1b720e),
	.w6(32'h3b30c52a),
	.w7(32'hbbbc12f9),
	.w8(32'hbc26a7d5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1ea30),
	.w1(32'hbbe58d3c),
	.w2(32'hbbb8c63b),
	.w3(32'hbb7f7a8b),
	.w4(32'hbb947049),
	.w5(32'hbc25cada),
	.w6(32'hba80d2bf),
	.w7(32'h3a24c984),
	.w8(32'hbb6862a8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba783300),
	.w1(32'h3afbbfd8),
	.w2(32'hbac19f3a),
	.w3(32'hbc504157),
	.w4(32'hba577c86),
	.w5(32'hbbae6e68),
	.w6(32'hbb1ef1f4),
	.w7(32'hbbe5fa74),
	.w8(32'h3a90140f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e5507),
	.w1(32'hb9e0ae9e),
	.w2(32'h3a386a09),
	.w3(32'hbb880492),
	.w4(32'hbbb3b5db),
	.w5(32'hbb533fc0),
	.w6(32'hba25ad29),
	.w7(32'h3bdf70c7),
	.w8(32'h3b3d4646),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa4a9f),
	.w1(32'hbbaae185),
	.w2(32'hbb1dc5eb),
	.w3(32'h3b1b513c),
	.w4(32'hbad92da6),
	.w5(32'hbb6fe333),
	.w6(32'hb9403506),
	.w7(32'h3b1f9aa9),
	.w8(32'h3a9d04c6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13edd),
	.w1(32'h3b74269d),
	.w2(32'hbb6c2c25),
	.w3(32'hbb239b77),
	.w4(32'h3b666259),
	.w5(32'hbb9f1e84),
	.w6(32'h3b4e7732),
	.w7(32'hba851e36),
	.w8(32'h3a6c62c8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3871495a),
	.w1(32'h3ad298f2),
	.w2(32'hb842d8dd),
	.w3(32'hbb49c7ec),
	.w4(32'h3b8a4ed5),
	.w5(32'h3b1a2b15),
	.w6(32'hbb0b20a0),
	.w7(32'hbb81979d),
	.w8(32'hbb094965),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1da0f),
	.w1(32'hba74a424),
	.w2(32'h3ba84743),
	.w3(32'h3b2456e4),
	.w4(32'hbbb23d46),
	.w5(32'hbb0e773c),
	.w6(32'hba9a1c08),
	.w7(32'h3a8e3adc),
	.w8(32'hbc0db8ff),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee8233),
	.w1(32'h3a823aa4),
	.w2(32'h3a8c77d4),
	.w3(32'hbc06b9d1),
	.w4(32'h3acf1757),
	.w5(32'h3b8842a3),
	.w6(32'hba1feeb0),
	.w7(32'hb87bed0c),
	.w8(32'h3c046be3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafe445),
	.w1(32'hba73530b),
	.w2(32'h3bea956a),
	.w3(32'hbb7d3e98),
	.w4(32'hbb6a0376),
	.w5(32'h39bef031),
	.w6(32'h3b30210e),
	.w7(32'h3b9cdc17),
	.w8(32'h3aafaefd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74b8ba),
	.w1(32'h3c73c428),
	.w2(32'h3c583c88),
	.w3(32'h3bede291),
	.w4(32'hbb0971e6),
	.w5(32'hbbc49add),
	.w6(32'h3bd6598e),
	.w7(32'h3c5a9d2b),
	.w8(32'h3b9819d9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c214f23),
	.w1(32'h3c0813b0),
	.w2(32'h3b6756d2),
	.w3(32'hbc93abd7),
	.w4(32'hba1502b9),
	.w5(32'hbb602fd3),
	.w6(32'hbb16ab90),
	.w7(32'hbbbd3d03),
	.w8(32'hbbf3ee8c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1665ec),
	.w1(32'h3b140003),
	.w2(32'hbacd2fb7),
	.w3(32'hbb078673),
	.w4(32'h3badc84e),
	.w5(32'h3c85972d),
	.w6(32'h3a8de77a),
	.w7(32'hbc2080f0),
	.w8(32'hba5d34d3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be064a2),
	.w1(32'h3b20cc99),
	.w2(32'h3c0f89a0),
	.w3(32'h3c2935b1),
	.w4(32'h3becb42e),
	.w5(32'h3a05fcd8),
	.w6(32'h3a87f909),
	.w7(32'hbbd3fb89),
	.w8(32'hbb97e9bc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9edd35),
	.w1(32'h3c8c847f),
	.w2(32'h3c98c2b5),
	.w3(32'hbbd38b8e),
	.w4(32'h3acd8341),
	.w5(32'hbbf71abb),
	.w6(32'hba97d0c6),
	.w7(32'h3b80b5f2),
	.w8(32'h3bb32e57),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978efe),
	.w1(32'h3a186613),
	.w2(32'h3b8b9816),
	.w3(32'hbbf56da1),
	.w4(32'h3bdd16b2),
	.w5(32'h3ad2eca7),
	.w6(32'h3acd98fc),
	.w7(32'hbbe42d92),
	.w8(32'hbb1d25bc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f94d4),
	.w1(32'h3b800ae1),
	.w2(32'h3c0df4f7),
	.w3(32'h3c119366),
	.w4(32'h3b2a98a2),
	.w5(32'hba4f5d52),
	.w6(32'h3b0a0b66),
	.w7(32'h3b859d69),
	.w8(32'h3c02b311),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2f49),
	.w1(32'h3c559a33),
	.w2(32'h3c89548d),
	.w3(32'hbc0a5ecd),
	.w4(32'hbb536c5c),
	.w5(32'hbb5303a4),
	.w6(32'hb997d2cf),
	.w7(32'hbb732dd3),
	.w8(32'hbb11f239),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23387d),
	.w1(32'h3a693e18),
	.w2(32'hb9d624a1),
	.w3(32'h395b7ea0),
	.w4(32'h39dc6c9d),
	.w5(32'hbb081e71),
	.w6(32'hbb20ed03),
	.w7(32'h3b7e471b),
	.w8(32'h3ba13e35),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf190d),
	.w1(32'h3cb250fe),
	.w2(32'h3caa1788),
	.w3(32'hbcf9873b),
	.w4(32'hb9131b0f),
	.w5(32'h3b0f01e1),
	.w6(32'h3c569fd0),
	.w7(32'hbb49cd73),
	.w8(32'hbd181b90),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09703d),
	.w1(32'h3bc5b32e),
	.w2(32'h3c0684e9),
	.w3(32'hbb9d1c67),
	.w4(32'h3bcf2d88),
	.w5(32'h3ae1e8f0),
	.w6(32'hbaf79b22),
	.w7(32'hbab7e2ca),
	.w8(32'h390f35df),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3917d6),
	.w1(32'hb799e826),
	.w2(32'hbab590d2),
	.w3(32'hba708ecd),
	.w4(32'hbbd58769),
	.w5(32'hbbfb5d02),
	.w6(32'hba0f2e7c),
	.w7(32'hbb968646),
	.w8(32'hbb0eb97e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1385a5),
	.w1(32'hbaf52d3f),
	.w2(32'hb9dd5843),
	.w3(32'hbc024150),
	.w4(32'h39fd51e7),
	.w5(32'h3a48e68e),
	.w6(32'h3b333e51),
	.w7(32'h3b74f0b3),
	.w8(32'h3be50377),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fb207),
	.w1(32'h3a9cc409),
	.w2(32'hbc162ae6),
	.w3(32'h3bab7f60),
	.w4(32'h3b171f37),
	.w5(32'h3b69db9f),
	.w6(32'hbae5a90e),
	.w7(32'hbc92d67d),
	.w8(32'hbbf918a9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabef20c),
	.w1(32'h3b81a758),
	.w2(32'h3b79dcae),
	.w3(32'h3bbeb825),
	.w4(32'hbb665166),
	.w5(32'hbb9ae158),
	.w6(32'h3c01d41e),
	.w7(32'h3c00dde0),
	.w8(32'h3b2d830c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa81f),
	.w1(32'h3b214519),
	.w2(32'hba473784),
	.w3(32'hbbe0dab3),
	.w4(32'hbaf72214),
	.w5(32'hbb192fa3),
	.w6(32'h3b8abdd0),
	.w7(32'hbc0c0901),
	.w8(32'hbbcce465),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf7ad6),
	.w1(32'hbb15e53b),
	.w2(32'hbb1cc56b),
	.w3(32'h3ac1b55d),
	.w4(32'hbb1d1c13),
	.w5(32'hbb160b22),
	.w6(32'h3a023bac),
	.w7(32'hbb3d07db),
	.w8(32'h3a8d25ed),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f10a0),
	.w1(32'hbaa191f4),
	.w2(32'hba2aaa1c),
	.w3(32'hbadaf767),
	.w4(32'h3bc4f2af),
	.w5(32'h3b9a77b3),
	.w6(32'h3b902975),
	.w7(32'hbb2f0ec3),
	.w8(32'h3b23cfcd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3b309),
	.w1(32'h3b73ab30),
	.w2(32'h3b50bcc1),
	.w3(32'hba42fcdd),
	.w4(32'h392d3126),
	.w5(32'hba4a8a09),
	.w6(32'h3afa86ed),
	.w7(32'h3b261d01),
	.w8(32'hbb015f1b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d104a),
	.w1(32'hba031c6f),
	.w2(32'hbb5959b2),
	.w3(32'hbbe48194),
	.w4(32'h3a3ebb28),
	.w5(32'h3ae6d653),
	.w6(32'hbb985f03),
	.w7(32'hbc25df7e),
	.w8(32'hbbd3d9ef),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbd8d3),
	.w1(32'h3aabb8a2),
	.w2(32'h3a1cf8f5),
	.w3(32'h3bc06853),
	.w4(32'h3c01a500),
	.w5(32'h3c1786e5),
	.w6(32'h3b0c22c1),
	.w7(32'h3b81605f),
	.w8(32'h3b534e48),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4fb50),
	.w1(32'h3b80b541),
	.w2(32'h3a8ef5e2),
	.w3(32'h3bea3cc6),
	.w4(32'h3b6cdb9a),
	.w5(32'h3b813794),
	.w6(32'hb9ebb2a8),
	.w7(32'hbc24a366),
	.w8(32'hbaa8f18d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f507e),
	.w1(32'hbb50cb5a),
	.w2(32'hba5216f8),
	.w3(32'hba2578c3),
	.w4(32'hbb4876bc),
	.w5(32'hbb1c4a97),
	.w6(32'hbbfd7b93),
	.w7(32'hbbabc38c),
	.w8(32'hbb9c97a3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64633d),
	.w1(32'h3be18b92),
	.w2(32'h3c19ee11),
	.w3(32'hb994b1bc),
	.w4(32'hbab183f8),
	.w5(32'h39fb4b0a),
	.w6(32'h3c01c69c),
	.w7(32'h3c20d2aa),
	.w8(32'hbb2f915d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec4af3),
	.w1(32'h3bafb920),
	.w2(32'h3c17029f),
	.w3(32'hbaabcc48),
	.w4(32'hbb3306fe),
	.w5(32'hbbaa847c),
	.w6(32'h3b03d2b9),
	.w7(32'h3c05e013),
	.w8(32'hbafb3f40),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed718),
	.w1(32'h3a957228),
	.w2(32'h3bf606d6),
	.w3(32'hbc03a22c),
	.w4(32'h3bb039ca),
	.w5(32'hba8ef46c),
	.w6(32'h3bb10585),
	.w7(32'h3c2ec6a3),
	.w8(32'h3b83b6db),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bddcb),
	.w1(32'h3b6734eb),
	.w2(32'h3b0932ad),
	.w3(32'hbb823651),
	.w4(32'hbbc999c5),
	.w5(32'hbc179321),
	.w6(32'hbb8a752f),
	.w7(32'hbbd1ce73),
	.w8(32'hbbb102d6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae59af1),
	.w1(32'h36db850c),
	.w2(32'hba48839d),
	.w3(32'hbc864a46),
	.w4(32'h3a650ed2),
	.w5(32'hbb5b3398),
	.w6(32'hb8dadab2),
	.w7(32'hba9309c2),
	.w8(32'hba1ad78c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc4181),
	.w1(32'h39d9239a),
	.w2(32'h3b82b5b9),
	.w3(32'hbad8483a),
	.w4(32'hba8a1fa2),
	.w5(32'h3a346df7),
	.w6(32'h3b59cd04),
	.w7(32'h3b96640f),
	.w8(32'h3af31608),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab00bc),
	.w1(32'h3b93442f),
	.w2(32'h3b065327),
	.w3(32'hbb4eb51a),
	.w4(32'hbb9455b5),
	.w5(32'h3bef406a),
	.w6(32'hbb2637e1),
	.w7(32'hba826e73),
	.w8(32'hbc0256cd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af857d1),
	.w1(32'h3ba82ea8),
	.w2(32'h3b9737d4),
	.w3(32'h3a338a48),
	.w4(32'h3a7ae7c9),
	.w5(32'h39c16b3d),
	.w6(32'h3ad91a9d),
	.w7(32'hbaa74fe6),
	.w8(32'h3b8c17c7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabf764),
	.w1(32'h3c314aa1),
	.w2(32'h3ae1d502),
	.w3(32'hbb0ab725),
	.w4(32'h395e95a4),
	.w5(32'hbb2010bc),
	.w6(32'h3c1d576a),
	.w7(32'h3bc131c1),
	.w8(32'hbbb848fb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa991b),
	.w1(32'hbbaa0d47),
	.w2(32'hbacbe1f6),
	.w3(32'hbade3bba),
	.w4(32'hbbce538f),
	.w5(32'hbbc6215d),
	.w6(32'hbb6eb158),
	.w7(32'hbb81ecc9),
	.w8(32'hbc00c896),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9f36c),
	.w1(32'h3c77a92d),
	.w2(32'h3c7ac866),
	.w3(32'h3b8f115a),
	.w4(32'h3c7581fa),
	.w5(32'h3c1d5da7),
	.w6(32'h3babd8f9),
	.w7(32'h3c476e6a),
	.w8(32'h3c2f8167),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f84f),
	.w1(32'h3c3357f7),
	.w2(32'h3b84c7f0),
	.w3(32'hbb8ed2b7),
	.w4(32'h3bd801a6),
	.w5(32'h3b22b5d9),
	.w6(32'h3a74ab18),
	.w7(32'hba8680f4),
	.w8(32'hb887cb74),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f1753),
	.w1(32'hbb15abff),
	.w2(32'h3abc1452),
	.w3(32'h3ba1a54e),
	.w4(32'hbb5c6e8f),
	.w5(32'h3b623595),
	.w6(32'hbb899f51),
	.w7(32'h3bcd3dd7),
	.w8(32'hbae0fb77),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb884c89),
	.w1(32'h3bd4ae75),
	.w2(32'h3c0d6cd6),
	.w3(32'hbb8f2cd5),
	.w4(32'h3b316ddf),
	.w5(32'hba84232f),
	.w6(32'hb9d27671),
	.w7(32'h3c4225d0),
	.w8(32'h3c0c559d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c719879),
	.w1(32'h3be79d51),
	.w2(32'h3bc05f78),
	.w3(32'hbac05f86),
	.w4(32'hbb0f54a7),
	.w5(32'hbb8c94d0),
	.w6(32'hbb194ce1),
	.w7(32'hbb713f57),
	.w8(32'hbc0f762d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd655),
	.w1(32'hbaf65439),
	.w2(32'hb97bf6c3),
	.w3(32'h3b5f0d9e),
	.w4(32'hbaa03d89),
	.w5(32'hbbf847e4),
	.w6(32'hbb0c982e),
	.w7(32'h3c622ce4),
	.w8(32'h3b148af7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb0686),
	.w1(32'h3b41432a),
	.w2(32'h3b1c50a5),
	.w3(32'hbbd24cfc),
	.w4(32'hbb2411b4),
	.w5(32'hbb61dccb),
	.w6(32'h3b125f7c),
	.w7(32'h3b97d288),
	.w8(32'h3b987ae6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba6df1),
	.w1(32'h3a2865cc),
	.w2(32'h3ac87ba9),
	.w3(32'hbc34cc62),
	.w4(32'hba99eb9e),
	.w5(32'hbb4e824a),
	.w6(32'hbaa5e181),
	.w7(32'h3ab12c41),
	.w8(32'h3b12eb51),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94020cf),
	.w1(32'h3c1ed955),
	.w2(32'h3bdcb09f),
	.w3(32'hbb5387eb),
	.w4(32'h3b1a81cd),
	.w5(32'h3b5971dd),
	.w6(32'hbb9790f9),
	.w7(32'h396da18f),
	.w8(32'hba97b14f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16aaa7),
	.w1(32'hbb9c0c93),
	.w2(32'hba46ac34),
	.w3(32'h3b6f82ab),
	.w4(32'hbb37d060),
	.w5(32'hbbefc5cb),
	.w6(32'hbb4ca2f5),
	.w7(32'h3bd6a330),
	.w8(32'hbab9e0db),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eaa0c),
	.w1(32'hbab00c00),
	.w2(32'h3bc42639),
	.w3(32'hbbc03289),
	.w4(32'h3bdadd78),
	.w5(32'h3c80f37d),
	.w6(32'hbc4dc8e4),
	.w7(32'hbc747dee),
	.w8(32'hbc38dd9a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132673),
	.w1(32'h3befb241),
	.w2(32'hbbbbb8aa),
	.w3(32'h3bcc46a9),
	.w4(32'h3c233fa5),
	.w5(32'h3c0ad3be),
	.w6(32'hbc148aff),
	.w7(32'hbcac5005),
	.w8(32'hbc94311d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb391e71),
	.w1(32'h3b73d3eb),
	.w2(32'h3b95a79f),
	.w3(32'h3c650d10),
	.w4(32'h3bc513fb),
	.w5(32'h39273d76),
	.w6(32'h3b587a3d),
	.w7(32'h3c167243),
	.w8(32'h3bd5e188),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42e706),
	.w1(32'h3b2e508b),
	.w2(32'h3b2fedca),
	.w3(32'h3aa74870),
	.w4(32'h3b3cc40a),
	.w5(32'hba1485ec),
	.w6(32'hbad33c01),
	.w7(32'hb98751da),
	.w8(32'h3aeee464),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3f2ea),
	.w1(32'hbaee74d3),
	.w2(32'hbb63b5d1),
	.w3(32'hb8327086),
	.w4(32'h3b28497b),
	.w5(32'h3b115821),
	.w6(32'hbbdbaa74),
	.w7(32'hbc4cfe85),
	.w8(32'hba2302b1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fe462),
	.w1(32'h3bba5493),
	.w2(32'h3c551040),
	.w3(32'hba2b67ac),
	.w4(32'hbbd59c3c),
	.w5(32'h3b6535db),
	.w6(32'h3bbd6193),
	.w7(32'h3aca2d80),
	.w8(32'hbbafe8c0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38abed),
	.w1(32'h3b4c57cc),
	.w2(32'h3be0446a),
	.w3(32'h3b89eedb),
	.w4(32'hbb5fb1a9),
	.w5(32'h3b80c460),
	.w6(32'hbbc09c85),
	.w7(32'hbbafcbb3),
	.w8(32'hbb77dac9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ac1a7),
	.w1(32'hbb907df8),
	.w2(32'h3a599c9b),
	.w3(32'h39ba54ce),
	.w4(32'hbbd897a2),
	.w5(32'hbb2cdc1c),
	.w6(32'h3af742e7),
	.w7(32'hba8d64e4),
	.w8(32'h3b72cb09),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb791dd),
	.w1(32'h3c07c4d4),
	.w2(32'h3c14e784),
	.w3(32'hbb098642),
	.w4(32'h3b62745b),
	.w5(32'hb9e43877),
	.w6(32'hba6df2ff),
	.w7(32'hb9dc8038),
	.w8(32'hbb1b0e98),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98c83c),
	.w1(32'hbaf2ab46),
	.w2(32'hbb8a7c2b),
	.w3(32'hbab94c35),
	.w4(32'h3a22ed98),
	.w5(32'h3b381b5d),
	.w6(32'hbb6fa60b),
	.w7(32'hbb2d2deb),
	.w8(32'h3ba59b6e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17c60a),
	.w1(32'h3be7bb12),
	.w2(32'h3bc4c1ab),
	.w3(32'h3af884d9),
	.w4(32'hb9e7a531),
	.w5(32'h3b3787ba),
	.w6(32'hbaed43f8),
	.w7(32'h3b099b99),
	.w8(32'h3ad913a4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b980764),
	.w1(32'h3bbe98a1),
	.w2(32'h3c53b97b),
	.w3(32'h3a137590),
	.w4(32'hb9db4a0d),
	.w5(32'h3b315d8f),
	.w6(32'h3bb332ea),
	.w7(32'h3be144c6),
	.w8(32'h3c0c61ad),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be898b6),
	.w1(32'h39a0071c),
	.w2(32'h3ad73252),
	.w3(32'h3aff09ff),
	.w4(32'hbab91917),
	.w5(32'hbbad5ed6),
	.w6(32'hbb9183d8),
	.w7(32'hba86aa90),
	.w8(32'h3a2e6721),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70ffc6),
	.w1(32'h39baf24c),
	.w2(32'h3c6bc029),
	.w3(32'h3acf3c80),
	.w4(32'h3a132fe2),
	.w5(32'h3bca55c1),
	.w6(32'hbb6c53c4),
	.w7(32'h3be98da2),
	.w8(32'h3be30729),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61f015),
	.w1(32'h3a986ba7),
	.w2(32'h3bbb8956),
	.w3(32'h3b9cf0d5),
	.w4(32'h3b542a26),
	.w5(32'h3b4adcdf),
	.w6(32'h3b26ab9a),
	.w7(32'hb9f9bb59),
	.w8(32'hbb1e2fa8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac0fc),
	.w1(32'hbb15b4ea),
	.w2(32'h3af37590),
	.w3(32'hbba76d0e),
	.w4(32'hbb93b761),
	.w5(32'hbbe29f1f),
	.w6(32'h3b1284bb),
	.w7(32'h3c0a7e82),
	.w8(32'h3b5a38c7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215763),
	.w1(32'h3c596047),
	.w2(32'h3c43935f),
	.w3(32'hbbbe5829),
	.w4(32'hba9e93c1),
	.w5(32'hbbcf179a),
	.w6(32'h3c34a132),
	.w7(32'h3c694e50),
	.w8(32'h3aec0c2b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6eeb26),
	.w1(32'h3ac3b604),
	.w2(32'h3a8df303),
	.w3(32'hbc270f15),
	.w4(32'hbb6f5050),
	.w5(32'hbc01e8b6),
	.w6(32'h3bd4fea6),
	.w7(32'h3bfaa252),
	.w8(32'h3bf40642),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c96ae),
	.w1(32'h39d55699),
	.w2(32'h3c085ed3),
	.w3(32'hbc45ca3e),
	.w4(32'hbaf38806),
	.w5(32'h3b990b81),
	.w6(32'h3b03631b),
	.w7(32'h3b64744c),
	.w8(32'h3b2aa555),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c022c30),
	.w1(32'h3b87c629),
	.w2(32'h3ade5a95),
	.w3(32'h3a54a8b2),
	.w4(32'h3b8e54ea),
	.w5(32'h3aa3d976),
	.w6(32'h3b385471),
	.w7(32'h3c00971f),
	.w8(32'h3c1c4ebb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec3603),
	.w1(32'h3ac35056),
	.w2(32'hba66d57b),
	.w3(32'hbab752f9),
	.w4(32'hbb64d342),
	.w5(32'h3bb00834),
	.w6(32'hbba6c5d5),
	.w7(32'hbbaf45d1),
	.w8(32'hbbf54097),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98701f9),
	.w1(32'h3a713ee5),
	.w2(32'h3b91d1f8),
	.w3(32'hbb12a953),
	.w4(32'h3b246446),
	.w5(32'hbba74d94),
	.w6(32'hbb8c8dfb),
	.w7(32'hbad4815c),
	.w8(32'hbb5e4401),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ed44d),
	.w1(32'h39edbcbf),
	.w2(32'h3c1eeeb7),
	.w3(32'hbbc73457),
	.w4(32'hbb666696),
	.w5(32'h3ae09852),
	.w6(32'hbafe83cf),
	.w7(32'h3c0fa652),
	.w8(32'h3bd07eb6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2ef0c),
	.w1(32'h3c6df2c7),
	.w2(32'h3c390f82),
	.w3(32'hbab3d8a8),
	.w4(32'h3aa82d77),
	.w5(32'hbb798413),
	.w6(32'hbb3c9e72),
	.w7(32'h38762d7b),
	.w8(32'hbba779a9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf3b4d),
	.w1(32'h3b72927a),
	.w2(32'hbb91d5b1),
	.w3(32'hba579ce7),
	.w4(32'h3aec4984),
	.w5(32'h3ba3058b),
	.w6(32'hbb87f92e),
	.w7(32'hbc275ca7),
	.w8(32'hbc066a9d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c298),
	.w1(32'hbba4a8a8),
	.w2(32'hbc2a0ef4),
	.w3(32'hb9a1c8eb),
	.w4(32'hbb313341),
	.w5(32'hbc084170),
	.w6(32'hb9e000c0),
	.w7(32'hbb309434),
	.w8(32'hbb01400a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe720d4),
	.w1(32'h3b27e4e7),
	.w2(32'h3b13f14f),
	.w3(32'hbba29645),
	.w4(32'h3b6d401f),
	.w5(32'hbb9fae1b),
	.w6(32'h3b9430ab),
	.w7(32'h3c60259b),
	.w8(32'h3c3ca4a2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24eb4),
	.w1(32'hb9db5838),
	.w2(32'hbb43bf25),
	.w3(32'hbc063c18),
	.w4(32'hbb0e0f45),
	.w5(32'hbb9b2c81),
	.w6(32'h3951ce5b),
	.w7(32'h3ac21241),
	.w8(32'h3b22fea0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66ce3e),
	.w1(32'hb9d7095e),
	.w2(32'h3b06d344),
	.w3(32'hbb3bdb21),
	.w4(32'hbbdd9e23),
	.w5(32'hbbd41a69),
	.w6(32'h3ae63483),
	.w7(32'h3bfa0c72),
	.w8(32'h3be4f862),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf43fc),
	.w1(32'h3ba3793d),
	.w2(32'h3b3ae31d),
	.w3(32'hbbedb16a),
	.w4(32'h3ba67f5f),
	.w5(32'h3be74b25),
	.w6(32'h3b2245a0),
	.w7(32'h3b844308),
	.w8(32'h3b2b5fe9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe044d),
	.w1(32'hb9c13d99),
	.w2(32'hba96013d),
	.w3(32'h3b8549ab),
	.w4(32'hbac75540),
	.w5(32'hbb22f8af),
	.w6(32'hbb3077c7),
	.w7(32'hbac2e415),
	.w8(32'h3a273509),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8c654),
	.w1(32'h3b172dcf),
	.w2(32'h3a405e7b),
	.w3(32'h3afbeb9c),
	.w4(32'h37c263fa),
	.w5(32'hbacbed1e),
	.w6(32'h3b8e34d1),
	.w7(32'h3bb63eb9),
	.w8(32'h3a8db44a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c77b3),
	.w1(32'h3b85ea4c),
	.w2(32'h3b8dafcd),
	.w3(32'hba55a88a),
	.w4(32'hb914cd32),
	.w5(32'hbb081986),
	.w6(32'h3b2d3eef),
	.w7(32'h3b89bda9),
	.w8(32'h3af56fa3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b0c76),
	.w1(32'h3b5c7b6a),
	.w2(32'h3b6dc0a4),
	.w3(32'hbbbc3795),
	.w4(32'hbb4f5e5e),
	.w5(32'hbc15a0f5),
	.w6(32'h3ba77afb),
	.w7(32'h3c01c77e),
	.w8(32'h3b94180d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e200),
	.w1(32'h3ad47856),
	.w2(32'hbb3816e6),
	.w3(32'hbc0384d5),
	.w4(32'hbaf6a36e),
	.w5(32'hbbc9a177),
	.w6(32'h3b91a0be),
	.w7(32'h3b332948),
	.w8(32'hbb407ca7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ba8b),
	.w1(32'h3c76a91e),
	.w2(32'h3ba8a58e),
	.w3(32'hbb8926f9),
	.w4(32'h3aa891f3),
	.w5(32'hb80a38f9),
	.w6(32'h3b34db31),
	.w7(32'h3b93313f),
	.w8(32'h3b5d64c6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a073d71),
	.w1(32'h3bdedd3a),
	.w2(32'h3c23c006),
	.w3(32'hba95cd8d),
	.w4(32'h3c110edf),
	.w5(32'h3be53903),
	.w6(32'h3a27151d),
	.w7(32'h3beaaef6),
	.w8(32'hba70bc30),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bf432),
	.w1(32'hba019bad),
	.w2(32'h3add223f),
	.w3(32'hbaf9f8c4),
	.w4(32'hbb9368d3),
	.w5(32'hbb96b542),
	.w6(32'h3a6b3d73),
	.w7(32'h3b9c4917),
	.w8(32'h3b6bdaa0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bc0ff),
	.w1(32'h3a7fc32f),
	.w2(32'h3b2fc922),
	.w3(32'h3b2be549),
	.w4(32'hbbd7b8cc),
	.w5(32'hbc231b5f),
	.w6(32'h391e98a3),
	.w7(32'h3baff21f),
	.w8(32'hbb16c145),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf50bd),
	.w1(32'hbb07eddc),
	.w2(32'hb90b0e21),
	.w3(32'hbc658a48),
	.w4(32'h3a53d6db),
	.w5(32'h3b46774d),
	.w6(32'hba13b31c),
	.w7(32'hbc24955a),
	.w8(32'hbb8b8fe3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43c2c6),
	.w1(32'h3ac89af8),
	.w2(32'h3bc912ce),
	.w3(32'hbb9ae25e),
	.w4(32'hbc5e4e3a),
	.w5(32'hbc8eb3cc),
	.w6(32'h3a80f485),
	.w7(32'h3c4cf307),
	.w8(32'h3b543255),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231639),
	.w1(32'h39710a18),
	.w2(32'h3ba91636),
	.w3(32'hbc554b00),
	.w4(32'h39aaaaab),
	.w5(32'h3809cbf6),
	.w6(32'hbb0fbe46),
	.w7(32'h3babe84d),
	.w8(32'h3b68d807),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd777e1),
	.w1(32'hba5c7e67),
	.w2(32'hba8c435d),
	.w3(32'h3a231dcb),
	.w4(32'hbb08bac4),
	.w5(32'hbbebcad0),
	.w6(32'hbbe453a4),
	.w7(32'hbbcb4248),
	.w8(32'hbc03de77),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1486a5),
	.w1(32'h3ba0bcbf),
	.w2(32'h3c0ef539),
	.w3(32'hbb138cf1),
	.w4(32'hbb8fbaa7),
	.w5(32'h3a1026b8),
	.w6(32'hbadb604e),
	.w7(32'h3befced7),
	.w8(32'h3bd168b5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b3098),
	.w1(32'h3c0c7ca6),
	.w2(32'h3a79caeb),
	.w3(32'hbb8537aa),
	.w4(32'h3b8a6abf),
	.w5(32'h398ce9c9),
	.w6(32'hbb4e2041),
	.w7(32'hbbbd086a),
	.w8(32'hbba4825d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a075767),
	.w1(32'hbb4eed21),
	.w2(32'hbc42b789),
	.w3(32'hbb411bdc),
	.w4(32'hbbc6809a),
	.w5(32'hbc850e4b),
	.w6(32'h3a7cd95a),
	.w7(32'h3b10140f),
	.w8(32'hbad38d34),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d1b9b),
	.w1(32'h3c3b0fb2),
	.w2(32'h3c5ede48),
	.w3(32'hbbffcf4f),
	.w4(32'h3b4a0599),
	.w5(32'hb919c99a),
	.w6(32'h3bb9d21c),
	.w7(32'h3c0cbf6f),
	.w8(32'h3b399b15),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e688),
	.w1(32'hbab1ed56),
	.w2(32'hbb95aa54),
	.w3(32'hbb7c90e1),
	.w4(32'hbaba2726),
	.w5(32'h3b9233e8),
	.w6(32'hbb328dd4),
	.w7(32'hbbddb4de),
	.w8(32'hbb734341),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5e6f5),
	.w1(32'h3b85f799),
	.w2(32'h3aaa0676),
	.w3(32'h3b811246),
	.w4(32'hba2632e6),
	.w5(32'hba63bfee),
	.w6(32'h3b0f2d17),
	.w7(32'hbb1f6d87),
	.w8(32'hbb4aa63f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e67c8),
	.w1(32'hbabed65c),
	.w2(32'hbb5176b2),
	.w3(32'h3ac8dcfa),
	.w4(32'hbba54b67),
	.w5(32'h3b142693),
	.w6(32'h3ad29706),
	.w7(32'hba467c1e),
	.w8(32'hba1c7283),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1d149),
	.w1(32'h3ac68e09),
	.w2(32'h3abe2b55),
	.w3(32'h3b8e37c3),
	.w4(32'hb7dd0a8b),
	.w5(32'hbacab2b4),
	.w6(32'h3b309ffa),
	.w7(32'h3af307b5),
	.w8(32'h3b9d91d7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2414d4),
	.w1(32'h3bba9daa),
	.w2(32'h3b989c78),
	.w3(32'hbb6550a9),
	.w4(32'hb98c0815),
	.w5(32'h3b752ace),
	.w6(32'h3bad9c9f),
	.w7(32'h3b86642a),
	.w8(32'h3aa08cc7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c056c22),
	.w1(32'h3c373920),
	.w2(32'h3c845fbb),
	.w3(32'h3b80212a),
	.w4(32'hbbdcfbfb),
	.w5(32'h3a159583),
	.w6(32'h3b92955b),
	.w7(32'h3c7c19e7),
	.w8(32'h3c432c34),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c1782),
	.w1(32'hbb1a4736),
	.w2(32'hbb3bec68),
	.w3(32'hbc1f43cf),
	.w4(32'hbb3f1d84),
	.w5(32'hbaf8b193),
	.w6(32'hbb29f2e5),
	.w7(32'hbb3f4bca),
	.w8(32'hbb71de52),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08118c),
	.w1(32'h3b7604a0),
	.w2(32'h3ae65b49),
	.w3(32'hbb2f3dae),
	.w4(32'h3ae2d6ea),
	.w5(32'h3999cedd),
	.w6(32'h3aeb218b),
	.w7(32'h3a58d5d3),
	.w8(32'h3acd352d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219f34),
	.w1(32'hbb8ce2d6),
	.w2(32'hbb8e78a2),
	.w3(32'h3adcccf2),
	.w4(32'hbbdb4b8d),
	.w5(32'hbbb6c804),
	.w6(32'hbb2ab973),
	.w7(32'hbb8e604f),
	.w8(32'hbc020810),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a7014),
	.w1(32'h3bc5fb7e),
	.w2(32'h3a89ee41),
	.w3(32'hbc179eba),
	.w4(32'h3b8e564a),
	.w5(32'hba84bda2),
	.w6(32'h3b23c5f3),
	.w7(32'hba958a37),
	.w8(32'h3afacfd4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee28e3),
	.w1(32'h3b671199),
	.w2(32'h3bbf05a7),
	.w3(32'hb9232291),
	.w4(32'hbbad9ed3),
	.w5(32'hbba1a3f3),
	.w6(32'h3c05c9e2),
	.w7(32'h3c535359),
	.w8(32'h3b7d5f72),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814757),
	.w1(32'hb9bd2041),
	.w2(32'h3b90d98c),
	.w3(32'hbbe8b4a2),
	.w4(32'hbb66042e),
	.w5(32'hbaf870e7),
	.w6(32'h3bad46ae),
	.w7(32'h3ba7be3f),
	.w8(32'h3b7b01e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e14f9),
	.w1(32'h3b35582a),
	.w2(32'h3ac638fb),
	.w3(32'hbb99f7d7),
	.w4(32'h3af41a8c),
	.w5(32'hbb873151),
	.w6(32'hba96adfc),
	.w7(32'h3c01f6d9),
	.w8(32'h3b4880ed),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b976814),
	.w1(32'hba548ad4),
	.w2(32'h3b8f4438),
	.w3(32'hbb42e407),
	.w4(32'hbb7fb1fd),
	.w5(32'hbbd865ef),
	.w6(32'hbadb301b),
	.w7(32'h3bc467a9),
	.w8(32'h3bae719c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a244b),
	.w1(32'hbac5221a),
	.w2(32'h39114beb),
	.w3(32'hbbb734aa),
	.w4(32'hbb47ec44),
	.w5(32'hbba760f4),
	.w6(32'h3b1d176b),
	.w7(32'h3b8f22f2),
	.w8(32'h3b558a99),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc861),
	.w1(32'h3ab839f5),
	.w2(32'h38ad848f),
	.w3(32'hbbbbedbe),
	.w4(32'h3bf846e4),
	.w5(32'h3b3413e3),
	.w6(32'h3bc80fb6),
	.w7(32'hba137d58),
	.w8(32'h3ab17392),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8533ae),
	.w1(32'h3b502845),
	.w2(32'h3b38e02e),
	.w3(32'h38a2b8ce),
	.w4(32'hbb44dc37),
	.w5(32'hbbc51887),
	.w6(32'h3b822053),
	.w7(32'h3b15d89b),
	.w8(32'h3b225fe4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5df29),
	.w1(32'h3b87030e),
	.w2(32'h3c213967),
	.w3(32'hbbcf2502),
	.w4(32'h3bed1146),
	.w5(32'h39c29f2a),
	.w6(32'h3b439db5),
	.w7(32'h3bc14a03),
	.w8(32'h3bc379e9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30440e),
	.w1(32'hba1b3918),
	.w2(32'hbb3ad390),
	.w3(32'h3bd5dddc),
	.w4(32'hbb27f942),
	.w5(32'hbb44d789),
	.w6(32'hbaebad6f),
	.w7(32'hbb455bb4),
	.w8(32'hbb8733d5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28fe01),
	.w1(32'hbc174588),
	.w2(32'h3a6def00),
	.w3(32'hbabc78c5),
	.w4(32'hbc35a9d2),
	.w5(32'h3b6b0ce4),
	.w6(32'hbc55ed8a),
	.w7(32'hbb73772b),
	.w8(32'hbb00c143),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule