module layer_10_featuremap_205(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51caf1),
	.w1(32'h3a6b1ee8),
	.w2(32'h3a6d12da),
	.w3(32'h3a25ebd3),
	.w4(32'hb8ee8203),
	.w5(32'h3ab7f2b1),
	.w6(32'h39114de7),
	.w7(32'hb9ea532d),
	.w8(32'h390698ab),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fef31),
	.w1(32'hb96371e6),
	.w2(32'hb9d819a0),
	.w3(32'h3a8f0d0d),
	.w4(32'h38c82744),
	.w5(32'hba616344),
	.w6(32'hb9d7b8d7),
	.w7(32'hb91de601),
	.w8(32'hba8c58ef),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad87395),
	.w1(32'hbad82928),
	.w2(32'hbac0b091),
	.w3(32'hbaf34b7f),
	.w4(32'hbab7eb14),
	.w5(32'hbacbb6fa),
	.w6(32'hba912f07),
	.w7(32'hbab74fd1),
	.w8(32'hbae0d320),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac943f1),
	.w1(32'hbaf48af1),
	.w2(32'hbab3af7b),
	.w3(32'hbb0058ad),
	.w4(32'hba80675c),
	.w5(32'hba72298c),
	.w6(32'hba20ab18),
	.w7(32'hba5a8f0e),
	.w8(32'hba9d664d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3ccaf),
	.w1(32'h3b10b459),
	.w2(32'h377cb565),
	.w3(32'hba7fd71b),
	.w4(32'h3b27ba59),
	.w5(32'h3ad617fd),
	.w6(32'h3b14c6c2),
	.w7(32'hb958ef4f),
	.w8(32'h38ba7a6d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebbb3a),
	.w1(32'hb931ab79),
	.w2(32'h3a8d4d3f),
	.w3(32'h3a7f0556),
	.w4(32'hb9945f54),
	.w5(32'h3a56d54f),
	.w6(32'h39a04a54),
	.w7(32'h3a75cdc3),
	.w8(32'h3a7d5d3d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6afc4),
	.w1(32'hbb03d695),
	.w2(32'hbaedfcaa),
	.w3(32'hb96cdada),
	.w4(32'hbac29595),
	.w5(32'hba6963dd),
	.w6(32'hb9cbe55e),
	.w7(32'hba08cf3a),
	.w8(32'h37b2aa80),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32315e),
	.w1(32'h3af91246),
	.w2(32'h3b070ce4),
	.w3(32'h3acbc9c5),
	.w4(32'h3b0a612e),
	.w5(32'h3b16370c),
	.w6(32'h3b216603),
	.w7(32'h3b042360),
	.w8(32'hb972a14f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a671ec9),
	.w1(32'h38ca2618),
	.w2(32'h398b38d7),
	.w3(32'h3a1d83b4),
	.w4(32'h39cb2cd5),
	.w5(32'h3a261ba1),
	.w6(32'h3999faca),
	.w7(32'h39737aa4),
	.w8(32'h35ed1522),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d8261),
	.w1(32'hba45badf),
	.w2(32'hb95bf187),
	.w3(32'h394f2b5f),
	.w4(32'hbaa16714),
	.w5(32'hba34bbd9),
	.w6(32'hbab58208),
	.w7(32'hbad254a4),
	.w8(32'hb7486a18),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0191),
	.w1(32'hbabe1379),
	.w2(32'hbaa6aa95),
	.w3(32'hbac514ad),
	.w4(32'hbb102522),
	.w5(32'hbb1b1c7c),
	.w6(32'hb919b184),
	.w7(32'hba917e23),
	.w8(32'hba420a90),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf264b),
	.w1(32'hbb8c3474),
	.w2(32'hbb13bed1),
	.w3(32'hbb118719),
	.w4(32'hbb66e46d),
	.w5(32'hbadcac34),
	.w6(32'h3aa31b8b),
	.w7(32'h3a2a28ef),
	.w8(32'h38d5eddf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba191ec1),
	.w1(32'hb7cbc7af),
	.w2(32'h3a339821),
	.w3(32'hba7b471e),
	.w4(32'hbadb8527),
	.w5(32'hb9383c00),
	.w6(32'hb9b82e4e),
	.w7(32'hba7a57b5),
	.w8(32'h39c89e13),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d574f),
	.w1(32'hb9ed3004),
	.w2(32'hba7293b5),
	.w3(32'hb9f937ba),
	.w4(32'hba1bdca8),
	.w5(32'hba4627d3),
	.w6(32'h39468c4f),
	.w7(32'h3a38c524),
	.w8(32'h39dacf74),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51fd88),
	.w1(32'hbadcc0ee),
	.w2(32'hbac63b89),
	.w3(32'hba222e8a),
	.w4(32'hbabfc33e),
	.w5(32'hba84ca16),
	.w6(32'hb9ae5f6e),
	.w7(32'h39254b6e),
	.w8(32'hba93b3bc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1462),
	.w1(32'h3a97014b),
	.w2(32'h3af16855),
	.w3(32'hb9e45232),
	.w4(32'h3a68bf18),
	.w5(32'h3aa3f981),
	.w6(32'h3a9a7373),
	.w7(32'h3ab32389),
	.w8(32'h3a3dd7c4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39096624),
	.w1(32'h38e84efb),
	.w2(32'h3a82129e),
	.w3(32'h3a000768),
	.w4(32'h3a35713c),
	.w5(32'hb86d88ee),
	.w6(32'h3a02c12b),
	.w7(32'h3a9ab241),
	.w8(32'h3a765159),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e9245),
	.w1(32'hbb1d9324),
	.w2(32'hba505a4a),
	.w3(32'h3b0829ed),
	.w4(32'hbaa3c5d8),
	.w5(32'h3a3e6a49),
	.w6(32'h3a9332f1),
	.w7(32'hbaba3180),
	.w8(32'hb9ced838),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1438c),
	.w1(32'hba7d8491),
	.w2(32'h391d5025),
	.w3(32'hbad5ae79),
	.w4(32'hba8a7fc2),
	.w5(32'h38fe6c10),
	.w6(32'h39ecdf85),
	.w7(32'hba2ce699),
	.w8(32'hb98ff3f4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ff2dc),
	.w1(32'h38e56f31),
	.w2(32'h39f5cf62),
	.w3(32'hba5dba4c),
	.w4(32'hb899c632),
	.w5(32'h38b46a81),
	.w6(32'h38b0d326),
	.w7(32'h393a85e9),
	.w8(32'h38a5fbd8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39680844),
	.w1(32'h38a5b9c4),
	.w2(32'h3a5511b9),
	.w3(32'h39254426),
	.w4(32'hb945542e),
	.w5(32'h3a22bf77),
	.w6(32'hba049ed4),
	.w7(32'hb928b0e0),
	.w8(32'hba1c6090),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8021c32),
	.w1(32'hbb2e9e01),
	.w2(32'hbb442cd3),
	.w3(32'hb9db38af),
	.w4(32'hbb4d36a9),
	.w5(32'hbae916d8),
	.w6(32'hbb382399),
	.w7(32'hbad50240),
	.w8(32'hbafea748),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53e112),
	.w1(32'hbb0082a7),
	.w2(32'h3b0aaaeb),
	.w3(32'hba31dbf8),
	.w4(32'hbac45657),
	.w5(32'hb85cc0a7),
	.w6(32'h3b58373b),
	.w7(32'h3b10c099),
	.w8(32'h3b0f9a45),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51e0ea),
	.w1(32'h3b0b522e),
	.w2(32'h3b1a6cbe),
	.w3(32'hb932732e),
	.w4(32'h3a2e3e99),
	.w5(32'h3a980417),
	.w6(32'h3a8619c1),
	.w7(32'h3aaa37ad),
	.w8(32'h3ab2063a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d5881),
	.w1(32'h3a219dfd),
	.w2(32'h3aa3c9f6),
	.w3(32'h39f85d96),
	.w4(32'hb9a71396),
	.w5(32'hb99e977e),
	.w6(32'hb9e2c195),
	.w7(32'hb8cc4391),
	.w8(32'hb9e501c1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba747b22),
	.w1(32'hb8a0155a),
	.w2(32'hb9de2b87),
	.w3(32'hba4363e1),
	.w4(32'hba33146c),
	.w5(32'hb9827c6f),
	.w6(32'h38348e7d),
	.w7(32'h3a8e3201),
	.w8(32'h3a701ccd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a942c29),
	.w1(32'hb98620cc),
	.w2(32'h399306df),
	.w3(32'h399524bd),
	.w4(32'hb9a05bcc),
	.w5(32'h391543a1),
	.w6(32'hb9995e36),
	.w7(32'hb8d8d682),
	.w8(32'hb97c47f1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c27ea),
	.w1(32'hbb843d5a),
	.w2(32'hbaae3d86),
	.w3(32'hbaa9a377),
	.w4(32'hbb682e53),
	.w5(32'hbaf8c2fe),
	.w6(32'hbb5ab834),
	.w7(32'hbb21c2ec),
	.w8(32'hbb3e5580),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24012),
	.w1(32'hbb22b7c4),
	.w2(32'hb9cc5e7d),
	.w3(32'hbabe5b4d),
	.w4(32'hbb18b53e),
	.w5(32'hba746b5b),
	.w6(32'hbb329c8c),
	.w7(32'hbab5deae),
	.w8(32'hba0f72a5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953fde6),
	.w1(32'hbad9e025),
	.w2(32'hbabcef79),
	.w3(32'hba2562b3),
	.w4(32'hba9de89a),
	.w5(32'hbaa37b87),
	.w6(32'hbaada053),
	.w7(32'hb9a1005f),
	.w8(32'h3a1e10a8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98900c2),
	.w1(32'hb91e7fbf),
	.w2(32'h39a81513),
	.w3(32'hb8b5f7a2),
	.w4(32'hb9122c31),
	.w5(32'h390a14a2),
	.w6(32'hba14f38c),
	.w7(32'hba05c371),
	.w8(32'hba3701ce),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae73eb),
	.w1(32'hba05f40b),
	.w2(32'hb9d3f7ed),
	.w3(32'hb91092a0),
	.w4(32'hba4f535d),
	.w5(32'hba08cb86),
	.w6(32'hba111f17),
	.w7(32'hba453821),
	.w8(32'hba52d206),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e108fa),
	.w1(32'h3982ba9b),
	.w2(32'hba1c0396),
	.w3(32'hba0bc911),
	.w4(32'hb86057d1),
	.w5(32'h37024354),
	.w6(32'h3a25b091),
	.w7(32'hba0521dd),
	.w8(32'hb9a18298),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6df78),
	.w1(32'h38878b32),
	.w2(32'h3a232214),
	.w3(32'hba91e385),
	.w4(32'hb8e4349f),
	.w5(32'h3a340c3a),
	.w6(32'h39dfe30e),
	.w7(32'h3a4f7bfe),
	.w8(32'h3ab6e01b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7395c6),
	.w1(32'hbaf74f73),
	.w2(32'hba82b74c),
	.w3(32'h39ed0d09),
	.w4(32'hba4677bf),
	.w5(32'hba8e4017),
	.w6(32'hbaf1fe28),
	.w7(32'hbb00b4c1),
	.w8(32'hba8deb52),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f982a),
	.w1(32'hba5ab46e),
	.w2(32'hb950497c),
	.w3(32'hba9bfe69),
	.w4(32'hbad1306f),
	.w5(32'hba37892a),
	.w6(32'hba1c2b0f),
	.w7(32'hba86a9c0),
	.w8(32'hba88a4c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4b95),
	.w1(32'hba2cd607),
	.w2(32'hbb113378),
	.w3(32'h3b978f3a),
	.w4(32'hba12a34f),
	.w5(32'hbbb26767),
	.w6(32'h3ba2b296),
	.w7(32'hbaeff638),
	.w8(32'hbb95d274),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4093b3),
	.w1(32'hba3dbaff),
	.w2(32'hba82610b),
	.w3(32'hbb589df1),
	.w4(32'hbaa7eca3),
	.w5(32'hbb048ac1),
	.w6(32'hba8fcedb),
	.w7(32'hba9edc5a),
	.w8(32'hbb128477),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48b449),
	.w1(32'hbad0f81c),
	.w2(32'hba86dcff),
	.w3(32'hbb309932),
	.w4(32'hbabd4651),
	.w5(32'hba0da74b),
	.w6(32'h3a0af0e7),
	.w7(32'h3aa885b7),
	.w8(32'h39c9d641),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fc991),
	.w1(32'hb985bc0f),
	.w2(32'hb9e5c679),
	.w3(32'h3a296dd1),
	.w4(32'hb736b491),
	.w5(32'hb9b1fcd8),
	.w6(32'hb922810a),
	.w7(32'hb9f73779),
	.w8(32'hba517a09),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43d576),
	.w1(32'hba0970d0),
	.w2(32'hbab712d7),
	.w3(32'hba65a596),
	.w4(32'hba131ab4),
	.w5(32'hba8ca481),
	.w6(32'hba2195db),
	.w7(32'hba8b984f),
	.w8(32'hb9e5f9d5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ee568),
	.w1(32'hbadd0c8f),
	.w2(32'hbae55955),
	.w3(32'hb9e386ec),
	.w4(32'hbaf65794),
	.w5(32'hbb1549f7),
	.w6(32'hba820f88),
	.w7(32'hba8fbfdd),
	.w8(32'hbad38ed5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9060),
	.w1(32'hbaaff88c),
	.w2(32'hba8982d9),
	.w3(32'hbb2aa7ee),
	.w4(32'hbaaef768),
	.w5(32'hba86b333),
	.w6(32'hba517a44),
	.w7(32'hba60bb6b),
	.w8(32'hba5a935e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c181d),
	.w1(32'hba913cf3),
	.w2(32'hbab52178),
	.w3(32'h3919e2d2),
	.w4(32'hb9db080a),
	.w5(32'h3892db8c),
	.w6(32'h3ac2f0ba),
	.w7(32'hba39fc29),
	.w8(32'h3afba362),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff334e),
	.w1(32'h3b09bbc5),
	.w2(32'h38e281d2),
	.w3(32'hba370b2d),
	.w4(32'h3af223c8),
	.w5(32'h3a272152),
	.w6(32'hb94bfa79),
	.w7(32'h38837a01),
	.w8(32'h3a185e9e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa16f70),
	.w1(32'h3af74ac2),
	.w2(32'h3b0d4f93),
	.w3(32'h382f69d1),
	.w4(32'h39a45e16),
	.w5(32'h3ab12b0b),
	.w6(32'h3a0000d2),
	.w7(32'h3a92bdbb),
	.w8(32'h3a42da02),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a462969),
	.w1(32'h3834ef68),
	.w2(32'hba99bd53),
	.w3(32'h3a83e87f),
	.w4(32'h3a02a088),
	.w5(32'h3a2a6b02),
	.w6(32'h3ae4f6f4),
	.w7(32'h3a5ee185),
	.w8(32'hb9b14881),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63dbfd),
	.w1(32'hbaf97789),
	.w2(32'h3a263c39),
	.w3(32'h3ad41e8d),
	.w4(32'hbb18a20e),
	.w5(32'h39bde373),
	.w6(32'h3ac6b3af),
	.w7(32'h39b0cf3d),
	.w8(32'h3a81605b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ed87f),
	.w1(32'hba042382),
	.w2(32'hb8f12a00),
	.w3(32'h3a4a43f5),
	.w4(32'hba28814b),
	.w5(32'hb961f209),
	.w6(32'hb9486743),
	.w7(32'hb912085f),
	.w8(32'h383a5706),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c8c63),
	.w1(32'h3a2478c9),
	.w2(32'h39c5b642),
	.w3(32'hb931f938),
	.w4(32'h39cad768),
	.w5(32'h398cd639),
	.w6(32'h3a5b4e4c),
	.w7(32'h3a452788),
	.w8(32'h39dbc577),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8d2a4),
	.w1(32'hb9ea1e7c),
	.w2(32'h38805c84),
	.w3(32'h3924e5f2),
	.w4(32'h3969a242),
	.w5(32'h39969f28),
	.w6(32'h38ee4aa1),
	.w7(32'h372b18d2),
	.w8(32'hba43bc0e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2f031),
	.w1(32'h3a1272fc),
	.w2(32'h3a956332),
	.w3(32'h39023eed),
	.w4(32'hba7431d3),
	.w5(32'h39094042),
	.w6(32'hb9e7a73f),
	.w7(32'hba87cfb4),
	.w8(32'hbac5d9be),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc50d8),
	.w1(32'hba3b0750),
	.w2(32'h39b22de9),
	.w3(32'hba73825b),
	.w4(32'hba2f371c),
	.w5(32'hb9321baa),
	.w6(32'hb91ea52e),
	.w7(32'hb98d4f75),
	.w8(32'hba11762b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e7861),
	.w1(32'hb99a1cd6),
	.w2(32'h3a1775a1),
	.w3(32'h3998a0f1),
	.w4(32'hba0adaa5),
	.w5(32'h3ac60d19),
	.w6(32'h3b083d11),
	.w7(32'hb8401a5d),
	.w8(32'h3ab4b97a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9756042),
	.w1(32'hb8746360),
	.w2(32'h39cc5d21),
	.w3(32'hb92262e6),
	.w4(32'h3964953c),
	.w5(32'h39a2856b),
	.w6(32'h39a1e359),
	.w7(32'h3a1220c2),
	.w8(32'h3a9b0b4a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50f04c),
	.w1(32'hba912973),
	.w2(32'hba682ba7),
	.w3(32'h39a69b0c),
	.w4(32'hba935e6c),
	.w5(32'hbaaf842f),
	.w6(32'hba1d3e59),
	.w7(32'hba494f0f),
	.w8(32'hba98fdd4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2c6a),
	.w1(32'hbac000a5),
	.w2(32'hba8dd8b9),
	.w3(32'hba1ecc03),
	.w4(32'hbaf026d4),
	.w5(32'hbacaf6db),
	.w6(32'hbaf46a57),
	.w7(32'hba9766eb),
	.w8(32'hbaac9382),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3718c),
	.w1(32'h3a568c35),
	.w2(32'h3a532fd8),
	.w3(32'hbb0194b1),
	.w4(32'h3a65dee7),
	.w5(32'h3a358598),
	.w6(32'h3ae1b7f5),
	.w7(32'h3a460543),
	.w8(32'hb8d53089),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c4c62),
	.w1(32'hba878643),
	.w2(32'hba8002bb),
	.w3(32'h39bc76ac),
	.w4(32'hba05c1ec),
	.w5(32'hba85b40d),
	.w6(32'hba6514bc),
	.w7(32'hba82c0c2),
	.w8(32'hbaa9cc47),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1d7f0),
	.w1(32'h3a056e3c),
	.w2(32'h3a34c587),
	.w3(32'hbac59b45),
	.w4(32'h39f7bc9b),
	.w5(32'h3a69f4e2),
	.w6(32'h3a86fd09),
	.w7(32'h3a7f6695),
	.w8(32'h3a7edecf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98c862),
	.w1(32'hba70e767),
	.w2(32'hb9d10186),
	.w3(32'h3a2cc907),
	.w4(32'hb95dd511),
	.w5(32'hb97b5a80),
	.w6(32'h3a350514),
	.w7(32'hb97ca4fa),
	.w8(32'hb939bf88),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab00ca3),
	.w1(32'h3a11747f),
	.w2(32'h3a2c5514),
	.w3(32'hba18a7fb),
	.w4(32'h3a57bdf2),
	.w5(32'h3a782943),
	.w6(32'h3a9f4fb7),
	.w7(32'h39a1606f),
	.w8(32'h38d1840b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f8203),
	.w1(32'h3b0592a3),
	.w2(32'hbada62a8),
	.w3(32'hb9243fab),
	.w4(32'h3aa87a5f),
	.w5(32'hb99ef8ba),
	.w6(32'h3996c45d),
	.w7(32'hbb19f39a),
	.w8(32'hba7660d0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc617),
	.w1(32'hba3b5821),
	.w2(32'hba8fd291),
	.w3(32'hbb171744),
	.w4(32'h38662f9d),
	.w5(32'hba304325),
	.w6(32'hb9fd954b),
	.w7(32'hba6ded4c),
	.w8(32'hb951f188),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d22e1),
	.w1(32'hba1f0c80),
	.w2(32'hb9995ad6),
	.w3(32'hb9b63c4f),
	.w4(32'hba356244),
	.w5(32'hb9edc50a),
	.w6(32'hba327394),
	.w7(32'hb98e311b),
	.w8(32'hba6888f1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba534972),
	.w1(32'h39a13a3f),
	.w2(32'h38a1efee),
	.w3(32'hbaa1e014),
	.w4(32'hb9ce9048),
	.w5(32'h3919ddfb),
	.w6(32'h3a655fcc),
	.w7(32'h39a84591),
	.w8(32'hba2f0be3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba596354),
	.w1(32'hba80494c),
	.w2(32'hb9bbbe5c),
	.w3(32'hba238fe4),
	.w4(32'hb9fc5884),
	.w5(32'hb9f43798),
	.w6(32'h3b051306),
	.w7(32'hb8a0efaa),
	.w8(32'h3b19928b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7fd95),
	.w1(32'h3ab7e90c),
	.w2(32'h3b0d2027),
	.w3(32'h3ab005a6),
	.w4(32'h3a403845),
	.w5(32'h3afdf48f),
	.w6(32'h3aab8b48),
	.w7(32'h3ae10e93),
	.w8(32'h3a8c97c0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9611836),
	.w1(32'hba6138be),
	.w2(32'h3a9c07ac),
	.w3(32'h38729e00),
	.w4(32'hb944dfa3),
	.w5(32'h3a9687a0),
	.w6(32'h3b00c2eb),
	.w7(32'h3a6a31ad),
	.w8(32'h3a9dad1d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06206e),
	.w1(32'h3ab8978b),
	.w2(32'h3aa7001f),
	.w3(32'h38d1c6c0),
	.w4(32'h3971b6dd),
	.w5(32'h3a1887ed),
	.w6(32'h3a8f3084),
	.w7(32'h3aaeb0a8),
	.w8(32'h39f87f32),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9603c),
	.w1(32'hbabde1e4),
	.w2(32'hbaaea18e),
	.w3(32'h3a3848c9),
	.w4(32'hba561165),
	.w5(32'hbab73c8b),
	.w6(32'hbac1493e),
	.w7(32'hbac70b0f),
	.w8(32'hbae831c1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc8333),
	.w1(32'h3a07027b),
	.w2(32'h3a4e517c),
	.w3(32'hbafaa614),
	.w4(32'h3a2c23f7),
	.w5(32'h3a38a16f),
	.w6(32'h3a08a489),
	.w7(32'h3a394611),
	.w8(32'h39f191d7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1385dc),
	.w1(32'h3a1967b6),
	.w2(32'h3a4aaa6b),
	.w3(32'h3a077698),
	.w4(32'h3a01b912),
	.w5(32'h3a4e6a3f),
	.w6(32'h3a211c05),
	.w7(32'h3a4e476f),
	.w8(32'h39cd8057),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31e780),
	.w1(32'hba49c8d3),
	.w2(32'h382b382b),
	.w3(32'h3a28973c),
	.w4(32'hba90021d),
	.w5(32'hb8f805b0),
	.w6(32'hba1499e8),
	.w7(32'hba0c271b),
	.w8(32'hba17b03b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e055d),
	.w1(32'hbac3fcf2),
	.w2(32'hba92e132),
	.w3(32'hba3c9004),
	.w4(32'hba77f87d),
	.w5(32'hbab7354f),
	.w6(32'hbab65f63),
	.w7(32'hbac3825c),
	.w8(32'hbb0596e7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dde81),
	.w1(32'hbaa520e7),
	.w2(32'hbaf32253),
	.w3(32'hba6a1863),
	.w4(32'hbb40abc5),
	.w5(32'hbb0ffa44),
	.w6(32'h3abc9b41),
	.w7(32'h3a7c41d9),
	.w8(32'hbada4fb1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab30df2),
	.w1(32'h38f62306),
	.w2(32'h38a9d40e),
	.w3(32'hba190ce5),
	.w4(32'hb90ffcf3),
	.w5(32'h3a573f83),
	.w6(32'h3b6cf061),
	.w7(32'h3a9d3a78),
	.w8(32'h3a43fcbd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c2ac9),
	.w1(32'h3a7bb4e5),
	.w2(32'hb8855946),
	.w3(32'hb85460c8),
	.w4(32'h39412f80),
	.w5(32'hba9d202b),
	.w6(32'hba7e7d44),
	.w7(32'hba9f886c),
	.w8(32'hbaa27fcc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae36a09),
	.w1(32'h39a2434d),
	.w2(32'h3a3dd823),
	.w3(32'hbac10809),
	.w4(32'h3a0b1bb1),
	.w5(32'h3931b19f),
	.w6(32'h3a8c41b9),
	.w7(32'h3a6fbe88),
	.w8(32'h3abfcc45),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de05c),
	.w1(32'hba31211f),
	.w2(32'h3a0da044),
	.w3(32'hb96b6c20),
	.w4(32'hb9f372e5),
	.w5(32'hb9e3bc15),
	.w6(32'hba2f676c),
	.w7(32'hba4904a8),
	.w8(32'hb82056a8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7ea17),
	.w1(32'h39315617),
	.w2(32'h3a86507b),
	.w3(32'hba028063),
	.w4(32'hba540e40),
	.w5(32'hb8df8fcf),
	.w6(32'hba995edc),
	.w7(32'hb9e3e978),
	.w8(32'hba463552),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6baffe),
	.w1(32'hb9a28f2d),
	.w2(32'hb7e5f8af),
	.w3(32'h39076d41),
	.w4(32'hba89f7de),
	.w5(32'hb923c507),
	.w6(32'hb81b2c3b),
	.w7(32'hba6f1701),
	.w8(32'hba5edd75),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b8301),
	.w1(32'hba9d0c14),
	.w2(32'hba4401da),
	.w3(32'hba95a248),
	.w4(32'hba93c688),
	.w5(32'hba886b2a),
	.w6(32'hba953982),
	.w7(32'hba5b3ec6),
	.w8(32'hba513c67),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bbab0),
	.w1(32'hb8c437fd),
	.w2(32'hb9f3fe43),
	.w3(32'hb9c521f6),
	.w4(32'hb98c7758),
	.w5(32'hba1a6d57),
	.w6(32'h37ab52a4),
	.w7(32'hb8e38a07),
	.w8(32'hba2481c8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a1ec5),
	.w1(32'hba227352),
	.w2(32'h3ab34129),
	.w3(32'hba9974da),
	.w4(32'hb9851270),
	.w5(32'h3a8dfe3b),
	.w6(32'h39c04994),
	.w7(32'h39252e53),
	.w8(32'h3a4f87f9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39070101),
	.w1(32'hb8e31645),
	.w2(32'hb83080e4),
	.w3(32'hb91a84be),
	.w4(32'hba1495bf),
	.w5(32'hb9c0386a),
	.w6(32'hba435ddf),
	.w7(32'hb9a883d9),
	.w8(32'hb9b3d560),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930c2b5),
	.w1(32'h3629623e),
	.w2(32'hba59d4f5),
	.w3(32'h3977a875),
	.w4(32'hb996a907),
	.w5(32'hbad26184),
	.w6(32'hba1e9363),
	.w7(32'hb939e814),
	.w8(32'hba9bb46c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11220b),
	.w1(32'hb90722f8),
	.w2(32'h3991625a),
	.w3(32'hba30625b),
	.w4(32'hb8f1f948),
	.w5(32'h379ddb07),
	.w6(32'hb9d427a1),
	.w7(32'hb9e44f88),
	.w8(32'hba28bdf6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a908d22),
	.w1(32'h3ac9d594),
	.w2(32'h3aaa15a8),
	.w3(32'h39ec0ecc),
	.w4(32'h3aa7fb65),
	.w5(32'h3a417207),
	.w6(32'h3ab27c8b),
	.w7(32'h3a8e5d39),
	.w8(32'h3ab52bb6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a6fe7),
	.w1(32'hb963ab00),
	.w2(32'h3a579787),
	.w3(32'h3b0f82cb),
	.w4(32'hb92d4114),
	.w5(32'h39c0215d),
	.w6(32'h3ab5994e),
	.w7(32'hb965eef1),
	.w8(32'hb9eda444),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa767ef),
	.w1(32'hbac8c63c),
	.w2(32'hba0cd9ca),
	.w3(32'hba6b9c4b),
	.w4(32'hbacdbe38),
	.w5(32'hba8dc32e),
	.w6(32'hba49a974),
	.w7(32'hba894b7f),
	.w8(32'hbaa4936b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a830a9e),
	.w1(32'hba9aab76),
	.w2(32'hbaed5987),
	.w3(32'h3aa89c55),
	.w4(32'hba52fe76),
	.w5(32'hbb28c1e3),
	.w6(32'h3adc6830),
	.w7(32'hb9d62c7b),
	.w8(32'hb95b2087),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48500e),
	.w1(32'hbafbb46d),
	.w2(32'hba8245ff),
	.w3(32'hbb65ee0b),
	.w4(32'hbb398a47),
	.w5(32'hbae97e81),
	.w6(32'hbb4cdeae),
	.w7(32'hbafe4b60),
	.w8(32'hba66564b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134af7),
	.w1(32'hba530d7c),
	.w2(32'h3aa18e37),
	.w3(32'hba760d50),
	.w4(32'hba059a19),
	.w5(32'h3a04a923),
	.w6(32'h3a418a66),
	.w7(32'h3a2ab750),
	.w8(32'h39d2f027),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a767c),
	.w1(32'h3a046332),
	.w2(32'h39ead7be),
	.w3(32'hb99e1aea),
	.w4(32'h38fc0bf6),
	.w5(32'hbaa0ef62),
	.w6(32'hb98b33d6),
	.w7(32'h387641e5),
	.w8(32'hb9a5801c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc1dc7),
	.w1(32'hba28af88),
	.w2(32'h389b5e0c),
	.w3(32'hbb1206f3),
	.w4(32'hba9a064c),
	.w5(32'hb98c7ed6),
	.w6(32'h39007386),
	.w7(32'h39ec5946),
	.w8(32'h38acdd97),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968d588),
	.w1(32'h37931c52),
	.w2(32'h3a437c63),
	.w3(32'h3969e5c9),
	.w4(32'hba5c274e),
	.w5(32'h398769d4),
	.w6(32'hb98d8dd5),
	.w7(32'h3a1605e0),
	.w8(32'hb9ba0abe),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9d448),
	.w1(32'hba9f4253),
	.w2(32'h3a7d5263),
	.w3(32'hb8a2cf37),
	.w4(32'hbab0597d),
	.w5(32'h3b127c6a),
	.w6(32'h3a1957b4),
	.w7(32'hba328d31),
	.w8(32'hb8d778be),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33ab6b),
	.w1(32'hb9ffd1e2),
	.w2(32'hb906d582),
	.w3(32'hbb0d70ed),
	.w4(32'hbaf94a32),
	.w5(32'hbad11cfd),
	.w6(32'h3a35aede),
	.w7(32'hba1fc375),
	.w8(32'h391aa410),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b745c5b),
	.w1(32'h3aa9925f),
	.w2(32'h3acae316),
	.w3(32'h3af677e4),
	.w4(32'h3aa695fa),
	.w5(32'h39f09b54),
	.w6(32'h3b8decd7),
	.w7(32'h395e21a7),
	.w8(32'hbab228b8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988babf),
	.w1(32'hb9572071),
	.w2(32'hba978d8c),
	.w3(32'hb97035a5),
	.w4(32'hbacc02f9),
	.w5(32'hbad00502),
	.w6(32'h3b27cf31),
	.w7(32'h3a647a94),
	.w8(32'hbad36cce),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4edbde),
	.w1(32'h3bb938e8),
	.w2(32'h3b86e364),
	.w3(32'hbad6a47d),
	.w4(32'h3b27bec8),
	.w5(32'h3b1be6fa),
	.w6(32'h3b56dfb6),
	.w7(32'h3b2bb2a1),
	.w8(32'hb9d558dc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b167646),
	.w1(32'hba801703),
	.w2(32'hba20d2f5),
	.w3(32'h3ae85d3f),
	.w4(32'hba5e433a),
	.w5(32'hba8d73b4),
	.w6(32'h3b9103ec),
	.w7(32'h3afd33db),
	.w8(32'h3b170c63),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cabd1),
	.w1(32'h393964b0),
	.w2(32'h3a25d369),
	.w3(32'h3a917421),
	.w4(32'h39d06acf),
	.w5(32'h3a398c7d),
	.w6(32'h3a11314f),
	.w7(32'h39ae0f8d),
	.w8(32'h3900a541),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcac0d0),
	.w1(32'h3b955ac3),
	.w2(32'h3aea4f8f),
	.w3(32'h3b99b401),
	.w4(32'h3b8d17c6),
	.w5(32'h3af2326c),
	.w6(32'h3be3c5ea),
	.w7(32'h3b621914),
	.w8(32'h3b05c4fb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7ae89),
	.w1(32'hbaa1b872),
	.w2(32'hba971f29),
	.w3(32'h3a72c197),
	.w4(32'hba8045a6),
	.w5(32'hbac14fd8),
	.w6(32'h3a4c14da),
	.w7(32'hba11edcf),
	.w8(32'hba0adbbb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912bfaa),
	.w1(32'hba90388e),
	.w2(32'hba6ef339),
	.w3(32'hb929cc49),
	.w4(32'hba708938),
	.w5(32'hba8868d0),
	.w6(32'hba17f812),
	.w7(32'hba6cb854),
	.w8(32'hba852917),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c806e),
	.w1(32'h3aaa3902),
	.w2(32'h3af7f587),
	.w3(32'hbadd5fe1),
	.w4(32'h3a2b8587),
	.w5(32'h3a4a13c2),
	.w6(32'hb9a896f7),
	.w7(32'hb947c375),
	.w8(32'hb9f09ab9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836301),
	.w1(32'h3963bb68),
	.w2(32'h398e6efa),
	.w3(32'h39aca6d7),
	.w4(32'hb9e6f70c),
	.w5(32'h3952d91f),
	.w6(32'h3ae946d8),
	.w7(32'h3a84eee3),
	.w8(32'h3ab646a1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f4fc),
	.w1(32'h3ae59673),
	.w2(32'h3a7a0b5b),
	.w3(32'h385c216f),
	.w4(32'h3ac78010),
	.w5(32'h3a7bf17a),
	.w6(32'h395173b2),
	.w7(32'h39f0d41c),
	.w8(32'h3a060300),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81c015),
	.w1(32'h38f90004),
	.w2(32'h3aaf126e),
	.w3(32'hba8ac926),
	.w4(32'hba3b66a6),
	.w5(32'h3a0068c1),
	.w6(32'h3919bf88),
	.w7(32'h3a6ed1b2),
	.w8(32'h3a258011),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5e80d),
	.w1(32'h3ba010be),
	.w2(32'hba9aa72b),
	.w3(32'h3a276ebc),
	.w4(32'h3b870114),
	.w5(32'h3a937e01),
	.w6(32'h3b156fbc),
	.w7(32'hba42a9a9),
	.w8(32'hb930443e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d3e2d),
	.w1(32'hb99b02d0),
	.w2(32'h38e67b65),
	.w3(32'h379fb296),
	.w4(32'hba39f4ef),
	.w5(32'hba2b1d63),
	.w6(32'h39c4f54b),
	.w7(32'h397b3538),
	.w8(32'hbad6a7ad),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ef9255),
	.w1(32'hba4fa6d6),
	.w2(32'hb8963fa1),
	.w3(32'h3a40e72d),
	.w4(32'hb8dc1968),
	.w5(32'hba0d4bb6),
	.w6(32'hb9dec88c),
	.w7(32'hba1937ed),
	.w8(32'hba5dc369),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa2789),
	.w1(32'h3a1b0bbf),
	.w2(32'h39cc314c),
	.w3(32'hba958628),
	.w4(32'h39c1cef0),
	.w5(32'h381328dd),
	.w6(32'hb8d5c977),
	.w7(32'h39672e4d),
	.w8(32'h3981180d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885df17),
	.w1(32'h3a5c3658),
	.w2(32'h39d559b4),
	.w3(32'hb9a2377e),
	.w4(32'h3a0c1390),
	.w5(32'h3a0d2176),
	.w6(32'h3a9f2cb6),
	.w7(32'h3a901596),
	.w8(32'h3a86d651),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a707cbc),
	.w1(32'h3a2f748a),
	.w2(32'h3a37c004),
	.w3(32'h3a8a3e68),
	.w4(32'h3a039421),
	.w5(32'h3a19795f),
	.w6(32'h3a82b40d),
	.w7(32'h3a663929),
	.w8(32'h3a03f29f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e0a0a),
	.w1(32'h39e2afc3),
	.w2(32'h3a4310b9),
	.w3(32'h39d55b5e),
	.w4(32'h3968764a),
	.w5(32'h3a2cc3f1),
	.w6(32'h3a426fff),
	.w7(32'h3a4b9893),
	.w8(32'h3a1e7dc0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a318012),
	.w1(32'hba323ffe),
	.w2(32'hbaa12d11),
	.w3(32'h3a01ab69),
	.w4(32'hba96945c),
	.w5(32'hb7bad821),
	.w6(32'hb967bbf2),
	.w7(32'hba26b8f4),
	.w8(32'hb7caea6b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64a5d2),
	.w1(32'h398a984f),
	.w2(32'h3a5b2336),
	.w3(32'hb64678ba),
	.w4(32'hba22ef03),
	.w5(32'hba488fdb),
	.w6(32'hba3a11a2),
	.w7(32'hb9b54cbb),
	.w8(32'hbb069a47),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb2342),
	.w1(32'hb74940c9),
	.w2(32'h3a6e5159),
	.w3(32'hbadece9e),
	.w4(32'hb86e8fad),
	.w5(32'h3a3408e9),
	.w6(32'h394fe906),
	.w7(32'h3986b646),
	.w8(32'hb9a42d8b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2484fe),
	.w1(32'hba40137c),
	.w2(32'h3a9c8e18),
	.w3(32'h39b28a71),
	.w4(32'hba9bedb6),
	.w5(32'h387b8cf7),
	.w6(32'h3a4c25f4),
	.w7(32'hb90f60ce),
	.w8(32'hba2eb219),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cff802),
	.w1(32'h3ade5655),
	.w2(32'h3afa8cf1),
	.w3(32'h3a2d1705),
	.w4(32'h3ab9aa24),
	.w5(32'h3ae38074),
	.w6(32'h3a851a52),
	.w7(32'h3af84042),
	.w8(32'h3ac4ca97),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a0b76),
	.w1(32'h3abec6e8),
	.w2(32'h3ab0266a),
	.w3(32'h39eff5e0),
	.w4(32'h3a812d12),
	.w5(32'h3b236432),
	.w6(32'h3b178971),
	.w7(32'h3b3d9e03),
	.w8(32'h3aeb1688),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae427dc),
	.w1(32'hbacb95f0),
	.w2(32'hb864eda4),
	.w3(32'h3b26e017),
	.w4(32'hba9cb79a),
	.w5(32'hb9c6d2bf),
	.w6(32'hba88a175),
	.w7(32'hba7d3f7b),
	.w8(32'hba88e295),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba125963),
	.w1(32'hb9dd2672),
	.w2(32'h3a359faa),
	.w3(32'hba5b0101),
	.w4(32'hb9f8a162),
	.w5(32'h38c354ca),
	.w6(32'hba856929),
	.w7(32'hba315b97),
	.w8(32'hba8bb773),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3b3a4),
	.w1(32'h3a124f1e),
	.w2(32'h3a9d429d),
	.w3(32'hb9c48bea),
	.w4(32'h393eec18),
	.w5(32'hb814e214),
	.w6(32'h3a81d831),
	.w7(32'h3a1c7b98),
	.w8(32'h39bf01ea),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8aa76),
	.w1(32'hb8ea8a28),
	.w2(32'h39b9857d),
	.w3(32'h3a5bcc90),
	.w4(32'h3a48ed07),
	.w5(32'h3acf5f29),
	.w6(32'h3a2b5885),
	.w7(32'h3aaad850),
	.w8(32'h3ad56e7a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6aa2d),
	.w1(32'hbb96da63),
	.w2(32'hbb75915f),
	.w3(32'hba10c4a6),
	.w4(32'hbb6205cc),
	.w5(32'hbb1536d8),
	.w6(32'hbb629290),
	.w7(32'hbb864528),
	.w8(32'hbb0f5546),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb379a87),
	.w1(32'hb8a6bc00),
	.w2(32'h39bad765),
	.w3(32'hbb4a073e),
	.w4(32'hb9e71732),
	.w5(32'h396610df),
	.w6(32'h39a20204),
	.w7(32'hb960d42f),
	.w8(32'h3992469c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f770f),
	.w1(32'hba19287c),
	.w2(32'hba3aa82b),
	.w3(32'h3ad01189),
	.w4(32'hb9cdb023),
	.w5(32'hb94bb587),
	.w6(32'h3950162a),
	.w7(32'hb98b7aa4),
	.w8(32'h39aa21f6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e7b90),
	.w1(32'hb97e049e),
	.w2(32'h3b7aeb8c),
	.w3(32'h399df989),
	.w4(32'hba4b4519),
	.w5(32'hbb64e50a),
	.w6(32'h39cf5e54),
	.w7(32'h39e3f0c0),
	.w8(32'h3a53bffe),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe39a),
	.w1(32'h37c70538),
	.w2(32'h375abf18),
	.w3(32'hbad84bb8),
	.w4(32'hb98c2fe8),
	.w5(32'h3a998672),
	.w6(32'hb981897d),
	.w7(32'hba7d0191),
	.w8(32'hba99e130),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6322d6),
	.w1(32'h3b1e5027),
	.w2(32'h3b503b2a),
	.w3(32'hb99f24b8),
	.w4(32'h3b094d2d),
	.w5(32'h3af07edd),
	.w6(32'h3aba1589),
	.w7(32'h3ae55587),
	.w8(32'h3a83e9de),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147784),
	.w1(32'hba4f2215),
	.w2(32'hb91eb248),
	.w3(32'h3b09f1d1),
	.w4(32'hbaa5476e),
	.w5(32'h397e31ff),
	.w6(32'h3adf6789),
	.w7(32'h3852d071),
	.w8(32'h3aa1f7ab),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f129c),
	.w1(32'hb89fe7ec),
	.w2(32'hb826db03),
	.w3(32'h3984eb32),
	.w4(32'h3909100c),
	.w5(32'hb91abad5),
	.w6(32'h389295d0),
	.w7(32'h3a14e2d4),
	.w8(32'h39a63f44),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c983f),
	.w1(32'hb8bc375c),
	.w2(32'h3a8ab8d5),
	.w3(32'hba82abb2),
	.w4(32'h385a072c),
	.w5(32'h3a2eb004),
	.w6(32'h39834830),
	.w7(32'hb98926bf),
	.w8(32'h3a54b06a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f55f2),
	.w1(32'hbb0c0225),
	.w2(32'hb9503595),
	.w3(32'h385a22e6),
	.w4(32'hbaaae9c0),
	.w5(32'h3a68c234),
	.w6(32'h3a6a1fa6),
	.w7(32'hba56df0f),
	.w8(32'h3a8fdb98),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba1b3),
	.w1(32'hb9a87fc8),
	.w2(32'h38d049c3),
	.w3(32'h3b56f5a8),
	.w4(32'h3a02453b),
	.w5(32'hb9fb37a9),
	.w6(32'h3a24a65a),
	.w7(32'h3ad6130d),
	.w8(32'h3a16ceb2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39034a70),
	.w1(32'h382affd0),
	.w2(32'h3b0495c1),
	.w3(32'hb8820c85),
	.w4(32'h3a52a090),
	.w5(32'hb92bc55b),
	.w6(32'h3b296d43),
	.w7(32'h3b3051f3),
	.w8(32'h3b3c043a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93678d),
	.w1(32'hb84b4c2c),
	.w2(32'h3928fd72),
	.w3(32'hb9dadadb),
	.w4(32'hba041d5f),
	.w5(32'hba2239b8),
	.w6(32'h3942c383),
	.w7(32'h39d9a714),
	.w8(32'h39c02708),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaeaba),
	.w1(32'hbb4dbf77),
	.w2(32'hbb104fe0),
	.w3(32'hba8a5df0),
	.w4(32'hbaaba824),
	.w5(32'hbaa422fd),
	.w6(32'hbac1b006),
	.w7(32'hba526af2),
	.w8(32'hba463e29),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43be75),
	.w1(32'hbb350ca9),
	.w2(32'h390663d9),
	.w3(32'hbaa8a802),
	.w4(32'hb9ffba35),
	.w5(32'hbaeaf876),
	.w6(32'h3a47a044),
	.w7(32'h3b017040),
	.w8(32'h3acb2224),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac40f09),
	.w1(32'hb9b24c03),
	.w2(32'h3904a84e),
	.w3(32'hbaaf04f1),
	.w4(32'hba15fdb7),
	.w5(32'hb950537d),
	.w6(32'hb9126ac7),
	.w7(32'hb9d704cf),
	.w8(32'hb9b5777c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9644716),
	.w1(32'hbb1fddba),
	.w2(32'hbacd807f),
	.w3(32'hb9ca1f30),
	.w4(32'hbac052ed),
	.w5(32'hb82f5dad),
	.w6(32'hba3d0f91),
	.w7(32'hba56b584),
	.w8(32'h3abefdf2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a508729),
	.w1(32'hba2d2730),
	.w2(32'hba1a278e),
	.w3(32'h3b28e70e),
	.w4(32'hb9ca94eb),
	.w5(32'hb9a760dc),
	.w6(32'hba222f6c),
	.w7(32'hbaa64109),
	.w8(32'hb9a276a2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910e29f),
	.w1(32'hb90f8429),
	.w2(32'hb9ebd917),
	.w3(32'h3a82cc6c),
	.w4(32'hb9e650a4),
	.w5(32'hba59478c),
	.w6(32'hb7ff40d6),
	.w7(32'hb983f491),
	.w8(32'hb9a87896),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35915377),
	.w1(32'hb83959c8),
	.w2(32'h3a2a9219),
	.w3(32'hba3208c6),
	.w4(32'hba4a3303),
	.w5(32'h39bea9e2),
	.w6(32'hba2f3e9a),
	.w7(32'hba3453cc),
	.w8(32'h3a23a012),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf1418),
	.w1(32'h3adbc8d0),
	.w2(32'h3b7933a0),
	.w3(32'hb9abdfeb),
	.w4(32'h3ac09a6c),
	.w5(32'h3aa07bba),
	.w6(32'h3afe148a),
	.w7(32'h3b1bdfe8),
	.w8(32'h3ad054d4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe132),
	.w1(32'hbb6669d6),
	.w2(32'hbb31bd35),
	.w3(32'h3aced845),
	.w4(32'hbb8728e5),
	.w5(32'hbb893745),
	.w6(32'hbab1e6a5),
	.w7(32'hba7c2146),
	.w8(32'hbaf4520c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e517),
	.w1(32'h3aaed446),
	.w2(32'h3b7ce77b),
	.w3(32'hbb8fb831),
	.w4(32'hb9a98168),
	.w5(32'h3a989e43),
	.w6(32'hba81cf56),
	.w7(32'hb9ecbc3c),
	.w8(32'h3a286228),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55e109),
	.w1(32'hba8c9c3a),
	.w2(32'h39f8d9f9),
	.w3(32'hb95411f1),
	.w4(32'hbb10a534),
	.w5(32'hba9af2a0),
	.w6(32'h3a814136),
	.w7(32'hba342986),
	.w8(32'h390bb010),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeae51),
	.w1(32'hba4d9265),
	.w2(32'h3a62804c),
	.w3(32'hbae51f65),
	.w4(32'hba196605),
	.w5(32'hba07701b),
	.w6(32'hba9cd331),
	.w7(32'hba97d43b),
	.w8(32'h3a62409e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7d1e),
	.w1(32'hbb2d4e2b),
	.w2(32'hbaf89957),
	.w3(32'h3aaa7a96),
	.w4(32'hba67c48f),
	.w5(32'hbabf61ce),
	.w6(32'h3ac8feeb),
	.w7(32'h3b03b0d7),
	.w8(32'h3b259c5f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d8134),
	.w1(32'hb9f989a4),
	.w2(32'h389b81f1),
	.w3(32'hb835eff0),
	.w4(32'hba0c279d),
	.w5(32'hb984ed30),
	.w6(32'h38a5db87),
	.w7(32'hb87b0ad0),
	.w8(32'hb98ecdb6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f458d),
	.w1(32'hbae3ff31),
	.w2(32'hba9cfd9d),
	.w3(32'hb9bfb6d9),
	.w4(32'hbb19f477),
	.w5(32'hbb21b24b),
	.w6(32'hbaa237a1),
	.w7(32'hbaf5b10a),
	.w8(32'hbab0749f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27b635),
	.w1(32'hba5a1563),
	.w2(32'h3af4abf2),
	.w3(32'hba983829),
	.w4(32'hbaab191a),
	.w5(32'hba48b890),
	.w6(32'hba93a118),
	.w7(32'hba9d2cbb),
	.w8(32'h3a987fb0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46c1ee),
	.w1(32'hba876264),
	.w2(32'hb9ffa6b5),
	.w3(32'h3a7c4b31),
	.w4(32'hb7814cd6),
	.w5(32'h3ad16696),
	.w6(32'hb9d9b768),
	.w7(32'hb9d325bf),
	.w8(32'h3b37b8f9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e2508),
	.w1(32'h3a20e23c),
	.w2(32'h3ada0cbf),
	.w3(32'h3bc08cea),
	.w4(32'h39ced041),
	.w5(32'h39fa0756),
	.w6(32'h3aac051b),
	.w7(32'h3a956bc7),
	.w8(32'h3a76d934),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca4feb),
	.w1(32'h396761b8),
	.w2(32'h3a8bc75b),
	.w3(32'h395f14ef),
	.w4(32'hb8a48216),
	.w5(32'h386fbd11),
	.w6(32'h3a281a26),
	.w7(32'h3a84da5d),
	.w8(32'h39c2b7a8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977ce88),
	.w1(32'hbb616d32),
	.w2(32'hba95f3d2),
	.w3(32'hba8539fe),
	.w4(32'hbb640c1b),
	.w5(32'hba8337b2),
	.w6(32'hbb13345d),
	.w7(32'hba75ddf5),
	.w8(32'hba4f4df0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae92e62),
	.w1(32'hbb05b7bb),
	.w2(32'hbb7247d2),
	.w3(32'hbab25b25),
	.w4(32'hbacbb0cb),
	.w5(32'hbb603033),
	.w6(32'hbb6b1332),
	.w7(32'hbb863127),
	.w8(32'hbb209b54),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168de6),
	.w1(32'h3914c634),
	.w2(32'h3a6af8c6),
	.w3(32'hbb1faae1),
	.w4(32'h3a022958),
	.w5(32'h3aa86639),
	.w6(32'hb8d16e85),
	.w7(32'h3850992d),
	.w8(32'h3a9fe34f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af579b3),
	.w1(32'hb933bd64),
	.w2(32'h3a97af7d),
	.w3(32'h3b25f3b7),
	.w4(32'hb8d88bbd),
	.w5(32'h3958539b),
	.w6(32'h3980e83d),
	.w7(32'h39f249db),
	.w8(32'h3998fe9b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d14df),
	.w1(32'hb9979808),
	.w2(32'h3ab5ed76),
	.w3(32'hba829710),
	.w4(32'h39be2b3f),
	.w5(32'h3b091ab8),
	.w6(32'h3a229101),
	.w7(32'h3a683937),
	.w8(32'h3b00bbf6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8f938),
	.w1(32'hb9088961),
	.w2(32'hb9a4ab8e),
	.w3(32'h3af6da7c),
	.w4(32'hb9457de1),
	.w5(32'h39794bfe),
	.w6(32'hb8fc08f0),
	.w7(32'hba23a0bd),
	.w8(32'h38341457),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfc0e6),
	.w1(32'h36930802),
	.w2(32'h3a18abdd),
	.w3(32'h3a5b28a3),
	.w4(32'hb71d1724),
	.w5(32'h388265d5),
	.w6(32'h3925e07e),
	.w7(32'h39c92b4b),
	.w8(32'h39eaf9db),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fd37a),
	.w1(32'h3954d44d),
	.w2(32'h3806abc8),
	.w3(32'hb7560c85),
	.w4(32'h382ff201),
	.w5(32'hb92a396e),
	.w6(32'h38d1bad2),
	.w7(32'h3944ef7b),
	.w8(32'h397fd2e6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad00f41),
	.w1(32'h397705a0),
	.w2(32'h3b3bb236),
	.w3(32'h3aba6069),
	.w4(32'h39013167),
	.w5(32'h3b735d18),
	.w6(32'h3b0e1464),
	.w7(32'h3b3ec955),
	.w8(32'h3bbf4fe4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02fe75),
	.w1(32'hba0c9d48),
	.w2(32'h39a38aae),
	.w3(32'h3be03acb),
	.w4(32'h3901f59e),
	.w5(32'h39ff0f0c),
	.w6(32'h39fdfe0e),
	.w7(32'h3a788983),
	.w8(32'h3a8d9654),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d58fdb),
	.w1(32'h3a327e78),
	.w2(32'h3a3eb80b),
	.w3(32'h39e9feb3),
	.w4(32'hb8abd9fd),
	.w5(32'hb9f75e23),
	.w6(32'h3923aa69),
	.w7(32'h3a32cf7c),
	.w8(32'h39faf3ea),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba529533),
	.w1(32'hbac82557),
	.w2(32'hba2ce163),
	.w3(32'hba48563b),
	.w4(32'hba8ffa82),
	.w5(32'h393eba4c),
	.w6(32'hbaf92fc4),
	.w7(32'hbb4e1e14),
	.w8(32'hbaac863c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34e39c),
	.w1(32'hbade754f),
	.w2(32'hba942088),
	.w3(32'h3b23e541),
	.w4(32'hbb57e748),
	.w5(32'hbb08c504),
	.w6(32'hba84b25f),
	.w7(32'hbb204a09),
	.w8(32'hba0c9d47),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6441),
	.w1(32'hba8d4876),
	.w2(32'hb9daff9f),
	.w3(32'hbab452ac),
	.w4(32'hbb0a5ce2),
	.w5(32'hba933a8f),
	.w6(32'h38761c44),
	.w7(32'hba32b5f9),
	.w8(32'h3953d7f2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24082f),
	.w1(32'hba5941ec),
	.w2(32'h3b05e986),
	.w3(32'hb929ff14),
	.w4(32'hbaa35d85),
	.w5(32'hbb49936f),
	.w6(32'h3afce985),
	.w7(32'h3b176574),
	.w8(32'h3ad9e94e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90d064),
	.w1(32'hba96d010),
	.w2(32'hbaaa235d),
	.w3(32'hbb2c24e8),
	.w4(32'hbaaca585),
	.w5(32'hbaef6c7a),
	.w6(32'hbae2bc4f),
	.w7(32'hbb81d9e5),
	.w8(32'h397d9475),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b457614),
	.w1(32'h39290f97),
	.w2(32'h3a89399c),
	.w3(32'h3b0867b1),
	.w4(32'hb90cc795),
	.w5(32'h395f2571),
	.w6(32'h3a187a71),
	.w7(32'h3a304126),
	.w8(32'h3a49995f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba574752),
	.w1(32'hba48384a),
	.w2(32'hb9a39085),
	.w3(32'hba468f49),
	.w4(32'hba2672fb),
	.w5(32'hba2d9f82),
	.w6(32'hba1bbae8),
	.w7(32'hb93b532a),
	.w8(32'hba017624),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9408c6),
	.w1(32'hbab90ec5),
	.w2(32'hba971ef8),
	.w3(32'hba8da3a5),
	.w4(32'hba997f3e),
	.w5(32'hba4588d1),
	.w6(32'hb96c3695),
	.w7(32'hb90c35a5),
	.w8(32'h3a8e889a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17bdbe),
	.w1(32'hbb64208d),
	.w2(32'hbb591c14),
	.w3(32'hba7a93bc),
	.w4(32'hbb2ab8b8),
	.w5(32'hbb4e978e),
	.w6(32'hbb5b3425),
	.w7(32'hbb67d98a),
	.w8(32'hba853f91),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf01d5),
	.w1(32'h3ae30971),
	.w2(32'h3b5761b5),
	.w3(32'hbb0446c5),
	.w4(32'h3950342b),
	.w5(32'h3a7b052d),
	.w6(32'h3adedf69),
	.w7(32'h3a8e7a2c),
	.w8(32'h3b0b749e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2923b8),
	.w1(32'h3a4cf87c),
	.w2(32'h3a11271f),
	.w3(32'h3abbf8d6),
	.w4(32'h3a165661),
	.w5(32'h3aff6fbb),
	.w6(32'h39cc5d61),
	.w7(32'h3a4185a0),
	.w8(32'hba4f1c5f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9c5fa),
	.w1(32'hba5e97bf),
	.w2(32'h3734036c),
	.w3(32'h3967b5c1),
	.w4(32'hba8bd39d),
	.w5(32'hba16d9eb),
	.w6(32'hb877772d),
	.w7(32'h383e0ac8),
	.w8(32'h3a699562),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acedf09),
	.w1(32'h3b6c488f),
	.w2(32'h3bdd38b1),
	.w3(32'h3a985116),
	.w4(32'h3af15887),
	.w5(32'h3bb106c6),
	.w6(32'h3a9f727a),
	.w7(32'h3b65bee4),
	.w8(32'h3b1bde35),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde0ac0),
	.w1(32'hbb174d16),
	.w2(32'hba740eba),
	.w3(32'h3b8ade2d),
	.w4(32'hbb0494ee),
	.w5(32'hbb1f145e),
	.w6(32'hb9c092a8),
	.w7(32'hba91c2be),
	.w8(32'h3a2ad127),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089fc5),
	.w1(32'hba87d5bc),
	.w2(32'hbb3c3600),
	.w3(32'h3aafd56b),
	.w4(32'hbade7643),
	.w5(32'hbb2dde1a),
	.w6(32'h39ddb515),
	.w7(32'hbac15ef1),
	.w8(32'hbaecc701),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab56f79),
	.w1(32'h3621588a),
	.w2(32'hba112bf5),
	.w3(32'hba449572),
	.w4(32'hba493d29),
	.w5(32'hba94286f),
	.w6(32'hb9cade57),
	.w7(32'hba885551),
	.w8(32'hb989b7f3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b8bbd),
	.w1(32'hba8bc5b5),
	.w2(32'h3ad4415f),
	.w3(32'hbad56911),
	.w4(32'hbb025e48),
	.w5(32'h3a336df2),
	.w6(32'h3971c85e),
	.w7(32'hba9a116a),
	.w8(32'h3af74975),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08be63),
	.w1(32'h3a666fb4),
	.w2(32'hb9549a09),
	.w3(32'h395a52ea),
	.w4(32'hb9632e78),
	.w5(32'hba7f26e5),
	.w6(32'hb8c77d6f),
	.w7(32'hb7c320eb),
	.w8(32'hba232844),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971a37c),
	.w1(32'hba832e33),
	.w2(32'hba12d8a5),
	.w3(32'hb6ee4efb),
	.w4(32'hba334a9c),
	.w5(32'hba62cfbf),
	.w6(32'hb9af7b03),
	.w7(32'hb9bdbd78),
	.w8(32'hb88f2032),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24d65a),
	.w1(32'hbb0d50d3),
	.w2(32'hbb1eaea6),
	.w3(32'hb9c26db6),
	.w4(32'hbaa301ce),
	.w5(32'hba153c21),
	.w6(32'hbb8b4098),
	.w7(32'hbb4f3fe1),
	.w8(32'hbb70c7e5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55c78e),
	.w1(32'hba6e77d2),
	.w2(32'hb98752e4),
	.w3(32'hbad35f2a),
	.w4(32'hba1a47f5),
	.w5(32'h39ce809c),
	.w6(32'hba69d61a),
	.w7(32'hbafca5c3),
	.w8(32'hba325ea2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac19196),
	.w1(32'hba2128f0),
	.w2(32'hb96bb2b9),
	.w3(32'h3b016ba8),
	.w4(32'hba6fddb1),
	.w5(32'hba87325b),
	.w6(32'hba532faa),
	.w7(32'hba941af8),
	.w8(32'hba5fb87d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ba7a2),
	.w1(32'hbb510283),
	.w2(32'hbb7aa5a7),
	.w3(32'hb9275fb1),
	.w4(32'hbb3e8435),
	.w5(32'hbb1bfec2),
	.w6(32'hbaf7bec1),
	.w7(32'hbb2c0ead),
	.w8(32'hbaf90d1b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3163b),
	.w1(32'h3b0b0703),
	.w2(32'h3b6c7e1a),
	.w3(32'hba5d8e75),
	.w4(32'h3b158dbf),
	.w5(32'h3b9a038c),
	.w6(32'h3ab113bb),
	.w7(32'h3afdd7d5),
	.w8(32'h3b9dead5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01b621),
	.w1(32'h3ae4de42),
	.w2(32'h3b33d336),
	.w3(32'h3c1799ec),
	.w4(32'hba09dcd6),
	.w5(32'hbab100f0),
	.w6(32'h3a674c77),
	.w7(32'hb9c59b42),
	.w8(32'h3b1a70f3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba652a9),
	.w1(32'h388d1100),
	.w2(32'h3a9d8404),
	.w3(32'h3b07cca1),
	.w4(32'hb956998f),
	.w5(32'hb83b4c96),
	.w6(32'h39e27ae3),
	.w7(32'h3a2f4603),
	.w8(32'h393ddc54),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a613f45),
	.w1(32'hbb4f418b),
	.w2(32'hbb223c5a),
	.w3(32'hba102dfe),
	.w4(32'hbb59ab25),
	.w5(32'hbaea5b4f),
	.w6(32'hbad509fe),
	.w7(32'hbb1b0fec),
	.w8(32'h37805b8d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936a39e),
	.w1(32'hb9811d40),
	.w2(32'hba01cbcf),
	.w3(32'hba22722c),
	.w4(32'hb984b40c),
	.w5(32'hb9b34186),
	.w6(32'hba04ce7b),
	.w7(32'hbaf3fe6a),
	.w8(32'hba8c3628),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5897c),
	.w1(32'hb99465b8),
	.w2(32'h3a373a78),
	.w3(32'h3a7dc740),
	.w4(32'hb9e8f77a),
	.w5(32'hb8befcf6),
	.w6(32'hb93fcf10),
	.w7(32'h39aa91e8),
	.w8(32'hb8ccde1e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5243d9),
	.w1(32'h3a2f0827),
	.w2(32'h39b3fc5c),
	.w3(32'h38b9088f),
	.w4(32'h3a2d9fbb),
	.w5(32'h38915dd6),
	.w6(32'h3a8964db),
	.w7(32'h3a2e02ee),
	.w8(32'h3a09e5f3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb822a7e9),
	.w1(32'h39178533),
	.w2(32'h3ad04f58),
	.w3(32'hb9aa35f4),
	.w4(32'hb8141978),
	.w5(32'h39391356),
	.w6(32'h3a54a91e),
	.w7(32'h3a9692bd),
	.w8(32'h3a0b6c4a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e9e6d),
	.w1(32'hba394fd7),
	.w2(32'hb9b25fdb),
	.w3(32'hba4302f3),
	.w4(32'hba8723ff),
	.w5(32'hba1f6aa3),
	.w6(32'h396338b2),
	.w7(32'hba806bd0),
	.w8(32'h3a134cad),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f29c3),
	.w1(32'hbacb47c4),
	.w2(32'h3a0a4556),
	.w3(32'hb920be1d),
	.w4(32'hba49ca70),
	.w5(32'hbb254d1b),
	.w6(32'h3a5a8454),
	.w7(32'h3b4510e8),
	.w8(32'h3ad21bdc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c9c68),
	.w1(32'hb9af2092),
	.w2(32'h3a0d2b96),
	.w3(32'hbaee5805),
	.w4(32'h3929fed3),
	.w5(32'h39b928cf),
	.w6(32'hba7bb9b2),
	.w7(32'hba104796),
	.w8(32'hb9876e88),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa93ac),
	.w1(32'hba8ef64d),
	.w2(32'hba8c99c6),
	.w3(32'h39bd1278),
	.w4(32'hba354f82),
	.w5(32'hba206f7f),
	.w6(32'hbac71756),
	.w7(32'hbac79c47),
	.w8(32'hba7a0fba),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c679b1),
	.w1(32'hbb17dacb),
	.w2(32'hba23377f),
	.w3(32'h3a64877c),
	.w4(32'hbb19faaf),
	.w5(32'hbafa7eb2),
	.w6(32'hbaa0855a),
	.w7(32'h3a243a15),
	.w8(32'h3a708e43),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc6803),
	.w1(32'h3ae0dcf2),
	.w2(32'h3b6e3f5e),
	.w3(32'h39bcbca6),
	.w4(32'h3ac2b4a8),
	.w5(32'h3ab9b217),
	.w6(32'h3b08bf67),
	.w7(32'h3b06ca52),
	.w8(32'h3ac925fd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30303b),
	.w1(32'h3b35c41d),
	.w2(32'h3bccd74b),
	.w3(32'hba2a82d3),
	.w4(32'hba13f021),
	.w5(32'h3adb5953),
	.w6(32'hb90fe72f),
	.w7(32'hb91fee7a),
	.w8(32'h3b3822e0),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0312be),
	.w1(32'hb9cf9d79),
	.w2(32'hb9c813cc),
	.w3(32'h3b926d74),
	.w4(32'hba4a1ab0),
	.w5(32'hba2642dd),
	.w6(32'hb99276bf),
	.w7(32'hba0e3f78),
	.w8(32'hb96e6579),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904e1fd),
	.w1(32'h3a8ec5ea),
	.w2(32'h3b21a6c0),
	.w3(32'hb903884f),
	.w4(32'h39de8359),
	.w5(32'h3aea5c92),
	.w6(32'h3959b18c),
	.w7(32'h39270d17),
	.w8(32'h3ab802f6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba23b80),
	.w1(32'h3a0bb667),
	.w2(32'h3943a166),
	.w3(32'h3b47c1b8),
	.w4(32'hb9c71abd),
	.w5(32'h38c452a1),
	.w6(32'h3a3097ee),
	.w7(32'hb9f600ce),
	.w8(32'h394a4217),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b9c7f),
	.w1(32'h3ad26a52),
	.w2(32'h3a99dd65),
	.w3(32'h3a369ebe),
	.w4(32'h39b23f1c),
	.w5(32'h39a68656),
	.w6(32'h3b254544),
	.w7(32'h3974e6f4),
	.w8(32'h3b4fa90d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30db12),
	.w1(32'h3b0c5592),
	.w2(32'h3b2594de),
	.w3(32'h3b15d0b5),
	.w4(32'h3a887bf1),
	.w5(32'h3afd0fb3),
	.w6(32'h39ffebab),
	.w7(32'h3a362177),
	.w8(32'h3a97cf99),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb4d51),
	.w1(32'hbb216c21),
	.w2(32'hbb2f1b96),
	.w3(32'h3b18bf3b),
	.w4(32'hbaae8ed0),
	.w5(32'hbb3d50e2),
	.w6(32'h39430964),
	.w7(32'hb926555c),
	.w8(32'h3a720f3e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8862f5),
	.w1(32'h3a539907),
	.w2(32'h3afba529),
	.w3(32'hbabc38b7),
	.w4(32'h3a627259),
	.w5(32'h3a47d5c3),
	.w6(32'h3a58f57c),
	.w7(32'h3a9e4e32),
	.w8(32'h3a5c4677),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a202e16),
	.w1(32'h3a01ceb5),
	.w2(32'h3a6788d4),
	.w3(32'h39d805ec),
	.w4(32'hb99e3dd1),
	.w5(32'hb8a251a6),
	.w6(32'h3a94801d),
	.w7(32'h3a4d436c),
	.w8(32'h3aa42d77),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8ab09),
	.w1(32'hb9c5a65b),
	.w2(32'hb99d09cd),
	.w3(32'h3b813750),
	.w4(32'hb9bb5a63),
	.w5(32'hba287778),
	.w6(32'h3b81f7ba),
	.w7(32'h3a9d2186),
	.w8(32'hb9bf04a6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ff6e2),
	.w1(32'hba0dbe48),
	.w2(32'h3b1bfc5f),
	.w3(32'h3908eb37),
	.w4(32'hbac8068c),
	.w5(32'h3a1a42db),
	.w6(32'h3acde61b),
	.w7(32'h39a9799e),
	.w8(32'h3ac69248),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b4fa4),
	.w1(32'hba8c3120),
	.w2(32'hbab8627d),
	.w3(32'h3adeefee),
	.w4(32'hba736afc),
	.w5(32'hb9e54fbf),
	.w6(32'h3b22e49f),
	.w7(32'hb878c4e9),
	.w8(32'hba30548b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dafa1),
	.w1(32'h39b192cc),
	.w2(32'h3a840a89),
	.w3(32'h3ad8d548),
	.w4(32'hb73f5980),
	.w5(32'h3a59829b),
	.w6(32'h39215fc7),
	.w7(32'hba611b8d),
	.w8(32'h39290660),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba584),
	.w1(32'h3b2edc8a),
	.w2(32'h3bcb20ae),
	.w3(32'h3b3bb7cf),
	.w4(32'h3a95ac25),
	.w5(32'h3ae2ff6b),
	.w6(32'h385d8b65),
	.w7(32'h3a1eddf0),
	.w8(32'h3acec692),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78f07),
	.w1(32'hba53fdab),
	.w2(32'hba7916c1),
	.w3(32'h3b3105e8),
	.w4(32'hba5b77e1),
	.w5(32'hba35cceb),
	.w6(32'hb8346f5f),
	.w7(32'hb96f6b3e),
	.w8(32'h39dbcf3f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98952e3),
	.w1(32'hb9e114a5),
	.w2(32'hb9ab0db5),
	.w3(32'hb88bad03),
	.w4(32'hbaa2eb10),
	.w5(32'hba9d4811),
	.w6(32'hba070a3c),
	.w7(32'hb97d86e0),
	.w8(32'hba44c164),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ffe3),
	.w1(32'hbaeba481),
	.w2(32'h39a8194d),
	.w3(32'hba9a6531),
	.w4(32'hbb21810f),
	.w5(32'hba3c107a),
	.w6(32'hbb092c4a),
	.w7(32'hb9791e17),
	.w8(32'h39e06d2d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c5507),
	.w1(32'hbb0c95f4),
	.w2(32'hbb5eaf1b),
	.w3(32'hba39c801),
	.w4(32'hba84f220),
	.w5(32'hbad297ac),
	.w6(32'hbb69d99b),
	.w7(32'hbb8756b4),
	.w8(32'hbb08beae),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba909062),
	.w1(32'hb9d07dca),
	.w2(32'hb841ea48),
	.w3(32'hba86e4bb),
	.w4(32'hba6e28ab),
	.w5(32'hb82523f1),
	.w6(32'hb848f128),
	.w7(32'hba447127),
	.w8(32'h39e76f34),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dc932),
	.w1(32'h3af75040),
	.w2(32'h3b63cfac),
	.w3(32'h3ad39960),
	.w4(32'h3b10142d),
	.w5(32'h3b3f42d6),
	.w6(32'h3b35aae3),
	.w7(32'hb907c916),
	.w8(32'h3b13fec2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5299bd),
	.w1(32'hbb682a42),
	.w2(32'hbb76c1f1),
	.w3(32'h3b4de282),
	.w4(32'hbb5ecaf1),
	.w5(32'hba9ee32d),
	.w6(32'hbb731735),
	.w7(32'hbaefa1d4),
	.w8(32'hbb06cc47),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23eb5e),
	.w1(32'hbae027bc),
	.w2(32'hbb0f5cc5),
	.w3(32'hbad86681),
	.w4(32'hbb5b7c18),
	.w5(32'hbad5ce11),
	.w6(32'hba5ba3fa),
	.w7(32'hb9a46e0d),
	.w8(32'hbb3f18d8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a575dd6),
	.w1(32'hbadcf06f),
	.w2(32'hba87ccb4),
	.w3(32'h3b273be6),
	.w4(32'hba8f6f97),
	.w5(32'hbab97d66),
	.w6(32'h3b2a6cd7),
	.w7(32'hba8c4d0d),
	.w8(32'hbb0a5942),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f7ae3),
	.w1(32'hb9cb3af8),
	.w2(32'h3a8883d8),
	.w3(32'h3a1c5d80),
	.w4(32'hba236fbd),
	.w5(32'h388d6028),
	.w6(32'h39a17643),
	.w7(32'h391ec3b9),
	.w8(32'h372e955e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d320a4),
	.w1(32'hba16d66c),
	.w2(32'h39423a77),
	.w3(32'hba2ff4b7),
	.w4(32'h376a3904),
	.w5(32'h399840a0),
	.w6(32'hba632922),
	.w7(32'hba36ccbd),
	.w8(32'hb9d0e0db),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e0d76),
	.w1(32'hba84e0f5),
	.w2(32'hb88fd10e),
	.w3(32'h39d9164a),
	.w4(32'hba420701),
	.w5(32'hb9093e2e),
	.w6(32'hb8274fa5),
	.w7(32'hb9c839f2),
	.w8(32'h397c521c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b141d),
	.w1(32'hba1f91eb),
	.w2(32'hb992e3c4),
	.w3(32'hb9de4989),
	.w4(32'hb98d2d48),
	.w5(32'hb9bf8042),
	.w6(32'hb59f1b9e),
	.w7(32'hb9275c64),
	.w8(32'h3a043c94),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6b4f8),
	.w1(32'h3ab48ca8),
	.w2(32'h3b525c8e),
	.w3(32'h3a336c59),
	.w4(32'h3a8488b3),
	.w5(32'h3a826aca),
	.w6(32'h3ad27de5),
	.w7(32'h3b07e8bd),
	.w8(32'h3abd4d40),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad174b4),
	.w1(32'hba203cc1),
	.w2(32'h38977a8a),
	.w3(32'h3a24ac9e),
	.w4(32'hb89d2c46),
	.w5(32'h395c769d),
	.w6(32'hba7912b2),
	.w7(32'hba407467),
	.w8(32'hb9f85bd5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972d6b8),
	.w1(32'h38a0e8e2),
	.w2(32'hb90ab709),
	.w3(32'h397641c6),
	.w4(32'hba48e419),
	.w5(32'hba4fee56),
	.w6(32'h3950be46),
	.w7(32'h395f3cea),
	.w8(32'hb96e7944),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ff62c),
	.w1(32'hb99e2186),
	.w2(32'h39d9bfdd),
	.w3(32'hba962f58),
	.w4(32'hb9e82dea),
	.w5(32'hb9cd0786),
	.w6(32'hb903af01),
	.w7(32'hb70aa7c2),
	.w8(32'h39574449),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b5b38),
	.w1(32'hb99d5061),
	.w2(32'hb9904b18),
	.w3(32'hb9215670),
	.w4(32'hbaa36d01),
	.w5(32'h38873bd1),
	.w6(32'hbaba4f93),
	.w7(32'hbaa65c92),
	.w8(32'h39e92362),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55d0d3),
	.w1(32'hba8f742d),
	.w2(32'h3a14a5c9),
	.w3(32'hba8db73b),
	.w4(32'hba8e06e3),
	.w5(32'hb8fbd779),
	.w6(32'h3a770bd2),
	.w7(32'hba12a48d),
	.w8(32'h3979fbc9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a638281),
	.w1(32'hb9fb6809),
	.w2(32'hb998b8c5),
	.w3(32'hba086ec7),
	.w4(32'hba879503),
	.w5(32'hba61be7d),
	.w6(32'h3ab4e1c4),
	.w7(32'h3a897e11),
	.w8(32'h3b3eec15),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce5f11),
	.w1(32'hba218a10),
	.w2(32'hb8915851),
	.w3(32'hba130d99),
	.w4(32'hba84de36),
	.w5(32'hba75afab),
	.w6(32'hb982c4c1),
	.w7(32'h382e1fea),
	.w8(32'h39114a3b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8189),
	.w1(32'hba5d0951),
	.w2(32'h396e1071),
	.w3(32'hba5ba8af),
	.w4(32'h3871ac54),
	.w5(32'h39e5a3a1),
	.w6(32'hbaabfb14),
	.w7(32'hba890a07),
	.w8(32'hba275be9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d872ad),
	.w1(32'hb884e473),
	.w2(32'h39a58b5e),
	.w3(32'h39ca207e),
	.w4(32'h39323c5c),
	.w5(32'h39918098),
	.w6(32'hb8b76224),
	.w7(32'h377b8d16),
	.w8(32'h38c2ef0d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38948950),
	.w1(32'hb81d24bb),
	.w2(32'h3a0e8fbd),
	.w3(32'h395316bb),
	.w4(32'h39ad224a),
	.w5(32'h3a1cf2f8),
	.w6(32'hb8c86a1e),
	.w7(32'hb8987b18),
	.w8(32'h386588ef),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc51b1),
	.w1(32'hbaa88404),
	.w2(32'h3a3b6d79),
	.w3(32'h3a52328b),
	.w4(32'hbab6131e),
	.w5(32'hb9ff63a3),
	.w6(32'h3aaa190c),
	.w7(32'h3ae07031),
	.w8(32'h3ad0a52e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67974a),
	.w1(32'hbb0d5697),
	.w2(32'hbb2574b4),
	.w3(32'hb9b4340a),
	.w4(32'hbb10e324),
	.w5(32'hba915fdd),
	.w6(32'hbaff5173),
	.w7(32'hbb322699),
	.w8(32'hba0b304a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5ff08),
	.w1(32'hb99fb4b8),
	.w2(32'h3a8da67e),
	.w3(32'h39ebc718),
	.w4(32'hba946818),
	.w5(32'hb989a013),
	.w6(32'h3a333893),
	.w7(32'h3a0639bf),
	.w8(32'hb96c6e58),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db472c),
	.w1(32'h397fe5c3),
	.w2(32'h3a2c45c8),
	.w3(32'hba02a1e3),
	.w4(32'hb9c39bd8),
	.w5(32'h39bb1778),
	.w6(32'h3a34c451),
	.w7(32'h39ecdc8f),
	.w8(32'h39be2210),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a241b92),
	.w1(32'hb9483ace),
	.w2(32'h39833cea),
	.w3(32'h390405f9),
	.w4(32'hb941b9ee),
	.w5(32'hb92939a4),
	.w6(32'hb812f67d),
	.w7(32'h399b2fb1),
	.w8(32'h39332ff2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af6751),
	.w1(32'hbae5d570),
	.w2(32'h38de940a),
	.w3(32'hba421da4),
	.w4(32'hbb117130),
	.w5(32'hbaef0202),
	.w6(32'h3a198f06),
	.w7(32'h3a9e5d7e),
	.w8(32'h3845754b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba156e46),
	.w1(32'h3ac4f0bf),
	.w2(32'h3b15bbbe),
	.w3(32'h3915aa27),
	.w4(32'h3a08f0bb),
	.w5(32'h3a81bbdf),
	.w6(32'h3a46ce36),
	.w7(32'hb9f764e4),
	.w8(32'h39504874),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af12b40),
	.w1(32'h3b4379d1),
	.w2(32'h3ba1178d),
	.w3(32'h3abd3dbc),
	.w4(32'h3b0bf45d),
	.w5(32'h3b1eb18d),
	.w6(32'h3b4c0d9e),
	.w7(32'h3b36ec2e),
	.w8(32'h3b1d4a11),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fbc6d),
	.w1(32'hb9972a5b),
	.w2(32'hb8aa4bea),
	.w3(32'h39e4bf8d),
	.w4(32'hb9d0eb81),
	.w5(32'hb9efc139),
	.w6(32'hb9fd3fca),
	.w7(32'hb94c418c),
	.w8(32'hb9b4c17e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a061027),
	.w1(32'h3abaa428),
	.w2(32'h3a2ae2ef),
	.w3(32'h3a0c798f),
	.w4(32'h3a91b181),
	.w5(32'h38c6f270),
	.w6(32'h3ab81a89),
	.w7(32'h39f5ac8f),
	.w8(32'hb9da4d73),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule