module layer_10_featuremap_494(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a7cc6),
	.w1(32'hba41d94b),
	.w2(32'hba29282c),
	.w3(32'hbab14c4e),
	.w4(32'hbb212a36),
	.w5(32'hbb150e59),
	.w6(32'h39e9323d),
	.w7(32'hba4ca7d3),
	.w8(32'h3a76a2ba),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b0fb1),
	.w1(32'h3b91862f),
	.w2(32'h3af195f7),
	.w3(32'h3a887c60),
	.w4(32'h3b3db841),
	.w5(32'hb8f71925),
	.w6(32'h3b1d3534),
	.w7(32'h3ad7a48a),
	.w8(32'h39040a93),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb825e63c),
	.w1(32'hbb3137e2),
	.w2(32'h3a551375),
	.w3(32'hb993a153),
	.w4(32'hbb2027b5),
	.w5(32'hbb289444),
	.w6(32'hba709f4d),
	.w7(32'hba36f6a2),
	.w8(32'h38a251a1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90ae96),
	.w1(32'hba73c573),
	.w2(32'hba947243),
	.w3(32'hb9c740d6),
	.w4(32'hbad28554),
	.w5(32'hb91c15f6),
	.w6(32'hba77fb8f),
	.w7(32'hbadabfe7),
	.w8(32'h391c69ab),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba4127),
	.w1(32'h3aa05c0d),
	.w2(32'h3a512e8c),
	.w3(32'h3b28fd83),
	.w4(32'h3a42ff19),
	.w5(32'hba5cc3f5),
	.w6(32'h3abaf7fe),
	.w7(32'hb89a176d),
	.w8(32'hba0740a6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05cc99),
	.w1(32'hbacf4de2),
	.w2(32'hba759e78),
	.w3(32'hb7750b09),
	.w4(32'h3aa64f2e),
	.w5(32'hba12306c),
	.w6(32'hbaa073d5),
	.w7(32'hb894ee3e),
	.w8(32'hbaa8dbb1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa66ac8),
	.w1(32'h3a34e629),
	.w2(32'h3aab6d4b),
	.w3(32'hba7367df),
	.w4(32'hb9d806dc),
	.w5(32'h39044eff),
	.w6(32'hba0fda36),
	.w7(32'hba4bfa8f),
	.w8(32'h3a10ab24),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dcf92),
	.w1(32'hbb97e0c1),
	.w2(32'hbb9f471c),
	.w3(32'hbbbe9ce1),
	.w4(32'hbbacf3d0),
	.w5(32'hbbcbfa0e),
	.w6(32'hbbd84dbd),
	.w7(32'hbb96951d),
	.w8(32'hbb60d667),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2353d4),
	.w1(32'hb9025c4e),
	.w2(32'h3921d706),
	.w3(32'h39fc6f0a),
	.w4(32'h3a589a08),
	.w5(32'h37c6efad),
	.w6(32'h3b0a2c0b),
	.w7(32'hbab0c086),
	.w8(32'hba8ceac4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39226),
	.w1(32'h3b730095),
	.w2(32'h3c0e3837),
	.w3(32'h3af9e6b7),
	.w4(32'h3ae8e5bd),
	.w5(32'h3be09c43),
	.w6(32'hb7986c8e),
	.w7(32'h3b1eabd2),
	.w8(32'h3b501be7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb3595),
	.w1(32'hbaa4ec02),
	.w2(32'hba6235fb),
	.w3(32'h3a1b39e5),
	.w4(32'hb9d8c607),
	.w5(32'hbaa5e0c9),
	.w6(32'h390e299f),
	.w7(32'h3a92d4f9),
	.w8(32'h3998870b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f5c70),
	.w1(32'hb99ab7d5),
	.w2(32'hbb213268),
	.w3(32'hbb089278),
	.w4(32'h3a75b8fb),
	.w5(32'hba03caea),
	.w6(32'hbb1ada33),
	.w7(32'hbab7a36c),
	.w8(32'hbaecc7d8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0929b6),
	.w1(32'h3ac8e72d),
	.w2(32'h3a9deff4),
	.w3(32'h3a9a1ef5),
	.w4(32'h3adb4a3e),
	.w5(32'h3b53aa68),
	.w6(32'h3a09d170),
	.w7(32'hb9b6c9b1),
	.w8(32'h3afb1f17),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c5624),
	.w1(32'h3908c0a3),
	.w2(32'h39efdd88),
	.w3(32'h3ac627c4),
	.w4(32'h39beb62c),
	.w5(32'hba4f6f2d),
	.w6(32'h3b03efc9),
	.w7(32'h3ac90ef5),
	.w8(32'hb98d3ca5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d0092),
	.w1(32'hba95a298),
	.w2(32'h3a86f32a),
	.w3(32'h3b2dfbe4),
	.w4(32'hb8efcf3e),
	.w5(32'hbac189d6),
	.w6(32'h3b2e0326),
	.w7(32'hb9c603db),
	.w8(32'hbac8f157),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807ae8e),
	.w1(32'hbaa35264),
	.w2(32'h3a61fa0a),
	.w3(32'hb9a8bf7e),
	.w4(32'hb9b7343f),
	.w5(32'h3b6e44e8),
	.w6(32'hbacf17ba),
	.w7(32'hbb6b5d53),
	.w8(32'h3aabc7fb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b5c80),
	.w1(32'hb8cadc6d),
	.w2(32'hb944c33c),
	.w3(32'h37ab6a0f),
	.w4(32'hba87f83b),
	.w5(32'hbaa5a563),
	.w6(32'hba29c42d),
	.w7(32'hba8e7cf2),
	.w8(32'hbabd6ff6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196a95),
	.w1(32'hbc54b68f),
	.w2(32'hbc6a612e),
	.w3(32'hbc812c07),
	.w4(32'hbc2ef740),
	.w5(32'hbc063805),
	.w6(32'hbc76411a),
	.w7(32'hbc1ed6c9),
	.w8(32'hbbdabbf0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba344cc0),
	.w1(32'hbb95056c),
	.w2(32'hbb928da9),
	.w3(32'hbb457041),
	.w4(32'hba880fca),
	.w5(32'hbaaa0f39),
	.w6(32'hbb9df34b),
	.w7(32'hbb20eb0d),
	.w8(32'hba55613e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae47a93),
	.w1(32'hbab78b1f),
	.w2(32'hbb8922d3),
	.w3(32'hba1ea61d),
	.w4(32'hb9de1e87),
	.w5(32'hba730094),
	.w6(32'hb8ccb0b3),
	.w7(32'hba0daa19),
	.w8(32'h3a0e7653),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3d0d),
	.w1(32'hbaadf885),
	.w2(32'hb981a590),
	.w3(32'hbb1bc3d5),
	.w4(32'h3ad0210c),
	.w5(32'hb9c9db79),
	.w6(32'hbaaa8e32),
	.w7(32'h3a993332),
	.w8(32'h39bce536),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5b95b),
	.w1(32'h3a950475),
	.w2(32'hbb1e6d7f),
	.w3(32'h3b2cd238),
	.w4(32'h3a21ccbd),
	.w5(32'hbb178c6e),
	.w6(32'h3b17d85a),
	.w7(32'h3a284208),
	.w8(32'hbb45d497),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2815b3),
	.w1(32'hbc94edb6),
	.w2(32'hbc704248),
	.w3(32'hbc41594e),
	.w4(32'hbc31072d),
	.w5(32'hbbd04d35),
	.w6(32'hbc8338d3),
	.w7(32'hbc06a129),
	.w8(32'hbc3730d1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3fe45),
	.w1(32'hb97d13ee),
	.w2(32'h3b201b5e),
	.w3(32'h3b85d4f3),
	.w4(32'h3a3277fb),
	.w5(32'h3b38a669),
	.w6(32'h3a5dbc50),
	.w7(32'hba0d09d3),
	.w8(32'hb932fe75),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe01ed),
	.w1(32'h3b6d4adb),
	.w2(32'h3b875ed2),
	.w3(32'h3b94edab),
	.w4(32'h3b73fbcd),
	.w5(32'h3b71c6fc),
	.w6(32'h3b168ac0),
	.w7(32'hba0b0722),
	.w8(32'h3a5a9edb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79844f),
	.w1(32'hbaec3713),
	.w2(32'hbb3cd215),
	.w3(32'hba8326cd),
	.w4(32'hb9c5f0e4),
	.w5(32'hbaf7e98f),
	.w6(32'hbb0bd407),
	.w7(32'hb707b83a),
	.w8(32'h39d453a3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40173),
	.w1(32'h3a87d055),
	.w2(32'h39796989),
	.w3(32'hbae93791),
	.w4(32'h3a675500),
	.w5(32'h3b6a858e),
	.w6(32'h39d0323d),
	.w7(32'h3ac0ba9e),
	.w8(32'h3b735b5b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf251e),
	.w1(32'h3b72eb53),
	.w2(32'h3b833bc1),
	.w3(32'h3c0a0121),
	.w4(32'h3b8088f3),
	.w5(32'h3a49db47),
	.w6(32'h3beaabdc),
	.w7(32'h3ac6f3d8),
	.w8(32'h38a7867e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c49cd),
	.w1(32'hbad54caf),
	.w2(32'hb90f48b4),
	.w3(32'h3aad5a93),
	.w4(32'hba44ef01),
	.w5(32'h3ad2b86b),
	.w6(32'hb99c9c10),
	.w7(32'h397dcfae),
	.w8(32'h3a007153),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5765a9),
	.w1(32'h3b9d2b3e),
	.w2(32'h3befaf45),
	.w3(32'h3bb3c23f),
	.w4(32'h3ba1ec18),
	.w5(32'h3b8c3f59),
	.w6(32'h3bb45234),
	.w7(32'h3b8a38d9),
	.w8(32'h3b741f78),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfdef2),
	.w1(32'hba205e2f),
	.w2(32'h3abaf735),
	.w3(32'h3aa006ce),
	.w4(32'hbaf25288),
	.w5(32'h3a7bc4ca),
	.w6(32'h3aef31e5),
	.w7(32'h3a2a3a32),
	.w8(32'hb8d60edd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dc7d1),
	.w1(32'h38ea96eb),
	.w2(32'h39cd0707),
	.w3(32'hb7bfc11e),
	.w4(32'h3a8b1d7e),
	.w5(32'h382812b3),
	.w6(32'hb99c343f),
	.w7(32'h3aaddadb),
	.w8(32'h3a2521b8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aece023),
	.w1(32'h3b4af5f2),
	.w2(32'h3b052ef6),
	.w3(32'h3b0ae538),
	.w4(32'h3a2cd667),
	.w5(32'h3b2c8cc5),
	.w6(32'h3ad06e27),
	.w7(32'h3af9a1cd),
	.w8(32'h3aeac14d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab71d3e),
	.w1(32'h3b610b6d),
	.w2(32'h3bbd4917),
	.w3(32'h3af18795),
	.w4(32'h3a8e1985),
	.w5(32'h3b377dc9),
	.w6(32'hb9f2b11d),
	.w7(32'h3a306d50),
	.w8(32'h3ade01fb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5d18b),
	.w1(32'h3b2cb3dc),
	.w2(32'h3aa94c17),
	.w3(32'h3a4d7f6e),
	.w4(32'h3af5ccb1),
	.w5(32'hba9a5c49),
	.w6(32'h3ac3f983),
	.w7(32'h3a9c6fd4),
	.w8(32'h3b0e2c76),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38209931),
	.w1(32'h3925ef86),
	.w2(32'h38c3ecdf),
	.w3(32'h39de80c6),
	.w4(32'hb96d3c7b),
	.w5(32'h3a0db9ef),
	.w6(32'hba69f2d6),
	.w7(32'hbb2c6283),
	.w8(32'hbaf3a74d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c6c7),
	.w1(32'hbb42bcdc),
	.w2(32'hbb33ea5c),
	.w3(32'hbaa6d52c),
	.w4(32'hbb65a791),
	.w5(32'hba609a22),
	.w6(32'hbb94cd6d),
	.w7(32'hb9bbfd27),
	.w8(32'h3956a04e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd8446),
	.w1(32'h3c5abef1),
	.w2(32'h3c0722cd),
	.w3(32'h3c451d45),
	.w4(32'h3c27b04d),
	.w5(32'h3ace7114),
	.w6(32'h3c154a07),
	.w7(32'h3bdbc5fe),
	.w8(32'h3b006124),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1393d7),
	.w1(32'h3c0d8220),
	.w2(32'h3bae1f8e),
	.w3(32'h3c3dbe4b),
	.w4(32'h3ba24ae2),
	.w5(32'hbb0e5441),
	.w6(32'h3c27beec),
	.w7(32'h3b0e278e),
	.w8(32'h3a6bf1f3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ace2a8),
	.w1(32'h3b254d85),
	.w2(32'h3ab59e4d),
	.w3(32'h3aaad4fa),
	.w4(32'h3ab68c2c),
	.w5(32'h3a808cc2),
	.w6(32'h3b039c8a),
	.w7(32'h3b0e3cac),
	.w8(32'h3a615ba9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abecdf5),
	.w1(32'h3af77502),
	.w2(32'hba926a2e),
	.w3(32'h3a9ee9c1),
	.w4(32'hba855431),
	.w5(32'h3b0be3f8),
	.w6(32'h3a918ab1),
	.w7(32'h3a965114),
	.w8(32'h3a809958),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a304c3b),
	.w1(32'hba4e2bff),
	.w2(32'hb9a2652c),
	.w3(32'h3a921393),
	.w4(32'h3adf1840),
	.w5(32'h3839a2f4),
	.w6(32'h3b036e26),
	.w7(32'h38c1f2f6),
	.w8(32'hba84d9ea),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0d524),
	.w1(32'hba0581fe),
	.w2(32'hbb3571b5),
	.w3(32'hba8904b4),
	.w4(32'hb9dd8222),
	.w5(32'hb95c5b5f),
	.w6(32'hba8ce06c),
	.w7(32'hbaee0449),
	.w8(32'hba2f971d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb271cb5),
	.w1(32'hbadce66f),
	.w2(32'hb974d49a),
	.w3(32'hba998207),
	.w4(32'hbb1e706c),
	.w5(32'h3a88816e),
	.w6(32'hbb6246de),
	.w7(32'hbab9024e),
	.w8(32'h3ae32c76),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb734),
	.w1(32'h3adfb6d6),
	.w2(32'h3b980656),
	.w3(32'h3b3bdc7e),
	.w4(32'h3b7fb34e),
	.w5(32'h3bc54d86),
	.w6(32'h3b6cbb0b),
	.w7(32'h3b52bc17),
	.w8(32'h3ae99724),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ad4db),
	.w1(32'hb9b6dbfb),
	.w2(32'h3bc9c966),
	.w3(32'h3b44c49b),
	.w4(32'hbae35bea),
	.w5(32'h3b750e60),
	.w6(32'h3b175e8d),
	.w7(32'hbb3d22c6),
	.w8(32'h3afdbb87),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad99f92),
	.w1(32'hbb20642d),
	.w2(32'hba410952),
	.w3(32'hb9c2ded3),
	.w4(32'hbb4e79b6),
	.w5(32'h3a808e7a),
	.w6(32'hbb92fd2e),
	.w7(32'hbb897e6c),
	.w8(32'hb9562dd1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8cec),
	.w1(32'hbc60f4f0),
	.w2(32'hbc831263),
	.w3(32'hbc621f8c),
	.w4(32'hbc1f6309),
	.w5(32'hbbe9097f),
	.w6(32'hbc80a520),
	.w7(32'hbbfb7d25),
	.w8(32'hbb680453),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d84f10),
	.w1(32'h3ab72467),
	.w2(32'h3a925dbe),
	.w3(32'hba89470d),
	.w4(32'h3ab202d8),
	.w5(32'h3a249142),
	.w6(32'hb90fce2a),
	.w7(32'h3a0ac7c9),
	.w8(32'hb8183206),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32a2c8),
	.w1(32'hba6d9254),
	.w2(32'hb98a9063),
	.w3(32'h3aebb54c),
	.w4(32'hb91ab0a7),
	.w5(32'h3a8435c7),
	.w6(32'hba5560f0),
	.w7(32'hbac272a4),
	.w8(32'hbabf6a90),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfcf79),
	.w1(32'hb7d14672),
	.w2(32'hba31fcf3),
	.w3(32'h3b4df1a8),
	.w4(32'h394ffff9),
	.w5(32'hb921f0e6),
	.w6(32'h3a5298a6),
	.w7(32'hba8536c6),
	.w8(32'hba3dd9cf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac98146),
	.w1(32'hb9c6e7ba),
	.w2(32'hba77a3cc),
	.w3(32'hb9133614),
	.w4(32'hbb471e72),
	.w5(32'hbb0704ea),
	.w6(32'hba5a93ce),
	.w7(32'hbb7387ab),
	.w8(32'hbadcb37b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ed24),
	.w1(32'hbac3ef8e),
	.w2(32'hba85378f),
	.w3(32'hba69521a),
	.w4(32'h39b76a02),
	.w5(32'hb99b888d),
	.w6(32'hbb3ae8b5),
	.w7(32'hb8c684d6),
	.w8(32'hba04670f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e8c4),
	.w1(32'hbbfe42b4),
	.w2(32'hbc016ad4),
	.w3(32'hbc17bf40),
	.w4(32'hbc0b0361),
	.w5(32'hbb3863aa),
	.w6(32'hbc1e0139),
	.w7(32'hbb925a27),
	.w8(32'hbaa351f3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba608fbf),
	.w1(32'h3ac00057),
	.w2(32'hbace1217),
	.w3(32'h39d0e8a1),
	.w4(32'h3b28da54),
	.w5(32'hbab07e10),
	.w6(32'hb941b05b),
	.w7(32'h3af2b55f),
	.w8(32'h3a1ed859),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a321a),
	.w1(32'h39b2f2c1),
	.w2(32'hbb1ddae5),
	.w3(32'h3aadcf50),
	.w4(32'h3a450ada),
	.w5(32'hbb21313f),
	.w6(32'h3ad0829c),
	.w7(32'hba6662ca),
	.w8(32'hbb6235a1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39143924),
	.w1(32'h39e0257b),
	.w2(32'h39b1fea1),
	.w3(32'h3a53f4f6),
	.w4(32'hba3a0fe8),
	.w5(32'hbad199ef),
	.w6(32'hbafda459),
	.w7(32'hbae7d69c),
	.w8(32'hba4f3b3f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9e5a7),
	.w1(32'hba95c87d),
	.w2(32'h3a99b57c),
	.w3(32'hbaa97c83),
	.w4(32'hb98346ac),
	.w5(32'h3a94fd06),
	.w6(32'hb8685c9c),
	.w7(32'h3906ff6a),
	.w8(32'h3a0a36bb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e400da),
	.w1(32'h3b1fa247),
	.w2(32'h3b007c43),
	.w3(32'h3a96d675),
	.w4(32'h3b33432d),
	.w5(32'h3b152591),
	.w6(32'hb8c473e5),
	.w7(32'h3af95473),
	.w8(32'h3b7f1590),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a900939),
	.w1(32'hba53bc00),
	.w2(32'h38f197e6),
	.w3(32'h3a36d8d2),
	.w4(32'hba3ca6da),
	.w5(32'hba4b3d30),
	.w6(32'h3a9f7fb4),
	.w7(32'hba88d332),
	.w8(32'h3ae2fb78),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb286467),
	.w1(32'hbbdf742a),
	.w2(32'hbbba1760),
	.w3(32'hbb966e58),
	.w4(32'hbb892cb8),
	.w5(32'hbb602da5),
	.w6(32'hbba44bce),
	.w7(32'hbb5158ba),
	.w8(32'hbb5f3f0b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16e2f),
	.w1(32'hbba69a53),
	.w2(32'hbb5a4840),
	.w3(32'hbbc78fbd),
	.w4(32'hbaf3ed20),
	.w5(32'hbb8ebed1),
	.w6(32'hbb91f2c2),
	.w7(32'hbb695140),
	.w8(32'hbb96b81f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f550f),
	.w1(32'h39acee00),
	.w2(32'hbb337d9f),
	.w3(32'h396d1518),
	.w4(32'h3a124e62),
	.w5(32'hbac17f53),
	.w6(32'hb9fedd0f),
	.w7(32'h3956a8b2),
	.w8(32'hba6f02e5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45140f),
	.w1(32'hba153b05),
	.w2(32'hba18da13),
	.w3(32'h3a6c09ab),
	.w4(32'hb9ef051d),
	.w5(32'hba349f63),
	.w6(32'hba2474d4),
	.w7(32'h3787ce44),
	.w8(32'h3a7c013c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82d38),
	.w1(32'h3b3ca7ac),
	.w2(32'h3b54b58c),
	.w3(32'hba99cf87),
	.w4(32'h3b58d6d7),
	.w5(32'h3b5339c5),
	.w6(32'hba401459),
	.w7(32'h3b8a2fe3),
	.w8(32'h3b652d51),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420f51),
	.w1(32'hb986c46a),
	.w2(32'h3997ed88),
	.w3(32'h3b6a1b3d),
	.w4(32'h3a8d38be),
	.w5(32'h3a8b4b53),
	.w6(32'h3b82b108),
	.w7(32'hb822caa5),
	.w8(32'h3a087036),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba878f49),
	.w1(32'hbb202f28),
	.w2(32'hbb25488c),
	.w3(32'hba81af91),
	.w4(32'hba65ffd1),
	.w5(32'hbb0c2928),
	.w6(32'hba94d9da),
	.w7(32'hba825dad),
	.w8(32'hbb68e1ca),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60cbd6),
	.w1(32'h3ab007b4),
	.w2(32'h3b8ff75f),
	.w3(32'h3b2b06b1),
	.w4(32'h3a4bd8b8),
	.w5(32'h3ad9a9fa),
	.w6(32'h3a00a70a),
	.w7(32'hbacea421),
	.w8(32'h3a601e04),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca714c),
	.w1(32'hbbdbf9e2),
	.w2(32'hbc10ff3f),
	.w3(32'hbb90d269),
	.w4(32'hbb34eebb),
	.w5(32'hbbcc4c3d),
	.w6(32'hbbd0b0e0),
	.w7(32'hbbc351a9),
	.w8(32'hbb991bc1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca849a),
	.w1(32'h3bced158),
	.w2(32'h3c50dbbe),
	.w3(32'h3be2e129),
	.w4(32'h3b81b6bc),
	.w5(32'h3be22606),
	.w6(32'h3ba9f599),
	.w7(32'h3b4c5171),
	.w8(32'h3bb6dbb1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a76bf),
	.w1(32'hbaafc620),
	.w2(32'hbac80f13),
	.w3(32'h395da45c),
	.w4(32'hb9b945e7),
	.w5(32'hba5103e4),
	.w6(32'hb9fdbd3f),
	.w7(32'hb9a577b1),
	.w8(32'hb8ca4938),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bc884),
	.w1(32'hbad5c5a5),
	.w2(32'hbaf8c657),
	.w3(32'hba5f128c),
	.w4(32'hbb627769),
	.w5(32'hbb6d3748),
	.w6(32'h3a2491b3),
	.w7(32'hbabe13a7),
	.w8(32'hba99e85c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c197c3),
	.w1(32'h39a975a5),
	.w2(32'h3a0913dc),
	.w3(32'hbad27c66),
	.w4(32'h3ac2124b),
	.w5(32'h3ab1271a),
	.w6(32'hba6e9583),
	.w7(32'h3a98751b),
	.w8(32'h3ab71754),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fe4a2),
	.w1(32'hba8b42c2),
	.w2(32'hbac7211e),
	.w3(32'hbadda231),
	.w4(32'hba338ffd),
	.w5(32'hb9b9834f),
	.w6(32'hba841db3),
	.w7(32'hba87d080),
	.w8(32'hba39b967),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39988513),
	.w1(32'hba5fd997),
	.w2(32'hb99caf52),
	.w3(32'h3a0ef9fe),
	.w4(32'hb934f0f0),
	.w5(32'hba9b9bed),
	.w6(32'h3a0e275a),
	.w7(32'h3911d130),
	.w8(32'hb9e53de1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a56c2),
	.w1(32'hbbe05a82),
	.w2(32'hbbc76c31),
	.w3(32'hbbf2ac2c),
	.w4(32'hbc0f27f4),
	.w5(32'hbb6ffb99),
	.w6(32'hbc356395),
	.w7(32'hbbc6d9fd),
	.w8(32'hbb6eb839),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839d5b),
	.w1(32'hbbfd6669),
	.w2(32'hbc26f54a),
	.w3(32'hbc19a7cd),
	.w4(32'hbc1f1a38),
	.w5(32'hbb450ae1),
	.w6(32'hbc5e7b7f),
	.w7(32'hbbca88df),
	.w8(32'hbb681d6e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6b44a),
	.w1(32'h3b899445),
	.w2(32'h3baeddcc),
	.w3(32'h3c091291),
	.w4(32'h3b743a78),
	.w5(32'h3bac839d),
	.w6(32'h3bf7d29f),
	.w7(32'h3ba81552),
	.w8(32'h3b964cc8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bb1c5),
	.w1(32'hbb75ab29),
	.w2(32'hbab72fbc),
	.w3(32'hba8e487c),
	.w4(32'hbaff5120),
	.w5(32'hba113cf3),
	.w6(32'hbb03aae8),
	.w7(32'hbafe5d05),
	.w8(32'hba98ac7a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98493fc),
	.w1(32'h3a84c076),
	.w2(32'hb96374d0),
	.w3(32'h3a7c42b3),
	.w4(32'h3aa9945b),
	.w5(32'h3b3c87c8),
	.w6(32'hbadedf1a),
	.w7(32'h3a1cf107),
	.w8(32'h3a88988b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8656395),
	.w1(32'h3aab59c5),
	.w2(32'h3b422cda),
	.w3(32'h39c52765),
	.w4(32'h3a8d26b7),
	.w5(32'h3a45a433),
	.w6(32'h3afe1451),
	.w7(32'h3a68a2a8),
	.w8(32'h3aa6ce31),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40d882),
	.w1(32'hbbf026ca),
	.w2(32'hbc02de1f),
	.w3(32'hbaf36141),
	.w4(32'hbba9a761),
	.w5(32'hbb4e8cef),
	.w6(32'hbb4b6b4f),
	.w7(32'hbb963fed),
	.w8(32'hbb335fbb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75b71b),
	.w1(32'h3a15a8ca),
	.w2(32'h3a4a4b6d),
	.w3(32'hba6f7735),
	.w4(32'hb8a2ac87),
	.w5(32'h394feaec),
	.w6(32'hba9071a7),
	.w7(32'h3a2af6d4),
	.w8(32'h3a9f5a5d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a911d10),
	.w1(32'hb9b86baa),
	.w2(32'h3a4cf8d1),
	.w3(32'h39ead41b),
	.w4(32'hb9300bce),
	.w5(32'h3aecbc6d),
	.w6(32'h3abb8573),
	.w7(32'h399287e4),
	.w8(32'hba28eab3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b601b0),
	.w1(32'hbae35168),
	.w2(32'hbac45691),
	.w3(32'hbadafc72),
	.w4(32'hbacab07a),
	.w5(32'hb9ac9f8d),
	.w6(32'hbafc01cf),
	.w7(32'hba43f762),
	.w8(32'hb9d51f2a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabdeb4),
	.w1(32'h395b6193),
	.w2(32'h3a9825ae),
	.w3(32'hbaea8765),
	.w4(32'hba62add5),
	.w5(32'hbad0659b),
	.w6(32'hba5b75c4),
	.w7(32'hba2337c2),
	.w8(32'hbafe4881),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b91d),
	.w1(32'h3b448f85),
	.w2(32'h3b8912c3),
	.w3(32'h3b5d09ad),
	.w4(32'h3b3b0330),
	.w5(32'h3b89684e),
	.w6(32'h3a9fcbe7),
	.w7(32'h3b4e590f),
	.w8(32'h3aae2ca7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7cf60),
	.w1(32'h3a72f0bd),
	.w2(32'hb860ba9d),
	.w3(32'h3a0a488b),
	.w4(32'h3aa17422),
	.w5(32'hb98a74fb),
	.w6(32'hb9ea6800),
	.w7(32'h3aaea813),
	.w8(32'hb873d76a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac578bc),
	.w1(32'hbae4620e),
	.w2(32'h3a1ee77a),
	.w3(32'hba48ecf7),
	.w4(32'h39fe33f4),
	.w5(32'h3b754bbb),
	.w6(32'h3a3e4df1),
	.w7(32'h3a22a7a2),
	.w8(32'h3b0ac0f4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ca8c),
	.w1(32'hbc47ae42),
	.w2(32'hbc2dce7e),
	.w3(32'hbc8134aa),
	.w4(32'hbc3c211e),
	.w5(32'hbb85da5e),
	.w6(32'hbca22113),
	.w7(32'hbc22ff38),
	.w8(32'hbbb17d14),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866b4f),
	.w1(32'hb8a751ca),
	.w2(32'hba82d695),
	.w3(32'h3ba54c30),
	.w4(32'h390b4b2c),
	.w5(32'h3a11c065),
	.w6(32'h3b48c7a1),
	.w7(32'h3a39d9e5),
	.w8(32'hba5798e6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e7aa),
	.w1(32'hbaaa3d28),
	.w2(32'hb9aa96f7),
	.w3(32'hbb48e15a),
	.w4(32'hba58364d),
	.w5(32'h3ad96fe3),
	.w6(32'hb96333d0),
	.w7(32'h3a9eb8c2),
	.w8(32'h39964233),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32f968),
	.w1(32'h3b8610de),
	.w2(32'h3b71576c),
	.w3(32'h3b68c377),
	.w4(32'h3b068211),
	.w5(32'h3aa99e94),
	.w6(32'h3b15e269),
	.w7(32'h3ac26cdc),
	.w8(32'h3aba7fbb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926972),
	.w1(32'hbb88ee9e),
	.w2(32'hb9ea919d),
	.w3(32'hbbb9b26e),
	.w4(32'hbb87e62e),
	.w5(32'hba0f0e28),
	.w6(32'hbb478282),
	.w7(32'hbbb03f3c),
	.w8(32'hbb63fc36),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7ae44),
	.w1(32'h3aa638e2),
	.w2(32'h3af884d4),
	.w3(32'h3a971b93),
	.w4(32'h3b0a3c2a),
	.w5(32'h3ad57b78),
	.w6(32'hb779393f),
	.w7(32'hb90ff0d5),
	.w8(32'hb899de71),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c4d34),
	.w1(32'h3b7f5cbd),
	.w2(32'h3b8a5af0),
	.w3(32'h3b362c59),
	.w4(32'h3b34f463),
	.w5(32'h3ba9633d),
	.w6(32'h3b39b7ed),
	.w7(32'h3ac6c8aa),
	.w8(32'h3b2d7b64),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab92cc2),
	.w1(32'h3a2d8ff0),
	.w2(32'hba4f90c6),
	.w3(32'h3a1164fd),
	.w4(32'h39f2efe9),
	.w5(32'h397ad90d),
	.w6(32'h3aefeccc),
	.w7(32'hb923298d),
	.w8(32'hb9c1f9f6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a3f7a),
	.w1(32'hba5f540e),
	.w2(32'h3b1c5e17),
	.w3(32'hbac1fc4c),
	.w4(32'hba4b7644),
	.w5(32'h3b5b12d7),
	.w6(32'hba47f3a0),
	.w7(32'hba6514a7),
	.w8(32'h3b0891bc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71f397),
	.w1(32'hba1f5596),
	.w2(32'h397d88d1),
	.w3(32'h3a802c2b),
	.w4(32'hb9516e53),
	.w5(32'h3ac2c3f7),
	.w6(32'hb7f964ec),
	.w7(32'hbaa71e63),
	.w8(32'hbb6eda3d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f24b),
	.w1(32'hbc544ecb),
	.w2(32'hbc44d4e9),
	.w3(32'hbc255650),
	.w4(32'hbc33a31b),
	.w5(32'hbb8a4b5c),
	.w6(32'hbc60d7ad),
	.w7(32'hbc04f2c1),
	.w8(32'hbb8e7a79),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e58c7),
	.w1(32'h3ba6a461),
	.w2(32'h3b3b33db),
	.w3(32'h3c1d0a4f),
	.w4(32'h3b8c1af7),
	.w5(32'h3ab8487a),
	.w6(32'h3c0f65ca),
	.w7(32'h3b5cc7bd),
	.w8(32'h3aa2fb0b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad9060),
	.w1(32'h3ba4717d),
	.w2(32'h3c04d3a7),
	.w3(32'h3bab038f),
	.w4(32'h3b408567),
	.w5(32'h3bee1418),
	.w6(32'h3b84e981),
	.w7(32'h3ab31c98),
	.w8(32'h3b97dc59),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09943),
	.w1(32'hbbdfec4b),
	.w2(32'hbc121ca7),
	.w3(32'hbbdb76d5),
	.w4(32'hbba654d3),
	.w5(32'hbbc7722d),
	.w6(32'hbba2b679),
	.w7(32'hbb50220c),
	.w8(32'hbb926774),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba224486),
	.w1(32'hbaa6cd08),
	.w2(32'hbac79c2b),
	.w3(32'hbab36d94),
	.w4(32'hbb097bb4),
	.w5(32'hbae1151a),
	.w6(32'hb9fa7f36),
	.w7(32'hba8a9372),
	.w8(32'hbaf75f05),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2af227),
	.w1(32'hbc97b647),
	.w2(32'hbc96c7f5),
	.w3(32'hbc5bfd24),
	.w4(32'hbc8ee001),
	.w5(32'hbc38b561),
	.w6(32'hbc9004ed),
	.w7(32'hbc6159e6),
	.w8(32'hbc0037e7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e6cdd),
	.w1(32'h3afea307),
	.w2(32'h3aae0e61),
	.w3(32'h3b85b2c8),
	.w4(32'hb9bb4dfa),
	.w5(32'hb9e87e52),
	.w6(32'h3baf4d2f),
	.w7(32'h3a6cb01a),
	.w8(32'hba624c6a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7ad0d),
	.w1(32'h3a4d31a6),
	.w2(32'h39b72b6d),
	.w3(32'h3a1e57ba),
	.w4(32'h3a9a3b46),
	.w5(32'h3a39d291),
	.w6(32'h3a40c58b),
	.w7(32'h3a0c1d8d),
	.w8(32'h39f530a0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46e2dc),
	.w1(32'h3aa4bc2a),
	.w2(32'h3b201edd),
	.w3(32'hba12fa4f),
	.w4(32'hb831651c),
	.w5(32'h39fc5149),
	.w6(32'hba5fd30a),
	.w7(32'hb88ced79),
	.w8(32'hb998423c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bda43),
	.w1(32'h3b1540ff),
	.w2(32'h3b2d1c53),
	.w3(32'h3ba91642),
	.w4(32'h39c4701c),
	.w5(32'h3b0fe4b9),
	.w6(32'h3b6e4314),
	.w7(32'h39c2a760),
	.w8(32'h3ae69060),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9043ae),
	.w1(32'h3b8c6862),
	.w2(32'h3c047f33),
	.w3(32'h3b2dc709),
	.w4(32'h3a8ced91),
	.w5(32'h3c0d208b),
	.w6(32'h3b450aa5),
	.w7(32'h3a363bff),
	.w8(32'h3b86f499),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4b67b),
	.w1(32'h3a53256b),
	.w2(32'h3b0adbe9),
	.w3(32'h38913c75),
	.w4(32'h3a29f452),
	.w5(32'h398b8e1a),
	.w6(32'h3b18fe8b),
	.w7(32'hba2c21f5),
	.w8(32'hba834c14),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24139f),
	.w1(32'hba697d6f),
	.w2(32'h3a5742ba),
	.w3(32'h3abcf6d5),
	.w4(32'hbaba2035),
	.w5(32'h3a684f26),
	.w6(32'h3939a67c),
	.w7(32'hba862bd0),
	.w8(32'h3a4b86de),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a697a0e),
	.w1(32'h39fa5202),
	.w2(32'hb9577501),
	.w3(32'h3970278e),
	.w4(32'h3a355b2e),
	.w5(32'h3aa039ff),
	.w6(32'h3a25adac),
	.w7(32'h38f0b491),
	.w8(32'h3a1b08b1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a6dc),
	.w1(32'hbb6d84c9),
	.w2(32'hba6475ee),
	.w3(32'hbaea6a8f),
	.w4(32'hbba794a3),
	.w5(32'hbac77e8e),
	.w6(32'hba3b478e),
	.w7(32'hbb96b7ab),
	.w8(32'hbb06138a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa243ff),
	.w1(32'h3b1736da),
	.w2(32'h3b8f5e5a),
	.w3(32'h3963fd01),
	.w4(32'h3b049411),
	.w5(32'h3b6f0abc),
	.w6(32'h39a3c39d),
	.w7(32'h3ab9c0dc),
	.w8(32'h3b19cbe0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89d59d),
	.w1(32'h392b4c22),
	.w2(32'hb9176bdc),
	.w3(32'h3a97ffd6),
	.w4(32'hb951b745),
	.w5(32'hba29b6b2),
	.w6(32'h3abd3d29),
	.w7(32'h394d56b6),
	.w8(32'hba0880a9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10587c),
	.w1(32'h3a4c9934),
	.w2(32'h3ae02d84),
	.w3(32'h3b1997b9),
	.w4(32'h39efc727),
	.w5(32'h3b36046d),
	.w6(32'h3b2fe5ea),
	.w7(32'h3908d76a),
	.w8(32'h3a1dd95c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ec31e),
	.w1(32'h3a01867f),
	.w2(32'h3942cd3e),
	.w3(32'h3a45ee74),
	.w4(32'hb9c7810d),
	.w5(32'h396ac78c),
	.w6(32'h3adfa6c7),
	.w7(32'hb922a43e),
	.w8(32'hb8f6b3d5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0a84),
	.w1(32'h3aa1a001),
	.w2(32'h3ac7ce51),
	.w3(32'h3a49c5d7),
	.w4(32'h3a89e4d5),
	.w5(32'hb9e11da9),
	.w6(32'h3a5a75c1),
	.w7(32'h3ac754bb),
	.w8(32'h3a5fb5d9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae55e98),
	.w1(32'h3aeeecf3),
	.w2(32'h3b66538b),
	.w3(32'h3b662044),
	.w4(32'h3abd0341),
	.w5(32'h3b64b246),
	.w6(32'h3b4dcb98),
	.w7(32'h3a8c8493),
	.w8(32'h3b344372),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef9e13),
	.w1(32'hba274cca),
	.w2(32'hb97770a6),
	.w3(32'h3a53d7eb),
	.w4(32'h3ab35749),
	.w5(32'h3b0c0f19),
	.w6(32'h3abcd58b),
	.w7(32'h3ab5819d),
	.w8(32'h3a6012b7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb377d9b),
	.w1(32'hbac0d1bf),
	.w2(32'hbb271a3b),
	.w3(32'hbafe704e),
	.w4(32'hbaa7570c),
	.w5(32'hbafe45da),
	.w6(32'hbb52ca93),
	.w7(32'hbb2fe108),
	.w8(32'hba380c90),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0558e),
	.w1(32'h3be50248),
	.w2(32'h3b9d1c65),
	.w3(32'h3bc6e5b6),
	.w4(32'h3bc0df09),
	.w5(32'h3a280dde),
	.w6(32'h3bbb73fe),
	.w7(32'h3b6a2088),
	.w8(32'hb9ba9b5f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab816e4),
	.w1(32'hb94197fe),
	.w2(32'hba4558bd),
	.w3(32'hbaf0f602),
	.w4(32'hba5ea368),
	.w5(32'hba2b545d),
	.w6(32'h39300d1a),
	.w7(32'hbafd2c7d),
	.w8(32'hba4d508a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393558de),
	.w1(32'hba453c9f),
	.w2(32'hba626980),
	.w3(32'hb983d495),
	.w4(32'hbb04eaa8),
	.w5(32'hbacb8c94),
	.w6(32'h39df7778),
	.w7(32'hba8f270f),
	.w8(32'hba4408fd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9883baf),
	.w1(32'h394476c2),
	.w2(32'hb943b4b6),
	.w3(32'hbb314365),
	.w4(32'hba329744),
	.w5(32'hbac376e2),
	.w6(32'hbaefc71e),
	.w7(32'hba8837c0),
	.w8(32'hbaabf945),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82f321),
	.w1(32'hbb1765c2),
	.w2(32'hbaefe417),
	.w3(32'h39fe4e9b),
	.w4(32'hbb2722ff),
	.w5(32'hba43e530),
	.w6(32'h39f21a72),
	.w7(32'hbad99bd8),
	.w8(32'hbafecf1c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6becaf),
	.w1(32'h38df2f43),
	.w2(32'hb8f7a1b2),
	.w3(32'hbb990b5d),
	.w4(32'h3a8f76bb),
	.w5(32'hb904f667),
	.w6(32'hbb81cf76),
	.w7(32'hba66e2c3),
	.w8(32'hbaaacb6d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3845a),
	.w1(32'hb9875c67),
	.w2(32'h3b0ca3d4),
	.w3(32'hbb4096f0),
	.w4(32'h3a403e53),
	.w5(32'h3b8de5a6),
	.w6(32'hbb54142d),
	.w7(32'h3920e92f),
	.w8(32'h3b5a719c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fd199),
	.w1(32'hbb25d888),
	.w2(32'hbb49fa7f),
	.w3(32'h3a4ec5c3),
	.w4(32'hbb179fc2),
	.w5(32'hbaf6f8e6),
	.w6(32'h39975345),
	.w7(32'hbac7e260),
	.w8(32'hbadd1d6e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0a68a),
	.w1(32'hbadbf253),
	.w2(32'hbad5093e),
	.w3(32'hba199df8),
	.w4(32'hba98aa37),
	.w5(32'hba8936b3),
	.w6(32'hba965769),
	.w7(32'hbad5724f),
	.w8(32'hbb1cfc40),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaba0d2),
	.w1(32'h3aa5754e),
	.w2(32'h3ae082b2),
	.w3(32'hb9595357),
	.w4(32'h3994c7a5),
	.w5(32'hba1f425e),
	.w6(32'hb90111f8),
	.w7(32'h3a0ea69e),
	.w8(32'h3a7af4b1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c2039),
	.w1(32'hba2ec91e),
	.w2(32'h3a27e0bd),
	.w3(32'hba46cd5e),
	.w4(32'hba58d799),
	.w5(32'h3aaf748f),
	.w6(32'hba76c6c2),
	.w7(32'hbaa2a42d),
	.w8(32'h3a695176),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab106a2),
	.w1(32'h3ae72510),
	.w2(32'h3ba3c3cc),
	.w3(32'hbb0e8d3f),
	.w4(32'h3b139fa9),
	.w5(32'h3b863d6b),
	.w6(32'hbabc0624),
	.w7(32'h3a6440d2),
	.w8(32'h3b16b0bf),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1e3c),
	.w1(32'hbbde1b08),
	.w2(32'hbbe3e77a),
	.w3(32'hbbea8b20),
	.w4(32'hbbcbba3f),
	.w5(32'hbb84186e),
	.w6(32'hbbf5b278),
	.w7(32'hbb9a47e6),
	.w8(32'hbb535adf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2e2d5),
	.w1(32'h3b3a5aa1),
	.w2(32'h3b57876e),
	.w3(32'h3b0515af),
	.w4(32'h3b047da9),
	.w5(32'h3acbd715),
	.w6(32'h3b31b028),
	.w7(32'h3b11027c),
	.w8(32'h3ab85094),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e916cb),
	.w1(32'hba854ecb),
	.w2(32'hb9d7f532),
	.w3(32'hba233c6b),
	.w4(32'hbb5bd623),
	.w5(32'hba6d2a85),
	.w6(32'hba120c30),
	.w7(32'hbb382dd9),
	.w8(32'hbb142a89),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd93095),
	.w1(32'hbbef890b),
	.w2(32'hbbba6c44),
	.w3(32'hbc00399e),
	.w4(32'hbbce932e),
	.w5(32'hbba1b871),
	.w6(32'hbbe73eb7),
	.w7(32'hbb480570),
	.w8(32'hbb669544),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994148e),
	.w1(32'h3a32e53c),
	.w2(32'h3a9950ac),
	.w3(32'hbac450a3),
	.w4(32'hba13f3d7),
	.w5(32'h3a45d4af),
	.w6(32'hbae0337b),
	.w7(32'hba2bda91),
	.w8(32'h3a18c367),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab93cd4),
	.w1(32'hbb5355ef),
	.w2(32'hbaa00e0e),
	.w3(32'hba948960),
	.w4(32'hbb3c3492),
	.w5(32'h3a6c3708),
	.w6(32'hb916224f),
	.w7(32'hbacf2b76),
	.w8(32'hba286bb0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb098ebc),
	.w1(32'hba834a73),
	.w2(32'h3a42e085),
	.w3(32'hba04d63f),
	.w4(32'hb8fb64dc),
	.w5(32'h3b15f6a0),
	.w6(32'hba501be3),
	.w7(32'h39e84dc0),
	.w8(32'h39a5067a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8fa9a),
	.w1(32'h3bbf9f4a),
	.w2(32'h3bac8792),
	.w3(32'h3c18a2d6),
	.w4(32'h3b6d7c3f),
	.w5(32'h3b850ef4),
	.w6(32'h3c2751bb),
	.w7(32'h3b6d43a3),
	.w8(32'h3b24aafe),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02eb5e),
	.w1(32'hbb28e2f4),
	.w2(32'hbb59a5b8),
	.w3(32'hbb28263d),
	.w4(32'hbb3b38e6),
	.w5(32'hbaa1d413),
	.w6(32'hbb2359fa),
	.w7(32'hbb28a4a1),
	.w8(32'hbb205994),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72e62f),
	.w1(32'hb98d9107),
	.w2(32'hb96b2c10),
	.w3(32'hbb1d8b4a),
	.w4(32'hba7861e9),
	.w5(32'h3a35a91c),
	.w6(32'hba9d8d51),
	.w7(32'hba0e080b),
	.w8(32'h38821056),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ffcf7),
	.w1(32'hbaadc811),
	.w2(32'hba8124d0),
	.w3(32'h3a25cad1),
	.w4(32'hba40201e),
	.w5(32'hba0256b3),
	.w6(32'h3a07e517),
	.w7(32'h3a1f3800),
	.w8(32'hb8a0293a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52fa37),
	.w1(32'h3b03fcb1),
	.w2(32'h3a944fb8),
	.w3(32'hb99faba8),
	.w4(32'h3ae45658),
	.w5(32'h3a460792),
	.w6(32'hb9a62420),
	.w7(32'h3af1a8d7),
	.w8(32'h3ada2fed),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cb31),
	.w1(32'h3aada472),
	.w2(32'hba68ab8c),
	.w3(32'h3b58b814),
	.w4(32'hb9d7b445),
	.w5(32'h3a3560a7),
	.w6(32'h3b20d422),
	.w7(32'hba94cd3d),
	.w8(32'hba23fa8d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beffb7),
	.w1(32'hba8b3eca),
	.w2(32'h3b22908c),
	.w3(32'h396f53de),
	.w4(32'h3a842cb7),
	.w5(32'h3bc708c0),
	.w6(32'h3a48cf30),
	.w7(32'h3a59ec21),
	.w8(32'h3adf056e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08eb2e),
	.w1(32'hb9a2230c),
	.w2(32'hb8ff8aba),
	.w3(32'h3a48a9bb),
	.w4(32'h399e0732),
	.w5(32'h3a42ed9f),
	.w6(32'h3a5699ae),
	.w7(32'h37968433),
	.w8(32'h3963f0ea),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72244),
	.w1(32'hba34d8f4),
	.w2(32'h3b3d1c11),
	.w3(32'h3a7aad64),
	.w4(32'hba18eea1),
	.w5(32'h3b465e23),
	.w6(32'h3a950b76),
	.w7(32'hba536656),
	.w8(32'h3ad71bd8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac22478),
	.w1(32'h3b8cd68f),
	.w2(32'h3bb22847),
	.w3(32'h3aefddb7),
	.w4(32'h3ae81ec4),
	.w5(32'h3b88afac),
	.w6(32'h3a9aa3d2),
	.w7(32'h3ada9fdb),
	.w8(32'h3b1fb901),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc0d7c),
	.w1(32'hbb85fb56),
	.w2(32'hbbc4817a),
	.w3(32'hbb069a7d),
	.w4(32'hbb94f6ee),
	.w5(32'hbb805549),
	.w6(32'hbb917f13),
	.w7(32'hbb7f1ddf),
	.w8(32'hbb274ea5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bfc52),
	.w1(32'h3999fa78),
	.w2(32'h3a900093),
	.w3(32'h3b17cc4a),
	.w4(32'hba313c55),
	.w5(32'h3b084a79),
	.w6(32'h3b6926a2),
	.w7(32'h3997595c),
	.w8(32'h3a20a0c0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf978b7),
	.w1(32'h3af71d75),
	.w2(32'h3b1ae11e),
	.w3(32'hbb356992),
	.w4(32'h3ae29f19),
	.w5(32'hbaa22a75),
	.w6(32'hba8d1379),
	.w7(32'h39bcdbb8),
	.w8(32'hb9b8eff6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5591ee),
	.w1(32'h3b38f195),
	.w2(32'h3aac39b8),
	.w3(32'h3b4c64a1),
	.w4(32'h3ae63d90),
	.w5(32'h38421991),
	.w6(32'h3a6d9592),
	.w7(32'h38bb3ed1),
	.w8(32'h3a3648c5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae8aae),
	.w1(32'h3a2a47dc),
	.w2(32'h3aa24c2e),
	.w3(32'h3b21d904),
	.w4(32'h3a97538d),
	.w5(32'h3a2a95f0),
	.w6(32'h3af6a89b),
	.w7(32'h3ac3c983),
	.w8(32'h3a992667),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a033138),
	.w1(32'h3ac735c8),
	.w2(32'hb9eea458),
	.w3(32'h3a4ff49f),
	.w4(32'h39d96b12),
	.w5(32'hb8a5a0f7),
	.w6(32'h3aff77a0),
	.w7(32'hb9858db2),
	.w8(32'hbacdbd8d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978fd7c),
	.w1(32'h3a931155),
	.w2(32'hb8dd0bb2),
	.w3(32'h3ab959d8),
	.w4(32'h3a50a45b),
	.w5(32'h3a65b604),
	.w6(32'hb7325b93),
	.w7(32'hb924a352),
	.w8(32'hb7a4c636),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42ff4),
	.w1(32'hbb80f20f),
	.w2(32'hbb168a58),
	.w3(32'hbb2d0cac),
	.w4(32'hbb183a71),
	.w5(32'h3aa2fc3e),
	.w6(32'hbb4babcd),
	.w7(32'hbaf2d7d3),
	.w8(32'hba2c243d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0968b),
	.w1(32'hbabc213a),
	.w2(32'hba5a1a4a),
	.w3(32'h3ae14e32),
	.w4(32'hba79a223),
	.w5(32'hba3c7744),
	.w6(32'h3a0e220a),
	.w7(32'hba46126d),
	.w8(32'hba054870),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd3887),
	.w1(32'hba7c168a),
	.w2(32'h3a77591b),
	.w3(32'hbae88414),
	.w4(32'h38f858a7),
	.w5(32'h3b2ee361),
	.w6(32'hbaab0729),
	.w7(32'h399c8de9),
	.w8(32'h3afda57e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a303e55),
	.w1(32'h3a655b66),
	.w2(32'h3a99e4a7),
	.w3(32'h3a04ce96),
	.w4(32'h3aa10551),
	.w5(32'hb9816d3d),
	.w6(32'h3a290c6f),
	.w7(32'h3ae00ee4),
	.w8(32'h3a936b87),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3abdb),
	.w1(32'hba26c84a),
	.w2(32'h3a8af400),
	.w3(32'h3aeae7e1),
	.w4(32'hb9df1370),
	.w5(32'hb9e4c95b),
	.w6(32'h3b110e89),
	.w7(32'h3a82efff),
	.w8(32'h3aa90e4d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba334fe9),
	.w1(32'hb9c607bb),
	.w2(32'hba4f7089),
	.w3(32'hb966f338),
	.w4(32'hb9b888aa),
	.w5(32'hbaaec73b),
	.w6(32'h3a2cfca8),
	.w7(32'h39e619a7),
	.w8(32'hb9cf3519),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afce6d0),
	.w1(32'h3b84d9f5),
	.w2(32'h3b6537a6),
	.w3(32'h3a76e71c),
	.w4(32'h3af2c27f),
	.w5(32'h3b4a9ac5),
	.w6(32'h3a2215de),
	.w7(32'h3ad968f0),
	.w8(32'h3a99adcb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953c1e3),
	.w1(32'hbb088c3e),
	.w2(32'h39217fb1),
	.w3(32'hb915842c),
	.w4(32'hbb06c5e4),
	.w5(32'h3a12105f),
	.w6(32'h3958fb77),
	.w7(32'hba17fe5c),
	.w8(32'hba2aa671),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aaeac),
	.w1(32'h3a0368c4),
	.w2(32'h3a317ded),
	.w3(32'h3a2c3749),
	.w4(32'hba6a43dd),
	.w5(32'h3b0fd0af),
	.w6(32'hba37d934),
	.w7(32'hb9a23023),
	.w8(32'h39b48792),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42a76),
	.w1(32'h3a396013),
	.w2(32'h3b1045dc),
	.w3(32'h3b716001),
	.w4(32'h3b47f5b9),
	.w5(32'h3aabbfe1),
	.w6(32'h3bc99614),
	.w7(32'h3b4fd5c2),
	.w8(32'h3a9445ea),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706a0a),
	.w1(32'hba565352),
	.w2(32'hbb7b4630),
	.w3(32'hbb95adcb),
	.w4(32'hbb5c24c2),
	.w5(32'hba3bd8f8),
	.w6(32'hbc1fd030),
	.w7(32'hbba49274),
	.w8(32'hba9232d0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b055073),
	.w1(32'h3b06ade1),
	.w2(32'h3a4d4377),
	.w3(32'h3ac0aeeb),
	.w4(32'h3aa2f1e2),
	.w5(32'h3a8d2f1c),
	.w6(32'h3a9a1b2c),
	.w7(32'h393d2d88),
	.w8(32'hb941ba19),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94166be),
	.w1(32'hba029b9d),
	.w2(32'h39f6d192),
	.w3(32'h3b32227a),
	.w4(32'h38ca12c0),
	.w5(32'h3a61abff),
	.w6(32'h3b736b8f),
	.w7(32'h3aabd1cc),
	.w8(32'h3aec1c47),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39c3e4),
	.w1(32'h39a205db),
	.w2(32'h3b0a8f26),
	.w3(32'h3a22bc35),
	.w4(32'h39f3cfca),
	.w5(32'h3b2a444a),
	.w6(32'hb89c5bc4),
	.w7(32'hba555cc6),
	.w8(32'h3a9a574d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b123613),
	.w1(32'h3adae626),
	.w2(32'h3ad1000b),
	.w3(32'h3b7bcd65),
	.w4(32'h3af05b7a),
	.w5(32'h3ad63f33),
	.w6(32'h3b1f383f),
	.w7(32'h3a9098ce),
	.w8(32'h3ad71282),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031104),
	.w1(32'hbb2e12f9),
	.w2(32'hbb0f899a),
	.w3(32'hbac11632),
	.w4(32'hbb5c6d5a),
	.w5(32'hba206cb2),
	.w6(32'hba8ccd38),
	.w7(32'hbb1f5954),
	.w8(32'hbac54e88),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd95807),
	.w1(32'hbae09e70),
	.w2(32'hb90c2bbe),
	.w3(32'hbbbdb5df),
	.w4(32'hbb27289a),
	.w5(32'h3b077246),
	.w6(32'hbbf6c445),
	.w7(32'hbb4166b0),
	.w8(32'h3939ea36),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2311fc),
	.w1(32'h39ad1f6e),
	.w2(32'h3a5dcfa4),
	.w3(32'h3a6aecdb),
	.w4(32'hb8e63e39),
	.w5(32'h3a7e7795),
	.w6(32'h3af23d73),
	.w7(32'h3a48ac42),
	.w8(32'h3a8ff356),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac718e8),
	.w1(32'hba8814c5),
	.w2(32'h3ad116a1),
	.w3(32'hbacca6e0),
	.w4(32'hb91020e7),
	.w5(32'h3b042df8),
	.w6(32'hbaa0771f),
	.w7(32'hbad7084c),
	.w8(32'h3ac198e4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d0244),
	.w1(32'h3a12d861),
	.w2(32'h3a2613c2),
	.w3(32'h3a92344f),
	.w4(32'h3a0adc6c),
	.w5(32'hb9aaab6b),
	.w6(32'h3ae58763),
	.w7(32'h394e25be),
	.w8(32'h3a6267e3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad60eaa),
	.w1(32'h3b1e5b5e),
	.w2(32'h3a4f0b0f),
	.w3(32'h3afbe7be),
	.w4(32'h3af025ad),
	.w5(32'h3a46b626),
	.w6(32'h3b13572d),
	.w7(32'h3aa07c72),
	.w8(32'h3a26222f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e9f60),
	.w1(32'hb938bec4),
	.w2(32'hb72c2078),
	.w3(32'hba290bc5),
	.w4(32'hba8a3e83),
	.w5(32'hb98fdcde),
	.w6(32'h38f194e3),
	.w7(32'h38c52c12),
	.w8(32'h3a2a07a7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa092f),
	.w1(32'h3b06b63e),
	.w2(32'h3ae82a18),
	.w3(32'h3a8c57a1),
	.w4(32'h3b26db1f),
	.w5(32'h3b0e3383),
	.w6(32'h3a1bd6fa),
	.w7(32'h3a9a268a),
	.w8(32'h3af3e883),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a455768),
	.w1(32'hba07958b),
	.w2(32'hba217410),
	.w3(32'h3aa6695f),
	.w4(32'h39fb39b1),
	.w5(32'hba85a63e),
	.w6(32'h3ac92c9f),
	.w7(32'h3a98049d),
	.w8(32'hb90c24a6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fed86),
	.w1(32'hbb0550ae),
	.w2(32'hba5135a1),
	.w3(32'hb91b610f),
	.w4(32'h3996e86b),
	.w5(32'h3a33dc3e),
	.w6(32'hb8cd2784),
	.w7(32'h3a904f8d),
	.w8(32'hb8960d56),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5cf53),
	.w1(32'hbac036e6),
	.w2(32'hb89e679b),
	.w3(32'h39e6b355),
	.w4(32'h3a014ad9),
	.w5(32'h3aa09a3a),
	.w6(32'hbab6b221),
	.w7(32'h3a47a442),
	.w8(32'h37030d7b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8455fd),
	.w1(32'h39da15cd),
	.w2(32'h3a6a425f),
	.w3(32'h3b0c5743),
	.w4(32'h39c9d081),
	.w5(32'h39e6d178),
	.w6(32'hb9a0f47c),
	.w7(32'hbadcf693),
	.w8(32'hbad2085c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7f425),
	.w1(32'h39a93981),
	.w2(32'h3a940ca7),
	.w3(32'hbb2bdb75),
	.w4(32'h3a17171f),
	.w5(32'h3b4bce2b),
	.w6(32'hbb1928ac),
	.w7(32'h3a11123d),
	.w8(32'h3ace6ae6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4acc9a),
	.w1(32'hba5873c7),
	.w2(32'hbb14c974),
	.w3(32'hb8e33080),
	.w4(32'h3882994e),
	.w5(32'hbb2a5969),
	.w6(32'h3a2a17e6),
	.w7(32'hb916516e),
	.w8(32'hbaf85f52),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf7e3c),
	.w1(32'hbbc3c773),
	.w2(32'hbac4a2c0),
	.w3(32'hbbeaedb2),
	.w4(32'hbbd4a06f),
	.w5(32'h3b056e51),
	.w6(32'hbbdf94b1),
	.w7(32'hbb197380),
	.w8(32'hbb213837),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b9d04),
	.w1(32'h3c08c377),
	.w2(32'h3c010336),
	.w3(32'h3bd1a6c5),
	.w4(32'h3bed5563),
	.w5(32'h3bb319ab),
	.w6(32'h3be53d97),
	.w7(32'h3b8d4e2c),
	.w8(32'h3af757bf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83f968),
	.w1(32'hb9f85518),
	.w2(32'hb946efe5),
	.w3(32'h3b44eb56),
	.w4(32'hba87d8eb),
	.w5(32'h39bb2f60),
	.w6(32'h3a6f0b1c),
	.w7(32'hba9db1ae),
	.w8(32'hbadeb55a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba169d81),
	.w1(32'h39a724f4),
	.w2(32'hbabf476d),
	.w3(32'hb9c3961c),
	.w4(32'hb9d172db),
	.w5(32'hba962fdc),
	.w6(32'h38d6c5c0),
	.w7(32'h3908788e),
	.w8(32'h39bc7122),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a92bf5),
	.w1(32'h39841bd9),
	.w2(32'hb9b7acc9),
	.w3(32'hb9f6f988),
	.w4(32'h3a135273),
	.w5(32'h3992375d),
	.w6(32'hba03aba7),
	.w7(32'hb988eb52),
	.w8(32'hb9e7b30a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38576a60),
	.w1(32'h3b1a1cfb),
	.w2(32'h3b092393),
	.w3(32'h3a33c735),
	.w4(32'h3af7a02d),
	.w5(32'h39ea32ee),
	.w6(32'h3a60aa41),
	.w7(32'h3b14cc51),
	.w8(32'h3ad58288),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075a71),
	.w1(32'h3ab5842f),
	.w2(32'h3aae40d9),
	.w3(32'h3a83fe6a),
	.w4(32'h390e8d25),
	.w5(32'h3ab9ed87),
	.w6(32'h3ad0f8be),
	.w7(32'hb943dac1),
	.w8(32'h3a8473b0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c62e99),
	.w1(32'hbb34ee3e),
	.w2(32'hbb3f85cb),
	.w3(32'hb9a144ce),
	.w4(32'hba5a7421),
	.w5(32'hbb143134),
	.w6(32'h3a89878f),
	.w7(32'hba34d200),
	.w8(32'hbb1f7d4a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a967890),
	.w1(32'h3b9d1bc6),
	.w2(32'h3bd82d14),
	.w3(32'h3b2bcad0),
	.w4(32'h3b85b150),
	.w5(32'h3bed7309),
	.w6(32'h3b81628a),
	.w7(32'h3b934c8d),
	.w8(32'h3bc24322),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995f1cc),
	.w1(32'hbaa0103a),
	.w2(32'hbaa67b7f),
	.w3(32'hb861c07c),
	.w4(32'hbab755af),
	.w5(32'h39dbaa7b),
	.w6(32'h38b06c06),
	.w7(32'hba915d26),
	.w8(32'hbaba0689),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277f92),
	.w1(32'h38d438f3),
	.w2(32'h3ba4ae36),
	.w3(32'hbacabcb2),
	.w4(32'hba825f6b),
	.w5(32'hb9f2f64f),
	.w6(32'hbac23873),
	.w7(32'hbae30d0e),
	.w8(32'h3aa3973d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e2bb4),
	.w1(32'h3a0d7c85),
	.w2(32'h39ffee7a),
	.w3(32'hbb946730),
	.w4(32'h3aa11e1b),
	.w5(32'h3afe5fb8),
	.w6(32'hbba7af0f),
	.w7(32'h3ae4d8e7),
	.w8(32'h39a80d2a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36421e),
	.w1(32'hbb851d9b),
	.w2(32'hbaff5639),
	.w3(32'hbb9cb340),
	.w4(32'hbb1677c9),
	.w5(32'h3b708d3b),
	.w6(32'hbb9be486),
	.w7(32'hbbba4211),
	.w8(32'h3babdad3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68fb11),
	.w1(32'hbb794ce2),
	.w2(32'hbb4124a7),
	.w3(32'hba952c55),
	.w4(32'hbbb428cd),
	.w5(32'hbb1622fc),
	.w6(32'hb914f5b7),
	.w7(32'hbbdb39ee),
	.w8(32'hba2fa746),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36920c),
	.w1(32'hba7de37c),
	.w2(32'hbb4b78c4),
	.w3(32'hbad6d732),
	.w4(32'hba92ce18),
	.w5(32'hbb183db4),
	.w6(32'hbac90eba),
	.w7(32'hbb1efa92),
	.w8(32'hbad3cead),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c194b),
	.w1(32'hbb106422),
	.w2(32'h3b4a7be6),
	.w3(32'hbbb86ad0),
	.w4(32'h3bbb00e4),
	.w5(32'hb902d690),
	.w6(32'hbb2b940d),
	.w7(32'h3baa33ad),
	.w8(32'hbab0f992),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a965a),
	.w1(32'h3a740019),
	.w2(32'h3a6d37cf),
	.w3(32'hbaa42fff),
	.w4(32'h3a8be0bc),
	.w5(32'h3b3d4458),
	.w6(32'h3997e5eb),
	.w7(32'hb9b071e0),
	.w8(32'hba045650),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98b11e),
	.w1(32'hba93b4ae),
	.w2(32'hbb9efb3a),
	.w3(32'h3b0feb97),
	.w4(32'hb90d4295),
	.w5(32'hbaf57436),
	.w6(32'h3b83f286),
	.w7(32'hbb07e5b1),
	.w8(32'hbb6892ab),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbccbf),
	.w1(32'h3b932a95),
	.w2(32'hbb4b93c1),
	.w3(32'hbbc09290),
	.w4(32'h3b48e186),
	.w5(32'h3ab3d88c),
	.w6(32'hbbf352fb),
	.w7(32'h3b345fe3),
	.w8(32'hbbeac087),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88df79),
	.w1(32'h39bfcd8e),
	.w2(32'h3b6154ed),
	.w3(32'hbb00f504),
	.w4(32'hb9996d3a),
	.w5(32'h3c0628d7),
	.w6(32'h3b0f159a),
	.w7(32'h3b2e4682),
	.w8(32'hba852a16),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb952351),
	.w1(32'h3b3acd84),
	.w2(32'hbad44f98),
	.w3(32'hba81208e),
	.w4(32'hb979453a),
	.w5(32'hbab14dff),
	.w6(32'hba0243bc),
	.w7(32'hb94dbbac),
	.w8(32'hbb05adaa),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03cf47),
	.w1(32'h3b1f19da),
	.w2(32'h3c1d5d01),
	.w3(32'hb9e850f2),
	.w4(32'h3999829e),
	.w5(32'h3bdaf410),
	.w6(32'hbacfcaa8),
	.w7(32'hbab1396e),
	.w8(32'h3bc65368),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b858bc6),
	.w1(32'h3ae4afdb),
	.w2(32'hbac7c43f),
	.w3(32'h3be750ab),
	.w4(32'h3b8b86b6),
	.w5(32'h3b3515cf),
	.w6(32'h3bcc7a9b),
	.w7(32'h3b00c08b),
	.w8(32'hba02df55),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9ff4),
	.w1(32'h3a27213a),
	.w2(32'h3b40e7c3),
	.w3(32'hbb7e972e),
	.w4(32'hbb58016f),
	.w5(32'h3bc3e22e),
	.w6(32'hbb3ce018),
	.w7(32'h3a0ab55f),
	.w8(32'h3be1654d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78d8b3),
	.w1(32'hbb05ac44),
	.w2(32'h3b801bd2),
	.w3(32'h3b9191d8),
	.w4(32'hbbd0023a),
	.w5(32'h3c6ecb05),
	.w6(32'h3b270478),
	.w7(32'hbad26d3e),
	.w8(32'h3c14db76),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf54351),
	.w1(32'hbbc6fe9d),
	.w2(32'hbb8b4a7f),
	.w3(32'hbc13eab4),
	.w4(32'hbbd1dcea),
	.w5(32'h3b41c76c),
	.w6(32'hbc6c8cf4),
	.w7(32'hbc3c891a),
	.w8(32'hbb17567a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86c580),
	.w1(32'hb90762c8),
	.w2(32'h3b64debf),
	.w3(32'hbae7993c),
	.w4(32'h3b2c92e8),
	.w5(32'h3b76de57),
	.w6(32'h3a3bcbd9),
	.w7(32'h3c076292),
	.w8(32'h3af7b49a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15e73e),
	.w1(32'h3ad4aa7b),
	.w2(32'hb93df7d0),
	.w3(32'h3ae0122c),
	.w4(32'hbb7a13dd),
	.w5(32'h3bbbecf3),
	.w6(32'h3aa8cea1),
	.w7(32'h3ac22cb4),
	.w8(32'hbb2a546e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2421b4),
	.w1(32'h3b1db3aa),
	.w2(32'hb8a63c13),
	.w3(32'h3a7eabc2),
	.w4(32'hb9b1eed3),
	.w5(32'h3b53d4d0),
	.w6(32'h3b08cc55),
	.w7(32'h3875549f),
	.w8(32'h3b3fdf53),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e7567),
	.w1(32'hbb2c818a),
	.w2(32'hbb0f46c6),
	.w3(32'hbad7fc16),
	.w4(32'h3a8a4294),
	.w5(32'h3a8673c6),
	.w6(32'hb9022c6f),
	.w7(32'hbaa60f17),
	.w8(32'h39ae6bd4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4604f6),
	.w1(32'hbb2a3b0c),
	.w2(32'hbb014d7f),
	.w3(32'hbc1325a8),
	.w4(32'h39871786),
	.w5(32'h3bdf8335),
	.w6(32'hbc33f2e3),
	.w7(32'h3a03c6b8),
	.w8(32'h3a327929),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2df4),
	.w1(32'hbc0855f6),
	.w2(32'hbb4d5ec0),
	.w3(32'hbc0a948c),
	.w4(32'hbb931fe9),
	.w5(32'h3b8014d4),
	.w6(32'hbc043067),
	.w7(32'hbbbd5c35),
	.w8(32'h3ae516fe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ec4f),
	.w1(32'hbc14bf10),
	.w2(32'hbbcf2be0),
	.w3(32'hbbb5ae93),
	.w4(32'hbbc3d84e),
	.w5(32'hbbc4f3f3),
	.w6(32'hbc096557),
	.w7(32'hbb5f8623),
	.w8(32'hbb319d08),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d8afb),
	.w1(32'hbb3d495a),
	.w2(32'h3bb3618d),
	.w3(32'hbbd51308),
	.w4(32'hbbc0b59d),
	.w5(32'h3b338d8c),
	.w6(32'hbadd1901),
	.w7(32'hbbc98d1e),
	.w8(32'h3bd6cb2d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5e70),
	.w1(32'hba743778),
	.w2(32'h3baca25c),
	.w3(32'h3b816278),
	.w4(32'hba9995a3),
	.w5(32'h3bb35107),
	.w6(32'h3b98487a),
	.w7(32'hbb011ebb),
	.w8(32'h3b9620fb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb47d8f),
	.w1(32'hba5a40a3),
	.w2(32'hba65b1c4),
	.w3(32'h3b94f8a8),
	.w4(32'hbac40304),
	.w5(32'h39e853a5),
	.w6(32'h3bb517b7),
	.w7(32'hbb05573d),
	.w8(32'h3aa8f987),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dacc3),
	.w1(32'hba1d182e),
	.w2(32'h39e59898),
	.w3(32'hbae1483b),
	.w4(32'hba9c1e18),
	.w5(32'h39f9d51a),
	.w6(32'hbb2fd8d4),
	.w7(32'hbb12d3b6),
	.w8(32'h3acebdb4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac957),
	.w1(32'h3a49204d),
	.w2(32'hbb8380f4),
	.w3(32'hbb8a645d),
	.w4(32'h3acbd2b8),
	.w5(32'hba8f2a87),
	.w6(32'hba4e6837),
	.w7(32'h3a352d76),
	.w8(32'hbabd9af9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04d083),
	.w1(32'h3c4121b4),
	.w2(32'h3b9f2f33),
	.w3(32'hbb6c7699),
	.w4(32'h3c8f1e3a),
	.w5(32'h3c39cbda),
	.w6(32'hba3c8414),
	.w7(32'h3c6b807c),
	.w8(32'h3bc0032a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1bbc),
	.w1(32'hbb043ad9),
	.w2(32'hbc03cec4),
	.w3(32'h3ae8adf0),
	.w4(32'h3b97eb67),
	.w5(32'hba9ed490),
	.w6(32'h3a1e1231),
	.w7(32'h3ab8762a),
	.w8(32'hbbd72089),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa421f),
	.w1(32'hba1f6e6e),
	.w2(32'hbab2eb9c),
	.w3(32'hbb489a38),
	.w4(32'h3bacbc2f),
	.w5(32'h3a8fe1e1),
	.w6(32'hbbb19af1),
	.w7(32'hbb630843),
	.w8(32'h3acaeab2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d198f),
	.w1(32'hb852d492),
	.w2(32'hbb2de856),
	.w3(32'hbb553b19),
	.w4(32'hb9816fb3),
	.w5(32'h3ace0635),
	.w6(32'h35b022f5),
	.w7(32'hba97eb81),
	.w8(32'hba3bbcd3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cf638),
	.w1(32'h3abfbe8e),
	.w2(32'h3b1e3da5),
	.w3(32'hbb54400e),
	.w4(32'hbb855d3d),
	.w5(32'h3b2d1075),
	.w6(32'hbb352e55),
	.w7(32'hbab40766),
	.w8(32'h3ac79429),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aab392),
	.w1(32'hbc204b55),
	.w2(32'hbc1a8438),
	.w3(32'hbbe6a61b),
	.w4(32'hbc2602e4),
	.w5(32'hbb3fe5c5),
	.w6(32'hbc05b4ef),
	.w7(32'hbc352354),
	.w8(32'hbb38785c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb2ba8),
	.w1(32'hbb4c31eb),
	.w2(32'h3b8486c1),
	.w3(32'hbb91fc83),
	.w4(32'hbbbecb9f),
	.w5(32'h3ba26b60),
	.w6(32'hbbfa280d),
	.w7(32'hbb115ce1),
	.w8(32'hba6b3d39),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d00c),
	.w1(32'hbb0f7c8c),
	.w2(32'h3a8b83d9),
	.w3(32'hbaa7f5b9),
	.w4(32'hbbab3456),
	.w5(32'h3b8ca7dc),
	.w6(32'hbade28be),
	.w7(32'hb996ca9c),
	.w8(32'h3adc2ecd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7b657),
	.w1(32'hbb8e1ed2),
	.w2(32'hbb53df3b),
	.w3(32'hbc347eac),
	.w4(32'hbb2ebafa),
	.w5(32'h398ef0c3),
	.w6(32'hbc303173),
	.w7(32'hba561f28),
	.w8(32'hbb03ea50),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2659a),
	.w1(32'h3b7d5f14),
	.w2(32'h3ac12a23),
	.w3(32'hb9bf199a),
	.w4(32'h3bbc5b19),
	.w5(32'h3ba43c30),
	.w6(32'h3a24b80b),
	.w7(32'h3b21501f),
	.w8(32'hbaea90b9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b65f0),
	.w1(32'hb895b40c),
	.w2(32'h3b57d689),
	.w3(32'hbbd3373f),
	.w4(32'h3962e877),
	.w5(32'h3b1ae2e5),
	.w6(32'hbb6f1917),
	.w7(32'hbb081d6b),
	.w8(32'h3b9eaa2e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92cb00),
	.w1(32'hba7a834c),
	.w2(32'h3b65059b),
	.w3(32'hbb13cd36),
	.w4(32'hbb7162a9),
	.w5(32'h3b74e9bf),
	.w6(32'hba6999c7),
	.w7(32'h3aeafc0e),
	.w8(32'h3ba93ee7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1801c2),
	.w1(32'hbb26d85f),
	.w2(32'hba49b9d6),
	.w3(32'h3907936c),
	.w4(32'hbb063706),
	.w5(32'hba79821d),
	.w6(32'hbb0a3afc),
	.w7(32'h3b126120),
	.w8(32'h3ad0b671),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba54d7d),
	.w1(32'hbb6aa709),
	.w2(32'h3ab05805),
	.w3(32'hbc08c63e),
	.w4(32'h3a1bab43),
	.w5(32'h3b8ddcfb),
	.w6(32'hbb8638da),
	.w7(32'hbaee7641),
	.w8(32'hbb15de2a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e63a),
	.w1(32'hbb6c9eef),
	.w2(32'h39a81fb4),
	.w3(32'hbaf988ff),
	.w4(32'hbb6d773b),
	.w5(32'h39a7b215),
	.w6(32'hba83e896),
	.w7(32'hbac4def0),
	.w8(32'hbaf596df),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2a003),
	.w1(32'hbb98a972),
	.w2(32'hba8f535f),
	.w3(32'hb9f55113),
	.w4(32'hbbda19dd),
	.w5(32'h3af91dd3),
	.w6(32'hbb25b4ab),
	.w7(32'hbb651aa5),
	.w8(32'h389d7369),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1587c),
	.w1(32'hbb715467),
	.w2(32'hbb9e6a4a),
	.w3(32'hbb8c0698),
	.w4(32'hb99cb10c),
	.w5(32'hba0290af),
	.w6(32'hbb5b5456),
	.w7(32'hba9266fc),
	.w8(32'h3a51ecef),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5083ee),
	.w1(32'hbb194dac),
	.w2(32'h3b623003),
	.w3(32'hbb60c91c),
	.w4(32'hbb968cea),
	.w5(32'h3b676d9d),
	.w6(32'hbbde1bcd),
	.w7(32'hbb1a0419),
	.w8(32'h3ba6ea10),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e4ae9),
	.w1(32'hbb739e78),
	.w2(32'hbb1cefab),
	.w3(32'h3ba4ace4),
	.w4(32'hbb6dc2b6),
	.w5(32'hb93e8e94),
	.w6(32'h3baf3267),
	.w7(32'hbb761fc7),
	.w8(32'hba2c6ff8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022cfa),
	.w1(32'hbb19aa65),
	.w2(32'h3b2f2581),
	.w3(32'hbb0189b7),
	.w4(32'h3a0cb8b0),
	.w5(32'h3bcfb046),
	.w6(32'hbb138944),
	.w7(32'hbb3202f9),
	.w8(32'h3bcdf260),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f7029),
	.w1(32'h3a9c0b8e),
	.w2(32'hbb78165c),
	.w3(32'h3b24b0f4),
	.w4(32'h3aba72e1),
	.w5(32'hbad7aeb1),
	.w6(32'h3b4e729f),
	.w7(32'h390e1ea6),
	.w8(32'hbac8a494),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba171f59),
	.w1(32'hb987ff29),
	.w2(32'h3ad6614c),
	.w3(32'hba154894),
	.w4(32'hba4dbf0b),
	.w5(32'h38d63ed8),
	.w6(32'hbb993a25),
	.w7(32'hba98ab5b),
	.w8(32'h39aea74f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf5e8d),
	.w1(32'h3b531894),
	.w2(32'h3bd873e4),
	.w3(32'hbbbf238c),
	.w4(32'hbb8adf42),
	.w5(32'h3c17a4c1),
	.w6(32'hbb8a352e),
	.w7(32'hbb66095f),
	.w8(32'h3bb48cdb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da6f5),
	.w1(32'hbb05af08),
	.w2(32'hbaac7669),
	.w3(32'h3b43608f),
	.w4(32'h38844c1f),
	.w5(32'h3b3792c5),
	.w6(32'h3bc74907),
	.w7(32'hbb1edcf8),
	.w8(32'hbacd1da4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ef5cb),
	.w1(32'hbb09f7cd),
	.w2(32'h3b16c5f2),
	.w3(32'hbb53bc0f),
	.w4(32'hbab317be),
	.w5(32'hbb7e73e7),
	.w6(32'hbbc91ac5),
	.w7(32'hbad343e0),
	.w8(32'h3a976036),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e2136),
	.w1(32'h3aa5385d),
	.w2(32'hbb560206),
	.w3(32'hbb11aeac),
	.w4(32'hba82aa34),
	.w5(32'hba661bd1),
	.w6(32'h38bc4836),
	.w7(32'h3accdf77),
	.w8(32'hbacd9556),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07fe81),
	.w1(32'h3aeeb802),
	.w2(32'hba6ec35b),
	.w3(32'hbb5971a0),
	.w4(32'hbb471ac7),
	.w5(32'hbaecb28d),
	.w6(32'hbaaa207b),
	.w7(32'hba58c44c),
	.w8(32'hba83e592),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d8e3b),
	.w1(32'h3a14d216),
	.w2(32'h3a076757),
	.w3(32'hbb078015),
	.w4(32'hb9de989d),
	.w5(32'h3a65b0f4),
	.w6(32'h3b02cd2a),
	.w7(32'hbb238485),
	.w8(32'h3ae48d6a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc008e1a),
	.w1(32'hbb95b29f),
	.w2(32'hbbbba0fc),
	.w3(32'hbbee8c34),
	.w4(32'hba2ae7d9),
	.w5(32'h3b2d56e6),
	.w6(32'hbbe17b51),
	.w7(32'hbaa1b117),
	.w8(32'h39a9d6f8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefd771),
	.w1(32'h3bbb063d),
	.w2(32'hbb90cade),
	.w3(32'hbbd0625b),
	.w4(32'h3b967d1c),
	.w5(32'hbc04fb4a),
	.w6(32'hbb6faa5c),
	.w7(32'h3bb41e43),
	.w8(32'hbbe097ba),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32fc20),
	.w1(32'hbbe8f4c3),
	.w2(32'hbb954798),
	.w3(32'hbbfce896),
	.w4(32'hbb3fe11e),
	.w5(32'hbb11f494),
	.w6(32'hbc2ab160),
	.w7(32'hbabfaf84),
	.w8(32'hbb8707aa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule