module layer_10_featuremap_344(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300b86),
	.w1(32'h3adc7a9f),
	.w2(32'h3ac043e6),
	.w3(32'hbb0a53d1),
	.w4(32'h3aa4d5cf),
	.w5(32'hbb8afea4),
	.w6(32'hb9bd2235),
	.w7(32'h3b0d510c),
	.w8(32'hbb3a4eb3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1eca),
	.w1(32'hbac32ffe),
	.w2(32'h3a62e972),
	.w3(32'hbb8c0f25),
	.w4(32'hba95a20f),
	.w5(32'hbb19c9d2),
	.w6(32'hbb8b0a2c),
	.w7(32'hbad1c515),
	.w8(32'hbac1ec50),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61241c),
	.w1(32'hbb8f2d17),
	.w2(32'h39950ee9),
	.w3(32'h3ac4abc5),
	.w4(32'hb8e6ab6c),
	.w5(32'hbb10a1ce),
	.w6(32'hbb1406da),
	.w7(32'hbab71a48),
	.w8(32'hbac3dd7c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e9369c),
	.w1(32'h3a740147),
	.w2(32'h3aefedfe),
	.w3(32'hb8f01017),
	.w4(32'h3b26caeb),
	.w5(32'hba759a8f),
	.w6(32'h3a310458),
	.w7(32'h3ac10079),
	.w8(32'hbb083a73),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9630e6e),
	.w1(32'hbb59c207),
	.w2(32'hbb413b38),
	.w3(32'hbb6f4eaa),
	.w4(32'hba975ebb),
	.w5(32'hbb5ce02d),
	.w6(32'hbb9f6b36),
	.w7(32'hbab72889),
	.w8(32'hbba9d1a1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96fa45),
	.w1(32'hbb002230),
	.w2(32'h38f86dbd),
	.w3(32'hbb30793b),
	.w4(32'hba3a3098),
	.w5(32'hba9960c0),
	.w6(32'hbb52a2d9),
	.w7(32'hb910acaa),
	.w8(32'hbaef02db),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d01f4),
	.w1(32'h3a17766e),
	.w2(32'h3b8e3a17),
	.w3(32'h3a680c8a),
	.w4(32'h3ad28b55),
	.w5(32'h3b9fadbb),
	.w6(32'hba267368),
	.w7(32'h3ae3b34b),
	.w8(32'h3c064356),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c46c5),
	.w1(32'h3b5b2d0b),
	.w2(32'h3a83f5ad),
	.w3(32'h3c2cb7f9),
	.w4(32'h3c32fb92),
	.w5(32'h3ab759a3),
	.w6(32'h3c37e3ed),
	.w7(32'h3bd67cb2),
	.w8(32'h3a8aa11c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3edde),
	.w1(32'h3935cfc8),
	.w2(32'hb815d1d6),
	.w3(32'hb91b7dfb),
	.w4(32'h3ad5f057),
	.w5(32'hbbd13b56),
	.w6(32'hba9e6d3e),
	.w7(32'h3b185e31),
	.w8(32'hbbe6b1d8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0feaa9),
	.w1(32'hbb955736),
	.w2(32'hba201ba1),
	.w3(32'hbbff1e37),
	.w4(32'hbb6f9b2b),
	.w5(32'hbaa4a758),
	.w6(32'hbc0c5596),
	.w7(32'hbb9986ca),
	.w8(32'hbb6287d4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb564348),
	.w1(32'hbb0b7139),
	.w2(32'hb8039eab),
	.w3(32'hbb57bc31),
	.w4(32'hb9cb09d6),
	.w5(32'h3b9697fa),
	.w6(32'hbb7f381e),
	.w7(32'hba45d942),
	.w8(32'h3bb967c6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b761403),
	.w1(32'h3ab69c51),
	.w2(32'h3af4b96d),
	.w3(32'h3bde0756),
	.w4(32'h3b32e9ae),
	.w5(32'hbaa0c881),
	.w6(32'h3baa2592),
	.w7(32'h3aed8986),
	.w8(32'h3b044a50),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff7ca5),
	.w1(32'hbab4e4f0),
	.w2(32'hbb74579b),
	.w3(32'hbb3755e6),
	.w4(32'hbb6cd2aa),
	.w5(32'h3b9751b6),
	.w6(32'h39fab5ca),
	.w7(32'hbb2a82da),
	.w8(32'h3b52b70f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c44c7),
	.w1(32'hba5752d6),
	.w2(32'hbafa78ef),
	.w3(32'hbb0cae8b),
	.w4(32'hbb9748f4),
	.w5(32'h3b426807),
	.w6(32'hbb1e6ac2),
	.w7(32'hbb871c19),
	.w8(32'h3b06021c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63d59e),
	.w1(32'h3ab23edd),
	.w2(32'h3a91f752),
	.w3(32'hbb063ce8),
	.w4(32'h38dfc485),
	.w5(32'hb9de2c34),
	.w6(32'hba95ecc3),
	.w7(32'h3ab268d7),
	.w8(32'hba6e0c8c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7792e5),
	.w1(32'hba47e42a),
	.w2(32'hbaba162a),
	.w3(32'hbb86c44f),
	.w4(32'hbae69052),
	.w5(32'hbb03d6c6),
	.w6(32'hbb994f4e),
	.w7(32'hba42509e),
	.w8(32'hbb000a69),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfd10d),
	.w1(32'h3ac36d39),
	.w2(32'h3b86ecda),
	.w3(32'hbaa91d19),
	.w4(32'hba7ed209),
	.w5(32'h39b0033e),
	.w6(32'hba967ada),
	.w7(32'h3ac71e95),
	.w8(32'h3a4b92ec),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc5dcb),
	.w1(32'h3965a1eb),
	.w2(32'h3a76666c),
	.w3(32'hbac72d75),
	.w4(32'hb98476d9),
	.w5(32'h399e87aa),
	.w6(32'hba9c84e2),
	.w7(32'h39870a66),
	.w8(32'hbb05a648),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5cf1b),
	.w1(32'hb92d4b5a),
	.w2(32'hba2fc70d),
	.w3(32'hbb8c9e65),
	.w4(32'hbab55457),
	.w5(32'hbb94e640),
	.w6(32'hbb11cedd),
	.w7(32'hba2fbe61),
	.w8(32'hbb917a5b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f3df),
	.w1(32'hba82eca4),
	.w2(32'h3a12d075),
	.w3(32'hbb08beec),
	.w4(32'hb7b82815),
	.w5(32'hbafb22f3),
	.w6(32'hbb3f12e0),
	.w7(32'hb90e00ed),
	.w8(32'hbb0bf54c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eea9d),
	.w1(32'h3aa81491),
	.w2(32'h3afdb319),
	.w3(32'hbb25183e),
	.w4(32'hbae2190a),
	.w5(32'h3b1c8ca4),
	.w6(32'hbb053325),
	.w7(32'hb795e52b),
	.w8(32'h3b20a5bc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4a6e9),
	.w1(32'h3b06ce0a),
	.w2(32'h3b5ce31e),
	.w3(32'h3b972e6a),
	.w4(32'h3b59b983),
	.w5(32'hba633d97),
	.w6(32'h3b9a3b58),
	.w7(32'h3b28b415),
	.w8(32'hba847a21),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c6c1d),
	.w1(32'hbb5d4925),
	.w2(32'hbbd217ab),
	.w3(32'hbb479254),
	.w4(32'hbb4dc5b9),
	.w5(32'hbb4d0a39),
	.w6(32'hbb44d788),
	.w7(32'hbb801786),
	.w8(32'hbab9541b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefdecf),
	.w1(32'h3ab7ea59),
	.w2(32'hbb9ceb25),
	.w3(32'hbb896373),
	.w4(32'h3af3f8e9),
	.w5(32'hbb69e4fc),
	.w6(32'h3aec128b),
	.w7(32'h3aa53e8b),
	.w8(32'hbb4b6081),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d182f),
	.w1(32'hb9acd3a4),
	.w2(32'hbb97bebf),
	.w3(32'h3ae86a6e),
	.w4(32'h391d9ff4),
	.w5(32'hb90f7b0c),
	.w6(32'h3ac5cf6e),
	.w7(32'hb9e75df2),
	.w8(32'hbb068aa5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73975e),
	.w1(32'h3b20db36),
	.w2(32'h3bda16db),
	.w3(32'h39473086),
	.w4(32'h3b154443),
	.w5(32'h3b093872),
	.w6(32'h3aa4a9e6),
	.w7(32'h3b7a8b3c),
	.w8(32'h3a8d6af4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914d6e8),
	.w1(32'hba1a2384),
	.w2(32'h3a1dc215),
	.w3(32'h3b40c62e),
	.w4(32'h3ac27951),
	.w5(32'hbb8eef33),
	.w6(32'h3ac9124e),
	.w7(32'h394dc869),
	.w8(32'hbbc8aee2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706f6d),
	.w1(32'hbae2ba54),
	.w2(32'h3a1367d8),
	.w3(32'hbad35c2b),
	.w4(32'hbacc80c7),
	.w5(32'h3b2965fe),
	.w6(32'hbb0ecf33),
	.w7(32'hba17cfec),
	.w8(32'h3b1505c2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cb946),
	.w1(32'h3836490d),
	.w2(32'h39d8da75),
	.w3(32'h3b5e2fa0),
	.w4(32'hbb0095fd),
	.w5(32'h3a9c50c7),
	.w6(32'h3b672325),
	.w7(32'h3b2ac817),
	.w8(32'h3b75c5ca),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcee2f0),
	.w1(32'hbb05b611),
	.w2(32'h3b479ac9),
	.w3(32'hbbb031b2),
	.w4(32'hba840fa4),
	.w5(32'hb94c5263),
	.w6(32'hbb9953f2),
	.w7(32'h39fb1735),
	.w8(32'hbaaab1a3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84674c),
	.w1(32'hbb419afb),
	.w2(32'hbbc2b28d),
	.w3(32'h3ad7aee5),
	.w4(32'h3b73bc77),
	.w5(32'hbb327580),
	.w6(32'hba0ed185),
	.w7(32'hbac861ef),
	.w8(32'hbb59babe),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7f740),
	.w1(32'hbb69e00f),
	.w2(32'hba7e926d),
	.w3(32'hbad79285),
	.w4(32'hbb011a17),
	.w5(32'h3b4d9536),
	.w6(32'hbb5ad634),
	.w7(32'hb943d7ac),
	.w8(32'h3aea800f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b9562),
	.w1(32'h3b41acbf),
	.w2(32'h3b21c1bc),
	.w3(32'h3a842d23),
	.w4(32'h3b8b20c4),
	.w5(32'h3b115cda),
	.w6(32'h3b72ec61),
	.w7(32'h3b8edad6),
	.w8(32'h3a8699c4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0adef),
	.w1(32'h39967f8f),
	.w2(32'hba4d98f3),
	.w3(32'hba76d818),
	.w4(32'h39161cc0),
	.w5(32'hbb564e51),
	.w6(32'hba8c3757),
	.w7(32'h39d6adad),
	.w8(32'hbb411e3a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba161ce1),
	.w1(32'hba40fb54),
	.w2(32'hbad45998),
	.w3(32'hbb35b7eb),
	.w4(32'hb9a9ae21),
	.w5(32'hbaf6e82c),
	.w6(32'hbb39b130),
	.w7(32'hb97e210e),
	.w8(32'hbb492211),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd1e77),
	.w1(32'h3aba7417),
	.w2(32'hb9ca51f4),
	.w3(32'hbb27e346),
	.w4(32'hbaf7ca5e),
	.w5(32'hbb60b357),
	.w6(32'hba33b5be),
	.w7(32'h3ae88e9b),
	.w8(32'hbb62ac6c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e315),
	.w1(32'hbb83e091),
	.w2(32'h3ae24379),
	.w3(32'hbc09a5dc),
	.w4(32'hbb896a4d),
	.w5(32'h3ace08c7),
	.w6(32'hbc041042),
	.w7(32'hbbf9488d),
	.w8(32'hb95fae44),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8bec),
	.w1(32'h3b211ba1),
	.w2(32'h3bc4a7dd),
	.w3(32'h3ac137eb),
	.w4(32'h3b20bf6a),
	.w5(32'h3a4362ec),
	.w6(32'hba3501af),
	.w7(32'h3b0ac36b),
	.w8(32'h3ac36c2d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fbcab),
	.w1(32'h3beefb3c),
	.w2(32'h3b4ff31a),
	.w3(32'h3bbe6d13),
	.w4(32'h3b86a8cc),
	.w5(32'hbae1f7d7),
	.w6(32'h3be5e79d),
	.w7(32'h3b9e5350),
	.w8(32'hbb818a42),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3caf5),
	.w1(32'h3ae28768),
	.w2(32'h3aeec848),
	.w3(32'hbab20112),
	.w4(32'hbb98f24b),
	.w5(32'h3bad4efd),
	.w6(32'hb8f04646),
	.w7(32'hbb82c087),
	.w8(32'h3beab19b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59fe80),
	.w1(32'hba16e932),
	.w2(32'hbaf19812),
	.w3(32'hbaa355b8),
	.w4(32'hbb307d58),
	.w5(32'hb7a8130d),
	.w6(32'hbadca0a1),
	.w7(32'hbb2c39f4),
	.w8(32'h396c387e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48e2f0),
	.w1(32'h3ac686e0),
	.w2(32'h3bbb22fe),
	.w3(32'h3b29a15b),
	.w4(32'h3afbf92e),
	.w5(32'hbbae284b),
	.w6(32'h3b4c5918),
	.w7(32'h3b24d04c),
	.w8(32'hbb912c4a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf953d7),
	.w1(32'hba64bfbb),
	.w2(32'h3af5c6eb),
	.w3(32'hbb8bc173),
	.w4(32'h37e2899f),
	.w5(32'hb9e5d063),
	.w6(32'hbb904e54),
	.w7(32'h3983fc28),
	.w8(32'hbb061fd9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0269d2),
	.w1(32'hbc426fba),
	.w2(32'hbc3574bf),
	.w3(32'hbbcde975),
	.w4(32'hbb582101),
	.w5(32'hbb900c9c),
	.w6(32'hbbfef391),
	.w7(32'h3adfc403),
	.w8(32'hbb318ceb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffe968),
	.w1(32'hbb97eb79),
	.w2(32'hbb931173),
	.w3(32'hbbbfda04),
	.w4(32'hbb804a9b),
	.w5(32'h3aed1a83),
	.w6(32'hbba9cdb6),
	.w7(32'hbb92f11d),
	.w8(32'h3b19b673),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01f3e8),
	.w1(32'hbabe20b0),
	.w2(32'hbae45898),
	.w3(32'hba8803a0),
	.w4(32'hbb03ae39),
	.w5(32'h3a90e6fc),
	.w6(32'hb88628b2),
	.w7(32'hb99b2968),
	.w8(32'h3a9707f5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a6cf),
	.w1(32'hbc1f6029),
	.w2(32'hbc345fc7),
	.w3(32'hbbdcc519),
	.w4(32'hbba70f13),
	.w5(32'hbb3f81e9),
	.w6(32'hbbc4fdc3),
	.w7(32'hbba38dc3),
	.w8(32'hbb22ee98),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa153ec),
	.w1(32'h3a68aaaa),
	.w2(32'hba0b3be5),
	.w3(32'h3b1289b1),
	.w4(32'h3b236193),
	.w5(32'hbb540a8e),
	.w6(32'h3b5628ee),
	.w7(32'h3ab3a8bc),
	.w8(32'hbabf5866),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a757888),
	.w1(32'hbb0d556e),
	.w2(32'hbbb6ca8b),
	.w3(32'h3986770a),
	.w4(32'h3a2c30e0),
	.w5(32'h39eb2a48),
	.w6(32'h3b5b930d),
	.w7(32'h3adfcf47),
	.w8(32'h3af2517c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a4acf),
	.w1(32'h3a4706bf),
	.w2(32'h3a783a7a),
	.w3(32'h3bb0b3d0),
	.w4(32'h3b9ba521),
	.w5(32'hbbb3fa18),
	.w6(32'h3b6d79c1),
	.w7(32'h3b2ef473),
	.w8(32'hbb51fb47),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af28234),
	.w1(32'hb9a09f78),
	.w2(32'h3aad9f91),
	.w3(32'h3b3312dd),
	.w4(32'h3b403641),
	.w5(32'hbb162d21),
	.w6(32'h3ad0d79f),
	.w7(32'h3b7c63c6),
	.w8(32'hbb5e87a5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198ac3),
	.w1(32'hba8254df),
	.w2(32'h398d4784),
	.w3(32'hbaee7fe1),
	.w4(32'hb85da0d5),
	.w5(32'h3b02652b),
	.w6(32'hbb18fed1),
	.w7(32'h39cfd2d1),
	.w8(32'h3b875396),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00400c),
	.w1(32'hbb5224a1),
	.w2(32'hbb9c94ff),
	.w3(32'hb959fd3b),
	.w4(32'hbb6ebc4a),
	.w5(32'h3ba1b02d),
	.w6(32'hbaf401a4),
	.w7(32'hbb41c05f),
	.w8(32'h3bf25a9a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a0a57),
	.w1(32'h3b1f25f3),
	.w2(32'hb9ca0d73),
	.w3(32'h3ac951ae),
	.w4(32'hbb6788d6),
	.w5(32'hbb52c689),
	.w6(32'h3b10d4fc),
	.w7(32'hbb3f9b03),
	.w8(32'hbae4708f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba1dbd),
	.w1(32'hba1f19b9),
	.w2(32'hbaa62f8b),
	.w3(32'hbb0c14d5),
	.w4(32'hbb185d3a),
	.w5(32'h393faa00),
	.w6(32'hbac955fe),
	.w7(32'hbaea83aa),
	.w8(32'hb96edcbc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f6ae7),
	.w1(32'hba87b8ca),
	.w2(32'hbabfa8cd),
	.w3(32'hbb4fb1c4),
	.w4(32'hbb5284c4),
	.w5(32'h3b34e367),
	.w6(32'hbb4aba32),
	.w7(32'hbadfea5b),
	.w8(32'h3b7ba896),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447af2),
	.w1(32'hba61420b),
	.w2(32'hbb623bec),
	.w3(32'hba69d46e),
	.w4(32'hbb1dc3ea),
	.w5(32'h3ae630cc),
	.w6(32'hbacfadbb),
	.w7(32'hbb15d828),
	.w8(32'h3b5d8a0f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed1a86),
	.w1(32'hba9ba8bb),
	.w2(32'hbb11f9bf),
	.w3(32'hbb0a6c67),
	.w4(32'hbb0a20b9),
	.w5(32'h3b302270),
	.w6(32'hbb489ced),
	.w7(32'hbb22aca9),
	.w8(32'h3b2908dc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acde732),
	.w1(32'h3b9aedd6),
	.w2(32'h3c0e5405),
	.w3(32'h3bcd83d3),
	.w4(32'h3be77d22),
	.w5(32'h3bcf395c),
	.w6(32'h3b884367),
	.w7(32'h3b8c7122),
	.w8(32'h3aca43de),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c76d4),
	.w1(32'hbb944c64),
	.w2(32'hbb2faa78),
	.w3(32'h3bde1677),
	.w4(32'h3ad5cef9),
	.w5(32'hba4472d5),
	.w6(32'h3b90c495),
	.w7(32'h39d44449),
	.w8(32'hb92e08ec),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78c3e5),
	.w1(32'h3a87325f),
	.w2(32'h39ec81e0),
	.w3(32'hbaf6fc2a),
	.w4(32'h3a806e08),
	.w5(32'hbad37703),
	.w6(32'h37c144b0),
	.w7(32'h3b6d78f9),
	.w8(32'hba07c9c4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911a33e),
	.w1(32'h3a800a3f),
	.w2(32'h3b2b405a),
	.w3(32'hbac6fd20),
	.w4(32'hba686afb),
	.w5(32'hbac4eb9e),
	.w6(32'hb9a62843),
	.w7(32'h3a7c7be8),
	.w8(32'hba366086),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7720),
	.w1(32'hba85cfbd),
	.w2(32'hbaf297e6),
	.w3(32'hba834774),
	.w4(32'hb915274b),
	.w5(32'h39c44ea7),
	.w6(32'hb9511e23),
	.w7(32'h3919618b),
	.w8(32'h3ac8fbda),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af99d33),
	.w1(32'hb944aef0),
	.w2(32'hbad924b6),
	.w3(32'hbb0aa411),
	.w4(32'hba8bbd9d),
	.w5(32'hbb83dcc0),
	.w6(32'hbb014d3c),
	.w7(32'hba9ec00c),
	.w8(32'hbb072ec2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb098b72),
	.w1(32'hbaea0ec9),
	.w2(32'hb9930a0b),
	.w3(32'hbb44bd30),
	.w4(32'hbac07237),
	.w5(32'hba956942),
	.w6(32'hbb42e462),
	.w7(32'hba16c0cf),
	.w8(32'hba4744c4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81c7a),
	.w1(32'hba77498a),
	.w2(32'hbab4da62),
	.w3(32'h398770ae),
	.w4(32'hba7dbfb4),
	.w5(32'h3b1ee061),
	.w6(32'hba984abf),
	.w7(32'hba892258),
	.w8(32'h3b137f13),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900b35),
	.w1(32'h3b3dd893),
	.w2(32'h3a79cfc2),
	.w3(32'h3b1f0d6d),
	.w4(32'h3b7482ee),
	.w5(32'h3a9af1e8),
	.w6(32'h3aa029bf),
	.w7(32'h3ac28cd5),
	.w8(32'h38e9808c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17ad0b),
	.w1(32'h3ac4b1d7),
	.w2(32'hb9dafaca),
	.w3(32'h399b7d2f),
	.w4(32'h3b2c7cea),
	.w5(32'hbb971a97),
	.w6(32'hba30d094),
	.w7(32'h3ab9b18e),
	.w8(32'hbb9a7cb2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf8097),
	.w1(32'hbb11ecd8),
	.w2(32'hbb12d2f0),
	.w3(32'hbad55707),
	.w4(32'h3a915abc),
	.w5(32'hbaf49eff),
	.w6(32'hbaf45e4e),
	.w7(32'h3972664b),
	.w8(32'hbb974414),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904d25),
	.w1(32'hbb74986b),
	.w2(32'hbb639914),
	.w3(32'hbb99c3b0),
	.w4(32'hbb532633),
	.w5(32'hbb68cbfc),
	.w6(32'hbb43ceaa),
	.w7(32'hba70d61c),
	.w8(32'hbb940d3c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38788a9b),
	.w1(32'h3a5b8781),
	.w2(32'h3a941382),
	.w3(32'hba9d3ebb),
	.w4(32'h3abf1362),
	.w5(32'hba701e23),
	.w6(32'hba4ea1ed),
	.w7(32'hb9a36428),
	.w8(32'h3b1448f1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0831),
	.w1(32'h3b6f1567),
	.w2(32'h3a1ad69a),
	.w3(32'h3b013775),
	.w4(32'h3a001d54),
	.w5(32'hbba61b79),
	.w6(32'h3b515077),
	.w7(32'h3b0352bb),
	.w8(32'hbb7c074f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95e633),
	.w1(32'hbad3ea96),
	.w2(32'h38c7e98c),
	.w3(32'hbb2fc4b6),
	.w4(32'hbb04947a),
	.w5(32'hbb45d713),
	.w6(32'hbb505388),
	.w7(32'h3a0ca9cf),
	.w8(32'hbadda5b6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb498553),
	.w1(32'hb816d117),
	.w2(32'h3b1b58c2),
	.w3(32'hbb57466d),
	.w4(32'hba8ebe99),
	.w5(32'hba7453ac),
	.w6(32'hbb47a312),
	.w7(32'h39a119a0),
	.w8(32'hbb4290eb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e945),
	.w1(32'h3a677fa1),
	.w2(32'h3a193fc7),
	.w3(32'hbb34fa01),
	.w4(32'hba4e1a6f),
	.w5(32'hbb49c106),
	.w6(32'hbb690c94),
	.w7(32'h3a83b60c),
	.w8(32'hbb243944),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2993c5),
	.w1(32'hbb19f96f),
	.w2(32'hbb520ae6),
	.w3(32'hbb8f0612),
	.w4(32'hbb907266),
	.w5(32'h38ddf10a),
	.w6(32'hbb006899),
	.w7(32'hbab1250b),
	.w8(32'h3b3beafa),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b080227),
	.w1(32'h39d04ac4),
	.w2(32'hbb000d47),
	.w3(32'hba7fd40c),
	.w4(32'hb97fb7c5),
	.w5(32'hbaa170dc),
	.w6(32'h3a94774d),
	.w7(32'hba464aaf),
	.w8(32'hbb0a5a08),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a18c),
	.w1(32'h399f2851),
	.w2(32'hb9fb34fa),
	.w3(32'hbb370b2c),
	.w4(32'hba4246ea),
	.w5(32'h398f143f),
	.w6(32'hbaefa6c0),
	.w7(32'hb93f91ca),
	.w8(32'h3b0a52cc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc7ff),
	.w1(32'hba429fc8),
	.w2(32'hbabb80c8),
	.w3(32'h3b21ce0b),
	.w4(32'h3b0c1d79),
	.w5(32'hba688979),
	.w6(32'h3b271b6c),
	.w7(32'hb8e8e0df),
	.w8(32'hbb0596a1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad59d97),
	.w1(32'h3a158076),
	.w2(32'h36768241),
	.w3(32'hba5417c3),
	.w4(32'hba5b429b),
	.w5(32'h3b534f04),
	.w6(32'hbad41768),
	.w7(32'hba2c9fd8),
	.w8(32'h3be639e2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13afe7),
	.w1(32'h3b772e37),
	.w2(32'h3af79ca0),
	.w3(32'h3bb5b2bc),
	.w4(32'h3b7ccc39),
	.w5(32'hbae60c85),
	.w6(32'h3c0416f4),
	.w7(32'h3b2b1068),
	.w8(32'hbb146fe8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386b34b7),
	.w1(32'h3a86126e),
	.w2(32'h3a676f95),
	.w3(32'hba39e361),
	.w4(32'h39c916e9),
	.w5(32'hbaa7110b),
	.w6(32'hba3a657a),
	.w7(32'h3aa2cdfa),
	.w8(32'hbaab9f39),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ed343),
	.w1(32'hbae04710),
	.w2(32'hbb0ee869),
	.w3(32'hbab99237),
	.w4(32'h39b56f8a),
	.w5(32'hbb32eff0),
	.w6(32'hba200331),
	.w7(32'hb9d38b56),
	.w8(32'hbb814301),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6ea57),
	.w1(32'hbb51024a),
	.w2(32'hbb503279),
	.w3(32'hbbbcaf88),
	.w4(32'hbb228bde),
	.w5(32'hbb135297),
	.w6(32'hbbb4f08c),
	.w7(32'hbb4b892b),
	.w8(32'hbb1047cb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c16d),
	.w1(32'hb93f132a),
	.w2(32'hb9ffa0a0),
	.w3(32'hbb0645bc),
	.w4(32'hba41cba5),
	.w5(32'hbada69a7),
	.w6(32'h3915f1cf),
	.w7(32'hba2cf27d),
	.w8(32'hbacc576f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940292f),
	.w1(32'hbb05f51c),
	.w2(32'hba6553a6),
	.w3(32'hbad237d3),
	.w4(32'h3a9dc57a),
	.w5(32'h3ae419f9),
	.w6(32'hba1dd66d),
	.w7(32'h3b2901b0),
	.w8(32'h3b5fda5d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fc73b),
	.w1(32'hb9496042),
	.w2(32'h3b3e1ae4),
	.w3(32'h3b2a816d),
	.w4(32'hba20f9cd),
	.w5(32'hbac1def8),
	.w6(32'hba22a36a),
	.w7(32'hba977403),
	.w8(32'hbab3c1f7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce8454),
	.w1(32'h3a0823c7),
	.w2(32'hba334b70),
	.w3(32'h39e8e888),
	.w4(32'h3a989fe4),
	.w5(32'h38cb609c),
	.w6(32'h39f9a32c),
	.w7(32'h3a9ccb53),
	.w8(32'hba7f0168),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae8289),
	.w1(32'h38bca9bd),
	.w2(32'h3b0779e1),
	.w3(32'hba76ca18),
	.w4(32'hba45c92d),
	.w5(32'h383502a9),
	.w6(32'hbaf20f6a),
	.w7(32'hba290f80),
	.w8(32'h3aaca7c1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06897e),
	.w1(32'h3a7925f4),
	.w2(32'h3a149fe6),
	.w3(32'h3b5fb0c7),
	.w4(32'h3ac6acf8),
	.w5(32'hba9997cf),
	.w6(32'h3b4d5ddf),
	.w7(32'hba3463cd),
	.w8(32'hbb54bdc0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b15cb),
	.w1(32'h3b579729),
	.w2(32'h3aa61f3b),
	.w3(32'hba83c1fc),
	.w4(32'hba35f62d),
	.w5(32'h3b3ff622),
	.w6(32'h3a26de6f),
	.w7(32'hba1bb9b5),
	.w8(32'h3b5c7d41),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba59c5),
	.w1(32'h3addc2c1),
	.w2(32'h3b454f19),
	.w3(32'hbac6c9b4),
	.w4(32'hbab828cc),
	.w5(32'hbaff4bd1),
	.w6(32'hbacbc2b7),
	.w7(32'h3a69ff36),
	.w8(32'hbb28c178),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ae134),
	.w1(32'hbb118b9d),
	.w2(32'h3a822778),
	.w3(32'hba1aad6b),
	.w4(32'h3945ff32),
	.w5(32'hbab93bdc),
	.w6(32'hbb5f9942),
	.w7(32'hba641586),
	.w8(32'hbabbf27f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb704b9b),
	.w1(32'hbb422aa5),
	.w2(32'hbb894eb1),
	.w3(32'hbb122937),
	.w4(32'hbaf34548),
	.w5(32'hbb9de582),
	.w6(32'hbb4bd55e),
	.w7(32'hbb309bcd),
	.w8(32'hbbb2e94c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819e9a),
	.w1(32'hba76f61d),
	.w2(32'hbacbd32e),
	.w3(32'hbb094dc1),
	.w4(32'h39e2c0c8),
	.w5(32'hbba378af),
	.w6(32'hbadbf8f8),
	.w7(32'hba30e633),
	.w8(32'hbbecc8c7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9613e),
	.w1(32'hbb28b15e),
	.w2(32'hba05801a),
	.w3(32'hbb3eaceb),
	.w4(32'h392fcab8),
	.w5(32'hbbaebed0),
	.w6(32'hbba7552f),
	.w7(32'h3b01fd8e),
	.w8(32'hba9e7040),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb809cc9),
	.w1(32'hbb83af6d),
	.w2(32'hbb7e09d9),
	.w3(32'h3a049f3d),
	.w4(32'h39e10d2b),
	.w5(32'h3b750470),
	.w6(32'hba5c7440),
	.w7(32'h3b0a95fd),
	.w8(32'h3b867982),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf5a34),
	.w1(32'hbb8b53fe),
	.w2(32'hbc4b965d),
	.w3(32'hb9ffad15),
	.w4(32'h3b2e8040),
	.w5(32'hbadc5e4b),
	.w6(32'hb9f4c78e),
	.w7(32'h3aec66f3),
	.w8(32'hbb49e6a3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2c9ed),
	.w1(32'h3b89ae5c),
	.w2(32'h3a0fd174),
	.w3(32'h3bb8e463),
	.w4(32'h3b77e450),
	.w5(32'hbb2ea284),
	.w6(32'h3b144a52),
	.w7(32'h3923072f),
	.w8(32'hbb7f7140),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb272722),
	.w1(32'hbaf3614e),
	.w2(32'hbb58f707),
	.w3(32'hbb233b94),
	.w4(32'hbb2502fe),
	.w5(32'h39fb53cb),
	.w6(32'hbb0e3c3b),
	.w7(32'hbb2d0f3c),
	.w8(32'h38ecfb7d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970686),
	.w1(32'hbab3e7df),
	.w2(32'hb98bc1f9),
	.w3(32'hbb1b9ad4),
	.w4(32'hba9696ce),
	.w5(32'h3b7ab6f0),
	.w6(32'hbb576d88),
	.w7(32'hbb596372),
	.w8(32'h3a2f6a17),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9019686),
	.w1(32'hbadd1bde),
	.w2(32'hbbc51fb5),
	.w3(32'h39ba919a),
	.w4(32'h3a46eeb9),
	.w5(32'hbaf2c9f7),
	.w6(32'hba93d06e),
	.w7(32'h3a8dc214),
	.w8(32'hbb4025ce),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38fd3a),
	.w1(32'hb996dceb),
	.w2(32'hb9518262),
	.w3(32'hbb33bb15),
	.w4(32'h3a8a6249),
	.w5(32'hba1ce893),
	.w6(32'hbb34e82d),
	.w7(32'h3a34ac44),
	.w8(32'hbad00ccf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8fe81),
	.w1(32'hbad3b521),
	.w2(32'hbb9c8354),
	.w3(32'h3baf3313),
	.w4(32'h3bcfa262),
	.w5(32'h3a287ae0),
	.w6(32'h3b32521f),
	.w7(32'h3b972dd7),
	.w8(32'hba838414),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48e1ab),
	.w1(32'hbb1b7b0b),
	.w2(32'hbb1d535d),
	.w3(32'hbb0e4831),
	.w4(32'hbaf7c660),
	.w5(32'hbb0d25ea),
	.w6(32'hbb375d41),
	.w7(32'hbb2d9625),
	.w8(32'hba71a505),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace5a80),
	.w1(32'hb935b1c4),
	.w2(32'hbadcdf2f),
	.w3(32'hbb1bf951),
	.w4(32'hbb1695e0),
	.w5(32'hba771de2),
	.w6(32'h3a5c42a7),
	.w7(32'h390a8078),
	.w8(32'hb9226380),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55f725),
	.w1(32'hba69a5b8),
	.w2(32'hbaae9b2d),
	.w3(32'hbabd4224),
	.w4(32'hbaf1d596),
	.w5(32'h39bdc63c),
	.w6(32'hba8bdfa1),
	.w7(32'hba743510),
	.w8(32'h3813f1c1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970f716),
	.w1(32'h3992d5b5),
	.w2(32'h3acceb42),
	.w3(32'h39e0d0f6),
	.w4(32'h3a433a66),
	.w5(32'h3b083cb2),
	.w6(32'hb9326053),
	.w7(32'h3a149714),
	.w8(32'h3a9389db),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5541ed),
	.w1(32'h3aebfa2d),
	.w2(32'hba7d2db9),
	.w3(32'h3b5df103),
	.w4(32'h3a857f82),
	.w5(32'h3aeb95bb),
	.w6(32'h3a4343d9),
	.w7(32'hba4a56ef),
	.w8(32'h3a0e1f48),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdd84e),
	.w1(32'h39121d9d),
	.w2(32'hbb86d653),
	.w3(32'h3b3a0746),
	.w4(32'h3b2b6bf3),
	.w5(32'hbb455e8e),
	.w6(32'h3a901a89),
	.w7(32'h3ad4c492),
	.w8(32'hbb397550),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011417),
	.w1(32'hbb143aae),
	.w2(32'hbb2eb10f),
	.w3(32'hbb21b8ad),
	.w4(32'hbb22faa5),
	.w5(32'h3a3565f3),
	.w6(32'hbae8efc0),
	.w7(32'hbaa8fa0b),
	.w8(32'h390a5c9f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e46a88),
	.w1(32'h3aa76917),
	.w2(32'h3a6ca27b),
	.w3(32'h3a51b01d),
	.w4(32'h3ab731f5),
	.w5(32'hb9e3d667),
	.w6(32'hbaaa9f93),
	.w7(32'h3964f492),
	.w8(32'hba92ad59),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2be4f),
	.w1(32'h39080087),
	.w2(32'h3a55456e),
	.w3(32'hb92f091f),
	.w4(32'h39ef7e30),
	.w5(32'h3a90c255),
	.w6(32'h3a0b3391),
	.w7(32'h3a0c3513),
	.w8(32'h3a20a541),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f6f9),
	.w1(32'hbb1e33d7),
	.w2(32'hb9b45a01),
	.w3(32'hbb820066),
	.w4(32'hbb4f9883),
	.w5(32'hbb0dee6e),
	.w6(32'hbb830301),
	.w7(32'hbaefb76e),
	.w8(32'hbb045733),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf52c4f),
	.w1(32'hbac46b68),
	.w2(32'hbb419c17),
	.w3(32'hbad29766),
	.w4(32'hbb0423da),
	.w5(32'hb99c2840),
	.w6(32'hbaacffac),
	.w7(32'hbb2b577e),
	.w8(32'hbab11461),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba255052),
	.w1(32'hba158070),
	.w2(32'hb986b9fe),
	.w3(32'hb8f120f2),
	.w4(32'hba32848d),
	.w5(32'h3943ae34),
	.w6(32'hbae439db),
	.w7(32'hb989ce55),
	.w8(32'h39b66042),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56da31),
	.w1(32'h3a2b7fe6),
	.w2(32'h39962ecf),
	.w3(32'h3a01173a),
	.w4(32'h39360b2d),
	.w5(32'hb9c64ed2),
	.w6(32'h3a80e949),
	.w7(32'h3a355f35),
	.w8(32'hba5c2f54),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2457),
	.w1(32'hbb1bf1a7),
	.w2(32'hbb00a934),
	.w3(32'hba461805),
	.w4(32'h38ba3840),
	.w5(32'h3ad40e96),
	.w6(32'hbaa9860b),
	.w7(32'hba737047),
	.w8(32'h3a99cfc8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabd1c0),
	.w1(32'h3ae9754c),
	.w2(32'h3af3af96),
	.w3(32'h3a89e3b9),
	.w4(32'h3af5cb20),
	.w5(32'h3a20a68d),
	.w6(32'h3a8de6f4),
	.w7(32'h3abefc71),
	.w8(32'hba68294b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cef0d0),
	.w1(32'hba814a4f),
	.w2(32'hba6d6dc1),
	.w3(32'hba814014),
	.w4(32'hba6fcb21),
	.w5(32'h3a1704a4),
	.w6(32'hbb08f266),
	.w7(32'hbac03965),
	.w8(32'h3a1410d9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cecc82),
	.w1(32'h38818579),
	.w2(32'h3a44b3c2),
	.w3(32'h388d39a2),
	.w4(32'h3a2c061f),
	.w5(32'hba1e5e78),
	.w6(32'hb99d42bc),
	.w7(32'h3a13d999),
	.w8(32'hba126270),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cec8b),
	.w1(32'hbaeab458),
	.w2(32'hba8d0f54),
	.w3(32'hbaf96525),
	.w4(32'hba7d9bab),
	.w5(32'hbad909e2),
	.w6(32'hbb1fcb3f),
	.w7(32'hbab9ec78),
	.w8(32'hb9d5acd6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a1e03a),
	.w1(32'hba120b15),
	.w2(32'hba41acf4),
	.w3(32'hbb0653d4),
	.w4(32'hba918844),
	.w5(32'hba8b4896),
	.w6(32'hbab28d8a),
	.w7(32'h397d5fcc),
	.w8(32'hba87641c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a1f4),
	.w1(32'hbafa7793),
	.w2(32'hba476874),
	.w3(32'hbaa2580d),
	.w4(32'hba1567ef),
	.w5(32'hba692dd1),
	.w6(32'hbb1de5c8),
	.w7(32'hba46fe62),
	.w8(32'hb9a66979),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff4aba),
	.w1(32'h3a306048),
	.w2(32'h3903e64f),
	.w3(32'hba1d0e68),
	.w4(32'hba4b66a9),
	.w5(32'hb788dc63),
	.w6(32'hbaabcc90),
	.w7(32'hba7565c9),
	.w8(32'hba8555fa),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa903f9),
	.w1(32'hb9717f11),
	.w2(32'h3a6d1509),
	.w3(32'h3a4e9240),
	.w4(32'h3a9e6c61),
	.w5(32'h392e3886),
	.w6(32'hba3eac0b),
	.w7(32'h399f3f88),
	.w8(32'h3a522abc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ef765),
	.w1(32'h3892c568),
	.w2(32'h3912fa83),
	.w3(32'h391ca781),
	.w4(32'hb7be48bb),
	.w5(32'hba4db734),
	.w6(32'h3992312b),
	.w7(32'h391c021b),
	.w8(32'hba34b91f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6015d4),
	.w1(32'hbab64ee0),
	.w2(32'hba8a1d27),
	.w3(32'hbaf300ff),
	.w4(32'hbae0a0b4),
	.w5(32'hba4a9826),
	.w6(32'hbaa716bd),
	.w7(32'hbaed21bb),
	.w8(32'hba99e53e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968a24),
	.w1(32'hba8b00a1),
	.w2(32'h3a0b1761),
	.w3(32'hba7cc231),
	.w4(32'h39e7ef1f),
	.w5(32'hbaaecb81),
	.w6(32'hbaa879e4),
	.w7(32'hb927f556),
	.w8(32'hba182728),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31c1d4),
	.w1(32'hba92db6f),
	.w2(32'hba59793c),
	.w3(32'hbab7859d),
	.w4(32'hba98d412),
	.w5(32'h3a5abe36),
	.w6(32'hba8110ce),
	.w7(32'hba3cb1ed),
	.w8(32'h3a6c2fcd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c699a8),
	.w1(32'h3ac1191d),
	.w2(32'h3ad3d67c),
	.w3(32'h3a121c17),
	.w4(32'h38ba1040),
	.w5(32'h3ab3564b),
	.w6(32'h39a374aa),
	.w7(32'h3a9ab923),
	.w8(32'h3aa01ffd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac13068),
	.w1(32'h3a7f4195),
	.w2(32'h3a2bbd45),
	.w3(32'h3a648298),
	.w4(32'h3a11012e),
	.w5(32'h3b096cb4),
	.w6(32'h3a52ba7a),
	.w7(32'h3a5b0593),
	.w8(32'h3a2a2e64),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1b244),
	.w1(32'h396f3445),
	.w2(32'h37a14c1a),
	.w3(32'h3b0b60db),
	.w4(32'h3b42ad55),
	.w5(32'hba00322f),
	.w6(32'h3a304c99),
	.w7(32'h3ae08a2f),
	.w8(32'hb943aa8a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e24c41),
	.w1(32'h398a11d5),
	.w2(32'h3a1c6605),
	.w3(32'hb9556850),
	.w4(32'h39a3ece3),
	.w5(32'h396b5b13),
	.w6(32'hba0999e3),
	.w7(32'h39ce27e5),
	.w8(32'h3a37dc29),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91363f1),
	.w1(32'hb9ec0ed1),
	.w2(32'hba6c4429),
	.w3(32'hba4f22fe),
	.w4(32'hb9fd6404),
	.w5(32'h39ea26bc),
	.w6(32'hb9cf1963),
	.w7(32'hb94e15ca),
	.w8(32'hb6dfc278),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88cd0cc),
	.w1(32'h3a2378ea),
	.w2(32'h3a01f9c6),
	.w3(32'h36b25c51),
	.w4(32'h39e75009),
	.w5(32'hba792386),
	.w6(32'hb77e588c),
	.w7(32'h39675572),
	.w8(32'hba923181),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02bd79),
	.w1(32'hba31400c),
	.w2(32'hba8cc4ec),
	.w3(32'hba0f8f13),
	.w4(32'h36e99e7c),
	.w5(32'hb9796f8f),
	.w6(32'hba83059f),
	.w7(32'hb93bcda7),
	.w8(32'hb871aa9f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddf6dc),
	.w1(32'h39a8b457),
	.w2(32'h3a1f10da),
	.w3(32'hb8bc0a23),
	.w4(32'h39e4b01e),
	.w5(32'h390aa133),
	.w6(32'hba1fb911),
	.w7(32'h39887cb4),
	.w8(32'h39cc7ceb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba1ac9),
	.w1(32'h39195efb),
	.w2(32'h3a22a559),
	.w3(32'hbaa2b3c1),
	.w4(32'hba198228),
	.w5(32'hbb124b84),
	.w6(32'hbad6090c),
	.w7(32'h3955cd78),
	.w8(32'hbab01d04),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34b9df),
	.w1(32'hbb141c97),
	.w2(32'hbaf9dae0),
	.w3(32'hbb2fa1b1),
	.w4(32'hbb221814),
	.w5(32'hbb48de75),
	.w6(32'hbb27503f),
	.w7(32'hbafc1c68),
	.w8(32'hbb40e85c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf86c0d),
	.w1(32'hba4e48f2),
	.w2(32'hbb05e2a4),
	.w3(32'hba7581b0),
	.w4(32'hba92a761),
	.w5(32'h39a91dda),
	.w6(32'hbac48653),
	.w7(32'hbb0e1bd9),
	.w8(32'hb94fd318),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad278b),
	.w1(32'h399c6fb5),
	.w2(32'hba5b6b69),
	.w3(32'hb883f0e1),
	.w4(32'hb8db1be5),
	.w5(32'hbb481a3d),
	.w6(32'hba0daa6d),
	.w7(32'hb9c56613),
	.w8(32'hbb1502c4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cb7e2),
	.w1(32'hba489de4),
	.w2(32'hbab0f0dd),
	.w3(32'hbac50cb1),
	.w4(32'hbace39de),
	.w5(32'hb9bb0442),
	.w6(32'hba55e4e6),
	.w7(32'hba836043),
	.w8(32'hba0bbc01),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39216bd0),
	.w1(32'h388f6052),
	.w2(32'h395078db),
	.w3(32'hba174f91),
	.w4(32'hb91d1870),
	.w5(32'hb991406f),
	.w6(32'hba749788),
	.w7(32'hba125cfe),
	.w8(32'h37550e45),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823313d),
	.w1(32'h38895884),
	.w2(32'h3a23603f),
	.w3(32'hb8c759cc),
	.w4(32'hb90e6045),
	.w5(32'hbaf1eef7),
	.w6(32'h350dd7f8),
	.w7(32'h38eae64b),
	.w8(32'hba9a4c31),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4fc4a),
	.w1(32'hba7e92d6),
	.w2(32'hbae45e47),
	.w3(32'hbaf3615d),
	.w4(32'hbaf52347),
	.w5(32'hbace41bd),
	.w6(32'hba38563d),
	.w7(32'hbae43e40),
	.w8(32'hbad4933d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28c192),
	.w1(32'hbb2da670),
	.w2(32'hbb593b20),
	.w3(32'hbaac0357),
	.w4(32'hbb0019a1),
	.w5(32'hba9f363b),
	.w6(32'hbaa26fdd),
	.w7(32'hbb17221f),
	.w8(32'hbab3f65d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee6ab3),
	.w1(32'hb9ae055f),
	.w2(32'hb9324a0a),
	.w3(32'hb968973e),
	.w4(32'hb8f77378),
	.w5(32'h384025ee),
	.w6(32'hba88970a),
	.w7(32'hba1da0bc),
	.w8(32'hb9a51f48),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a539f84),
	.w1(32'h3a8c9877),
	.w2(32'h3a1861db),
	.w3(32'h3a2852f8),
	.w4(32'h394fa916),
	.w5(32'h3a6a876e),
	.w6(32'h39ce7b53),
	.w7(32'h39e819ce),
	.w8(32'h3a8c2ce0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960c477),
	.w1(32'h39090a98),
	.w2(32'hba78157b),
	.w3(32'hba16f945),
	.w4(32'h387bcd05),
	.w5(32'h38a118c1),
	.w6(32'hba1601a6),
	.w7(32'hb89c490a),
	.w8(32'hb9a45894),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3836bc),
	.w1(32'h39f27c58),
	.w2(32'hbb4c0ff8),
	.w3(32'h3adfd18d),
	.w4(32'h3a5dd140),
	.w5(32'hbb52a3cd),
	.w6(32'h3b1baccd),
	.w7(32'hb958fa0d),
	.w8(32'hbb9401bf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65b503),
	.w1(32'hbae72495),
	.w2(32'hba475f73),
	.w3(32'hbb8dad73),
	.w4(32'hbb2eb680),
	.w5(32'hbb7790b6),
	.w6(32'hbba1cbd6),
	.w7(32'hbb5dd8a4),
	.w8(32'hbb7a6d87),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa08761),
	.w1(32'hba2543e7),
	.w2(32'hba972c06),
	.w3(32'hba8d71f2),
	.w4(32'hba5768e1),
	.w5(32'h397f508e),
	.w6(32'hbac36e50),
	.w7(32'hba153f22),
	.w8(32'hb4d32a58),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f5489),
	.w1(32'h3b21d74b),
	.w2(32'h3a70a9c4),
	.w3(32'h3b6e7b19),
	.w4(32'h3b0868dd),
	.w5(32'h3a80ea52),
	.w6(32'h3b060ca5),
	.w7(32'h3a7a2799),
	.w8(32'hb99e1bb4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba702),
	.w1(32'h3a366888),
	.w2(32'hbb57b651),
	.w3(32'h3bf45bfc),
	.w4(32'h3b9f3398),
	.w5(32'h3b2434bd),
	.w6(32'h3b9f32af),
	.w7(32'h3b810052),
	.w8(32'h3b30aecc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad441),
	.w1(32'hbb888fa3),
	.w2(32'hbb89cd94),
	.w3(32'hbc0399c6),
	.w4(32'hbb50e35e),
	.w5(32'hbb533e9e),
	.w6(32'hbbcf3653),
	.w7(32'hbb105c72),
	.w8(32'hbac2d175),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba624c14),
	.w1(32'hba4e9628),
	.w2(32'hb81d6b0f),
	.w3(32'hb92b9632),
	.w4(32'h3a49173e),
	.w5(32'hba4c2b83),
	.w6(32'hba6ef2ca),
	.w7(32'h39bb0781),
	.w8(32'hba16938f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57bf0d),
	.w1(32'h3926e5c3),
	.w2(32'h3add2f17),
	.w3(32'hb997f00b),
	.w4(32'h3a81ddfa),
	.w5(32'h37f11432),
	.w6(32'hba33c01c),
	.w7(32'h3a0218b2),
	.w8(32'hba001b16),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c0188),
	.w1(32'hba367402),
	.w2(32'hbac20914),
	.w3(32'hba1abcf4),
	.w4(32'hba38a6df),
	.w5(32'hba072e79),
	.w6(32'hba9d8c11),
	.w7(32'hbabc574f),
	.w8(32'h398bef74),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3876739e),
	.w1(32'hb7adc6a6),
	.w2(32'hb64a6c35),
	.w3(32'h38a2cde2),
	.w4(32'hba78b743),
	.w5(32'hba6dbcfa),
	.w6(32'h3962e617),
	.w7(32'h39a83436),
	.w8(32'hbac30944),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab41221),
	.w1(32'hbae36529),
	.w2(32'hbb57cdc7),
	.w3(32'hbaaea4a1),
	.w4(32'hbb0cc85f),
	.w5(32'hbafbd973),
	.w6(32'hbad93639),
	.w7(32'hbb3e3c92),
	.w8(32'hbad4e216),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab13960),
	.w1(32'hba5929e2),
	.w2(32'hba61802b),
	.w3(32'hbadf0895),
	.w4(32'hba205bb1),
	.w5(32'hb9343302),
	.w6(32'hba0ae326),
	.w7(32'hba1dc519),
	.w8(32'h39f5aee4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cf4a4c),
	.w1(32'h387a0b25),
	.w2(32'hb96e4b5b),
	.w3(32'hbad5c885),
	.w4(32'h3925767b),
	.w5(32'hb99691ba),
	.w6(32'hba735ee5),
	.w7(32'h3a9fcbcb),
	.w8(32'h3a0dd694),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9960470),
	.w1(32'h3ac5433f),
	.w2(32'hb9f0593c),
	.w3(32'hba62aa00),
	.w4(32'hba5b317b),
	.w5(32'h3884eafe),
	.w6(32'hb93d9579),
	.w7(32'h38825283),
	.w8(32'h3a2b2c17),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1adb3),
	.w1(32'hba27f0ab),
	.w2(32'hbb034216),
	.w3(32'h3b4385a8),
	.w4(32'h3ac7ac2b),
	.w5(32'hb8835840),
	.w6(32'h3b06fd6a),
	.w7(32'hb973850e),
	.w8(32'h385e8645),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979154d),
	.w1(32'hb916da2e),
	.w2(32'hb9fdc85d),
	.w3(32'h3a1a2e8c),
	.w4(32'h39e065bd),
	.w5(32'h3a207eff),
	.w6(32'h3a14346c),
	.w7(32'h3a19e24d),
	.w8(32'hb9d55dce),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f9eca),
	.w1(32'hba8bc3f9),
	.w2(32'hba0fd470),
	.w3(32'h3a5c7625),
	.w4(32'h3a447f01),
	.w5(32'h3b135ccc),
	.w6(32'hba2587a3),
	.w7(32'hba0d3460),
	.w8(32'h3aefd2d2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fbb53),
	.w1(32'hba0d4162),
	.w2(32'hba3acb17),
	.w3(32'hbb0133f3),
	.w4(32'h3ac8015b),
	.w5(32'hb9aebd26),
	.w6(32'hbb1daaf1),
	.w7(32'hba06ee79),
	.w8(32'h39263e8d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6b4c3),
	.w1(32'hbb9535ef),
	.w2(32'hbb681348),
	.w3(32'hbba7aa9b),
	.w4(32'hbae910cc),
	.w5(32'hba1470ee),
	.w6(32'hbbb5b17c),
	.w7(32'hbb01024d),
	.w8(32'hba48be57),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971a73),
	.w1(32'h3b1d61e4),
	.w2(32'h3ab7a086),
	.w3(32'h3b90ff5f),
	.w4(32'h3aefa129),
	.w5(32'hba93c0ef),
	.w6(32'h3b9d5afd),
	.w7(32'h3b511820),
	.w8(32'h3a572d5b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a561541),
	.w1(32'h3a9d033e),
	.w2(32'h3a54cba6),
	.w3(32'h3aa98ae3),
	.w4(32'h3a0c3db4),
	.w5(32'hb8b7cf84),
	.w6(32'h39ffb323),
	.w7(32'hb9f43b88),
	.w8(32'hba0271b2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad348f8),
	.w1(32'hbaa5bbcf),
	.w2(32'hbad7a38f),
	.w3(32'hbaafb2da),
	.w4(32'hbb3a2f8d),
	.w5(32'h3acfa78a),
	.w6(32'hbadaacf5),
	.w7(32'hbb0692bd),
	.w8(32'h3a91af8c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392982d3),
	.w1(32'h3a6a7079),
	.w2(32'h3ac97856),
	.w3(32'hb9cbf9c4),
	.w4(32'h397a51c9),
	.w5(32'h3820f8ed),
	.w6(32'hb9fa05d8),
	.w7(32'hba386f4a),
	.w8(32'hb91a37cb),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85b086),
	.w1(32'hbab5b05d),
	.w2(32'hbb30c267),
	.w3(32'h38a4fbba),
	.w4(32'h39c5c914),
	.w5(32'hbb318a6a),
	.w6(32'hba921734),
	.w7(32'hba82bf8a),
	.w8(32'hbb48d7e9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1373e),
	.w1(32'hbb7367a0),
	.w2(32'hbb8ab21a),
	.w3(32'hbb80d91a),
	.w4(32'hbb171eb7),
	.w5(32'hba93e5b6),
	.w6(32'hbbcd6132),
	.w7(32'hbb8c4331),
	.w8(32'hbaf3c358),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1183c9),
	.w1(32'h3ade01f1),
	.w2(32'h3ac620c2),
	.w3(32'h3b2295b8),
	.w4(32'h3b42698e),
	.w5(32'h39c3aec4),
	.w6(32'h3b169df7),
	.w7(32'h3b7902eb),
	.w8(32'h3b05f052),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58287c),
	.w1(32'hbac041b4),
	.w2(32'hbb0f7835),
	.w3(32'hbb7108f2),
	.w4(32'hbb239446),
	.w5(32'hb7d2926c),
	.w6(32'hbb4ae36e),
	.w7(32'hbb2c460b),
	.w8(32'hb9049d43),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985b27),
	.w1(32'h3a0ace9e),
	.w2(32'h386119d3),
	.w3(32'h39dd67b4),
	.w4(32'hb90a9087),
	.w5(32'h3af32e96),
	.w6(32'h3a4721a5),
	.w7(32'hb896dd6c),
	.w8(32'h39fbfd4e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982f12),
	.w1(32'hba92fe83),
	.w2(32'hb908d949),
	.w3(32'h3a361162),
	.w4(32'h39cfbe33),
	.w5(32'hba4696ba),
	.w6(32'hbabcb2cf),
	.w7(32'hb916a7b8),
	.w8(32'hb9cccf71),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e0739),
	.w1(32'hba3fa0f4),
	.w2(32'hba62cf55),
	.w3(32'hba5da565),
	.w4(32'hba7efaca),
	.w5(32'h349fbdf8),
	.w6(32'hb7ddaf94),
	.w7(32'hba95c1f5),
	.w8(32'h3a165ae8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395239fa),
	.w1(32'h378e9281),
	.w2(32'h3998f7bc),
	.w3(32'hb9f819f6),
	.w4(32'hba49e349),
	.w5(32'hba2aabd1),
	.w6(32'hba7ed94a),
	.w7(32'hb9dbc5d0),
	.w8(32'hba6d0d66),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9deb8f3),
	.w1(32'hbaa13fd1),
	.w2(32'hb940ad9d),
	.w3(32'hbaec6ec2),
	.w4(32'hba33ee02),
	.w5(32'hba05a987),
	.w6(32'hba2d1b27),
	.w7(32'hba717062),
	.w8(32'hb9a1d656),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de0b7c),
	.w1(32'hb7eeaba8),
	.w2(32'hba105a8e),
	.w3(32'hb9d08414),
	.w4(32'hba78d404),
	.w5(32'h398be907),
	.w6(32'hba02751a),
	.w7(32'hb9db650b),
	.w8(32'h3a2d9ff5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a373a61),
	.w1(32'h39e827ce),
	.w2(32'h3a11732d),
	.w3(32'h3907086e),
	.w4(32'h3a3fdf10),
	.w5(32'hba6212e6),
	.w6(32'h37c2540a),
	.w7(32'h3a2498b7),
	.w8(32'hb9bd8829),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f30618),
	.w1(32'hb9df5374),
	.w2(32'h37fcb0df),
	.w3(32'h39900fca),
	.w4(32'h388c1549),
	.w5(32'h3942a8ba),
	.w6(32'h38b44dc2),
	.w7(32'h38fd4d2a),
	.w8(32'hb9c9b247),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77c4b15),
	.w1(32'h3849f070),
	.w2(32'h3a1bdb66),
	.w3(32'hb9c854be),
	.w4(32'h3a118ff8),
	.w5(32'h3a5bfb4d),
	.w6(32'hb97411f6),
	.w7(32'h3a37119e),
	.w8(32'h3a75d688),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1399f),
	.w1(32'h39d00385),
	.w2(32'hb96e480a),
	.w3(32'h3a0ff055),
	.w4(32'hb9efef06),
	.w5(32'h39ef3c8e),
	.w6(32'h3aa8d884),
	.w7(32'h390ef8e1),
	.w8(32'h3a7efdd7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce3b83),
	.w1(32'hba92f68b),
	.w2(32'hbba1fe04),
	.w3(32'h3b7acde5),
	.w4(32'h3b1cfd21),
	.w5(32'hbb768438),
	.w6(32'h39f2396a),
	.w7(32'h3ab5645c),
	.w8(32'hbb4cf9ce),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56ae1),
	.w1(32'hbb5f5ed7),
	.w2(32'hbb3c8a94),
	.w3(32'hbb56618a),
	.w4(32'hba8ea258),
	.w5(32'hbaa62ece),
	.w6(32'hbbad2172),
	.w7(32'hbb32fb17),
	.w8(32'hbab3ef78),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3607eb),
	.w1(32'h39b3f62c),
	.w2(32'h396d7b84),
	.w3(32'h3a46d901),
	.w4(32'h3a702c08),
	.w5(32'h3a4d5e4b),
	.w6(32'h3ad79588),
	.w7(32'h3ae4b82b),
	.w8(32'h3a9e3d86),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5b2c9),
	.w1(32'h39e34ee1),
	.w2(32'h39d87f41),
	.w3(32'hb9651a2e),
	.w4(32'hb8d9d43d),
	.w5(32'hba92331a),
	.w6(32'hba0c0ad8),
	.w7(32'h38c7c3a9),
	.w8(32'hba938ecb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb085590),
	.w1(32'hbad4691a),
	.w2(32'hba4fcc7d),
	.w3(32'hba9f078c),
	.w4(32'h3a0571c9),
	.w5(32'hb9414b0b),
	.w6(32'hbaa36771),
	.w7(32'hb73bad30),
	.w8(32'hb8d982dc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40d5bb),
	.w1(32'hb8093f56),
	.w2(32'h39d28b64),
	.w3(32'hb992afb9),
	.w4(32'h39ac7e5e),
	.w5(32'hb99559a4),
	.w6(32'hb98dbc2e),
	.w7(32'h39826cf3),
	.w8(32'h3836220b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f46cc7),
	.w1(32'hb9732173),
	.w2(32'hb8b985da),
	.w3(32'hba39cd20),
	.w4(32'hba68241e),
	.w5(32'h3a07472c),
	.w6(32'hba8b43a7),
	.w7(32'hb9e9601c),
	.w8(32'h39ef4211),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4652fd),
	.w1(32'hb9163ce3),
	.w2(32'h3acfd5aa),
	.w3(32'h3a90ec51),
	.w4(32'h3ac42c24),
	.w5(32'h3b17e1ad),
	.w6(32'h3a948924),
	.w7(32'h3b25dddb),
	.w8(32'h3b22f497),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c7ab9),
	.w1(32'h3b0fbf96),
	.w2(32'h3aae310b),
	.w3(32'h3b18fa8e),
	.w4(32'h3af42dbc),
	.w5(32'h3a466cd8),
	.w6(32'h3ac161f9),
	.w7(32'h3b08134a),
	.w8(32'h3a7d43cb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91c198),
	.w1(32'hb9760a12),
	.w2(32'h3a8b4ffb),
	.w3(32'hb9d1fee3),
	.w4(32'hb964dc5f),
	.w5(32'hba9816ca),
	.w6(32'hba805dd3),
	.w7(32'h38abbd37),
	.w8(32'hb9f333fc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba081bf8),
	.w1(32'hbaafa6b2),
	.w2(32'hbb78e154),
	.w3(32'hba880ffc),
	.w4(32'hbb30d217),
	.w5(32'hba9902bb),
	.w6(32'h3af2a986),
	.w7(32'hbb020a69),
	.w8(32'hba4b8fcf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05a0e8),
	.w1(32'hba364561),
	.w2(32'hba8a8d74),
	.w3(32'hba0d6647),
	.w4(32'hbad36989),
	.w5(32'h39bccb4a),
	.w6(32'hb9095100),
	.w7(32'hbad11a0d),
	.w8(32'h38fb627a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1abc54),
	.w1(32'h3a563cf4),
	.w2(32'h38039841),
	.w3(32'h3a587d9a),
	.w4(32'h39ee3eed),
	.w5(32'hba489a00),
	.w6(32'h39f4829a),
	.w7(32'h3990ad7b),
	.w8(32'h39aabebc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ad312),
	.w1(32'hbaacb990),
	.w2(32'hba3c2ed5),
	.w3(32'hbaa9b0d3),
	.w4(32'hba66bf0c),
	.w5(32'hba987d0f),
	.w6(32'h3a163ad4),
	.w7(32'h397b82db),
	.w8(32'hba1975cc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a6125),
	.w1(32'hbac267a4),
	.w2(32'hba9c4cf2),
	.w3(32'hbadd4ea0),
	.w4(32'hbaac7fa5),
	.w5(32'hb91a30ea),
	.w6(32'hb9e0c031),
	.w7(32'hb9f2d0d7),
	.w8(32'hb7ecb2c3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e684a8),
	.w1(32'h39c48ad5),
	.w2(32'h3aced3e5),
	.w3(32'h39810b35),
	.w4(32'h3a66eee3),
	.w5(32'hbb38e951),
	.w6(32'hb94691c8),
	.w7(32'h3aade22c),
	.w8(32'hbb1ce3bf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb396e5d),
	.w1(32'hbb00055d),
	.w2(32'hbb40aa65),
	.w3(32'hbb2dfd68),
	.w4(32'hbb497ec5),
	.w5(32'hbaa91485),
	.w6(32'hbb127336),
	.w7(32'hbb25195b),
	.w8(32'hbb2e6278),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6dcdb),
	.w1(32'hb9cbf40e),
	.w2(32'hba8714e5),
	.w3(32'hb85d7bcc),
	.w4(32'h38f414d2),
	.w5(32'hbab6606d),
	.w6(32'hbabc8762),
	.w7(32'hb92be6d7),
	.w8(32'hbb14bd9d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eeee4),
	.w1(32'hba95d7cf),
	.w2(32'hbac46dde),
	.w3(32'hbad18aa2),
	.w4(32'hba97ca55),
	.w5(32'h3a0df2aa),
	.w6(32'hbada6ae9),
	.w7(32'hbaff8788),
	.w8(32'hba5032cd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3da05),
	.w1(32'h3a19c984),
	.w2(32'h3ac7ce16),
	.w3(32'h392fe79f),
	.w4(32'h3ae28af0),
	.w5(32'hb9561a71),
	.w6(32'hbaa35861),
	.w7(32'h3a2669af),
	.w8(32'hba0bc8ab),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec2aae),
	.w1(32'hba80ff74),
	.w2(32'hbb03e9aa),
	.w3(32'hba0aaa65),
	.w4(32'hb751c6c3),
	.w5(32'hba93d784),
	.w6(32'hba530588),
	.w7(32'h3984d30d),
	.w8(32'h39dbecd6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3862418e),
	.w1(32'h3a3de321),
	.w2(32'h39f0bdb9),
	.w3(32'hbb29739a),
	.w4(32'hba4c44ed),
	.w5(32'hbb3b126b),
	.w6(32'hbb1e652a),
	.w7(32'hba5392f6),
	.w8(32'hbb4c161f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d24b2),
	.w1(32'hbad83597),
	.w2(32'hbb13c197),
	.w3(32'hbab48fc5),
	.w4(32'hbae846cf),
	.w5(32'h39f36bc7),
	.w6(32'h37b6709e),
	.w7(32'hba9fa341),
	.w8(32'h386b8fc0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6ed49),
	.w1(32'hb9babe0f),
	.w2(32'hb99b3d30),
	.w3(32'hb9b91dc2),
	.w4(32'h38654225),
	.w5(32'h3b3898c1),
	.w6(32'hba1ea4e3),
	.w7(32'h39d7ec8f),
	.w8(32'h3b083709),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf68e5),
	.w1(32'h3858f99c),
	.w2(32'hb9a7b34b),
	.w3(32'h3aa8e698),
	.w4(32'h3a910a1e),
	.w5(32'hb991ca85),
	.w6(32'hba6f0f5b),
	.w7(32'h388b5ecc),
	.w8(32'hba893ce5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad75f8d),
	.w1(32'hbac6a3aa),
	.w2(32'hbab2c2d6),
	.w3(32'hbad97d01),
	.w4(32'hbaba2e81),
	.w5(32'hba47af45),
	.w6(32'hbb17eae3),
	.w7(32'hbab61c3b),
	.w8(32'hba5ed286),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe24f8),
	.w1(32'hbb089089),
	.w2(32'hbb76776d),
	.w3(32'hbb25e242),
	.w4(32'hbafe7a3d),
	.w5(32'hbb53ee62),
	.w6(32'hbb36ae70),
	.w7(32'hbae42ef6),
	.w8(32'hbb78eb99),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f094ed),
	.w1(32'h3847a6d0),
	.w2(32'hb9927722),
	.w3(32'hb9cefed9),
	.w4(32'hbab221b2),
	.w5(32'h39d14aef),
	.w6(32'h396c069e),
	.w7(32'hbac39058),
	.w8(32'hba959425),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7035a8),
	.w1(32'hb9f3668b),
	.w2(32'hb747fd95),
	.w3(32'h3a822e05),
	.w4(32'h3a8d25d9),
	.w5(32'hba8202ea),
	.w6(32'hba9b8457),
	.w7(32'hb9d9f630),
	.w8(32'hba24ffe9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41c196),
	.w1(32'hba2a708f),
	.w2(32'hba235e2f),
	.w3(32'hbab8f509),
	.w4(32'hba9628b8),
	.w5(32'h3a2d40e1),
	.w6(32'hba51e2c2),
	.w7(32'hba2cdb4d),
	.w8(32'h3990905d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66089c),
	.w1(32'h3a4eb734),
	.w2(32'h3b22f50d),
	.w3(32'h39a37269),
	.w4(32'h3b0314f4),
	.w5(32'hb903114e),
	.w6(32'hb988de55),
	.w7(32'h3af9b4bf),
	.w8(32'h39dc7bbe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07247e),
	.w1(32'hbac601ab),
	.w2(32'hba1ccb3c),
	.w3(32'hbb0632a4),
	.w4(32'hba7b6cd5),
	.w5(32'hb91010cf),
	.w6(32'hbaa421af),
	.w7(32'hba9eb3f1),
	.w8(32'hba02c67c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b728e2),
	.w1(32'hb9b2ad9d),
	.w2(32'h3accb5a6),
	.w3(32'hba423a3e),
	.w4(32'h3ac2af8b),
	.w5(32'hb8db70a6),
	.w6(32'hba462fa8),
	.w7(32'h3a6a0f2f),
	.w8(32'hb9e47741),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6104a4),
	.w1(32'hba8d8cec),
	.w2(32'hb9b5f789),
	.w3(32'h37be398e),
	.w4(32'h379b6137),
	.w5(32'h39d3e1e0),
	.w6(32'hb9d676a8),
	.w7(32'hb9855965),
	.w8(32'h3993d6fc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba297687),
	.w1(32'h39527fc9),
	.w2(32'h3acc267d),
	.w3(32'hba8ba291),
	.w4(32'h3ababea2),
	.w5(32'hba9202d3),
	.w6(32'hbab7d914),
	.w7(32'h3aad2c6b),
	.w8(32'hbad5a4bc),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88221ac),
	.w1(32'h39aaf8de),
	.w2(32'h389cd06c),
	.w3(32'h39d804a5),
	.w4(32'h3a4c29b9),
	.w5(32'hb9f77302),
	.w6(32'h396e32d4),
	.w7(32'h393fe2da),
	.w8(32'h38f01072),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c6d73),
	.w1(32'hba29d02f),
	.w2(32'hba1735ca),
	.w3(32'hba78821a),
	.w4(32'hbafd6019),
	.w5(32'h3a877e7f),
	.w6(32'hba2ebe23),
	.w7(32'hbab0559f),
	.w8(32'hba00ff20),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f7c5d),
	.w1(32'h3ab4bb98),
	.w2(32'h3b1d5bf7),
	.w3(32'h3b00bf35),
	.w4(32'h3b611557),
	.w5(32'h38f7abbc),
	.w6(32'hb9f63dcd),
	.w7(32'h3b07e32d),
	.w8(32'hba54d3f3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39898d87),
	.w1(32'h39da9a0b),
	.w2(32'h3a9ee804),
	.w3(32'hb9c5c7f9),
	.w4(32'h3a2668ad),
	.w5(32'h3ad4abab),
	.w6(32'hb9ec6859),
	.w7(32'h3a5e2ae3),
	.w8(32'h3adb4cfc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1de3),
	.w1(32'h3a631302),
	.w2(32'h3b239f28),
	.w3(32'h39bdc711),
	.w4(32'h3ae32bae),
	.w5(32'hba8aede2),
	.w6(32'hb986ce1f),
	.w7(32'h3ab7404b),
	.w8(32'hbab8fc4d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268da5),
	.w1(32'hbb6c81f0),
	.w2(32'hbb2b4caf),
	.w3(32'hbbc5bb75),
	.w4(32'hbbbe18da),
	.w5(32'h3b617725),
	.w6(32'hbba0adf9),
	.w7(32'hbb9c401f),
	.w8(32'hba48cd1c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e0812),
	.w1(32'h3a707f27),
	.w2(32'h3b158f22),
	.w3(32'h3a87b939),
	.w4(32'hb9bd9f7f),
	.w5(32'hbb374929),
	.w6(32'hbaab7085),
	.w7(32'h3a036a0a),
	.w8(32'hba1c1426),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba454689),
	.w1(32'hbb60908a),
	.w2(32'hba8d9d5b),
	.w3(32'hbb8c3c78),
	.w4(32'hbb9157b2),
	.w5(32'h3a8c09f5),
	.w6(32'hbb1d1fe8),
	.w7(32'hb98434f3),
	.w8(32'h3a928392),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48df1a),
	.w1(32'hbb5ae672),
	.w2(32'hbb28b137),
	.w3(32'hbb8469ab),
	.w4(32'hbadd2e8c),
	.w5(32'hba71fc52),
	.w6(32'hbb63da9a),
	.w7(32'hbb132100),
	.w8(32'h37a49678),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0bc9b),
	.w1(32'hb9842731),
	.w2(32'hbaa03a84),
	.w3(32'hba9dbf04),
	.w4(32'hbb2f4eef),
	.w5(32'hba841895),
	.w6(32'hba92831a),
	.w7(32'hbb0b7676),
	.w8(32'hbb1b130a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb75d4),
	.w1(32'hbb0df9d5),
	.w2(32'hbb8a521d),
	.w3(32'hbad64ab0),
	.w4(32'hbba6818c),
	.w5(32'hbace7399),
	.w6(32'h3ae99046),
	.w7(32'hbb241cb5),
	.w8(32'hba7ffd2c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c6f7),
	.w1(32'hbb065409),
	.w2(32'hbae61cea),
	.w3(32'hbaa1b655),
	.w4(32'hba946d72),
	.w5(32'hbace439e),
	.w6(32'hba540b0b),
	.w7(32'hba1f0cf8),
	.w8(32'hbb0f9d44),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dfff1),
	.w1(32'h3b1d3c50),
	.w2(32'hbaab0aff),
	.w3(32'hbb52c6f7),
	.w4(32'hbb01ce07),
	.w5(32'hba3c91fa),
	.w6(32'hbb87d7c0),
	.w7(32'hbb53d80a),
	.w8(32'hbb36621a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76f783),
	.w1(32'hbb24dc3d),
	.w2(32'hbb02c0c8),
	.w3(32'hbb8872c3),
	.w4(32'hbb4f1664),
	.w5(32'h39ec501b),
	.w6(32'hbb86ac6a),
	.w7(32'h389eb178),
	.w8(32'h3b0a46ee),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3cefb),
	.w1(32'h3ab184cc),
	.w2(32'h3b2d10c2),
	.w3(32'hba71aedb),
	.w4(32'hb9552881),
	.w5(32'hba950557),
	.w6(32'hb9acea6f),
	.w7(32'h3a1946b1),
	.w8(32'h3b2bfab6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fbba0),
	.w1(32'h3b39e4cd),
	.w2(32'h3a915954),
	.w3(32'hb99053e1),
	.w4(32'h391261bc),
	.w5(32'h3892c3a5),
	.w6(32'h3b3995e0),
	.w7(32'h3b529463),
	.w8(32'hb98f3b8d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39450825),
	.w1(32'h3a06b6c3),
	.w2(32'h3a9de73f),
	.w3(32'h3a024dda),
	.w4(32'h3b21e399),
	.w5(32'hbae315cd),
	.w6(32'h39744c0c),
	.w7(32'h3b2b8684),
	.w8(32'h3a64515e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964013),
	.w1(32'hba08c1e9),
	.w2(32'hba9c071d),
	.w3(32'hbbb0ce81),
	.w4(32'hbbc57203),
	.w5(32'hbaaebc9a),
	.w6(32'hbb5d1448),
	.w7(32'hbb92a07a),
	.w8(32'hba934fc2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9516e5),
	.w1(32'h3b434360),
	.w2(32'hba690d2e),
	.w3(32'h3b2763d0),
	.w4(32'h3b662a56),
	.w5(32'hbb9bc84b),
	.w6(32'h3b3d0da0),
	.w7(32'h3accd22e),
	.w8(32'hbb82bf82),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed83bb),
	.w1(32'hbb4fa864),
	.w2(32'hbb59badb),
	.w3(32'hbba42a91),
	.w4(32'hbaf8e08c),
	.w5(32'hbb6408a8),
	.w6(32'hbb59098f),
	.w7(32'hbb084895),
	.w8(32'hbad47f32),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a514a2),
	.w1(32'hbab801e2),
	.w2(32'hba41f1e6),
	.w3(32'hbbb24560),
	.w4(32'hbb875ea4),
	.w5(32'hbb14c3b5),
	.w6(32'hbb21cb27),
	.w7(32'hbb2f85bf),
	.w8(32'h3a23ec7f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6fe7f),
	.w1(32'hbac0e71d),
	.w2(32'hb9c1f78e),
	.w3(32'hbb60cc98),
	.w4(32'hbb4942c7),
	.w5(32'h3b82c9f6),
	.w6(32'hbb02308c),
	.w7(32'hbaa63dc8),
	.w8(32'h3b73357b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f042e),
	.w1(32'hba163919),
	.w2(32'h3b2dd3bc),
	.w3(32'h3be0ac88),
	.w4(32'h3bf83e95),
	.w5(32'hbb77aeec),
	.w6(32'h3b36c00f),
	.w7(32'h3baf7093),
	.w8(32'hbb8bc866),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de6c0),
	.w1(32'hbb8a98d2),
	.w2(32'hba9687ea),
	.w3(32'hbad02780),
	.w4(32'hbb5758e4),
	.w5(32'hb988362d),
	.w6(32'h3b20004a),
	.w7(32'h3ab14ee5),
	.w8(32'hba14623e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac96058),
	.w1(32'h388dbae1),
	.w2(32'h3ac82679),
	.w3(32'h3a3b3f79),
	.w4(32'h3ad50ecb),
	.w5(32'hbb850d1f),
	.w6(32'hb9827ea6),
	.w7(32'h3abef85c),
	.w8(32'hbaebd793),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94d2db),
	.w1(32'hbb898295),
	.w2(32'hbaff2c04),
	.w3(32'hbbad72fd),
	.w4(32'hbb364534),
	.w5(32'hbb506727),
	.w6(32'hbbde35ec),
	.w7(32'hbb800d4b),
	.w8(32'hbafe6414),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0d338),
	.w1(32'hbb2c476c),
	.w2(32'hbb69b641),
	.w3(32'h38ee2444),
	.w4(32'hba638a31),
	.w5(32'hbb533460),
	.w6(32'h3aafc6d4),
	.w7(32'hba98ddf0),
	.w8(32'hbb6336b6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb777ea3),
	.w1(32'h3b03333c),
	.w2(32'h3ad03197),
	.w3(32'hba4a6685),
	.w4(32'hbb151c20),
	.w5(32'h3a933bef),
	.w6(32'hbb09bbf7),
	.w7(32'hba240663),
	.w8(32'hba8b8ab4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801268),
	.w1(32'hbb44eae4),
	.w2(32'hbba415e0),
	.w3(32'hbb1cc157),
	.w4(32'hb9d39507),
	.w5(32'hba64acba),
	.w6(32'hb94019a1),
	.w7(32'h3a2ce172),
	.w8(32'hba8fe438),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf5aa5),
	.w1(32'h3a4af9ca),
	.w2(32'hbb57b66d),
	.w3(32'hba2e895c),
	.w4(32'hbb2b1b03),
	.w5(32'hb903909e),
	.w6(32'hbb029498),
	.w7(32'hbb7d607b),
	.w8(32'h3986eae6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec20b0),
	.w1(32'hbb3f1e4c),
	.w2(32'hbb585db9),
	.w3(32'hbaa9766e),
	.w4(32'hb9f28025),
	.w5(32'hbb9d03df),
	.w6(32'h3ab8e1b3),
	.w7(32'h3af0fca1),
	.w8(32'hbb1b3b1f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc8d7f),
	.w1(32'hbb580ae2),
	.w2(32'hbb68d81d),
	.w3(32'hbc008c39),
	.w4(32'hbbfba03a),
	.w5(32'hba28ed45),
	.w6(32'hbbb60f05),
	.w7(32'hbb9f8422),
	.w8(32'hbb38c9dc),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2ddf),
	.w1(32'hbab99a21),
	.w2(32'hb9a6d219),
	.w3(32'hb9e14cb3),
	.w4(32'hbae4f360),
	.w5(32'hb9939dce),
	.w6(32'h3a9cc94e),
	.w7(32'h3a59043a),
	.w8(32'h39c1e69f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06a801),
	.w1(32'hb9c27307),
	.w2(32'h39f70bde),
	.w3(32'hbb28163e),
	.w4(32'hb93bbe8e),
	.w5(32'hb800ad1f),
	.w6(32'hbac15bb0),
	.w7(32'hba5ee0d2),
	.w8(32'h3afa4e23),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule