module layer_8_featuremap_112(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14bfd4),
	.w1(32'hbc2c2655),
	.w2(32'hbc85c10c),
	.w3(32'h3c408f07),
	.w4(32'h3c09db51),
	.w5(32'hbb859ecb),
	.w6(32'hbc651cef),
	.w7(32'hbb980f14),
	.w8(32'hbbb5ff0e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b1f9d),
	.w1(32'hbade6a39),
	.w2(32'hb8055177),
	.w3(32'hbc0766ec),
	.w4(32'h3a8c4001),
	.w5(32'hbb40fd18),
	.w6(32'hbc1b1128),
	.w7(32'hbc3f0038),
	.w8(32'hbc56cd68),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb39c),
	.w1(32'hbc201ea2),
	.w2(32'hbbf65c79),
	.w3(32'hbbd8daf7),
	.w4(32'hbb8be4c4),
	.w5(32'h3a8bbac2),
	.w6(32'hbc43ca9d),
	.w7(32'hbc24bdcc),
	.w8(32'hbc3bd4eb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf2fec),
	.w1(32'hbc368197),
	.w2(32'hbc9bafd8),
	.w3(32'hbc4ff966),
	.w4(32'hbc176d06),
	.w5(32'h3ab002a2),
	.w6(32'hbc19329d),
	.w7(32'hbbef0744),
	.w8(32'h3cc885ae),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc322c44),
	.w1(32'hb9f80ddb),
	.w2(32'hbc95aedb),
	.w3(32'hbb450ed2),
	.w4(32'hbca04153),
	.w5(32'hbc64d860),
	.w6(32'hba1042e1),
	.w7(32'hbc5a3392),
	.w8(32'h3b961b90),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc088d0d),
	.w1(32'h3c6677b3),
	.w2(32'h3c5642db),
	.w3(32'h3a4472de),
	.w4(32'h3bb72d83),
	.w5(32'hbb80634f),
	.w6(32'h3c37225c),
	.w7(32'h3b098e81),
	.w8(32'hbc0a646c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5e4e),
	.w1(32'h3b3d9f14),
	.w2(32'hbb12305c),
	.w3(32'hbb8297aa),
	.w4(32'hb90217a1),
	.w5(32'hbb8162f9),
	.w6(32'hbb9ee9bb),
	.w7(32'h3b4d8dae),
	.w8(32'h3b2c0d84),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b878e),
	.w1(32'hba2bb08f),
	.w2(32'hbbd320c5),
	.w3(32'hbb0e4d8e),
	.w4(32'hbbb5f05e),
	.w5(32'hbc77c3aa),
	.w6(32'hbc2c7d4e),
	.w7(32'hbbc4587f),
	.w8(32'hbbc82e39),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39807d34),
	.w1(32'hbbcdca0b),
	.w2(32'hba8c3408),
	.w3(32'h3a1da259),
	.w4(32'h3ba02b17),
	.w5(32'h3ba23b28),
	.w6(32'hbb922618),
	.w7(32'h3c15e70a),
	.w8(32'h3c74f274),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29f68e),
	.w1(32'hbca053a9),
	.w2(32'hbc96e79f),
	.w3(32'hbb568b6c),
	.w4(32'hba90dc2d),
	.w5(32'hbbff156b),
	.w6(32'hba72da61),
	.w7(32'hbc471698),
	.w8(32'hb9a2f370),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1d56c),
	.w1(32'h3b451115),
	.w2(32'hbbc4882c),
	.w3(32'h3c0803f0),
	.w4(32'hbc75fcce),
	.w5(32'hbcb7cbe5),
	.w6(32'h3b9ca24e),
	.w7(32'h3b0a9794),
	.w8(32'hb9c138db),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89dc99),
	.w1(32'hbc80dc94),
	.w2(32'hbc8856c4),
	.w3(32'hbc87b2a5),
	.w4(32'hbb973078),
	.w5(32'hbc229aa7),
	.w6(32'h3beb0535),
	.w7(32'hbc34cce7),
	.w8(32'hbb976855),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6af6c7),
	.w1(32'hbc261ae4),
	.w2(32'hbb656043),
	.w3(32'h3b8d5fc2),
	.w4(32'hb996213b),
	.w5(32'h3c0d0e6c),
	.w6(32'hbb23d860),
	.w7(32'hbb8b5bd9),
	.w8(32'h3b12ebc4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39442e3f),
	.w1(32'hb9989c52),
	.w2(32'hbb3531ad),
	.w3(32'h3b3d2e95),
	.w4(32'hb98c9619),
	.w5(32'hba3a2da6),
	.w6(32'h3b4a8df0),
	.w7(32'hbb154e36),
	.w8(32'hba8a6664),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd258),
	.w1(32'hba251584),
	.w2(32'hbb27523d),
	.w3(32'hba826fb8),
	.w4(32'hba51ccdc),
	.w5(32'hba85e427),
	.w6(32'h382f5d36),
	.w7(32'hbb0c8635),
	.w8(32'hbada7791),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6a3b),
	.w1(32'hbac47a57),
	.w2(32'hbb24bb59),
	.w3(32'hba458feb),
	.w4(32'hbb6b2363),
	.w5(32'hbbd59dd6),
	.w6(32'hb9ae0b04),
	.w7(32'hbbc06e9d),
	.w8(32'hbbea2a00),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e3ba),
	.w1(32'hbb7adfef),
	.w2(32'hbc9854f5),
	.w3(32'hbb4c464e),
	.w4(32'hbc05a8f1),
	.w5(32'hbc82c669),
	.w6(32'hbb0e034f),
	.w7(32'hbc7a1f7c),
	.w8(32'hbca655cf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c0d4b),
	.w1(32'hbc9bb0f5),
	.w2(32'hbc8081c1),
	.w3(32'hbc477943),
	.w4(32'hbab0b8c8),
	.w5(32'h3ab8cf29),
	.w6(32'hbc551582),
	.w7(32'hbad27224),
	.w8(32'hbb9da258),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0d989),
	.w1(32'hbce7d247),
	.w2(32'hbd4cf051),
	.w3(32'h3c946c0d),
	.w4(32'h3c4e789c),
	.w5(32'hbb6dd1a0),
	.w6(32'h3cc65f4a),
	.w7(32'h3cb9f655),
	.w8(32'h3bf1d022),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd5bb0),
	.w1(32'hbbc73afa),
	.w2(32'hbad90b52),
	.w3(32'h3bfef2ca),
	.w4(32'h3b1f8952),
	.w5(32'h3c030b51),
	.w6(32'hbb96635d),
	.w7(32'hbc512cd8),
	.w8(32'hbbb04dbe),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb5f38),
	.w1(32'hbb8010e2),
	.w2(32'hbbd2f787),
	.w3(32'h39038e93),
	.w4(32'h3c5249f4),
	.w5(32'h3bcbf628),
	.w6(32'h3b0e9b03),
	.w7(32'h3bbb9c50),
	.w8(32'h3be0a03d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132e9b),
	.w1(32'h3c2c87e7),
	.w2(32'hbbe24c6f),
	.w3(32'hbb92b46b),
	.w4(32'hbc21228f),
	.w5(32'hbc05daad),
	.w6(32'hbb6bd222),
	.w7(32'hbc71c5ab),
	.w8(32'hbc538288),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cfda4),
	.w1(32'hbd007899),
	.w2(32'hbd0bbc77),
	.w3(32'h3ce70635),
	.w4(32'h3b7599c2),
	.w5(32'hbbb16dd9),
	.w6(32'h3c71af03),
	.w7(32'h3c6c3be2),
	.w8(32'h3bf2852f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad462ea),
	.w1(32'hbb7868e6),
	.w2(32'h3b03997a),
	.w3(32'h3c1bd0db),
	.w4(32'hbb76e4bc),
	.w5(32'h3bd69dab),
	.w6(32'h3b591fff),
	.w7(32'hbb9208ed),
	.w8(32'h3b69351a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf89246),
	.w1(32'hbb6c8f7c),
	.w2(32'hba84880b),
	.w3(32'h3a4abe69),
	.w4(32'h3bd7fda3),
	.w5(32'hbb26dfc6),
	.w6(32'hbacc00a7),
	.w7(32'h3a64f268),
	.w8(32'hbbed958d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2299e),
	.w1(32'hbbd61dd2),
	.w2(32'hbc894379),
	.w3(32'h3c0d4250),
	.w4(32'hbc612a40),
	.w5(32'hbc512f8a),
	.w6(32'h3c4140ba),
	.w7(32'hbb4a4043),
	.w8(32'hbaf0b19e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb713),
	.w1(32'hbc123396),
	.w2(32'h3bb6381a),
	.w3(32'hbb3c2213),
	.w4(32'hbb4dc15d),
	.w5(32'h3a7f76e2),
	.w6(32'h3b0c4ec3),
	.w7(32'h3b51d724),
	.w8(32'h3b6dbf10),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66e1a6),
	.w1(32'hbd90361f),
	.w2(32'hbcc670ff),
	.w3(32'h3cea9fad),
	.w4(32'hbd5f09ac),
	.w5(32'h3c95eef1),
	.w6(32'h3dbef901),
	.w7(32'h3b422cda),
	.w8(32'h3d425c8e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac6c2f),
	.w1(32'hbb787428),
	.w2(32'hbc8eea67),
	.w3(32'h3cb1caf1),
	.w4(32'hba8d3ebb),
	.w5(32'hbc013f4a),
	.w6(32'h3c699aa7),
	.w7(32'hb8f47ea4),
	.w8(32'hbb159f32),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88476c),
	.w1(32'hba35290d),
	.w2(32'hbbd60aae),
	.w3(32'hb9ce693b),
	.w4(32'hba5f3e19),
	.w5(32'hba750bd3),
	.w6(32'h3a1ff44c),
	.w7(32'hbb9c1db1),
	.w8(32'h3c24e124),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcb95c),
	.w1(32'hbb23e08b),
	.w2(32'hbbb60a1d),
	.w3(32'hbc1f5b61),
	.w4(32'hbae4f054),
	.w5(32'hbb3b6a77),
	.w6(32'h3b730ca8),
	.w7(32'hbab50115),
	.w8(32'hba3c1938),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b128907),
	.w1(32'h3ba9762a),
	.w2(32'h3b379df2),
	.w3(32'h3a97a1bd),
	.w4(32'h3b2136b2),
	.w5(32'hbbc16393),
	.w6(32'h3b598504),
	.w7(32'h3bb9cb67),
	.w8(32'h3aae516f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30a913),
	.w1(32'hbb9d585d),
	.w2(32'hbc985499),
	.w3(32'hbc245e09),
	.w4(32'hbb904d1e),
	.w5(32'hbc859cd1),
	.w6(32'hbc02b224),
	.w7(32'h3b0bcf4f),
	.w8(32'hbbe97d3b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67ddc7),
	.w1(32'hbb1f1512),
	.w2(32'hbb843f41),
	.w3(32'hbc4db2fa),
	.w4(32'h3b68dcd7),
	.w5(32'hba639c93),
	.w6(32'h3b77d7d9),
	.w7(32'hbb43209f),
	.w8(32'hbc22d656),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0eb74),
	.w1(32'hb8cc18ad),
	.w2(32'h3b8fb922),
	.w3(32'hbc8288de),
	.w4(32'hbb213b48),
	.w5(32'h3b9025f2),
	.w6(32'hbcade5cb),
	.w7(32'hbbfdefe6),
	.w8(32'hba6f642e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba314d76),
	.w1(32'hbbe4b2b7),
	.w2(32'hbb90aa7e),
	.w3(32'h3becd6ed),
	.w4(32'h3ab5833d),
	.w5(32'hbb9d7e4d),
	.w6(32'h3c0cea18),
	.w7(32'h3cf11eec),
	.w8(32'h3cc15255),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926fc3),
	.w1(32'h3ba1a662),
	.w2(32'hbc24c623),
	.w3(32'h3ca1d4cc),
	.w4(32'hbb8e5567),
	.w5(32'hbc134953),
	.w6(32'h3cd6be3f),
	.w7(32'h3ab070ff),
	.w8(32'hbbca415f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c1453),
	.w1(32'hbb8a7c34),
	.w2(32'h3b1a4fe3),
	.w3(32'hbc166d13),
	.w4(32'h3be82106),
	.w5(32'hba5f64e2),
	.w6(32'hbb8c5a95),
	.w7(32'h3baba3b7),
	.w8(32'hbb080cb8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f249),
	.w1(32'h3ba56689),
	.w2(32'hbbb7a305),
	.w3(32'hbbc017ef),
	.w4(32'hb855a494),
	.w5(32'hbba10e3d),
	.w6(32'hba990d2d),
	.w7(32'hbbb94ba5),
	.w8(32'hbc5619ec),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dd17c),
	.w1(32'hbbc98e87),
	.w2(32'hbb2ed218),
	.w3(32'hbbb45fcc),
	.w4(32'hb9333639),
	.w5(32'hbb87a125),
	.w6(32'hbc31c4bf),
	.w7(32'hbbfa793d),
	.w8(32'hbc2d71da),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3621),
	.w1(32'hbcb8927e),
	.w2(32'hbc93e3f7),
	.w3(32'h3c6f8926),
	.w4(32'hbc8e7a96),
	.w5(32'h3b841f50),
	.w6(32'hba8e8b33),
	.w7(32'hbc6ba362),
	.w8(32'h3c5886fa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5293),
	.w1(32'hbc0e4e82),
	.w2(32'hbc24ccb6),
	.w3(32'hbba65d68),
	.w4(32'hbc3a3c6e),
	.w5(32'hba538f18),
	.w6(32'h3b69af41),
	.w7(32'hbb99e332),
	.w8(32'h3b7467ec),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb129b98),
	.w1(32'hbc88b5df),
	.w2(32'h39fe07c4),
	.w3(32'h3aa4a2b2),
	.w4(32'h3a437584),
	.w5(32'hb93f503e),
	.w6(32'h3b47aa26),
	.w7(32'h3a72a73a),
	.w8(32'h3b4d0404),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcc4ae),
	.w1(32'h3c3ca165),
	.w2(32'hbbdd281f),
	.w3(32'h3c7f470a),
	.w4(32'h3b51e8d9),
	.w5(32'h3bc3e3a7),
	.w6(32'h3c647783),
	.w7(32'h3b1df34c),
	.w8(32'h3becccb1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa56ef),
	.w1(32'hbc00c266),
	.w2(32'hbcc2026f),
	.w3(32'h3c88e0bf),
	.w4(32'h39db9958),
	.w5(32'hbc47b756),
	.w6(32'h3c7b6c2d),
	.w7(32'h3b701dcc),
	.w8(32'hb9551962),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba299af),
	.w1(32'hbc0b0778),
	.w2(32'hbcaab081),
	.w3(32'h39dc4e76),
	.w4(32'hbc94c531),
	.w5(32'hbc33d048),
	.w6(32'h3ae4fb60),
	.w7(32'hbb553aa5),
	.w8(32'h3ac83957),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a4c44),
	.w1(32'hbc96dcf6),
	.w2(32'hbbef431c),
	.w3(32'h38ca60e7),
	.w4(32'hbaa4ad6d),
	.w5(32'h3b6d3ee1),
	.w6(32'hbb9b0520),
	.w7(32'hbc21d156),
	.w8(32'hbb36bb64),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb274791),
	.w1(32'hbab09e2c),
	.w2(32'hbca8ef7d),
	.w3(32'h3c31a793),
	.w4(32'hbb9a13e8),
	.w5(32'hbc6c216f),
	.w6(32'h3c0fefd6),
	.w7(32'h3b0b8074),
	.w8(32'hbbcb2976),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c9cff),
	.w1(32'hbc3cbf0e),
	.w2(32'hbbb74616),
	.w3(32'h3a097522),
	.w4(32'hba09f1b6),
	.w5(32'hbb5cabeb),
	.w6(32'h3abf6de2),
	.w7(32'h3baa3e5b),
	.w8(32'h39022cb4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dd6aa),
	.w1(32'hbc564529),
	.w2(32'hbccb3008),
	.w3(32'hbbb2ff41),
	.w4(32'hbb65a6a6),
	.w5(32'hbc6a675d),
	.w6(32'h3c43f8d9),
	.w7(32'hbb8e8d51),
	.w8(32'hbc42ab9c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc866628),
	.w1(32'hbc11a5ef),
	.w2(32'h3b75feed),
	.w3(32'hbc54b960),
	.w4(32'hbc56f66a),
	.w5(32'h3c0dde4d),
	.w6(32'hbc837e35),
	.w7(32'hbb01063f),
	.w8(32'h3c78d0e1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f00ac),
	.w1(32'hbd026619),
	.w2(32'hbd3c312c),
	.w3(32'h3caeed38),
	.w4(32'hbcda4b17),
	.w5(32'hbd302d40),
	.w6(32'h3cf59fec),
	.w7(32'hbc9e2aca),
	.w8(32'hbcb2c1d0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f3422),
	.w1(32'hbc666742),
	.w2(32'hba867596),
	.w3(32'hbca4d45a),
	.w4(32'h3a959b6b),
	.w5(32'hbb92b235),
	.w6(32'hbca7456c),
	.w7(32'h3b314fb7),
	.w8(32'hbb1c6770),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc421d18),
	.w1(32'hbc8b7e84),
	.w2(32'hbcc9e017),
	.w3(32'h3c4b9fe3),
	.w4(32'h3c767764),
	.w5(32'h3bc3ee54),
	.w6(32'hbb0a15e9),
	.w7(32'h3b79ae64),
	.w8(32'hbad57eef),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972b03a),
	.w1(32'h39179e72),
	.w2(32'hba8ee092),
	.w3(32'h3b0ccd36),
	.w4(32'hbc181ca3),
	.w5(32'hbb671e16),
	.w6(32'h3b0f5ee6),
	.w7(32'hba9db748),
	.w8(32'hbb123bb8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcf70f),
	.w1(32'hbc5c6548),
	.w2(32'hbd05e4e9),
	.w3(32'h3cd52c5d),
	.w4(32'h3ca29de2),
	.w5(32'h3c088414),
	.w6(32'h3be2ad76),
	.w7(32'h3c4f850b),
	.w8(32'h3c0efc33),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1886c5),
	.w1(32'hbc0cfaee),
	.w2(32'hbb9d036e),
	.w3(32'h3bb36a88),
	.w4(32'h3bc72002),
	.w5(32'h3b65822b),
	.w6(32'h39f72794),
	.w7(32'hbb03a75b),
	.w8(32'hbc1f4914),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2caadc),
	.w1(32'hbc25c414),
	.w2(32'hbb2864d6),
	.w3(32'h3b7e4bc6),
	.w4(32'hbbbb98eb),
	.w5(32'h3c2ea46e),
	.w6(32'h3be0ca34),
	.w7(32'h3a6231b3),
	.w8(32'h3cc4e969),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe84c4),
	.w1(32'h3c0e2b8d),
	.w2(32'hbbd1d7d0),
	.w3(32'h3cfcbed7),
	.w4(32'h3aab7062),
	.w5(32'h3b65136f),
	.w6(32'h3cba7bea),
	.w7(32'h3b213c81),
	.w8(32'h3af857fb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb548a3d),
	.w1(32'hbadf7ee1),
	.w2(32'h3adbcef5),
	.w3(32'h3c15cc38),
	.w4(32'h3b6acd9b),
	.w5(32'hbbec1261),
	.w6(32'h3bb12c38),
	.w7(32'h3bbf822e),
	.w8(32'hb9d14513),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff04cf),
	.w1(32'h3bbbc4f3),
	.w2(32'h3bacd4ee),
	.w3(32'hbbc4a8b4),
	.w4(32'hbc4626aa),
	.w5(32'h3b778643),
	.w6(32'hbb70be94),
	.w7(32'h3a00500b),
	.w8(32'h3c6bc8d6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbba4f8),
	.w1(32'h3ba872e3),
	.w2(32'hba2016eb),
	.w3(32'h3babe7af),
	.w4(32'hb9470b8b),
	.w5(32'hbabaef68),
	.w6(32'h3c4e96f9),
	.w7(32'hba1f48a7),
	.w8(32'hbb2cd805),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8903),
	.w1(32'hbccb3fb5),
	.w2(32'hbc95451a),
	.w3(32'h3c3299e7),
	.w4(32'hba9ef38b),
	.w5(32'h3b5dfe4f),
	.w6(32'h3be142b9),
	.w7(32'h3a9efdf9),
	.w8(32'h3c31b0f8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32afe2),
	.w1(32'hb947db39),
	.w2(32'hba6c1c34),
	.w3(32'hbb333453),
	.w4(32'h3aaa2861),
	.w5(32'hbaaf1696),
	.w6(32'hbb8e2152),
	.w7(32'hbb2f93b9),
	.w8(32'hbb216496),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a902a),
	.w1(32'h3b6345b1),
	.w2(32'hbb463935),
	.w3(32'hba4ddd01),
	.w4(32'hbb718eb4),
	.w5(32'hbb80d2d4),
	.w6(32'hb8a4e4c4),
	.w7(32'hbbb93544),
	.w8(32'hbbdb84c0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8909),
	.w1(32'hbc11c41b),
	.w2(32'hbbe9ec29),
	.w3(32'hbb2e2847),
	.w4(32'hbb1a0890),
	.w5(32'hbb977fc1),
	.w6(32'hbbb7ed6c),
	.w7(32'hba77fedf),
	.w8(32'hbbaf637b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc2550),
	.w1(32'hbaff2d32),
	.w2(32'h3b09abf7),
	.w3(32'h3b273e9f),
	.w4(32'h3a1d0179),
	.w5(32'hba810a90),
	.w6(32'hba3db565),
	.w7(32'h3ae8603d),
	.w8(32'hbb833f93),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb96b85),
	.w1(32'hbc083567),
	.w2(32'hbc68de2e),
	.w3(32'hb925dcd7),
	.w4(32'hbbb0a12a),
	.w5(32'hbc0e75b6),
	.w6(32'hbab8291f),
	.w7(32'h3bac2368),
	.w8(32'h39ff7030),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8a71b),
	.w1(32'hbbd5f9e5),
	.w2(32'hbc37d30f),
	.w3(32'hbc2a37b0),
	.w4(32'hbb7fa0e2),
	.w5(32'hbb804e9a),
	.w6(32'hbc14ccf9),
	.w7(32'hbb66ff4d),
	.w8(32'hbbb2a308),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15a695),
	.w1(32'h3bc7f8bf),
	.w2(32'hbbec8124),
	.w3(32'h3c8a76c6),
	.w4(32'h3c976135),
	.w5(32'hbb6a0b62),
	.w6(32'h3c297a1c),
	.w7(32'h3c86d07d),
	.w8(32'h3bb07374),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1986a3),
	.w1(32'h3c678581),
	.w2(32'h399f5383),
	.w3(32'hb9710c39),
	.w4(32'hbb0aef51),
	.w5(32'h39c35891),
	.w6(32'h3c4cf6ae),
	.w7(32'h3acbafab),
	.w8(32'h3bd35895),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8487aaf),
	.w1(32'hbbfb1527),
	.w2(32'hbc4f0c73),
	.w3(32'h3b3f30e8),
	.w4(32'hbc6aa237),
	.w5(32'hbca0cb49),
	.w6(32'h3bd7d833),
	.w7(32'hbbe43886),
	.w8(32'hbc28a093),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e599cc),
	.w1(32'h3ad0d7d8),
	.w2(32'hbb419318),
	.w3(32'hbc0d21d4),
	.w4(32'hbb40e0ed),
	.w5(32'hbb830036),
	.w6(32'h3adfc6a7),
	.w7(32'hbb9703be),
	.w8(32'hbbde4159),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38ebf4),
	.w1(32'hbca0d6d2),
	.w2(32'hbc26b102),
	.w3(32'hba422849),
	.w4(32'h3bfbf429),
	.w5(32'h3c446e31),
	.w6(32'hbb77d892),
	.w7(32'h3c1b2604),
	.w8(32'h3c6e9bca),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a2302),
	.w1(32'h3b8b0cdf),
	.w2(32'hbc04c384),
	.w3(32'h3aa549b0),
	.w4(32'hbb6bff4b),
	.w5(32'hbb44c381),
	.w6(32'h3ad2e9b8),
	.w7(32'hbb138586),
	.w8(32'h3b7a40bb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034d23),
	.w1(32'hbc26e326),
	.w2(32'hbc593171),
	.w3(32'hbc007cc0),
	.w4(32'hbc108f6e),
	.w5(32'hbc6f3118),
	.w6(32'h3a48c8dc),
	.w7(32'hbbdb52ed),
	.w8(32'hbc1e6c4e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc063a7f),
	.w1(32'hbb3ac3b5),
	.w2(32'h37c1a2eb),
	.w3(32'hbb18b79f),
	.w4(32'h37763cec),
	.w5(32'h38076505),
	.w6(32'hb9d1b053),
	.w7(32'h388284e1),
	.w8(32'h38818560),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f626f),
	.w1(32'hbbbaf821),
	.w2(32'hbc71b055),
	.w3(32'h3c27db2e),
	.w4(32'hbb039723),
	.w5(32'hbbc447d9),
	.w6(32'h3c0613af),
	.w7(32'h3bd861d3),
	.w8(32'h3ac19baf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e75f4),
	.w1(32'hbc5289e8),
	.w2(32'hbc904734),
	.w3(32'h3bd52f9e),
	.w4(32'hbb499728),
	.w5(32'hbb94c646),
	.w6(32'h3c23dd03),
	.w7(32'h3b54a5c1),
	.w8(32'h3a53b114),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973449e),
	.w1(32'h39863eab),
	.w2(32'h3998e584),
	.w3(32'h38fb1968),
	.w4(32'h392c3f16),
	.w5(32'h39b9dc95),
	.w6(32'h38428840),
	.w7(32'hb6a68008),
	.w8(32'h39817aaf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6908f29),
	.w1(32'h376449d2),
	.w2(32'hb664133e),
	.w3(32'h387e6d3b),
	.w4(32'h38e21b25),
	.w5(32'h386e4e56),
	.w6(32'h38a6447c),
	.w7(32'h390e0964),
	.w8(32'h390a34ae),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6737),
	.w1(32'hbb86306c),
	.w2(32'hbb3cb904),
	.w3(32'h3bd557f0),
	.w4(32'h3b9853d4),
	.w5(32'hbb5b4ff6),
	.w6(32'h3ba87b35),
	.w7(32'h3ac063e8),
	.w8(32'hbbdd43ce),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc16856),
	.w1(32'hbb69f981),
	.w2(32'hbc08f37b),
	.w3(32'h3c6a9308),
	.w4(32'h3b98511e),
	.w5(32'h3b415631),
	.w6(32'h3c4618b1),
	.w7(32'h3bf5176a),
	.w8(32'h3bd9471c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc372090),
	.w1(32'hbd1e1f8a),
	.w2(32'hbcfcd15d),
	.w3(32'h3be589b9),
	.w4(32'hbcda5a29),
	.w5(32'hba5ec23e),
	.w6(32'hb9daf05d),
	.w7(32'hbbeb54fd),
	.w8(32'h3c57a2d5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e6174),
	.w1(32'hbc6e5ff9),
	.w2(32'hbcb4421f),
	.w3(32'h3ce999d5),
	.w4(32'h3c29e69e),
	.w5(32'h3ae022e8),
	.w6(32'h3caa1446),
	.w7(32'h3c84f99e),
	.w8(32'h3c94d6ef),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17051),
	.w1(32'hbc34b9ec),
	.w2(32'hbb849dd6),
	.w3(32'h3b3ca3b0),
	.w4(32'hbb0fe2b5),
	.w5(32'hb9c6eb81),
	.w6(32'h3ac4f484),
	.w7(32'hbaf42629),
	.w8(32'hbb67530e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c63122),
	.w1(32'h37da7672),
	.w2(32'hb8a7f0e8),
	.w3(32'hb9cb0b35),
	.w4(32'hb809b21a),
	.w5(32'hb88e44d4),
	.w6(32'hb9b91cbf),
	.w7(32'hb9478fa6),
	.w8(32'hb933146e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e58427),
	.w1(32'hb7ca8645),
	.w2(32'hb7cac8a1),
	.w3(32'hb80b3140),
	.w4(32'h37fad78c),
	.w5(32'h37fc7837),
	.w6(32'hb67d3402),
	.w7(32'h386ced41),
	.w8(32'h37c240e9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c2cab),
	.w1(32'hb8baab5b),
	.w2(32'h381eeb1a),
	.w3(32'hb9372d2e),
	.w4(32'hb98dcfa1),
	.w5(32'hb93ee97d),
	.w6(32'hb94224a7),
	.w7(32'hb97f02dd),
	.w8(32'hb910db4c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d6d8f),
	.w1(32'h3ab27e8e),
	.w2(32'h3a040510),
	.w3(32'h3ab5f688),
	.w4(32'h3a83db74),
	.w5(32'hb812f939),
	.w6(32'h3ac08851),
	.w7(32'h3aa55a99),
	.w8(32'hb8de421e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1698),
	.w1(32'hbc0076df),
	.w2(32'hbb46379a),
	.w3(32'h3bd8ac31),
	.w4(32'h39fbb3d3),
	.w5(32'h3a5e0b6a),
	.w6(32'h3b784078),
	.w7(32'hba879df0),
	.w8(32'hb9b86803),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39814b23),
	.w1(32'h3768dd64),
	.w2(32'hb92e56e9),
	.w3(32'h38be9e02),
	.w4(32'hb82a93e4),
	.w5(32'hb95b2c09),
	.w6(32'h3a3a7b1f),
	.w7(32'h3985fc6c),
	.w8(32'h39c18f04),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e62fe),
	.w1(32'hba353eed),
	.w2(32'h3b50d902),
	.w3(32'h3aec94b1),
	.w4(32'h39bceef4),
	.w5(32'h3b530b3d),
	.w6(32'hba95f7b1),
	.w7(32'hbb90ca20),
	.w8(32'hbb314377),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0f29c),
	.w1(32'hbbe0eabe),
	.w2(32'hbbf76ad2),
	.w3(32'h3ba2abce),
	.w4(32'hba9f8d3d),
	.w5(32'hbb0c95a2),
	.w6(32'h3b9c57da),
	.w7(32'h3952d3c6),
	.w8(32'h3a4db1be),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a5e36),
	.w1(32'hbb1b0c34),
	.w2(32'hbb7955ba),
	.w3(32'h3b909b43),
	.w4(32'h3b161959),
	.w5(32'h3a6ef805),
	.w6(32'h3a52a7d3),
	.w7(32'h39b9fb82),
	.w8(32'h3b3a3df3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea7f9f),
	.w1(32'hbb62aa34),
	.w2(32'hbc41716b),
	.w3(32'h3c1777b1),
	.w4(32'h3b59e34c),
	.w5(32'hbbe082b3),
	.w6(32'h3c04f11d),
	.w7(32'h3b78e9c4),
	.w8(32'hbb94813a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce89a1),
	.w1(32'hbc077062),
	.w2(32'hbc1a4c06),
	.w3(32'h3bc02a01),
	.w4(32'hbb4621a3),
	.w5(32'hbba36baa),
	.w6(32'h3c2ae94e),
	.w7(32'h3b98cff1),
	.w8(32'h3a81ea75),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f52f3),
	.w1(32'hb7df17e0),
	.w2(32'hb8b51d03),
	.w3(32'h3924e3d0),
	.w4(32'h39250706),
	.w5(32'hb79208fd),
	.w6(32'hb5b82968),
	.w7(32'h38eb176e),
	.w8(32'hb8a52183),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b372fa),
	.w1(32'h39027380),
	.w2(32'h38f685a7),
	.w3(32'hb88fcbbb),
	.w4(32'h3860dc7e),
	.w5(32'h3825322a),
	.w6(32'hb939c9b6),
	.w7(32'hb868a61e),
	.w8(32'hb89af364),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917f226),
	.w1(32'h378f3568),
	.w2(32'h38a96ade),
	.w3(32'hb8bb33d2),
	.w4(32'h38db4efe),
	.w5(32'h38b47752),
	.w6(32'hb922ee44),
	.w7(32'h381d2c78),
	.w8(32'hb8a74090),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fecb22),
	.w1(32'h3a28e7f2),
	.w2(32'h3a2ff4a2),
	.w3(32'h39989667),
	.w4(32'h39de7eed),
	.w5(32'h3a086c82),
	.w6(32'h39c9ce3f),
	.w7(32'h39ebed67),
	.w8(32'h39e49011),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01c974),
	.w1(32'h39cad20a),
	.w2(32'h3abd4d1e),
	.w3(32'h3ab3d7bd),
	.w4(32'h3b0976d3),
	.w5(32'h3af2072a),
	.w6(32'h3a4b36d4),
	.w7(32'h3a81b0c2),
	.w8(32'hb8bcb2c5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb9142),
	.w1(32'h3a4265ea),
	.w2(32'h3a7d3b97),
	.w3(32'h3aab367c),
	.w4(32'h3a4ae071),
	.w5(32'h3a0d1e49),
	.w6(32'h3abeca1a),
	.w7(32'h39fc73c2),
	.w8(32'hb735c7b5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a7692),
	.w1(32'hbb2c0cba),
	.w2(32'h3bad0d67),
	.w3(32'h3ad55848),
	.w4(32'h3a7df9a7),
	.w5(32'h3bc285d0),
	.w6(32'hbb87ef8b),
	.w7(32'hbb586506),
	.w8(32'hbb140a30),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7794ae),
	.w1(32'hb9c0e3fe),
	.w2(32'h3ab06b6b),
	.w3(32'hbb17e7b3),
	.w4(32'hbad92109),
	.w5(32'h39993bb3),
	.w6(32'hbb2c3c17),
	.w7(32'hbb219dc4),
	.w8(32'hba58d77d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f276),
	.w1(32'hbb03df65),
	.w2(32'hbbeefde9),
	.w3(32'h3c608f91),
	.w4(32'h3b8d84b9),
	.w5(32'hbb2cd4cc),
	.w6(32'h3c63a60e),
	.w7(32'h3c2477a4),
	.w8(32'h3bcbbcdd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a984dfc),
	.w1(32'h3a48a5b8),
	.w2(32'h3a1c3675),
	.w3(32'h3a5c4776),
	.w4(32'h39bbb567),
	.w5(32'h39a63944),
	.w6(32'h3aa47819),
	.w7(32'h3a82fc48),
	.w8(32'h3a23bf50),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab538d1),
	.w1(32'h3ac6cd3e),
	.w2(32'h3afc3890),
	.w3(32'hbb63be77),
	.w4(32'hba47ef2b),
	.w5(32'hb95e116b),
	.w6(32'hbb66a6d0),
	.w7(32'hbb38fa63),
	.w8(32'hbb09316d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a6306),
	.w1(32'h382d6f5a),
	.w2(32'h3a04d46a),
	.w3(32'hbad849e7),
	.w4(32'hba2d5144),
	.w5(32'h3613d676),
	.w6(32'hbacbfb06),
	.w7(32'hba8dcfbb),
	.w8(32'hba562b25),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68cc5),
	.w1(32'hbacea025),
	.w2(32'hba6ab63e),
	.w3(32'hb9412bc1),
	.w4(32'hbaa25438),
	.w5(32'hb90df510),
	.w6(32'hb9783e1b),
	.w7(32'h3a39da84),
	.w8(32'hb9bd6e93),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab75a9),
	.w1(32'hbb8d9001),
	.w2(32'hbb9725b7),
	.w3(32'h3b3b66c8),
	.w4(32'hb8a70708),
	.w5(32'h3a8f93c9),
	.w6(32'h3b0214b8),
	.w7(32'h3ae95ab0),
	.w8(32'h3aefe0de),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c4f0),
	.w1(32'hbb19888a),
	.w2(32'hbb0b7112),
	.w3(32'hb9c21917),
	.w4(32'hbb068b79),
	.w5(32'h3a3cf63c),
	.w6(32'h3b2cb46e),
	.w7(32'h3a255013),
	.w8(32'h3b364f6c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a149),
	.w1(32'hba2d0700),
	.w2(32'h3b04cf2b),
	.w3(32'hbb8d70ff),
	.w4(32'hbb048936),
	.w5(32'h3a2318b5),
	.w6(32'hbbb8c15f),
	.w7(32'hbb699501),
	.w8(32'hba4b1b70),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab2ba5),
	.w1(32'h36eebd38),
	.w2(32'h3947874e),
	.w3(32'hb85930b7),
	.w4(32'h38b918c9),
	.w5(32'h398380fd),
	.w6(32'hb8870dc4),
	.w7(32'h3991aeb7),
	.w8(32'h39ab20ec),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad65841),
	.w1(32'hbb81b6b2),
	.w2(32'hbbd007b4),
	.w3(32'hbb112d1b),
	.w4(32'hbb4a0437),
	.w5(32'hbba4793e),
	.w6(32'hba7461b8),
	.w7(32'hbb2dabf5),
	.w8(32'hbb375046),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e8668),
	.w1(32'h396426ea),
	.w2(32'h39122a9d),
	.w3(32'h39d12ce4),
	.w4(32'h38510e5e),
	.w5(32'hb8331aab),
	.w6(32'h3a5ff0ae),
	.w7(32'h39e19ae1),
	.w8(32'h39a1f396),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4b004),
	.w1(32'hbb44b2f3),
	.w2(32'hbb545550),
	.w3(32'h39650f40),
	.w4(32'hbb189804),
	.w5(32'hbb64edf9),
	.w6(32'h392b7c03),
	.w7(32'hbb01500c),
	.w8(32'hbb58a48b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a4aa0),
	.w1(32'hba85f582),
	.w2(32'hbbe5cc4c),
	.w3(32'h3c033196),
	.w4(32'h3b35f07d),
	.w5(32'hba95be69),
	.w6(32'h3bea6fe0),
	.w7(32'h3b859dc4),
	.w8(32'h3b9aec2e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83474d9),
	.w1(32'h37304dd0),
	.w2(32'hb62a22f5),
	.w3(32'hb896f02e),
	.w4(32'hb68fda67),
	.w5(32'h378117cc),
	.w6(32'hb8a6b643),
	.w7(32'hb7fee37a),
	.w8(32'h37996471),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8130b),
	.w1(32'hba1fca31),
	.w2(32'hbadb9c5e),
	.w3(32'h3b0abbec),
	.w4(32'h3a1b61cf),
	.w5(32'hb9c3fbb5),
	.w6(32'h3ae8a4a2),
	.w7(32'h3a2537ea),
	.w8(32'h3a0bc244),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f8d4),
	.w1(32'hbbf3ef14),
	.w2(32'hbb9ffdc6),
	.w3(32'h3c481275),
	.w4(32'h3c0ab334),
	.w5(32'h3bb705d3),
	.w6(32'hbaddad51),
	.w7(32'hbbd2a375),
	.w8(32'hbbea3986),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf121a2),
	.w1(32'hbbbc6c30),
	.w2(32'hbb20475a),
	.w3(32'hbb8759cb),
	.w4(32'hbb9aa022),
	.w5(32'hba72735d),
	.w6(32'hb6fe9c34),
	.w7(32'h3a96dbb7),
	.w8(32'h3b140ef3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84cc785),
	.w1(32'h390edd34),
	.w2(32'hb78da35e),
	.w3(32'hb99062b7),
	.w4(32'h384198a3),
	.w5(32'h3974b7ba),
	.w6(32'hb8cd14c9),
	.w7(32'h3904d602),
	.w8(32'h38bc0206),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8423c7),
	.w1(32'hba2789e0),
	.w2(32'hb9df8f91),
	.w3(32'hba87b055),
	.w4(32'hb9e9beff),
	.w5(32'hb9baeb21),
	.w6(32'hbac2d60f),
	.w7(32'hba902c01),
	.w8(32'hba8be905),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6b78),
	.w1(32'h3a4fb9c7),
	.w2(32'h3a846b78),
	.w3(32'h3a2de40f),
	.w4(32'h3a30e892),
	.w5(32'h3a51cfc6),
	.w6(32'h3a7db364),
	.w7(32'h3a33d0f2),
	.w8(32'h3a24f027),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca1dfc),
	.w1(32'h3b7b4e38),
	.w2(32'hbb167400),
	.w3(32'h3b81c615),
	.w4(32'h3bd51a10),
	.w5(32'h3a3f4dc3),
	.w6(32'h3b7b14d3),
	.w7(32'h3b8cc0a8),
	.w8(32'h39feb8de),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6f34),
	.w1(32'hbbd59afd),
	.w2(32'hbbdf7296),
	.w3(32'h3b71bfdf),
	.w4(32'hba388f1a),
	.w5(32'hbaa3bb46),
	.w6(32'h3aef224b),
	.w7(32'hba54e665),
	.w8(32'hb854c4f6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b9d8),
	.w1(32'h3ae1a030),
	.w2(32'hbbf7deb3),
	.w3(32'h3b6d252f),
	.w4(32'h3b245583),
	.w5(32'hbc0ed479),
	.w6(32'h3bab0d3b),
	.w7(32'h3acb5ad6),
	.w8(32'hbbbbd521),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule