module layer_10_featuremap_199(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990901d),
	.w1(32'h3ac02c1b),
	.w2(32'h3aef3eb8),
	.w3(32'hb95bf39b),
	.w4(32'h3b2bfe51),
	.w5(32'h3a80002e),
	.w6(32'h3a377d24),
	.w7(32'h3ad5df11),
	.w8(32'hba26591a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf8702),
	.w1(32'hba3065e1),
	.w2(32'h3985e9cc),
	.w3(32'h3b571221),
	.w4(32'hbb63c7dc),
	.w5(32'hbb72d5c0),
	.w6(32'h3b47c182),
	.w7(32'h39505b64),
	.w8(32'hba251755),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352a7682),
	.w1(32'hb9913e05),
	.w2(32'h3a824679),
	.w3(32'hb9ba37ac),
	.w4(32'h397db176),
	.w5(32'hb9caf887),
	.w6(32'hba5a95cf),
	.w7(32'hba0c1ade),
	.w8(32'hb9af3335),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985f95),
	.w1(32'hbb0dcd48),
	.w2(32'hbb4aa758),
	.w3(32'hba2e7806),
	.w4(32'hbae50d05),
	.w5(32'hba4c0ce5),
	.w6(32'h3b0213c2),
	.w7(32'h3b149338),
	.w8(32'h3b2b1284),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f310),
	.w1(32'h3a38ca43),
	.w2(32'h37e903b4),
	.w3(32'hba82c838),
	.w4(32'h3a85dafa),
	.w5(32'h3a83d0cc),
	.w6(32'h3a1f210a),
	.w7(32'hb934c26d),
	.w8(32'hb90a5b56),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a673a93),
	.w1(32'h3aa0293c),
	.w2(32'h39d5990f),
	.w3(32'h3a38532e),
	.w4(32'h3a883c23),
	.w5(32'h3a610f8b),
	.w6(32'h3951dc69),
	.w7(32'hb8b0f28d),
	.w8(32'hba2b069a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93215b),
	.w1(32'h3a20f1a8),
	.w2(32'h3b44e211),
	.w3(32'h3a4e501a),
	.w4(32'h3b175377),
	.w5(32'h3b823706),
	.w6(32'h3a633383),
	.w7(32'h3b2c5262),
	.w8(32'h3b1b6890),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7e89),
	.w1(32'h3b874465),
	.w2(32'h3b486da3),
	.w3(32'h3b60daa6),
	.w4(32'h3bee1f17),
	.w5(32'h3b871cca),
	.w6(32'h3b31bbf1),
	.w7(32'h3b6e4233),
	.w8(32'h3b222beb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7745a3),
	.w1(32'h3a833348),
	.w2(32'h3aa0e925),
	.w3(32'h38cb53e4),
	.w4(32'hb926c135),
	.w5(32'h3a05ed71),
	.w6(32'h3ac87db5),
	.w7(32'h3a2fbc43),
	.w8(32'h3a8ebe5f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe935d4),
	.w1(32'hbac478ec),
	.w2(32'h3c81b6f7),
	.w3(32'hbb4688b3),
	.w4(32'h3ac7a6bd),
	.w5(32'h3c815743),
	.w6(32'h3b976ded),
	.w7(32'h3beb3045),
	.w8(32'h3c5b9447),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af69156),
	.w1(32'h3ad33267),
	.w2(32'h3b6dbda5),
	.w3(32'h3ae401c7),
	.w4(32'hb9e52a2e),
	.w5(32'h3acb9e01),
	.w6(32'h3a234f27),
	.w7(32'hbae60503),
	.w8(32'hb9cee907),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba35bb),
	.w1(32'hbad562c5),
	.w2(32'h3c2bd059),
	.w3(32'hbaa98c58),
	.w4(32'h3ae41b42),
	.w5(32'h3c5533f9),
	.w6(32'h3adefebe),
	.w7(32'h3b361155),
	.w8(32'h3c28582c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf38026),
	.w1(32'hbb35e2ca),
	.w2(32'h3c6d8564),
	.w3(32'hbb39760f),
	.w4(32'h3b225fe8),
	.w5(32'h3c99136d),
	.w6(32'hbafcb370),
	.w7(32'h3b93f166),
	.w8(32'h3c663486),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d627),
	.w1(32'hbb911442),
	.w2(32'h3a5f512f),
	.w3(32'hbb107599),
	.w4(32'hbb784442),
	.w5(32'h3a5f373c),
	.w6(32'hbaeb7d7a),
	.w7(32'hbb816a72),
	.w8(32'hba7f1b5d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fb602),
	.w1(32'hbb04a482),
	.w2(32'hb94abae8),
	.w3(32'hbb6a69eb),
	.w4(32'hbb832297),
	.w5(32'hb6407bba),
	.w6(32'h3bb73e83),
	.w7(32'h3b98acdb),
	.w8(32'h3b6c2d58),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb980a0b),
	.w1(32'hbaee8bc3),
	.w2(32'h3bc63eb9),
	.w3(32'hbb400d7c),
	.w4(32'hbad388b0),
	.w5(32'h3baed2cb),
	.w6(32'h3aeb684d),
	.w7(32'h3b450d6e),
	.w8(32'h3c174622),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c6944),
	.w1(32'hbb0493ee),
	.w2(32'h3a8a25a3),
	.w3(32'h38d9b4a3),
	.w4(32'hbac481fb),
	.w5(32'hbac28dd6),
	.w6(32'hba731009),
	.w7(32'hbb58a960),
	.w8(32'hba92a63f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e0d83),
	.w1(32'hbaa0412a),
	.w2(32'h3bf43df3),
	.w3(32'hbbb0b7a3),
	.w4(32'h3b16f080),
	.w5(32'h3c49c669),
	.w6(32'h3c02cc89),
	.w7(32'h3c1bec70),
	.w8(32'h3c1936ff),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba914c55),
	.w1(32'hbb1d0128),
	.w2(32'h3bdc177c),
	.w3(32'hbba53bed),
	.w4(32'hb9e96ec8),
	.w5(32'h3be4b701),
	.w6(32'h3afca1b5),
	.w7(32'h3bac5d2a),
	.w8(32'h3ba9ed00),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b42c83),
	.w1(32'h3a15c720),
	.w2(32'h3a0da36e),
	.w3(32'hba09358c),
	.w4(32'hb9157969),
	.w5(32'hb9d2c492),
	.w6(32'h3a1683ce),
	.w7(32'h39e50186),
	.w8(32'h3948450b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923217a),
	.w1(32'hbadf9c55),
	.w2(32'hbab8e143),
	.w3(32'hb9a03eea),
	.w4(32'hbadbd090),
	.w5(32'hbaedd4ca),
	.w6(32'hbb09aca3),
	.w7(32'hbaddde9a),
	.w8(32'hbb249c8e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb726bcb),
	.w1(32'hba077211),
	.w2(32'h3bc9b4a5),
	.w3(32'hbba2e0e6),
	.w4(32'h383c4ef0),
	.w5(32'h3b1b7be3),
	.w6(32'hba1ac344),
	.w7(32'h3abcf184),
	.w8(32'h3b689d2e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34f32e),
	.w1(32'h3b9f979a),
	.w2(32'h3cc3bcb6),
	.w3(32'hbb80dfc1),
	.w4(32'hbbb05a4f),
	.w5(32'h3cb0a9c4),
	.w6(32'h3c7c1426),
	.w7(32'h3ca17888),
	.w8(32'h3d0b4cda),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5a66),
	.w1(32'hbb814160),
	.w2(32'h3c3ceb5f),
	.w3(32'hbbc9bfbd),
	.w4(32'hbbd6ccfd),
	.w5(32'h3bf82988),
	.w6(32'h3b169474),
	.w7(32'h3ab010ff),
	.w8(32'h3c33de7c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39521957),
	.w1(32'hba755cb8),
	.w2(32'h3c13f52f),
	.w3(32'hbb6f6a32),
	.w4(32'hbbc11f5e),
	.w5(32'h3b17e092),
	.w6(32'h3c153fbb),
	.w7(32'h3c02df72),
	.w8(32'h3c745fbd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20f368),
	.w1(32'h37ae706b),
	.w2(32'h3ab3b772),
	.w3(32'hba8b208b),
	.w4(32'hb9d78bd5),
	.w5(32'h3a873422),
	.w6(32'h38327cae),
	.w7(32'hb82c5f7d),
	.w8(32'h3a0dd108),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a323b05),
	.w1(32'h39d40485),
	.w2(32'h39510320),
	.w3(32'hbae5f779),
	.w4(32'hb9bc6cb9),
	.w5(32'hba52f7c2),
	.w6(32'hb8195504),
	.w7(32'hb8cb100e),
	.w8(32'hba39a5d1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4454),
	.w1(32'hba04e98e),
	.w2(32'h3ada9646),
	.w3(32'hbba4dd55),
	.w4(32'hba845036),
	.w5(32'hba3fc4c0),
	.w6(32'hb9a810cf),
	.w7(32'h3b7249b7),
	.w8(32'h3b64125f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb32a),
	.w1(32'hbb02d012),
	.w2(32'h3c2d7954),
	.w3(32'hbc0f02ee),
	.w4(32'hbbc09cd2),
	.w5(32'h3be4b0e2),
	.w6(32'hbc0330cd),
	.w7(32'hbb3ebdd1),
	.w8(32'h3bae23ce),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52684),
	.w1(32'hbc01be56),
	.w2(32'h3b0b2c97),
	.w3(32'hbbdbffc3),
	.w4(32'hbbff80b8),
	.w5(32'h38ab6a38),
	.w6(32'hbb05f1c1),
	.w7(32'hbb02f3de),
	.w8(32'h3bd38e85),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32f42a),
	.w1(32'hba5eeaa3),
	.w2(32'hb9e43f2c),
	.w3(32'h38d9330d),
	.w4(32'hba769880),
	.w5(32'hba861fac),
	.w6(32'hba90764a),
	.w7(32'hbaa7f5a1),
	.w8(32'hbad0e71e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c6c4b),
	.w1(32'hba05d822),
	.w2(32'h390ae435),
	.w3(32'hbaac73ff),
	.w4(32'hbaa5ec50),
	.w5(32'hb9fd09be),
	.w6(32'hba3cb58d),
	.w7(32'hba8ccc61),
	.w8(32'hba784c49),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee00c2),
	.w1(32'hbaff7f7d),
	.w2(32'h3b975254),
	.w3(32'hbb2ed800),
	.w4(32'hbb567439),
	.w5(32'h3afc4f7a),
	.w6(32'h3ac25512),
	.w7(32'h3aada6c2),
	.w8(32'h3b9dc9cf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c2c7),
	.w1(32'h3b27c65e),
	.w2(32'h3bced1c7),
	.w3(32'h38f805f4),
	.w4(32'h3a0fc5ef),
	.w5(32'h3b9e1cfc),
	.w6(32'h3ad4eb3b),
	.w7(32'h3b851a0a),
	.w8(32'h3b96eff0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ea864),
	.w1(32'h3a9928e2),
	.w2(32'h3af80515),
	.w3(32'h39b462cb),
	.w4(32'h3ac4f217),
	.w5(32'h3b75babb),
	.w6(32'hb815f3b3),
	.w7(32'h3a759bf2),
	.w8(32'h3acb7e14),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0dab2),
	.w1(32'h3aadc507),
	.w2(32'h3b10b0c9),
	.w3(32'h3a5ad76e),
	.w4(32'h3990ef59),
	.w5(32'h3b02cc8c),
	.w6(32'h3a18a0d0),
	.w7(32'h3a4de501),
	.w8(32'h3a7e8e82),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0011d0),
	.w1(32'hbae71844),
	.w2(32'h3c0095c6),
	.w3(32'h3ac3712a),
	.w4(32'hbbb223db),
	.w5(32'h3b5cf41d),
	.w6(32'h3b0f6f62),
	.w7(32'h3a0a40c3),
	.w8(32'h3bd9cd11),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1ce71),
	.w1(32'h39c2fa84),
	.w2(32'h3c478875),
	.w3(32'hbc14c118),
	.w4(32'hbc4ccbc6),
	.w5(32'hbbbbd2d6),
	.w6(32'h3c0a8824),
	.w7(32'h3a9470d5),
	.w8(32'h3c30579b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb28d),
	.w1(32'h3b683fed),
	.w2(32'h3cb87103),
	.w3(32'hbc4c5764),
	.w4(32'hbb8e5345),
	.w5(32'h3c7227cf),
	.w6(32'h3b359e01),
	.w7(32'h3ba2a6c1),
	.w8(32'h3ccb959e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39c092),
	.w1(32'hbac9fb5e),
	.w2(32'hbb455e1b),
	.w3(32'h39943542),
	.w4(32'hbb509000),
	.w5(32'hbbaea601),
	.w6(32'h3b75c25d),
	.w7(32'hb8b4b62e),
	.w8(32'hbb1f8eab),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b04b0),
	.w1(32'hb9907d3f),
	.w2(32'hbac02218),
	.w3(32'h3a77db4b),
	.w4(32'hb9f79a9a),
	.w5(32'hbaea3b3f),
	.w6(32'hb8bde48e),
	.w7(32'hba50c033),
	.w8(32'hba2f9a77),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38d8fd),
	.w1(32'hbac8b125),
	.w2(32'hba2bb012),
	.w3(32'hbaa262e0),
	.w4(32'hbad5397b),
	.w5(32'hbafefbb1),
	.w6(32'hb9860dfd),
	.w7(32'hb90b6bfd),
	.w8(32'hba962ed5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ebbc),
	.w1(32'hbbf5f283),
	.w2(32'h3ab4a846),
	.w3(32'hbba71ddf),
	.w4(32'hbbd0df2d),
	.w5(32'h3b9eab5f),
	.w6(32'hbb70d68e),
	.w7(32'hbbd7f29c),
	.w8(32'h3b69157f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01927e),
	.w1(32'hbba634eb),
	.w2(32'h3c1c894f),
	.w3(32'hbc59c16d),
	.w4(32'hbb5301de),
	.w5(32'h3c515a75),
	.w6(32'hb82e77d5),
	.w7(32'h3b929320),
	.w8(32'h3c5097e3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64c6ab),
	.w1(32'hbae6e40f),
	.w2(32'h3c407629),
	.w3(32'hbb12a300),
	.w4(32'hbbbeb97d),
	.w5(32'h3ba37898),
	.w6(32'h3b75e75e),
	.w7(32'h3b0df73c),
	.w8(32'h3c4a349f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33270e),
	.w1(32'hba160bcb),
	.w2(32'h3c66145c),
	.w3(32'hbbaac5fe),
	.w4(32'hbbb886d6),
	.w5(32'h3c0a7087),
	.w6(32'h3bcad73c),
	.w7(32'h3be26372),
	.w8(32'h3c8927f1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1b994),
	.w1(32'h3b47bab5),
	.w2(32'h3bb30de3),
	.w3(32'h3b6b1d1d),
	.w4(32'h39d34d59),
	.w5(32'h3bee0f2d),
	.w6(32'h3c553501),
	.w7(32'h3c123fbd),
	.w8(32'h3c343453),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afad19c),
	.w1(32'h3b69f834),
	.w2(32'h3c8ef577),
	.w3(32'h3aabad6d),
	.w4(32'h3c09a599),
	.w5(32'h3cc3bfa5),
	.w6(32'h3b946bd0),
	.w7(32'h3c4d691b),
	.w8(32'h3c8aab2f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add4b4e),
	.w1(32'h3949d103),
	.w2(32'h39d23adc),
	.w3(32'hba766fbe),
	.w4(32'hb9dae136),
	.w5(32'h38d1bcdc),
	.w6(32'hba6bb9c2),
	.w7(32'hb8207c58),
	.w8(32'hb7637c45),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f4dfb),
	.w1(32'hbae9c8a5),
	.w2(32'hbabeaeb0),
	.w3(32'h39ded539),
	.w4(32'hb9a3b8e8),
	.w5(32'hb983db08),
	.w6(32'hbac917af),
	.w7(32'hba784c42),
	.w8(32'hba17926d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dfa2b),
	.w1(32'hba2a7eff),
	.w2(32'h3a5d05bc),
	.w3(32'hbb4f9def),
	.w4(32'h398c9063),
	.w5(32'h3a8c1685),
	.w6(32'hbb0e8d6a),
	.w7(32'hb95ca7dd),
	.w8(32'h390a9591),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff2260),
	.w1(32'h3b30ce18),
	.w2(32'h3bd3192c),
	.w3(32'hbb20e029),
	.w4(32'h39d901d7),
	.w5(32'h3be50619),
	.w6(32'h3b76db4c),
	.w7(32'h3b0c3b4e),
	.w8(32'h3bda3dc2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39909008),
	.w1(32'h3b0eea6d),
	.w2(32'h3b01d757),
	.w3(32'hba160d63),
	.w4(32'h3abf65af),
	.w5(32'h3abfef1a),
	.w6(32'h3b0fc22c),
	.w7(32'h3b0c8281),
	.w8(32'h3ad23079),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd523f8),
	.w1(32'hba91a504),
	.w2(32'h3ba04882),
	.w3(32'hbb6c68e5),
	.w4(32'h3b246996),
	.w5(32'h3bf22bfe),
	.w6(32'h3bdbc95b),
	.w7(32'h3c0cc227),
	.w8(32'h3bd6a91e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbef6b),
	.w1(32'h3b0e40e2),
	.w2(32'h3b11a497),
	.w3(32'hb8bd8bdf),
	.w4(32'h382d84be),
	.w5(32'h3a9ff50c),
	.w6(32'h3a63d924),
	.w7(32'h3ae8cdbd),
	.w8(32'h3b17e689),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2f885),
	.w1(32'hbaf5c478),
	.w2(32'hb9af2e73),
	.w3(32'hb9ec843c),
	.w4(32'hbab7f3eb),
	.w5(32'hbabd7cfd),
	.w6(32'hbab56fc5),
	.w7(32'hbb0bd4ec),
	.w8(32'hba58a832),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66923b),
	.w1(32'hb9b69466),
	.w2(32'hbafab680),
	.w3(32'hba63c3a5),
	.w4(32'hba2a041a),
	.w5(32'hbaf8de26),
	.w6(32'hba42803a),
	.w7(32'hba896eab),
	.w8(32'hba95f709),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a87ef),
	.w1(32'h38c3e406),
	.w2(32'hb9e11c4e),
	.w3(32'hbabd8a09),
	.w4(32'h3aa3caef),
	.w5(32'h3a9dc561),
	.w6(32'h3a1ace88),
	.w7(32'h39bcf511),
	.w8(32'hba10511e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91021d),
	.w1(32'hbb2225ca),
	.w2(32'h3ab5a2b9),
	.w3(32'hba20baeb),
	.w4(32'hbb18b5bb),
	.w5(32'h3a16b543),
	.w6(32'hb9b0cde8),
	.w7(32'hbae5aac3),
	.w8(32'h3a806928),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2abfbb),
	.w1(32'hbb0e5dbe),
	.w2(32'hba7a5a7f),
	.w3(32'hba4aea33),
	.w4(32'hbb2faf9f),
	.w5(32'hbaa5b904),
	.w6(32'hba166fea),
	.w7(32'hbb1cf4d8),
	.w8(32'hbacd3063),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb447),
	.w1(32'hbb144425),
	.w2(32'h3a5f38ff),
	.w3(32'hbbdb0332),
	.w4(32'hbb5919c3),
	.w5(32'h3b54b562),
	.w6(32'hbb3ffce4),
	.w7(32'hbad18c38),
	.w8(32'h3b7eed71),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199534),
	.w1(32'h3845300a),
	.w2(32'h3b3095df),
	.w3(32'hba48255f),
	.w4(32'h3978b5b9),
	.w5(32'h3b34765b),
	.w6(32'h3b0a91de),
	.w7(32'h3a1bef77),
	.w8(32'h3ad1245d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba753c9c),
	.w1(32'h39665fcf),
	.w2(32'hba3533b7),
	.w3(32'hbaa815df),
	.w4(32'h3a2af0ff),
	.w5(32'hbaadb155),
	.w6(32'h3ac5bd67),
	.w7(32'hba92deb6),
	.w8(32'h3a841a20),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1b86b),
	.w1(32'h3a2ea8e5),
	.w2(32'h3a6361d7),
	.w3(32'hb7354c8f),
	.w4(32'h3aff1c81),
	.w5(32'h3b02d277),
	.w6(32'h399c5e6c),
	.w7(32'h3a867253),
	.w8(32'h3965cf4b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bf66f),
	.w1(32'hba82d07a),
	.w2(32'hba38f700),
	.w3(32'h3ad8bf9a),
	.w4(32'hbb001502),
	.w5(32'hba8e0eab),
	.w6(32'hba2cf173),
	.w7(32'hb9171cbc),
	.w8(32'hba9dba06),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd7f6),
	.w1(32'hbaac7c0a),
	.w2(32'hba1559ec),
	.w3(32'hb9a70245),
	.w4(32'hb91d05f6),
	.w5(32'h39972166),
	.w6(32'hba2865fe),
	.w7(32'hb99638d6),
	.w8(32'hba7b437a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa41b8),
	.w1(32'hbb98d2a0),
	.w2(32'hbb9edbbd),
	.w3(32'h3b872fbb),
	.w4(32'h3aa12e6b),
	.w5(32'hb9df0202),
	.w6(32'h3b877824),
	.w7(32'h3b5d6e0d),
	.w8(32'h3b01052d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a877e6d),
	.w1(32'h3b834247),
	.w2(32'h3c82bc52),
	.w3(32'hbbeb3c42),
	.w4(32'hbbca70b3),
	.w5(32'h3c1772aa),
	.w6(32'h3be9b0a9),
	.w7(32'h3bd37201),
	.w8(32'h3c95b9e3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e7b5c),
	.w1(32'h3bed691b),
	.w2(32'h3c8ccad0),
	.w3(32'hbb755b21),
	.w4(32'hb9b53566),
	.w5(32'h3c353f29),
	.w6(32'h3c181a47),
	.w7(32'h3bf65fb1),
	.w8(32'h3c827e0c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba398e44),
	.w1(32'h39b5b32c),
	.w2(32'h3ca39304),
	.w3(32'hbba892cf),
	.w4(32'hbbbf0550),
	.w5(32'h3c381c52),
	.w6(32'h3c3f5892),
	.w7(32'h3c3153d9),
	.w8(32'h3cbba7e2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35b9c5),
	.w1(32'h39809b9d),
	.w2(32'hb90414f1),
	.w3(32'h3a00a8d5),
	.w4(32'h38f43ff4),
	.w5(32'hb989351c),
	.w6(32'hb92e7b30),
	.w7(32'h38bbd36c),
	.w8(32'hba4b4ae4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390698ca),
	.w1(32'hb9b7a210),
	.w2(32'hba60b88f),
	.w3(32'hb9def062),
	.w4(32'hb988a847),
	.w5(32'hba68dc51),
	.w6(32'hb9c79295),
	.w7(32'hba20297a),
	.w8(32'hbac0eef4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aae0d),
	.w1(32'hba05694d),
	.w2(32'hba8c8136),
	.w3(32'hba7411e3),
	.w4(32'hb9c5d971),
	.w5(32'hba77f392),
	.w6(32'hb9ce62a4),
	.w7(32'hba350f51),
	.w8(32'hbac46407),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6dc16),
	.w1(32'hbab79d06),
	.w2(32'h3a198663),
	.w3(32'hba96bedf),
	.w4(32'hb8fe8fb8),
	.w5(32'h3ae43c48),
	.w6(32'h3892aa90),
	.w7(32'h3a1f40f9),
	.w8(32'h3a278d63),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba288e30),
	.w1(32'hba8081b2),
	.w2(32'hba4291fa),
	.w3(32'hba8eecd8),
	.w4(32'hba41f8a0),
	.w5(32'hba609226),
	.w6(32'hb8dd341c),
	.w7(32'h39ae96a2),
	.w8(32'hba193eeb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57fd2a),
	.w1(32'hb9a12e62),
	.w2(32'hbba788c2),
	.w3(32'h39e42164),
	.w4(32'h3ada26fd),
	.w5(32'h3ae3f280),
	.w6(32'h3b5d2420),
	.w7(32'h3b5a0796),
	.w8(32'hbb061783),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61996e),
	.w1(32'hbb51cb25),
	.w2(32'h3b9c1d8a),
	.w3(32'hbbd0aadf),
	.w4(32'hbb80535b),
	.w5(32'h3b84e9ee),
	.w6(32'h3955aaf3),
	.w7(32'hb933f4d1),
	.w8(32'h3b81bf6f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51ab7f),
	.w1(32'h3ae157d3),
	.w2(32'h3c2b7ad6),
	.w3(32'hbafacc80),
	.w4(32'h3b105099),
	.w5(32'h3c1b1bcf),
	.w6(32'hba322f5d),
	.w7(32'h3b861434),
	.w8(32'h3c411f30),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50a829),
	.w1(32'h3aa7830c),
	.w2(32'h3b540607),
	.w3(32'hbb57fda5),
	.w4(32'hba9d9fa0),
	.w5(32'h3b5e9e0f),
	.w6(32'h3b0899ec),
	.w7(32'h3a878dcd),
	.w8(32'h3bdb5b76),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd1150),
	.w1(32'hbb864c19),
	.w2(32'hb932ef3e),
	.w3(32'h3a037a89),
	.w4(32'hbb2cee07),
	.w5(32'h3acc5719),
	.w6(32'hbaf32326),
	.w7(32'hb97fecaf),
	.w8(32'h3a6dbfe3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587b67),
	.w1(32'hba7672ab),
	.w2(32'h3bc4108f),
	.w3(32'hbb7bb778),
	.w4(32'hbb1381fa),
	.w5(32'h3b873cc6),
	.w6(32'hbacf2b5e),
	.w7(32'hba761646),
	.w8(32'h3baa2601),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada1085),
	.w1(32'h3a155f0e),
	.w2(32'h3bdaefd4),
	.w3(32'hba105820),
	.w4(32'h3a098aa3),
	.w5(32'h3bd9c86f),
	.w6(32'h3a5948ab),
	.w7(32'h3b186c77),
	.w8(32'h3bb754a3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16c580),
	.w1(32'hb95671b7),
	.w2(32'h3a132bb6),
	.w3(32'h3a343578),
	.w4(32'hba4357a0),
	.w5(32'hba125519),
	.w6(32'hb9875cfc),
	.w7(32'hb9a129fa),
	.w8(32'hba330b27),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef6719),
	.w1(32'hb9dfc139),
	.w2(32'h39205bb0),
	.w3(32'hba9a4d0b),
	.w4(32'hba2c7515),
	.w5(32'hba657dcd),
	.w6(32'hb8037698),
	.w7(32'h3991fae5),
	.w8(32'h368b0314),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96128d),
	.w1(32'h3a10a276),
	.w2(32'h3ad01469),
	.w3(32'h392d0c10),
	.w4(32'hba972b56),
	.w5(32'hb8f7e9f1),
	.w6(32'hba5e20f7),
	.w7(32'hba9daea7),
	.w8(32'hb8caa347),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69af39),
	.w1(32'hba6946ab),
	.w2(32'hba5a64e9),
	.w3(32'hb8e072c8),
	.w4(32'hba05db28),
	.w5(32'hba1b1ba9),
	.w6(32'hb8244f7d),
	.w7(32'hba109213),
	.w8(32'hb9a25f0e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2e98),
	.w1(32'hbab3e6f8),
	.w2(32'hbae73348),
	.w3(32'h3a63392f),
	.w4(32'hbba58ad2),
	.w5(32'hbbd737b2),
	.w6(32'h3c026ca7),
	.w7(32'hba8cf5b6),
	.w8(32'h39f46b35),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898c4ce),
	.w1(32'hbb536b1a),
	.w2(32'h3a34cfaa),
	.w3(32'hb989f3e9),
	.w4(32'hbb444f34),
	.w5(32'h393de4e2),
	.w6(32'hb812ae38),
	.w7(32'hbb107e4f),
	.w8(32'h39dd0ac3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2ece),
	.w1(32'hbab0aa68),
	.w2(32'h3a93dda4),
	.w3(32'hbb2c3a14),
	.w4(32'hbbc1ad66),
	.w5(32'hbb5e4c3a),
	.w6(32'h3b959356),
	.w7(32'h3a91648a),
	.w8(32'hba200ecb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecb416),
	.w1(32'hba92a8c8),
	.w2(32'h3b6e8afa),
	.w3(32'hba1a5081),
	.w4(32'hbb1ed5d8),
	.w5(32'h3b86f72f),
	.w6(32'h3be0edce),
	.w7(32'h3b82e37d),
	.w8(32'h3bf06c6c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886e2e),
	.w1(32'hbb09fb89),
	.w2(32'h3b4fc97f),
	.w3(32'hbbd1b11d),
	.w4(32'hbb9f9297),
	.w5(32'hb4d39ae0),
	.w6(32'hba0a6c02),
	.w7(32'hbad14290),
	.w8(32'h3b5d9fef),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c854f),
	.w1(32'h3aca8ff0),
	.w2(32'h3bb215da),
	.w3(32'hbae32350),
	.w4(32'hbb221a80),
	.w5(32'h3ae9c935),
	.w6(32'h398d173a),
	.w7(32'h395ad6a4),
	.w8(32'h3b98fb66),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba910c2a),
	.w1(32'hbb9af959),
	.w2(32'h3a9b739c),
	.w3(32'hbae5e132),
	.w4(32'hbbf0de6a),
	.w5(32'hbb1cacc0),
	.w6(32'h3b2207c9),
	.w7(32'hbad3b44a),
	.w8(32'h3abec544),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6ce7),
	.w1(32'hbb28450b),
	.w2(32'h3b4b75f1),
	.w3(32'hbba9e817),
	.w4(32'hbbbcc48e),
	.w5(32'hbb068a51),
	.w6(32'h3b58c5bc),
	.w7(32'h3a9b6441),
	.w8(32'h3b4218b6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0827f7),
	.w1(32'hbb37302f),
	.w2(32'hbb02986d),
	.w3(32'hb8e091f6),
	.w4(32'hbb891381),
	.w5(32'hbbb86995),
	.w6(32'h3bbb5a9b),
	.w7(32'h37f26d3f),
	.w8(32'hbaee79ee),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee1519),
	.w1(32'hbaeeaf27),
	.w2(32'h3a80bb82),
	.w3(32'hbb8a5128),
	.w4(32'hbbc0cf66),
	.w5(32'hbb76300d),
	.w6(32'h3bd93e87),
	.w7(32'h3a59250f),
	.w8(32'h3abbe6d1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d343e6),
	.w1(32'hbb50ced1),
	.w2(32'hba9a1c1d),
	.w3(32'hbacb3c34),
	.w4(32'hbb836059),
	.w5(32'hbb16d3ca),
	.w6(32'hbb19b20e),
	.w7(32'hbb2d64d6),
	.w8(32'hbb33f5e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba94cd1),
	.w1(32'hbb54e17c),
	.w2(32'h3c20d448),
	.w3(32'hbb9a294c),
	.w4(32'hba2880f9),
	.w5(32'h3c255719),
	.w6(32'h3b8e6d1f),
	.w7(32'h3c0e5950),
	.w8(32'h3c6abf05),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbecf0),
	.w1(32'hbadf188c),
	.w2(32'h3ae96d6a),
	.w3(32'h3bb39edf),
	.w4(32'hb98a2c6d),
	.w5(32'h3ba8c51d),
	.w6(32'h3c52c623),
	.w7(32'h3c2821e8),
	.w8(32'h3c3e1f21),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be23c71),
	.w1(32'h3ae82d50),
	.w2(32'h3be7f62a),
	.w3(32'h3b88c37f),
	.w4(32'h3b904e89),
	.w5(32'h3c05caa5),
	.w6(32'h3c39cae5),
	.w7(32'h3c22fb47),
	.w8(32'h3c5b484d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c171ae8),
	.w1(32'h3bd61629),
	.w2(32'h3c1a2499),
	.w3(32'hb9db9b3c),
	.w4(32'hbbca9929),
	.w5(32'hbb513db7),
	.w6(32'h3c69c5e3),
	.w7(32'h3b83e1e0),
	.w8(32'h3c26c0fd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a0d9),
	.w1(32'hbbdd1f2d),
	.w2(32'h3bba7a0a),
	.w3(32'hbbd44496),
	.w4(32'hbafedbba),
	.w5(32'h3c006e13),
	.w6(32'h3b1e86fc),
	.w7(32'h3b43db92),
	.w8(32'h3c44ce6d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ebda),
	.w1(32'h3ab12133),
	.w2(32'h3bc0c503),
	.w3(32'h3ba689f8),
	.w4(32'h3971b69a),
	.w5(32'h3b907c27),
	.w6(32'h3babede8),
	.w7(32'h3b645cbf),
	.w8(32'h3aeb1546),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c1e60),
	.w1(32'hba16b57a),
	.w2(32'hba05aa9b),
	.w3(32'hbb383d08),
	.w4(32'hba1f8b70),
	.w5(32'hba07cf6b),
	.w6(32'hba9bd9de),
	.w7(32'hbac743db),
	.w8(32'hbb1dd0a2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc4dda),
	.w1(32'h3b688089),
	.w2(32'h3b9d88bf),
	.w3(32'h3b87370d),
	.w4(32'hba475bba),
	.w5(32'h3b4d5a71),
	.w6(32'h3bb0a639),
	.w7(32'h3b63dd88),
	.w8(32'h3baf10a9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca95b),
	.w1(32'hba9cb9e3),
	.w2(32'h3b29a797),
	.w3(32'hba516053),
	.w4(32'h3b1608d6),
	.w5(32'h3b989c0a),
	.w6(32'hbafe190d),
	.w7(32'h3b2f7832),
	.w8(32'h3bc724e7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924db9c),
	.w1(32'hb95698c2),
	.w2(32'h3ae13614),
	.w3(32'hba5072d6),
	.w4(32'hba4302d8),
	.w5(32'hb8cde1ed),
	.w6(32'hba1cd65e),
	.w7(32'hb9e8cb79),
	.w8(32'h38b987f6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20cbfc),
	.w1(32'hba1c3222),
	.w2(32'h38027a9f),
	.w3(32'h39d298c0),
	.w4(32'hba692e14),
	.w5(32'hba73c4dc),
	.w6(32'hb89b8ecf),
	.w7(32'hbaa99361),
	.w8(32'hba9f0247),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06237f),
	.w1(32'hbb9be84d),
	.w2(32'h3b8acfff),
	.w3(32'hbc24d57f),
	.w4(32'hbacbfaca),
	.w5(32'h3c004d99),
	.w6(32'hbba851fe),
	.w7(32'h3a875465),
	.w8(32'h3bb95ad4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf917c2),
	.w1(32'hbbcc1d67),
	.w2(32'h3b7b48fe),
	.w3(32'hbc0d8ce0),
	.w4(32'hbbc5c51b),
	.w5(32'h3b403372),
	.w6(32'hbb3d21c7),
	.w7(32'hba18e2c2),
	.w8(32'h3bf0e35b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cecc6),
	.w1(32'h39979fdd),
	.w2(32'h3af6b583),
	.w3(32'hba75566d),
	.w4(32'hbaee6ccf),
	.w5(32'hba5177f3),
	.w6(32'h3b8004e9),
	.w7(32'h3b9be2e5),
	.w8(32'h3b561d3a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70927c),
	.w1(32'h3aca51e1),
	.w2(32'hb9cb9d52),
	.w3(32'hbad25e5b),
	.w4(32'h381c9fb9),
	.w5(32'h3b09767a),
	.w6(32'h3bbdbe35),
	.w7(32'h3b5fa6e7),
	.w8(32'h3bfd9aa3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd93dd5),
	.w1(32'h3b89ecca),
	.w2(32'h3c1d60b5),
	.w3(32'h39b96823),
	.w4(32'hbabb83e3),
	.w5(32'h3b841b91),
	.w6(32'h3b056b5d),
	.w7(32'h3a62a1fa),
	.w8(32'h3be5e6fd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba715474),
	.w1(32'hbad25783),
	.w2(32'h3b4d7518),
	.w3(32'hbb21fdc6),
	.w4(32'hbb25fa4d),
	.w5(32'h39f29ac9),
	.w6(32'hb849a999),
	.w7(32'hb89e62f5),
	.w8(32'h3b703a86),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c619e),
	.w1(32'hbb2c5191),
	.w2(32'h3b45cae2),
	.w3(32'hbb7c61fe),
	.w4(32'hbb5a3c63),
	.w5(32'h3b1fa483),
	.w6(32'hb9f6e3d2),
	.w7(32'h390ddf47),
	.w8(32'h3ba0c9c2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94703ab),
	.w1(32'hba6c200f),
	.w2(32'hba7f0a1e),
	.w3(32'hba9e9e96),
	.w4(32'hb99ac7e1),
	.w5(32'hb9ee95ba),
	.w6(32'hbab98b3a),
	.w7(32'hbad358fb),
	.w8(32'hbb24b8d2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffd9d3),
	.w1(32'h3927dabc),
	.w2(32'hb9e5ac22),
	.w3(32'hbab3d8b3),
	.w4(32'hb91f5805),
	.w5(32'hb9d3e23e),
	.w6(32'hb9572e61),
	.w7(32'hba2412bc),
	.w8(32'hba70dacc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c53a5),
	.w1(32'hb8f9483a),
	.w2(32'hb9401954),
	.w3(32'hb82d85da),
	.w4(32'h3962f300),
	.w5(32'hb81590a7),
	.w6(32'hb891377e),
	.w7(32'hba354ca1),
	.w8(32'hba81b143),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba122f15),
	.w1(32'h3a933fad),
	.w2(32'h3ae64b89),
	.w3(32'hba19d7fb),
	.w4(32'h3afd11f7),
	.w5(32'h3ab2a767),
	.w6(32'h3a36c8b1),
	.w7(32'h3a866720),
	.w8(32'h3a60783a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3a598),
	.w1(32'hbb878b11),
	.w2(32'h3be29b08),
	.w3(32'hbb0ce681),
	.w4(32'hbba986cd),
	.w5(32'h3b85a8d0),
	.w6(32'hb7d7c6d5),
	.w7(32'hba1ccbd0),
	.w8(32'h3bbd7ab7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38634839),
	.w1(32'h3b1264d9),
	.w2(32'h3b331235),
	.w3(32'hba9750f1),
	.w4(32'h3a62b5b3),
	.w5(32'h3aaea44a),
	.w6(32'h3abe70a4),
	.w7(32'h3a94282e),
	.w8(32'h3a903856),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3a5b),
	.w1(32'h3b1aa17d),
	.w2(32'h3baad9aa),
	.w3(32'h3a900473),
	.w4(32'h3b430074),
	.w5(32'h3b36ce25),
	.w6(32'h3b5deb4e),
	.w7(32'h3b995a92),
	.w8(32'h3b62b8f4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238f13),
	.w1(32'hba875bd2),
	.w2(32'h3b155f33),
	.w3(32'hbb12e157),
	.w4(32'hbb327aea),
	.w5(32'hb92362c9),
	.w6(32'h3b8d9ab8),
	.w7(32'h3b3336c7),
	.w8(32'h3bd0f3a2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab58031),
	.w1(32'h3ae5df0e),
	.w2(32'h3b1f72da),
	.w3(32'hbab56102),
	.w4(32'h3b8858cd),
	.w5(32'h3b009c80),
	.w6(32'h3aac7bf2),
	.w7(32'h3b10feca),
	.w8(32'h3b0c2457),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeac4cd),
	.w1(32'h3b160994),
	.w2(32'h3adaa040),
	.w3(32'h3b3d0b86),
	.w4(32'h3abf19e3),
	.w5(32'h3a955f54),
	.w6(32'h39ca69f8),
	.w7(32'h39fa803b),
	.w8(32'h39f4e652),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a392ce),
	.w1(32'hba5af8be),
	.w2(32'hba82c943),
	.w3(32'h39e77257),
	.w4(32'hba9e41ea),
	.w5(32'hbabe360f),
	.w6(32'hbab1ca22),
	.w7(32'hbaf14f59),
	.w8(32'hbad0daa2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975ab48),
	.w1(32'h39832292),
	.w2(32'hba26f2c9),
	.w3(32'hba019451),
	.w4(32'h3aa75921),
	.w5(32'hb97d95f6),
	.w6(32'h3b228174),
	.w7(32'h3a478fee),
	.w8(32'h39ec3bd6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60a9b0),
	.w1(32'h3b738133),
	.w2(32'h3c0444ce),
	.w3(32'hbb393410),
	.w4(32'h39253335),
	.w5(32'h3be85704),
	.w6(32'h3a86b577),
	.w7(32'h3abf821c),
	.w8(32'h3bd52128),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef467a),
	.w1(32'hbbfbb3a1),
	.w2(32'hb9e07625),
	.w3(32'hbba3fe8a),
	.w4(32'hbb98224c),
	.w5(32'hbadf8db7),
	.w6(32'h39889233),
	.w7(32'h3843f341),
	.w8(32'hba476a0f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8f0ba),
	.w1(32'h3957dec3),
	.w2(32'h3a89aa75),
	.w3(32'hbab03aac),
	.w4(32'hb98ee84e),
	.w5(32'h3a09eb1b),
	.w6(32'h38240a49),
	.w7(32'h39f281e8),
	.w8(32'h3a526e79),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8787e9),
	.w1(32'h3aa42b85),
	.w2(32'h3b17c2fe),
	.w3(32'hbacf3155),
	.w4(32'hb9d9cf42),
	.w5(32'h3ad79847),
	.w6(32'h3a43d930),
	.w7(32'h3a31b8eb),
	.w8(32'h3a8e1878),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aaaef),
	.w1(32'h38ab2b46),
	.w2(32'h3844e3a2),
	.w3(32'h391be1ad),
	.w4(32'hb9a800f1),
	.w5(32'hba528d76),
	.w6(32'h3ad7e775),
	.w7(32'h39ce0ef0),
	.w8(32'h3a5ffb5d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bd124),
	.w1(32'hba63549f),
	.w2(32'h3b1f03fe),
	.w3(32'hbb541d55),
	.w4(32'hbad65baa),
	.w5(32'h3b16bbcf),
	.w6(32'hbaa896a1),
	.w7(32'h38b9f723),
	.w8(32'h3b4c337f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad34c59),
	.w1(32'h3ae17653),
	.w2(32'hb98b8e8f),
	.w3(32'h39dbb751),
	.w4(32'hba4fb71d),
	.w5(32'hbba4e31b),
	.w6(32'h3bd3eca2),
	.w7(32'h3ae06577),
	.w8(32'h3939220d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6c688),
	.w1(32'hba06942f),
	.w2(32'h3b812e33),
	.w3(32'h3aa9405b),
	.w4(32'h3b25f828),
	.w5(32'h3c17ccd5),
	.w6(32'h3bab5510),
	.w7(32'h3c08f473),
	.w8(32'h3c26f0dc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb126674),
	.w1(32'hbaf28f90),
	.w2(32'h3b6e6818),
	.w3(32'hbb27c986),
	.w4(32'hbb595cbf),
	.w5(32'h3931b3d7),
	.w6(32'h3b4d49b6),
	.w7(32'h3a10e3d7),
	.w8(32'h3b01d0d0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01fed7),
	.w1(32'h3b38164d),
	.w2(32'h3b78074d),
	.w3(32'hbb4c7cc9),
	.w4(32'hbb4e1bb0),
	.w5(32'h3a7a5f20),
	.w6(32'h3c0619fa),
	.w7(32'h3b16e5e7),
	.w8(32'h3b503afe),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b79f73),
	.w1(32'hbb131f38),
	.w2(32'h3b879a08),
	.w3(32'h3aa05b4e),
	.w4(32'hbb337f98),
	.w5(32'h3b66dc93),
	.w6(32'h3b40d34b),
	.w7(32'h3b5424db),
	.w8(32'h3b62a036),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4ae62),
	.w1(32'h3a079789),
	.w2(32'h3ad2f650),
	.w3(32'hbad5a60f),
	.w4(32'hb8f2cc76),
	.w5(32'h3b015176),
	.w6(32'h3b2d49f5),
	.w7(32'h3a2e26e0),
	.w8(32'h3ae13210),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5629),
	.w1(32'hbb8abdf3),
	.w2(32'h3a943aa0),
	.w3(32'hb9be7c5a),
	.w4(32'hbb190b25),
	.w5(32'h3b6e71fa),
	.w6(32'h3ab56097),
	.w7(32'h3a2b564b),
	.w8(32'h3aceab85),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f068),
	.w1(32'hb9d9798e),
	.w2(32'h3b051fcb),
	.w3(32'hbabec5c8),
	.w4(32'hb9828361),
	.w5(32'h3b1210ed),
	.w6(32'h3933be8f),
	.w7(32'h3880f11b),
	.w8(32'h3b190ba2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34d98c),
	.w1(32'hb9d606e5),
	.w2(32'h3b9093dc),
	.w3(32'hbb746d99),
	.w4(32'hbb888da5),
	.w5(32'h3b5bda34),
	.w6(32'h3bd70c11),
	.w7(32'h3b8ee6f5),
	.w8(32'h3c00f720),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba17ba8),
	.w1(32'hba8274de),
	.w2(32'hbba36f6f),
	.w3(32'h3b90807b),
	.w4(32'hbb0ecee2),
	.w5(32'hbbf20473),
	.w6(32'h3bdf844d),
	.w7(32'h3abeb5f9),
	.w8(32'hbb8b038f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c8ecf),
	.w1(32'h3a5c2daf),
	.w2(32'h37eb9b1b),
	.w3(32'hbad57671),
	.w4(32'h3a221b95),
	.w5(32'hb7f9ba83),
	.w6(32'h3a84c120),
	.w7(32'h39a86353),
	.w8(32'h38a1f558),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec6382),
	.w1(32'h3a6ca478),
	.w2(32'h3b5fc481),
	.w3(32'hb821b028),
	.w4(32'h3a063a66),
	.w5(32'h3b1526a1),
	.w6(32'hb8d548d0),
	.w7(32'h3ab607bd),
	.w8(32'hba29db49),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1a89b),
	.w1(32'hbb006141),
	.w2(32'h3a9d6a48),
	.w3(32'h39be21b0),
	.w4(32'hba502d8d),
	.w5(32'h3a597447),
	.w6(32'h39a637c4),
	.w7(32'h3ab25e13),
	.w8(32'h3b197b6b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65a3f4),
	.w1(32'h39e750fd),
	.w2(32'h3b2cc647),
	.w3(32'h3adcfcf1),
	.w4(32'hba9d1b0a),
	.w5(32'hbb61d56b),
	.w6(32'h3c102b4c),
	.w7(32'h3b88ea26),
	.w8(32'h383af998),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca5c54),
	.w1(32'hb9aabd41),
	.w2(32'h3c36d031),
	.w3(32'hbbfc5e12),
	.w4(32'h3b5ce4a3),
	.w5(32'h3c594097),
	.w6(32'hbb176c28),
	.w7(32'h3baa0267),
	.w8(32'h3c425c11),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921b0a5),
	.w1(32'h3a16ed9e),
	.w2(32'hba4e40ca),
	.w3(32'hb8f12b8e),
	.w4(32'h3aa50f94),
	.w5(32'hb94d1b7d),
	.w6(32'h3b07195c),
	.w7(32'h398f5582),
	.w8(32'h3a2cf6ca),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3d807),
	.w1(32'hbb0d0e72),
	.w2(32'h3bd1f9fc),
	.w3(32'hbb614641),
	.w4(32'hba5cadda),
	.w5(32'h3c00f936),
	.w6(32'h3a4eb3ec),
	.w7(32'h3b879f2f),
	.w8(32'h3c0d4336),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba825c20),
	.w1(32'h3a0d9fd3),
	.w2(32'h3b6bc564),
	.w3(32'h38489cd6),
	.w4(32'h3b25f791),
	.w5(32'h3b0de57c),
	.w6(32'h3bec823d),
	.w7(32'h3be8aeee),
	.w8(32'h3ba419b6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dce39),
	.w1(32'h3b7efce0),
	.w2(32'h3be32855),
	.w3(32'h3b25bbc7),
	.w4(32'h3ba035be),
	.w5(32'h3c15ab56),
	.w6(32'h3a1b8b86),
	.w7(32'h3b68ce8c),
	.w8(32'h3c078fc2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88332a9),
	.w1(32'h3aedf220),
	.w2(32'h3bc2d245),
	.w3(32'hbab3a2dd),
	.w4(32'hb8952448),
	.w5(32'h3b600cef),
	.w6(32'h3b9daee3),
	.w7(32'h3bd0b14e),
	.w8(32'h3c2e6c4e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b923499),
	.w1(32'h3b34bf27),
	.w2(32'hb93c1654),
	.w3(32'h3bbf1ad3),
	.w4(32'h3b1b5312),
	.w5(32'hbac6e0ed),
	.w6(32'h3bc78e55),
	.w7(32'h3bb06b9a),
	.w8(32'h3a4a914a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a0d2d),
	.w1(32'hbb628cf0),
	.w2(32'hbae3c277),
	.w3(32'hbafff8b2),
	.w4(32'hbab23508),
	.w5(32'hba729085),
	.w6(32'hbb56e4db),
	.w7(32'hbb66fc15),
	.w8(32'hbb039697),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d6ba4),
	.w1(32'h3a8cfcf0),
	.w2(32'h3c0265c0),
	.w3(32'hbba2eacf),
	.w4(32'hba8ec39a),
	.w5(32'h3bca638b),
	.w6(32'hbb3a1176),
	.w7(32'hba9e03ca),
	.w8(32'h3bfd7faf),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53570a),
	.w1(32'h3b965ad2),
	.w2(32'hbb5903b1),
	.w3(32'h3bbb77ac),
	.w4(32'h3b77c6dc),
	.w5(32'hbbec9da4),
	.w6(32'h3c9ce842),
	.w7(32'h3c1282eb),
	.w8(32'hbb6bef68),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66e3cd),
	.w1(32'hba74f7c1),
	.w2(32'h3ba683b8),
	.w3(32'hbab6068c),
	.w4(32'hbb2861a9),
	.w5(32'h3b1f1488),
	.w6(32'h3a79bd76),
	.w7(32'h39d147f3),
	.w8(32'h3bcc538d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55df65),
	.w1(32'h3a766dee),
	.w2(32'h393c2c94),
	.w3(32'h399cd114),
	.w4(32'h39a0fe93),
	.w5(32'h36ca4e17),
	.w6(32'h3aefbc11),
	.w7(32'h3a613dde),
	.w8(32'h3a733836),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d8db3),
	.w1(32'h39814b8f),
	.w2(32'hba092c66),
	.w3(32'hb9a4d4ec),
	.w4(32'h3a35f7d4),
	.w5(32'hb91729a6),
	.w6(32'h3a2af1fc),
	.w7(32'hb8946fde),
	.w8(32'h376d1d2f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba682d2d),
	.w1(32'h3a2ee82a),
	.w2(32'h3b61897e),
	.w3(32'hba8c23bc),
	.w4(32'hbaae5e70),
	.w5(32'h3b6b6345),
	.w6(32'h3bb9dcef),
	.w7(32'h3b84a2f1),
	.w8(32'h3b7474d9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35ce19),
	.w1(32'h3a8c42d3),
	.w2(32'h3ae13133),
	.w3(32'h3a3665aa),
	.w4(32'h3a3f74ed),
	.w5(32'h3ab29237),
	.w6(32'h3ab97ffb),
	.w7(32'h3a74f21c),
	.w8(32'h3af5d219),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71fcffc),
	.w1(32'hbb690cf6),
	.w2(32'h3b9683c6),
	.w3(32'hbacb5031),
	.w4(32'hbb990b78),
	.w5(32'h3aeef871),
	.w6(32'hbac17670),
	.w7(32'hba945faa),
	.w8(32'h3b066aec),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c1ca9),
	.w1(32'h3a87c45e),
	.w2(32'h3ab8440b),
	.w3(32'hba384a81),
	.w4(32'h39d1e62b),
	.w5(32'h3a9968bd),
	.w6(32'hb9894141),
	.w7(32'hba83629e),
	.w8(32'h38a6644a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0958),
	.w1(32'hbaad096a),
	.w2(32'h3c48ef0b),
	.w3(32'hbb840aa3),
	.w4(32'hbab49b47),
	.w5(32'h3c67c967),
	.w6(32'hbb5ad18e),
	.w7(32'h3aa94af6),
	.w8(32'h3c86b277),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d08583),
	.w1(32'hb9c9d579),
	.w2(32'h3a287418),
	.w3(32'hba648f16),
	.w4(32'hba66a7b0),
	.w5(32'h39185531),
	.w6(32'hba21933a),
	.w7(32'h395e1f1b),
	.w8(32'h39d7c3ee),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396765bd),
	.w1(32'h39b90a49),
	.w2(32'h3a32bbdd),
	.w3(32'h39676293),
	.w4(32'h3a93fa85),
	.w5(32'h3a92925a),
	.w6(32'h3a80a8cf),
	.w7(32'h39715530),
	.w8(32'h3aa17bf4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba870748),
	.w1(32'hbaffe774),
	.w2(32'hba185c57),
	.w3(32'hbadcb0f4),
	.w4(32'hbb8513a5),
	.w5(32'hbba45014),
	.w6(32'h3ac12b16),
	.w7(32'hba3dbfd6),
	.w8(32'hbb95f426),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2267a6),
	.w1(32'hbb4a590b),
	.w2(32'h3bbf24ef),
	.w3(32'hbb3244c8),
	.w4(32'hbbc88379),
	.w5(32'h3b9d2efc),
	.w6(32'h3be1638d),
	.w7(32'h3b8bd232),
	.w8(32'h3c39f98c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f90a1),
	.w1(32'hbae2b017),
	.w2(32'h3be06bc5),
	.w3(32'hbb5220b0),
	.w4(32'hbb0c0c16),
	.w5(32'h3be019e3),
	.w6(32'hbb4f7f3d),
	.w7(32'hbac5f639),
	.w8(32'h3b9e3d75),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92920b),
	.w1(32'hbb70009f),
	.w2(32'h3b9d60cf),
	.w3(32'hbb4375a8),
	.w4(32'hbb1a378f),
	.w5(32'h3b85c74a),
	.w6(32'h3a5723c3),
	.w7(32'h39856ffa),
	.w8(32'h3be4e464),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba435fc7),
	.w1(32'hbb85cc25),
	.w2(32'hba51ef13),
	.w3(32'h39fffe86),
	.w4(32'hbb8f9618),
	.w5(32'hbb1e9ae3),
	.w6(32'hbb071201),
	.w7(32'h3a526740),
	.w8(32'h3a7b8482),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69438c),
	.w1(32'hbae72509),
	.w2(32'h3ba279e6),
	.w3(32'hbc02668e),
	.w4(32'hba2eca28),
	.w5(32'h3bd1ebfb),
	.w6(32'h3bf6f28b),
	.w7(32'h3c32e7a8),
	.w8(32'h3c2a7a2e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad2b5c),
	.w1(32'h3ae04a4e),
	.w2(32'h3c275c4a),
	.w3(32'hbacd7f25),
	.w4(32'hbac51320),
	.w5(32'h3bc5d537),
	.w6(32'h3b7c1df9),
	.w7(32'h3b92d670),
	.w8(32'h3c20b0d4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306771),
	.w1(32'hbb2bf904),
	.w2(32'h3b852c72),
	.w3(32'hba4aed1a),
	.w4(32'hbae7bb6b),
	.w5(32'h3b7bae7d),
	.w6(32'h3a6e29e9),
	.w7(32'h3ab3810a),
	.w8(32'h3b91f242),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451d42),
	.w1(32'hbacd5c58),
	.w2(32'h3a1f7049),
	.w3(32'hbb8e29c3),
	.w4(32'hbaaa3b10),
	.w5(32'h39fb156c),
	.w6(32'hbae17113),
	.w7(32'hb93d9a16),
	.w8(32'hbaf09ba4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd38a),
	.w1(32'h3ae613d1),
	.w2(32'hbb009baf),
	.w3(32'h39a66a54),
	.w4(32'h39680ffc),
	.w5(32'hbb941335),
	.w6(32'h3b6a883b),
	.w7(32'h3a5f1020),
	.w8(32'hbb8ffa30),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0451ae),
	.w1(32'hb9152315),
	.w2(32'hba8a6e12),
	.w3(32'h3a141ed1),
	.w4(32'h39585d54),
	.w5(32'hba19bb53),
	.w6(32'h3997bb97),
	.w7(32'hb9a4bc28),
	.w8(32'hb9e9424c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8de47),
	.w1(32'hbb5331e5),
	.w2(32'hba6fb03a),
	.w3(32'hbacf16c1),
	.w4(32'hbb4ec567),
	.w5(32'h3aa001e7),
	.w6(32'hbb111c26),
	.w7(32'hbabaad71),
	.w8(32'h3b32afa9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b22971),
	.w1(32'hb969fa36),
	.w2(32'hbb4910d4),
	.w3(32'hb9c48799),
	.w4(32'hbabc2c19),
	.w5(32'hbb1b39f1),
	.w6(32'h3a512824),
	.w7(32'hbabcd416),
	.w8(32'hb99523e5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab07180),
	.w1(32'h3bae234a),
	.w2(32'h3bd3cd67),
	.w3(32'hbb38a439),
	.w4(32'h3bab14de),
	.w5(32'h3c069d24),
	.w6(32'h3b9ae344),
	.w7(32'h3c004d70),
	.w8(32'h3c2863b2),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a8643),
	.w1(32'hba6abf57),
	.w2(32'hba51e2bf),
	.w3(32'h394e3046),
	.w4(32'hba7971a9),
	.w5(32'hb9c969f9),
	.w6(32'hba83ea12),
	.w7(32'hb8d6fec8),
	.w8(32'hb9e15d55),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcee34),
	.w1(32'h3b377bba),
	.w2(32'h3b6b0199),
	.w3(32'hba40bfef),
	.w4(32'h3ace1fe3),
	.w5(32'h3b1308cd),
	.w6(32'h3afcb5b7),
	.w7(32'h3b122952),
	.w8(32'h3ae788de),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fcc75),
	.w1(32'h3b70e85a),
	.w2(32'h3b8de110),
	.w3(32'h3a2004d5),
	.w4(32'h3a704a59),
	.w5(32'h3a549e9f),
	.w6(32'h3ba595a9),
	.w7(32'h3bb24572),
	.w8(32'h3becf249),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b168071),
	.w1(32'h3ac74156),
	.w2(32'h3c086e41),
	.w3(32'hba126c1f),
	.w4(32'hba50ed87),
	.w5(32'h3be616cc),
	.w6(32'h3bced21b),
	.w7(32'h3bb4dd2c),
	.w8(32'h3c294485),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5da9ac),
	.w1(32'hbaf4f908),
	.w2(32'h3906da96),
	.w3(32'h3a2ca7fa),
	.w4(32'hba0255f1),
	.w5(32'hb97d3695),
	.w6(32'hb9b6b09d),
	.w7(32'hbaf6825e),
	.w8(32'hb9cca961),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720dfe),
	.w1(32'h3a54b6d6),
	.w2(32'h3a79978f),
	.w3(32'hbac4394b),
	.w4(32'h399a71f8),
	.w5(32'h3a8f6526),
	.w6(32'h3a37b566),
	.w7(32'h3a9b459a),
	.w8(32'h3ab0a501),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab02e4),
	.w1(32'hbc3f1e28),
	.w2(32'h3c2cd1b7),
	.w3(32'hbc83f6e0),
	.w4(32'hbba52783),
	.w5(32'h3c90fd9c),
	.w6(32'hbc43dbde),
	.w7(32'hbbd6fbf1),
	.w8(32'h3c1b8b2e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a799dbb),
	.w1(32'hbaeeec00),
	.w2(32'hbbde46d9),
	.w3(32'h3a77ce26),
	.w4(32'hbc1debe2),
	.w5(32'hbc85de45),
	.w6(32'h3c137d11),
	.w7(32'hbbb87920),
	.w8(32'hbc2ffb87),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2e98),
	.w1(32'hbaf23db4),
	.w2(32'h387c3230),
	.w3(32'hbac39f6a),
	.w4(32'hba469e15),
	.w5(32'h3a9b8c39),
	.w6(32'hba54eec0),
	.w7(32'hb92c2289),
	.w8(32'h3ac7f9b9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05589c),
	.w1(32'h3a73e832),
	.w2(32'h3949eac0),
	.w3(32'hb91447f2),
	.w4(32'h3974cb56),
	.w5(32'h39afb192),
	.w6(32'h38b22cc4),
	.w7(32'h3a1e2957),
	.w8(32'h38018a3b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fc56e),
	.w1(32'hbb23bba9),
	.w2(32'hb90abde8),
	.w3(32'h3a2a900f),
	.w4(32'hbb2b7393),
	.w5(32'hba5c45e2),
	.w6(32'hba967077),
	.w7(32'h3a127070),
	.w8(32'h3a8c7a60),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbf099),
	.w1(32'h39b474e6),
	.w2(32'hb9cb3b4e),
	.w3(32'hba22d8a6),
	.w4(32'h39dae1cf),
	.w5(32'h3955394f),
	.w6(32'hb96e693a),
	.w7(32'hba0182ca),
	.w8(32'hba18bb94),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75af74),
	.w1(32'hb9b6146d),
	.w2(32'h39a1eedc),
	.w3(32'h396047ee),
	.w4(32'h3a37cdca),
	.w5(32'h3aa23d2b),
	.w6(32'h3a64803c),
	.w7(32'h3b0239b7),
	.w8(32'h3a1006e2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981160c),
	.w1(32'hbb5d93f9),
	.w2(32'hbb41afe9),
	.w3(32'h3a4e187c),
	.w4(32'hbbcef4fc),
	.w5(32'hbb1bb860),
	.w6(32'h3bd3d72d),
	.w7(32'h3bbcc4db),
	.w8(32'h3ba93fb8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc66b7),
	.w1(32'hbb4c165e),
	.w2(32'h3b711117),
	.w3(32'hbbbc98a6),
	.w4(32'hbae18da2),
	.w5(32'h3ab699fa),
	.w6(32'h3c01fb42),
	.w7(32'h3ba502fe),
	.w8(32'h3c03274e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15515d),
	.w1(32'h39c45a49),
	.w2(32'h3b2f08a2),
	.w3(32'hb99cd1fa),
	.w4(32'hba871580),
	.w5(32'h3a7f09f8),
	.w6(32'h3ab02fe0),
	.w7(32'hba4cd041),
	.w8(32'h3b0a93e6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147076),
	.w1(32'hbaca5df5),
	.w2(32'h3c23c9d2),
	.w3(32'hbb1dcf49),
	.w4(32'h3b242c63),
	.w5(32'h3c8216a5),
	.w6(32'hba25bf64),
	.w7(32'h3bb79a6a),
	.w8(32'h3c6e8893),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fcf64),
	.w1(32'h3b31f312),
	.w2(32'h3b708ff8),
	.w3(32'hbb0557d6),
	.w4(32'h3b1b5b36),
	.w5(32'h3b8c58ab),
	.w6(32'hb9562be9),
	.w7(32'h3b804a15),
	.w8(32'h3bc0af85),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999493a),
	.w1(32'h39dc0b2c),
	.w2(32'hb9feefed),
	.w3(32'hb88443a9),
	.w4(32'h3a8817f3),
	.w5(32'hb8013ca1),
	.w6(32'h3a1d9599),
	.w7(32'hb84fe8d3),
	.w8(32'hb986d292),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a97cb6),
	.w1(32'h3a8c0428),
	.w2(32'hba115d85),
	.w3(32'h3a385add),
	.w4(32'h3a933456),
	.w5(32'hba230f02),
	.w6(32'h3a812c03),
	.w7(32'hb9cf872f),
	.w8(32'hba2ec604),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0c5e6),
	.w1(32'h384c4e32),
	.w2(32'hbab7622d),
	.w3(32'h390b9c51),
	.w4(32'h3a63ce58),
	.w5(32'hb9e5d60f),
	.w6(32'h3a1c8f08),
	.w7(32'hb9d27369),
	.w8(32'hba50969c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0add9f),
	.w1(32'hba3d8e8e),
	.w2(32'h3be53c84),
	.w3(32'hbb287e06),
	.w4(32'hbb46e5c4),
	.w5(32'h3bda2c67),
	.w6(32'h3b4d08c1),
	.w7(32'h3b4f39e2),
	.w8(32'h3c24dcec),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd97b00),
	.w1(32'hb9e0ed26),
	.w2(32'hba2faf64),
	.w3(32'h3b5ade0a),
	.w4(32'hbbe5c066),
	.w5(32'hbc1d0f86),
	.w6(32'h3c10efc7),
	.w7(32'hb953d558),
	.w8(32'hba655e04),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68696e),
	.w1(32'hba045aac),
	.w2(32'h3be267c3),
	.w3(32'hbb25cf0a),
	.w4(32'hbb0f4d3d),
	.w5(32'h3b5dc3a8),
	.w6(32'h3b9b9930),
	.w7(32'h3b57a1b4),
	.w8(32'h3c02f348),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba557dec),
	.w1(32'h3aa14b4e),
	.w2(32'h3b8e955d),
	.w3(32'hba85d442),
	.w4(32'h3a5d43dc),
	.w5(32'h3b82ac5c),
	.w6(32'hb9083d69),
	.w7(32'h3a82e418),
	.w8(32'h3b5152ab),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31a4b9),
	.w1(32'h3b624cd0),
	.w2(32'h3c081973),
	.w3(32'hbba4530c),
	.w4(32'hbb32b6bd),
	.w5(32'h3a56323c),
	.w6(32'h3bd9acbc),
	.w7(32'h3be6a12c),
	.w8(32'h3be8e9b3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4255),
	.w1(32'hbb1129c1),
	.w2(32'h3af74b3e),
	.w3(32'hba9056c1),
	.w4(32'hb95ff608),
	.w5(32'h3b4aa53e),
	.w6(32'h3ad51aa3),
	.w7(32'h3a24fca4),
	.w8(32'h3b5a3d37),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6de020),
	.w1(32'h3b38c3a5),
	.w2(32'h3c5ebc1c),
	.w3(32'hbb34b011),
	.w4(32'h3c00bf3e),
	.w5(32'h3c877317),
	.w6(32'h3c2027ad),
	.w7(32'h3c70a946),
	.w8(32'h3cb042ea),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989307f),
	.w1(32'h39c8c412),
	.w2(32'h3a3399fe),
	.w3(32'hb82d31dc),
	.w4(32'hb466bdc9),
	.w5(32'h3a15dc13),
	.w6(32'hb8f64636),
	.w7(32'h39fd362d),
	.w8(32'h39fc7ebc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33537b),
	.w1(32'h3a54d8a4),
	.w2(32'h3ad7e40a),
	.w3(32'h39dc6684),
	.w4(32'h3a2bc3d1),
	.w5(32'h3abf838e),
	.w6(32'h3aa06805),
	.w7(32'h3ad32206),
	.w8(32'h3a90d59f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a6d6),
	.w1(32'h3b444fcb),
	.w2(32'h3c349937),
	.w3(32'hbb0ef563),
	.w4(32'hbba425ec),
	.w5(32'h3ba7c3cd),
	.w6(32'h3bd64112),
	.w7(32'h3bb2fc9a),
	.w8(32'h3c39b983),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f585),
	.w1(32'hbb254f8a),
	.w2(32'h3c499326),
	.w3(32'hbbd74c73),
	.w4(32'hbb846aaa),
	.w5(32'h3c1ef6b0),
	.w6(32'h3bbbe911),
	.w7(32'h3ba69bcb),
	.w8(32'h3c5e5664),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfe76a),
	.w1(32'h39f7aff4),
	.w2(32'h3c0d8d9f),
	.w3(32'h3a3168bb),
	.w4(32'hbb6eadb2),
	.w5(32'h3b4c9aff),
	.w6(32'h3bd6f52d),
	.w7(32'h3bb04e9b),
	.w8(32'h3c036f72),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0ebd),
	.w1(32'hbbaebec3),
	.w2(32'hbb1d928a),
	.w3(32'hbac787d7),
	.w4(32'hbaa5c596),
	.w5(32'h3abb1a2f),
	.w6(32'hbb11453e),
	.w7(32'h39e1e7fc),
	.w8(32'h3a90aaab),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988f34e),
	.w1(32'h3977c598),
	.w2(32'hba6c0dc1),
	.w3(32'hb99315ae),
	.w4(32'h3a18d487),
	.w5(32'hba0f2393),
	.w6(32'h3aa2104c),
	.w7(32'h3969e1df),
	.w8(32'hb8f6768e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba449277),
	.w1(32'h3b21ba86),
	.w2(32'h3b57c9fa),
	.w3(32'hb9f26e06),
	.w4(32'h3a7cb2bb),
	.w5(32'h3b00b793),
	.w6(32'h3aff2a83),
	.w7(32'h3b09e705),
	.w8(32'h3ae12549),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b569d),
	.w1(32'hbb6e43a1),
	.w2(32'h3b7dc700),
	.w3(32'h3999af2c),
	.w4(32'hbb5c08aa),
	.w5(32'h3b841f8e),
	.w6(32'h38c81fe2),
	.w7(32'hbaab0213),
	.w8(32'h3b8c1c18),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7dba),
	.w1(32'hbb968299),
	.w2(32'h3c003154),
	.w3(32'hbb971ae9),
	.w4(32'hbad0d55b),
	.w5(32'h3c21f07b),
	.w6(32'h3a58a8e0),
	.w7(32'h3bdf44f0),
	.w8(32'h3c61f191),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc57df3),
	.w1(32'h3add727f),
	.w2(32'h3b1e02b6),
	.w3(32'h3a648aa3),
	.w4(32'hbb452dac),
	.w5(32'h3b27f371),
	.w6(32'h3b22b0ed),
	.w7(32'h3b49f1cd),
	.w8(32'h3b20a86a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256d8d),
	.w1(32'h3a941784),
	.w2(32'h3b5d1b53),
	.w3(32'hbae1df97),
	.w4(32'hbb73c18e),
	.w5(32'hbb456c9d),
	.w6(32'h3be0d972),
	.w7(32'h3b7274a7),
	.w8(32'h3b340325),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8778d0a),
	.w1(32'h3b41afdd),
	.w2(32'h3c1e068f),
	.w3(32'hbb5032d6),
	.w4(32'h39ae8563),
	.w5(32'h3bba9e68),
	.w6(32'h3be853c6),
	.w7(32'h3bb5bb97),
	.w8(32'h3c368f7f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958b065),
	.w1(32'h397d9845),
	.w2(32'h39f0f665),
	.w3(32'h38354b50),
	.w4(32'h39a7edb8),
	.w5(32'h39c0e412),
	.w6(32'h3784241a),
	.w7(32'hb8acf0fe),
	.w8(32'hb9908278),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb53d1),
	.w1(32'hb9c8fc4a),
	.w2(32'hba8164b8),
	.w3(32'h38712933),
	.w4(32'h38e66b15),
	.w5(32'hb9c413e0),
	.w6(32'h395d548b),
	.w7(32'hb5db655d),
	.w8(32'hba53478f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd1f8),
	.w1(32'h3aae57d5),
	.w2(32'h3a42ca16),
	.w3(32'hbaa0f43f),
	.w4(32'h3a9d720f),
	.w5(32'hb970eead),
	.w6(32'h3af7f86d),
	.w7(32'h3a7f6a92),
	.w8(32'h39979bfe),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da04d6),
	.w1(32'h39cec2bb),
	.w2(32'hbab06258),
	.w3(32'hbaba4e2e),
	.w4(32'h3a51ca9d),
	.w5(32'hba9812b3),
	.w6(32'h39c3fa3d),
	.w7(32'hba8b7e68),
	.w8(32'hb99b0c8e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f4e67),
	.w1(32'h3a8182b2),
	.w2(32'h3b4b8fa1),
	.w3(32'h39c0ab28),
	.w4(32'h3a750099),
	.w5(32'h3b52f602),
	.w6(32'h39266480),
	.w7(32'h3b146782),
	.w8(32'h3b2dbec6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88af088),
	.w1(32'h3b2dfec2),
	.w2(32'h3c288a87),
	.w3(32'hba35b615),
	.w4(32'hba45ee5e),
	.w5(32'h3be15042),
	.w6(32'h3bb5ec04),
	.w7(32'h3ba4a250),
	.w8(32'h3c15a806),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c200c),
	.w1(32'hba9006f7),
	.w2(32'h3acc821a),
	.w3(32'hbab2d996),
	.w4(32'hbb3d51dc),
	.w5(32'h3ad23665),
	.w6(32'h3ad7d5a3),
	.w7(32'h3aaa351a),
	.w8(32'h3b73329b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3849ea63),
	.w1(32'hba872b81),
	.w2(32'hbb1d7591),
	.w3(32'hba3128f2),
	.w4(32'hba9d31ca),
	.w5(32'hbaf7afd8),
	.w6(32'hba8ef629),
	.w7(32'hb97dc3e3),
	.w8(32'hbaf5dbb3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba57aed),
	.w1(32'h3b912204),
	.w2(32'h3bfd401a),
	.w3(32'h3b2c1981),
	.w4(32'h3ba5944a),
	.w5(32'h3c3759f9),
	.w6(32'h3b9a906b),
	.w7(32'h3beeb6cf),
	.w8(32'h3c53c930),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8fa7d),
	.w1(32'h3a2e054a),
	.w2(32'h3acb7fb6),
	.w3(32'hba8aba9d),
	.w4(32'h3a60daf8),
	.w5(32'h3af32be5),
	.w6(32'h3ae71510),
	.w7(32'h3ab98904),
	.w8(32'h3b1380d7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9930f49),
	.w1(32'h36e3bfa5),
	.w2(32'hba38eddf),
	.w3(32'h39983eba),
	.w4(32'h39bf92c7),
	.w5(32'hba0c948b),
	.w6(32'h3a662565),
	.w7(32'h39c93b02),
	.w8(32'h39688c9a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba950944),
	.w1(32'hb944bfb8),
	.w2(32'h3b95c0d3),
	.w3(32'hbadaedd6),
	.w4(32'h3a3afc33),
	.w5(32'h3bcdcc1f),
	.w6(32'h3a555172),
	.w7(32'h3b0c40c4),
	.w8(32'h3b972a95),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18f787),
	.w1(32'hb9ab8724),
	.w2(32'h38b7243c),
	.w3(32'hb9c1b5ec),
	.w4(32'h399829c3),
	.w5(32'h3a7bac29),
	.w6(32'hb81b7eac),
	.w7(32'hb9a8dab0),
	.w8(32'hb997b293),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a844e87),
	.w1(32'h39479bc6),
	.w2(32'hba90789b),
	.w3(32'h3a941e13),
	.w4(32'h3a2fa00c),
	.w5(32'hba3e1fb7),
	.w6(32'h3af3693d),
	.w7(32'hb463ac33),
	.w8(32'h39e90fde),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7aaeb),
	.w1(32'h3897d99a),
	.w2(32'hb9ca1c9f),
	.w3(32'hb9c96203),
	.w4(32'h39bea9d1),
	.w5(32'hb9b178eb),
	.w6(32'h3a49fc2c),
	.w7(32'h39bd59a9),
	.w8(32'h3986beed),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc8e31),
	.w1(32'hba96fcbf),
	.w2(32'hba2fefa8),
	.w3(32'hb9d12ad9),
	.w4(32'hba925be2),
	.w5(32'hba4226a0),
	.w6(32'hbaa80712),
	.w7(32'hbaa0522b),
	.w8(32'hbaa16c76),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd0eb1),
	.w1(32'h3b628c4c),
	.w2(32'h3b85bd8f),
	.w3(32'h3ac4e8ab),
	.w4(32'h3b1c7da1),
	.w5(32'h3b1dda2b),
	.w6(32'h3ba3811a),
	.w7(32'h3b84f1ea),
	.w8(32'h3b635d78),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe782d1),
	.w1(32'hbb46c028),
	.w2(32'h3bc1ca09),
	.w3(32'hbafbfcf2),
	.w4(32'hba97c87e),
	.w5(32'h3bc7a9bd),
	.w6(32'h3b3c273d),
	.w7(32'h3b6f4b06),
	.w8(32'h3c0e1afb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e42c),
	.w1(32'hbaf98cbe),
	.w2(32'h3b6a2512),
	.w3(32'hbb8fcede),
	.w4(32'hba9c93f2),
	.w5(32'h3b6595d4),
	.w6(32'hb9b4ba7c),
	.w7(32'hba2b2040),
	.w8(32'h3b050447),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51468),
	.w1(32'hbb82df88),
	.w2(32'h3a1b8d54),
	.w3(32'hbb8be670),
	.w4(32'hbab49b3b),
	.w5(32'h3b84f0a3),
	.w6(32'hba906f3e),
	.w7(32'h3aaab812),
	.w8(32'h3b3f7b20),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba598125),
	.w1(32'hbaa58dcb),
	.w2(32'hb831f5a6),
	.w3(32'hba2baea2),
	.w4(32'hbabd2db9),
	.w5(32'hba825a84),
	.w6(32'hba010ba0),
	.w7(32'hba53558f),
	.w8(32'hb9888981),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c637d9),
	.w1(32'h39cba4f8),
	.w2(32'hb9275c33),
	.w3(32'hb9e36394),
	.w4(32'h3a5721fb),
	.w5(32'hb98aa4ce),
	.w6(32'h3a96f572),
	.w7(32'h3a39183d),
	.w8(32'h3a36a79d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9e864),
	.w1(32'h3980f01b),
	.w2(32'hb9d0c027),
	.w3(32'hba05d505),
	.w4(32'h3a44889e),
	.w5(32'h36dd632c),
	.w6(32'h3a1f0145),
	.w7(32'h37691ca7),
	.w8(32'hb94ddf26),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cf5b0),
	.w1(32'h39a24ee4),
	.w2(32'hb99db2e4),
	.w3(32'hb93052cc),
	.w4(32'h3a5c6ca7),
	.w5(32'hb5836fa7),
	.w6(32'h3a4187d6),
	.w7(32'h3999cbfa),
	.w8(32'hb7e55ec9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e161d),
	.w1(32'h3b222105),
	.w2(32'h3b21df44),
	.w3(32'h3b0a92fa),
	.w4(32'h3aa064bf),
	.w5(32'h3aeb4b2a),
	.w6(32'h3bfaa3c8),
	.w7(32'h3baf3821),
	.w8(32'h3ada954a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa26229),
	.w1(32'h3a488e48),
	.w2(32'h3a559777),
	.w3(32'h3b3c2290),
	.w4(32'h3aa41eb2),
	.w5(32'h3aa1b7ec),
	.w6(32'h3a120f0a),
	.w7(32'h3a23d8d3),
	.w8(32'hba164974),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab102b9),
	.w1(32'hba838b5d),
	.w2(32'h3b386b96),
	.w3(32'hbb136110),
	.w4(32'hbaa02501),
	.w5(32'h3b1c1ea7),
	.w6(32'hb9bd0b2c),
	.w7(32'hbadad380),
	.w8(32'h3b081a12),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8deec87),
	.w1(32'h3ab5cd10),
	.w2(32'h3b1353a6),
	.w3(32'hb96638d8),
	.w4(32'h3a9290e3),
	.w5(32'h3ac6b3c8),
	.w6(32'h39407972),
	.w7(32'h38d9489a),
	.w8(32'h3aaf66bd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f99f0),
	.w1(32'h399be577),
	.w2(32'hba0f8a16),
	.w3(32'hba0705c0),
	.w4(32'h3a66f739),
	.w5(32'h3866eb27),
	.w6(32'h3a088b58),
	.w7(32'hb942057c),
	.w8(32'hb8d30006),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ae295),
	.w1(32'hbb557524),
	.w2(32'hb9ddb502),
	.w3(32'h399fae20),
	.w4(32'hbaad18f3),
	.w5(32'h39266ade),
	.w6(32'h3ad9aff2),
	.w7(32'h3af147a3),
	.w8(32'h3a838c80),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba909743),
	.w1(32'h3b1a236d),
	.w2(32'h3ad34357),
	.w3(32'hba06ebea),
	.w4(32'h3afc817e),
	.w5(32'h3a480c29),
	.w6(32'h3b2f71b4),
	.w7(32'h3adfb407),
	.w8(32'h3a98f0a1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a536b),
	.w1(32'h3ad53529),
	.w2(32'h3931395e),
	.w3(32'hbaa57775),
	.w4(32'hb9da4b7a),
	.w5(32'hbb1133b6),
	.w6(32'h3bc98b5b),
	.w7(32'h3b01ddc1),
	.w8(32'h3a8956f2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba872ec4),
	.w1(32'hba30a988),
	.w2(32'hba7edc43),
	.w3(32'hb8be1432),
	.w4(32'hb98ce464),
	.w5(32'hba0c2c36),
	.w6(32'hb9612439),
	.w7(32'hb9a001b6),
	.w8(32'hb6a212ae),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10f904),
	.w1(32'h3ac9b170),
	.w2(32'h3b5307a1),
	.w3(32'hbc02325f),
	.w4(32'hbb8512c7),
	.w5(32'hbc103416),
	.w6(32'h3b8deb7a),
	.w7(32'h3b87cbe3),
	.w8(32'hb9c02e8e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule