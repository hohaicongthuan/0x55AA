module layer_10_featuremap_79(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba26265),
	.w1(32'h3b96deee),
	.w2(32'hbb284376),
	.w3(32'hba1f4178),
	.w4(32'h3b1e070c),
	.w5(32'h3b7f45a4),
	.w6(32'h3c42edb7),
	.w7(32'hbb0ff526),
	.w8(32'h38f876cf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd6456),
	.w1(32'hbb898397),
	.w2(32'h3b0b5814),
	.w3(32'hbb5041eb),
	.w4(32'h3b90a605),
	.w5(32'hbbc531a2),
	.w6(32'hbb993e91),
	.w7(32'hbc1bc668),
	.w8(32'h3b81b013),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb951ace),
	.w1(32'h3a07fa1f),
	.w2(32'h3b696363),
	.w3(32'hba631f4e),
	.w4(32'hbc2343db),
	.w5(32'h3b84441b),
	.w6(32'hbd10dca7),
	.w7(32'hbc047c44),
	.w8(32'hbb9c89d3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8002c5d),
	.w1(32'h398b94dd),
	.w2(32'hbb0038ba),
	.w3(32'h3c4555ac),
	.w4(32'hbc422583),
	.w5(32'hbb95dee6),
	.w6(32'hbb4b3d0c),
	.w7(32'hbb4be21f),
	.w8(32'hbb93d905),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d35b1),
	.w1(32'hbba47457),
	.w2(32'h3b63a618),
	.w3(32'hbbf8ae97),
	.w4(32'hbbaea9ba),
	.w5(32'h39b57b7c),
	.w6(32'h3b4433d3),
	.w7(32'hbb09c16d),
	.w8(32'hbd93b243),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5105),
	.w1(32'hbb41530e),
	.w2(32'hbbb78ee3),
	.w3(32'h3bd11dd4),
	.w4(32'hba9621dd),
	.w5(32'h3c13e79c),
	.w6(32'h3b1e33e9),
	.w7(32'hba24665b),
	.w8(32'hb9490897),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab50c8),
	.w1(32'hba654342),
	.w2(32'h3bd3bf19),
	.w3(32'h3c0dadc2),
	.w4(32'h3c5e5b96),
	.w5(32'h3aa59a66),
	.w6(32'hbac06ecd),
	.w7(32'h383b9473),
	.w8(32'hbc093913),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e760),
	.w1(32'hbba48d7d),
	.w2(32'h3ab29760),
	.w3(32'h3a0d63a4),
	.w4(32'hba30fcfb),
	.w5(32'h3993342e),
	.w6(32'hbbcebb38),
	.w7(32'h3b0dbeeb),
	.w8(32'hba7eac3d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0ab60),
	.w1(32'h3bee0b40),
	.w2(32'hbba7d57d),
	.w3(32'h3a320c06),
	.w4(32'h3b9a7ad2),
	.w5(32'h3bfc03f2),
	.w6(32'hbc271baf),
	.w7(32'hba1879e0),
	.w8(32'h38c09748),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c778ad2),
	.w1(32'hb9cded14),
	.w2(32'hbc28cf3c),
	.w3(32'h3b8972b5),
	.w4(32'h3b25cf3e),
	.w5(32'hbac607a4),
	.w6(32'hbcf5affa),
	.w7(32'hbbcbd6ef),
	.w8(32'hba703dbf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c3d78),
	.w1(32'hbbf3064b),
	.w2(32'h3bb14537),
	.w3(32'h3a4f0bf6),
	.w4(32'hbc6d8927),
	.w5(32'h3aa0fa81),
	.w6(32'hba11cf04),
	.w7(32'h3be954e1),
	.w8(32'h3aa440c0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39970a9a),
	.w1(32'h3bae2761),
	.w2(32'hbc2ff436),
	.w3(32'h3a8590ca),
	.w4(32'hbb9dc70c),
	.w5(32'hb93f668c),
	.w6(32'h3a839f68),
	.w7(32'hbb01e4bc),
	.w8(32'h3b6df443),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a464),
	.w1(32'hbb17aee1),
	.w2(32'hbb16253e),
	.w3(32'hbbc555d3),
	.w4(32'hbb5736b6),
	.w5(32'hbb635c49),
	.w6(32'h3c29b5c8),
	.w7(32'hbabd11d8),
	.w8(32'hbb07725d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfbb0d),
	.w1(32'h3b5672dd),
	.w2(32'h3aab4c24),
	.w3(32'h3bbc5c53),
	.w4(32'hbcf4a6b5),
	.w5(32'h3b247f62),
	.w6(32'h3c27c9de),
	.w7(32'hb9dc7e66),
	.w8(32'hbb3506ee),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6fd0b),
	.w1(32'hbb855eef),
	.w2(32'h3c21b497),
	.w3(32'h3afc150c),
	.w4(32'hbb425983),
	.w5(32'h3aa88f89),
	.w6(32'hba172499),
	.w7(32'hbbad258a),
	.w8(32'h3b875bcc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd3c3a),
	.w1(32'h3aacf5b1),
	.w2(32'hba820e67),
	.w3(32'h3b9af8e8),
	.w4(32'hbb5c3b37),
	.w5(32'hbb5987f4),
	.w6(32'hbbe05c16),
	.w7(32'hbc15f5ca),
	.w8(32'h3caf47a7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada8a77),
	.w1(32'hbaed5d0f),
	.w2(32'h3b056170),
	.w3(32'hba875e3c),
	.w4(32'h37e1fa74),
	.w5(32'h3970acf7),
	.w6(32'h3a09d23e),
	.w7(32'hba8feb3a),
	.w8(32'h3b19024c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc25875),
	.w1(32'hbceb5105),
	.w2(32'hbc9d550b),
	.w3(32'hbae78342),
	.w4(32'hbbaa322d),
	.w5(32'hba547b44),
	.w6(32'hbbd0e1be),
	.w7(32'hbd739de1),
	.w8(32'hbbe18c06),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56b85f),
	.w1(32'hbb7e6f36),
	.w2(32'h3c09c3be),
	.w3(32'hbb7f7b35),
	.w4(32'hbadc9a46),
	.w5(32'hba49eb56),
	.w6(32'hbbe7ee27),
	.w7(32'hbc08f6e0),
	.w8(32'hb9ad0a6e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24704e),
	.w1(32'hbb360c83),
	.w2(32'hbbe30616),
	.w3(32'hbb792682),
	.w4(32'h3c9c8a1d),
	.w5(32'hb9fe9326),
	.w6(32'hbafa11da),
	.w7(32'h3bc2b95b),
	.w8(32'h3b5cc8de),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b603710),
	.w1(32'h39bbaea7),
	.w2(32'h3cbb5963),
	.w3(32'h3b2dd471),
	.w4(32'h3b862e22),
	.w5(32'hbb0ef5a9),
	.w6(32'h3bef24eb),
	.w7(32'hbb150b10),
	.w8(32'h3b41a86a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7184e),
	.w1(32'hbb2d1a8b),
	.w2(32'h3a839aa8),
	.w3(32'h39cdbc38),
	.w4(32'hba8d588a),
	.w5(32'hb92dcbbf),
	.w6(32'hbadf309a),
	.w7(32'hb8a392b1),
	.w8(32'hbacea96f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5ac10),
	.w1(32'hbb82a1c7),
	.w2(32'h3cccc356),
	.w3(32'hbc182fa5),
	.w4(32'h3b4e3c33),
	.w5(32'h3c2c5e69),
	.w6(32'hbb126ea4),
	.w7(32'hbbf637cb),
	.w8(32'h3be32fa9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf10cc1),
	.w1(32'h3a355cc7),
	.w2(32'h3b886c3b),
	.w3(32'h3b185fe2),
	.w4(32'h3a6f6fc6),
	.w5(32'hbb162c9c),
	.w6(32'hbaa88946),
	.w7(32'hbbcc6aaa),
	.w8(32'h3b262b33),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee217),
	.w1(32'h3a7d6351),
	.w2(32'h3acf5e23),
	.w3(32'h3bf72dc9),
	.w4(32'h3c27779b),
	.w5(32'hbab7aef5),
	.w6(32'h39c31060),
	.w7(32'h3b022663),
	.w8(32'hbc740be7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc928377),
	.w1(32'h3aebeb5f),
	.w2(32'h3c3f1280),
	.w3(32'hbb9c80e6),
	.w4(32'hbc1bc84e),
	.w5(32'h3b991a12),
	.w6(32'hbbbc2711),
	.w7(32'hbbdd902f),
	.w8(32'h39794bae),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce2844),
	.w1(32'h3b520a52),
	.w2(32'hbbbcf4b3),
	.w3(32'h3bd970c7),
	.w4(32'hbad7ffa2),
	.w5(32'h3c0330e1),
	.w6(32'hbb144f64),
	.w7(32'h3bf175cf),
	.w8(32'hbbb03ca6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb328a17),
	.w1(32'hba8ac887),
	.w2(32'h3b075c6b),
	.w3(32'hbab4e9de),
	.w4(32'hba38f2d7),
	.w5(32'h3c4cc1f7),
	.w6(32'hbadeaac3),
	.w7(32'hbd27569a),
	.w8(32'h3a16157a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb923416),
	.w1(32'hbb1202b8),
	.w2(32'hbadbecc4),
	.w3(32'hbb77f8bf),
	.w4(32'hbb1a6293),
	.w5(32'h3aa84588),
	.w6(32'hbb9e5131),
	.w7(32'h3ad8a94d),
	.w8(32'hb9b69aee),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87348da),
	.w1(32'h3ae78385),
	.w2(32'h3b29277c),
	.w3(32'hba907806),
	.w4(32'h3c906440),
	.w5(32'hbb184d8c),
	.w6(32'hbb89c39f),
	.w7(32'h3b84aa2e),
	.w8(32'h3bab7d0e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea5bef),
	.w1(32'hba7bf37e),
	.w2(32'hbbc07454),
	.w3(32'h3b74ba8d),
	.w4(32'h3abdc609),
	.w5(32'hbb3d8773),
	.w6(32'hbb33efdf),
	.w7(32'hbb1dff87),
	.w8(32'hbb2e6ef1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a936),
	.w1(32'hbb8626bc),
	.w2(32'hbb8131e1),
	.w3(32'hbaeb6174),
	.w4(32'hba3c9356),
	.w5(32'hba925a36),
	.w6(32'hbb199b32),
	.w7(32'h3bfc2998),
	.w8(32'h3ab191fa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b54c4),
	.w1(32'h3b9c84b6),
	.w2(32'h3afdcae6),
	.w3(32'hbb660a1b),
	.w4(32'h3bdb20fd),
	.w5(32'hbb287983),
	.w6(32'h3bf11b2a),
	.w7(32'hbba591de),
	.w8(32'hbb2b98fa),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef6a13),
	.w1(32'hbc482f75),
	.w2(32'h3bb28d47),
	.w3(32'h3b02bd4b),
	.w4(32'hbbdc6bb5),
	.w5(32'hbb66afa3),
	.w6(32'h39b48434),
	.w7(32'hbb88e9af),
	.w8(32'h3bed2edb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11dfc3),
	.w1(32'hbbb0ea47),
	.w2(32'hbb4fbabc),
	.w3(32'hbacc4987),
	.w4(32'hb9eca72d),
	.w5(32'hbb084d8a),
	.w6(32'hbb82df0b),
	.w7(32'hbab77796),
	.w8(32'h3b984533),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b602b85),
	.w1(32'h3b10d083),
	.w2(32'hbc0aa7e7),
	.w3(32'hba84bff7),
	.w4(32'h3c13a18b),
	.w5(32'hbb2db3dd),
	.w6(32'h3da588ce),
	.w7(32'hbbddabb8),
	.w8(32'hbb1682f0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb7a54),
	.w1(32'hb9e86c23),
	.w2(32'hbbbaba1b),
	.w3(32'hbb0133d0),
	.w4(32'hbbd201df),
	.w5(32'h3d000e63),
	.w6(32'hba09b840),
	.w7(32'hbbd0217a),
	.w8(32'hbbefb994),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b703e6e),
	.w1(32'h3a05da5d),
	.w2(32'hbb691ccf),
	.w3(32'h3bade7dd),
	.w4(32'hbb59686a),
	.w5(32'h3b2dc5be),
	.w6(32'h3aa085e0),
	.w7(32'h3ba7230c),
	.w8(32'h3b29628b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd6701),
	.w1(32'hbc04f200),
	.w2(32'h3b58d96c),
	.w3(32'h3b302936),
	.w4(32'h3b334084),
	.w5(32'hba7ac1eb),
	.w6(32'hbb1cb65d),
	.w7(32'hbc330687),
	.w8(32'hbbdb1d77),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb537dff),
	.w1(32'h3aff5435),
	.w2(32'h3ad40006),
	.w3(32'hbb7b6234),
	.w4(32'h39989e12),
	.w5(32'h3bbce62f),
	.w6(32'hbbcd940f),
	.w7(32'hbbb513b2),
	.w8(32'h3bc281d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3425d448),
	.w1(32'hbb9ddcc1),
	.w2(32'h3a04eb12),
	.w3(32'h3a062274),
	.w4(32'hbc038d78),
	.w5(32'hbb60be59),
	.w6(32'h39c97237),
	.w7(32'hbb90a620),
	.w8(32'hbb319b4d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa50882),
	.w1(32'h3b1016d7),
	.w2(32'hbb648652),
	.w3(32'hba470d6a),
	.w4(32'h3ccd87a4),
	.w5(32'h3abcb8db),
	.w6(32'hbc0f96d2),
	.w7(32'hbb69befc),
	.w8(32'hb7d374e1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61e40b),
	.w1(32'hbc1212bc),
	.w2(32'hbbaea8ec),
	.w3(32'hb99cd810),
	.w4(32'hb917047b),
	.w5(32'hbc24fae1),
	.w6(32'h3b4a16c9),
	.w7(32'hbbc1cf6f),
	.w8(32'h3ad6d84b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c2ac8),
	.w1(32'h3c23661c),
	.w2(32'hbb50b1ef),
	.w3(32'hbb3b63b8),
	.w4(32'hbc19016c),
	.w5(32'hbb748116),
	.w6(32'hba09043c),
	.w7(32'h3d899d2c),
	.w8(32'h3b0a7f85),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5319c1),
	.w1(32'h3c19ae79),
	.w2(32'h39a50cb5),
	.w3(32'h3b1a7552),
	.w4(32'hbba39aa1),
	.w5(32'h3cee3f92),
	.w6(32'h3bbaf754),
	.w7(32'hb9cbbedb),
	.w8(32'h3af87883),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c506f),
	.w1(32'hbb4443aa),
	.w2(32'hbb05e8fa),
	.w3(32'hba0fabbe),
	.w4(32'hbb3a32cd),
	.w5(32'h3b3449cf),
	.w6(32'hbcdee312),
	.w7(32'hbab86f9f),
	.w8(32'h3b5a9685),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a856a),
	.w1(32'hbaf06525),
	.w2(32'hbb916314),
	.w3(32'h3b8b7fa4),
	.w4(32'h3b84ce6f),
	.w5(32'h3c3bd757),
	.w6(32'h3a9d12c4),
	.w7(32'hbb55c7fc),
	.w8(32'h3b1e01ae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca5aa),
	.w1(32'hbc0dd126),
	.w2(32'hbc0629f5),
	.w3(32'hbca01450),
	.w4(32'hbb5e65ab),
	.w5(32'hbc0ad330),
	.w6(32'hbbb62e17),
	.w7(32'hbc5ef071),
	.w8(32'h3bc7539b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e275),
	.w1(32'hbb66a739),
	.w2(32'h3d344252),
	.w3(32'hbb79b017),
	.w4(32'h389d7d22),
	.w5(32'hbc391921),
	.w6(32'h3aa4367a),
	.w7(32'hbbeb03e7),
	.w8(32'hb9eeaf70),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b1210),
	.w1(32'hbaf36afa),
	.w2(32'h3b0d1b01),
	.w3(32'h3b8e9c2e),
	.w4(32'hbb077d8b),
	.w5(32'h3bd20f9c),
	.w6(32'h39adcef6),
	.w7(32'h39c1b205),
	.w8(32'hba87c8a9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1b654),
	.w1(32'hbb179b6a),
	.w2(32'hbb4fdd2d),
	.w3(32'hbb1a79bb),
	.w4(32'hbba32a75),
	.w5(32'h38376ea9),
	.w6(32'hbb0cdaea),
	.w7(32'hbaa2289c),
	.w8(32'hbb5a0ba0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9693e8),
	.w1(32'hbb3c79c5),
	.w2(32'hbaa0c135),
	.w3(32'hbcf4f72e),
	.w4(32'hbb993fe9),
	.w5(32'h3be2f230),
	.w6(32'hbc24b405),
	.w7(32'hbb8966e7),
	.w8(32'hbb6da804),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4cd06),
	.w1(32'hbbd4372c),
	.w2(32'hbb83df3c),
	.w3(32'h3b04d39d),
	.w4(32'h3a90d63c),
	.w5(32'hbbace418),
	.w6(32'hbb7525ac),
	.w7(32'h39a738ab),
	.w8(32'h3ba03a09),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf88769),
	.w1(32'hbb249bbc),
	.w2(32'hbc8648b9),
	.w3(32'hbac8503d),
	.w4(32'hbb978b17),
	.w5(32'h3b3415b8),
	.w6(32'hbbc7b413),
	.w7(32'hbb648138),
	.w8(32'h3c1eadfe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55290f),
	.w1(32'hbaa0f7a6),
	.w2(32'hbb60791b),
	.w3(32'hbbcd5202),
	.w4(32'h3befb266),
	.w5(32'h3ae2f5cd),
	.w6(32'hbb27794d),
	.w7(32'hbb4a94a9),
	.w8(32'h3a7384d4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8163b),
	.w1(32'h3ae4577e),
	.w2(32'hbb6b00a7),
	.w3(32'hbbf90d64),
	.w4(32'hbb250bc3),
	.w5(32'hbbd45497),
	.w6(32'h3aa7b120),
	.w7(32'h3aae23ce),
	.w8(32'hbb9bb103),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c431b80),
	.w1(32'hbb36348d),
	.w2(32'hbb39e328),
	.w3(32'h3728b79b),
	.w4(32'h3ab12ce7),
	.w5(32'h3ae816dd),
	.w6(32'hbc990cfa),
	.w7(32'hbb8441b4),
	.w8(32'h3b31566c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9838a3),
	.w1(32'h3bb51bfa),
	.w2(32'hba780ce0),
	.w3(32'h3cb1e596),
	.w4(32'h3b76bf1c),
	.w5(32'hba490f67),
	.w6(32'hbb152a09),
	.w7(32'hbae893b9),
	.w8(32'h3d3a2b2b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33837d),
	.w1(32'hba9b0eb7),
	.w2(32'hbacd0d73),
	.w3(32'hb919c783),
	.w4(32'hb9be3fa1),
	.w5(32'h3b079f9e),
	.w6(32'h3a9d4bb0),
	.w7(32'hbaa8c370),
	.w8(32'h3b96d513),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9476ae6),
	.w1(32'h3c4be29f),
	.w2(32'h3b16a58f),
	.w3(32'hbafb1246),
	.w4(32'hbaa860fe),
	.w5(32'h3a3cd9ff),
	.w6(32'hba7726da),
	.w7(32'h3bf79b35),
	.w8(32'h39fc484a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2791),
	.w1(32'h3c15ba04),
	.w2(32'h3a65a75d),
	.w3(32'hbbb4be63),
	.w4(32'h3a222aa9),
	.w5(32'h3b2d4d64),
	.w6(32'hbac63aff),
	.w7(32'hbb5d2e5f),
	.w8(32'hbb906a1f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14898a),
	.w1(32'hbb330e8d),
	.w2(32'hbafc7502),
	.w3(32'hbb53974f),
	.w4(32'h3a506dd4),
	.w5(32'hbc7d64d1),
	.w6(32'hbb644198),
	.w7(32'h394a0f44),
	.w8(32'h3ab8b5e2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a445227),
	.w1(32'h3b0d0cf5),
	.w2(32'h3c45df7c),
	.w3(32'h3a64f637),
	.w4(32'h3a9b38e9),
	.w5(32'h3b06a63f),
	.w6(32'hbb270e02),
	.w7(32'h3b4bad66),
	.w8(32'h392d809e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b1f2b),
	.w1(32'h3c00a186),
	.w2(32'hbadcf2e0),
	.w3(32'hbab3cb93),
	.w4(32'hbbebeb9a),
	.w5(32'hbb925bcf),
	.w6(32'hbabf07c5),
	.w7(32'hbb81173e),
	.w8(32'hbbe21bab),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aeffd),
	.w1(32'h3a1795ab),
	.w2(32'hba9b0094),
	.w3(32'hbb3df95c),
	.w4(32'hbb29edf9),
	.w5(32'h3ba0d156),
	.w6(32'h3b3c4597),
	.w7(32'h3b923a41),
	.w8(32'h3c3c8fe4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba978542),
	.w1(32'h3b2481de),
	.w2(32'hbb0a414f),
	.w3(32'hbb5998b4),
	.w4(32'hb9fcd727),
	.w5(32'hb78204d5),
	.w6(32'hbc839b43),
	.w7(32'h3a892373),
	.w8(32'hbbb0c046),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d7056),
	.w1(32'h3af8d233),
	.w2(32'hbb109f84),
	.w3(32'hbb0a2cf5),
	.w4(32'h3c624a82),
	.w5(32'hbb2b1264),
	.w6(32'hba65b6ea),
	.w7(32'h3b1847aa),
	.w8(32'h3b03cbfd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60aaf0),
	.w1(32'hbc2232b8),
	.w2(32'h3cd6eb92),
	.w3(32'hbad9fa4a),
	.w4(32'h3b2dfd82),
	.w5(32'hbbb424df),
	.w6(32'h3a25a2d2),
	.w7(32'hb8b95217),
	.w8(32'h3cc6a619),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba049118),
	.w1(32'hbb475927),
	.w2(32'hb7d18011),
	.w3(32'hbafd4c34),
	.w4(32'hba0e53d6),
	.w5(32'h3c33efa6),
	.w6(32'hbb057ae6),
	.w7(32'hbbf52a98),
	.w8(32'hba951f95),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f40e8),
	.w1(32'h3a7f9f7a),
	.w2(32'h3bb3ffa8),
	.w3(32'hbb0b07c8),
	.w4(32'h3bc8488c),
	.w5(32'hba93b70a),
	.w6(32'h3a8e204e),
	.w7(32'h3bd69129),
	.w8(32'hbcf42ddc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f8bdb),
	.w1(32'h3bea95fe),
	.w2(32'h3a3eead3),
	.w3(32'h3ba12048),
	.w4(32'hbcd84cae),
	.w5(32'h3a49c8af),
	.w6(32'hbb64c16b),
	.w7(32'h3b86cfb0),
	.w8(32'h3a22a373),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4c333),
	.w1(32'h3b03230c),
	.w2(32'hba91293c),
	.w3(32'h3ac5c263),
	.w4(32'hbbf8eeb7),
	.w5(32'hbb06b631),
	.w6(32'hbb1bad3a),
	.w7(32'hbab593dd),
	.w8(32'hb9a31542),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5072c9),
	.w1(32'hbafe88b8),
	.w2(32'hbae5b680),
	.w3(32'h3ac326ea),
	.w4(32'hbb2f4f14),
	.w5(32'hbd00199e),
	.w6(32'h3b317811),
	.w7(32'h3b08ad18),
	.w8(32'h390d51af),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb539cec),
	.w1(32'hba4a1c0d),
	.w2(32'h3c1d34a1),
	.w3(32'hb969350e),
	.w4(32'hbb40a41b),
	.w5(32'hbb9a2fad),
	.w6(32'hbc9ed43e),
	.w7(32'h3b803191),
	.w8(32'hb9a7b66e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252ad6),
	.w1(32'h3af359b0),
	.w2(32'hb6d3ed35),
	.w3(32'h3abea735),
	.w4(32'hbcb8dd5b),
	.w5(32'h3a788523),
	.w6(32'h3d1f92f9),
	.w7(32'h3c6ac290),
	.w8(32'hba4a2ce4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3526),
	.w1(32'hba64d71a),
	.w2(32'h3b159ea7),
	.w3(32'hbad38802),
	.w4(32'hbb33af38),
	.w5(32'h3ac5c8b3),
	.w6(32'h3c4c9afd),
	.w7(32'hba1f243f),
	.w8(32'h3c9c5623),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948b3a),
	.w1(32'h3c528bb0),
	.w2(32'hba01ddac),
	.w3(32'hbb983b6b),
	.w4(32'hbb8e01a9),
	.w5(32'hbb17efff),
	.w6(32'hbbf445f6),
	.w7(32'hbbbb2504),
	.w8(32'hbc171d25),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93076f),
	.w1(32'hbb73cb0c),
	.w2(32'hba6687a2),
	.w3(32'hbc14a036),
	.w4(32'h396153f5),
	.w5(32'hb9a632eb),
	.w6(32'h3af93da4),
	.w7(32'h3c3f8fc9),
	.w8(32'hba93c5ec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39729c80),
	.w1(32'hba20f0cc),
	.w2(32'h39abed91),
	.w3(32'hb9740af8),
	.w4(32'h39f04659),
	.w5(32'hbb0b6775),
	.w6(32'h3b0d18b1),
	.w7(32'h3aee8ab9),
	.w8(32'h3b1d2c25),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1ffe1),
	.w1(32'hbb3213aa),
	.w2(32'h3c78b2d3),
	.w3(32'hba562aad),
	.w4(32'h3b8cda26),
	.w5(32'hbb34272b),
	.w6(32'hb9807158),
	.w7(32'hbc3f7a2d),
	.w8(32'hbbb12888),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7da5c),
	.w1(32'h3a9ffa1f),
	.w2(32'h3b20479f),
	.w3(32'hbc0dbaed),
	.w4(32'hbb02329c),
	.w5(32'hbb5020ba),
	.w6(32'hbb688941),
	.w7(32'hba5ce962),
	.w8(32'hb9e0a637),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba06a80),
	.w1(32'h3ad1ceac),
	.w2(32'hbb38f3ad),
	.w3(32'h39223219),
	.w4(32'hba6b956e),
	.w5(32'h3a388233),
	.w6(32'hbb0c607f),
	.w7(32'hbb1d0e13),
	.w8(32'hb9cccb9f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b639212),
	.w1(32'hbc4b8cce),
	.w2(32'hb93468c4),
	.w3(32'hbc09a677),
	.w4(32'hb96173ae),
	.w5(32'h398d7203),
	.w6(32'h3b97d229),
	.w7(32'h39be7fd7),
	.w8(32'h3b3f713f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed5f6),
	.w1(32'h3a8b5445),
	.w2(32'h3af1b58b),
	.w3(32'hbb12c82e),
	.w4(32'h3a8980ef),
	.w5(32'hb70082d8),
	.w6(32'hbb15c783),
	.w7(32'hba7808ab),
	.w8(32'hbb042698),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ef4f),
	.w1(32'h3ab5734e),
	.w2(32'h3cea221f),
	.w3(32'hb9dce4f0),
	.w4(32'hbbc2d5c5),
	.w5(32'hba428aed),
	.w6(32'hbba0a2cd),
	.w7(32'hbaaf7ad8),
	.w8(32'hbac6be13),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877620),
	.w1(32'hb87c772e),
	.w2(32'hba2c3b83),
	.w3(32'hbb369297),
	.w4(32'hbabb6437),
	.w5(32'h3aec1faa),
	.w6(32'hb81e06e6),
	.w7(32'hbcad1e87),
	.w8(32'h3a691f3a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2059f5),
	.w1(32'hbcc12f6c),
	.w2(32'h3b2c9498),
	.w3(32'hb94a604e),
	.w4(32'h3a4a0c45),
	.w5(32'h3afd2f4f),
	.w6(32'h3b378346),
	.w7(32'h3a04b5c7),
	.w8(32'h3aa2c80e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0813f),
	.w1(32'h3b5ec857),
	.w2(32'h395cd948),
	.w3(32'hba32bc3c),
	.w4(32'h3a3a6033),
	.w5(32'hbb7aacfa),
	.w6(32'hba9cab39),
	.w7(32'hbc09c48b),
	.w8(32'hbba0345a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3324),
	.w1(32'h3907940f),
	.w2(32'h39018245),
	.w3(32'h39b818a4),
	.w4(32'hbb980ced),
	.w5(32'hbaad2be3),
	.w6(32'hba02f394),
	.w7(32'h3a8341fc),
	.w8(32'h3b4552af),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995fdc),
	.w1(32'h3ac25058),
	.w2(32'hbabfbc0b),
	.w3(32'hbb7f93b6),
	.w4(32'hbad11d96),
	.w5(32'hb8b1e8e6),
	.w6(32'hbbf0981e),
	.w7(32'hbb36083a),
	.w8(32'hbbad2822),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fcf451),
	.w1(32'h3aabff8f),
	.w2(32'hba9c816c),
	.w3(32'h3a80b925),
	.w4(32'h3acf5081),
	.w5(32'hba3879eb),
	.w6(32'hbc056220),
	.w7(32'hbc072fb5),
	.w8(32'hb9cb0785),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4df3f),
	.w1(32'hba451f9a),
	.w2(32'hbb6eda4f),
	.w3(32'h3b8e9ab0),
	.w4(32'h3b82dc84),
	.w5(32'h3b5db45d),
	.w6(32'hba979b64),
	.w7(32'hbb887d25),
	.w8(32'hbb026f7b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abec828),
	.w1(32'hb99a5850),
	.w2(32'h3b418829),
	.w3(32'h3c4e1b52),
	.w4(32'hbb08e2bc),
	.w5(32'hbadf0aeb),
	.w6(32'h3c0e9cd0),
	.w7(32'h3ab92f3e),
	.w8(32'h3b4f7d5c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da0fe),
	.w1(32'hbc0c759a),
	.w2(32'h3ca7b5a5),
	.w3(32'h3ad41e0a),
	.w4(32'h3a4fefa1),
	.w5(32'hba8e4081),
	.w6(32'h3ac7cb3d),
	.w7(32'hbb19c28d),
	.w8(32'h3ac58f96),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4d32f),
	.w1(32'h3a8a74f0),
	.w2(32'h395c5bcb),
	.w3(32'h3b12faee),
	.w4(32'h3ab92488),
	.w5(32'h3acdb820),
	.w6(32'h3aff40af),
	.w7(32'h3b81b89b),
	.w8(32'hbb9bf81c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977f6b2),
	.w1(32'h3aabd029),
	.w2(32'h3a1786e9),
	.w3(32'h39f78116),
	.w4(32'h395edee8),
	.w5(32'h3ba78233),
	.w6(32'hba9f5cf7),
	.w7(32'h3a78bc3a),
	.w8(32'h38f91f6a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87b307),
	.w1(32'hbca4f847),
	.w2(32'h3a8fd0d7),
	.w3(32'hbd02de3d),
	.w4(32'h39993d25),
	.w5(32'h3bbf915b),
	.w6(32'hb92e5b09),
	.w7(32'h3973e4ac),
	.w8(32'hb7a11761),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab87a80),
	.w1(32'h3b094b57),
	.w2(32'hba7df25e),
	.w3(32'hb981d8e4),
	.w4(32'hbaf1c537),
	.w5(32'hb9b33164),
	.w6(32'h3a0a2707),
	.w7(32'hba487b44),
	.w8(32'h3ba66da2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22925c),
	.w1(32'h3d0955ca),
	.w2(32'hba429f74),
	.w3(32'h3be390e3),
	.w4(32'h3a11926f),
	.w5(32'hbc05b488),
	.w6(32'h3a87e6cd),
	.w7(32'h3b207bab),
	.w8(32'h3cad2049),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1d5a),
	.w1(32'hbbc01af4),
	.w2(32'hbbf6af5b),
	.w3(32'hbbb69929),
	.w4(32'hbaf14dfc),
	.w5(32'h3a90e4d4),
	.w6(32'hbbf73e20),
	.w7(32'hbb56f4a9),
	.w8(32'hbb53b8ad),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84877b),
	.w1(32'hbb597298),
	.w2(32'h3ac35bdf),
	.w3(32'h3c0ab142),
	.w4(32'h3bb3f720),
	.w5(32'h3af7306f),
	.w6(32'h3bb57dcc),
	.w7(32'h3b7d1223),
	.w8(32'h3b1183eb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90954e),
	.w1(32'hbadafb6c),
	.w2(32'h3d01d0a4),
	.w3(32'h3b25d217),
	.w4(32'hbb416915),
	.w5(32'hb9607874),
	.w6(32'h3cdad867),
	.w7(32'h3b4634f9),
	.w8(32'hb96e8dab),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82ba08),
	.w1(32'hbb2577f8),
	.w2(32'hbcf48a86),
	.w3(32'hbc578e15),
	.w4(32'h3b2ee145),
	.w5(32'hbaaf0619),
	.w6(32'h3a806362),
	.w7(32'h3ac7fca6),
	.w8(32'hbc0f7aa5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc891fee),
	.w1(32'h3b850cfa),
	.w2(32'hbc4a52c4),
	.w3(32'hb7ab0d3b),
	.w4(32'h39fc9e4e),
	.w5(32'h3b0826fa),
	.w6(32'hb8f82455),
	.w7(32'hbad6597e),
	.w8(32'hbad9c922),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44d8e2),
	.w1(32'hbcbb6f38),
	.w2(32'hbbbdf6f1),
	.w3(32'hbb07180f),
	.w4(32'hba5db7f3),
	.w5(32'h3affcf51),
	.w6(32'hbbe9cdc6),
	.w7(32'hbbd9dc5e),
	.w8(32'hbbdb7981),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a06b1),
	.w1(32'hbb6f24fe),
	.w2(32'hbae26bab),
	.w3(32'h3a771968),
	.w4(32'hb9d8db03),
	.w5(32'h3adebd3c),
	.w6(32'hba225c2d),
	.w7(32'hbb411452),
	.w8(32'h3a1f84dd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4cab),
	.w1(32'h3c01dd88),
	.w2(32'hbae16fac),
	.w3(32'h3a147ec8),
	.w4(32'h38b8854a),
	.w5(32'h39894444),
	.w6(32'h3a93cb26),
	.w7(32'hba9e37d9),
	.w8(32'hb949166a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018a23),
	.w1(32'hbaa892ad),
	.w2(32'h39dac077),
	.w3(32'hb9c145cd),
	.w4(32'h3a8bb1e8),
	.w5(32'hba8d1039),
	.w6(32'h39a9b498),
	.w7(32'hbabd755a),
	.w8(32'h3b80cd28),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f127f),
	.w1(32'hbb452805),
	.w2(32'h3b01c272),
	.w3(32'hbc960c58),
	.w4(32'hba9ec15c),
	.w5(32'hbb50b395),
	.w6(32'hb973a88e),
	.w7(32'hbaae655a),
	.w8(32'hba890f31),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990b81e),
	.w1(32'h3812d74c),
	.w2(32'hb9cef101),
	.w3(32'h387eb3fd),
	.w4(32'hbaeaa97b),
	.w5(32'hba84499b),
	.w6(32'hba38c50a),
	.w7(32'h3a80614f),
	.w8(32'h3a0bc138),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a107489),
	.w1(32'h3a30c803),
	.w2(32'hbb1c0408),
	.w3(32'h3a816a94),
	.w4(32'h3adcd599),
	.w5(32'hba43c049),
	.w6(32'hba85e714),
	.w7(32'h3a723504),
	.w8(32'hbb4e7283),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56041f),
	.w1(32'h3a4ae460),
	.w2(32'h3b10cf04),
	.w3(32'h3af5a64a),
	.w4(32'h3a1f9c57),
	.w5(32'hb994519f),
	.w6(32'h3b1b4081),
	.w7(32'h3a9cf76f),
	.w8(32'hb929bfe9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0a4e),
	.w1(32'h3b6efc97),
	.w2(32'hba946eaf),
	.w3(32'h3ae47798),
	.w4(32'h38112ca5),
	.w5(32'hbb435549),
	.w6(32'hba865e41),
	.w7(32'hb9ffbd3f),
	.w8(32'hbc56bf1c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919eb1),
	.w1(32'hbaa2166f),
	.w2(32'h38421e66),
	.w3(32'h3b8a1867),
	.w4(32'hbb3b50d5),
	.w5(32'h386178ed),
	.w6(32'hbaf74810),
	.w7(32'hba0930b8),
	.w8(32'h3a4f8fe5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e350c9),
	.w1(32'hbb990874),
	.w2(32'h3afafb19),
	.w3(32'h3b3f956c),
	.w4(32'hbac99134),
	.w5(32'h3a2d0ef3),
	.w6(32'h3bd5ce94),
	.w7(32'hba8e8ff4),
	.w8(32'h3ba1fa7e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943af53),
	.w1(32'h3ba7da4c),
	.w2(32'h3bfd625a),
	.w3(32'hb961def6),
	.w4(32'hb83c43c2),
	.w5(32'hba457c33),
	.w6(32'hbb2c73d1),
	.w7(32'h3985c1aa),
	.w8(32'hba9982bb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b10c4),
	.w1(32'h3a02c556),
	.w2(32'h3b4a230d),
	.w3(32'h3b582a93),
	.w4(32'h3b9a23e4),
	.w5(32'h3aa37c7a),
	.w6(32'h3bc2bc50),
	.w7(32'h3af4e801),
	.w8(32'hbb2b1e01),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7ceef),
	.w1(32'hba942f40),
	.w2(32'hbb81c100),
	.w3(32'h3c020b77),
	.w4(32'hbb2ff456),
	.w5(32'h3b4dc056),
	.w6(32'hbabcdc03),
	.w7(32'hbb0991fe),
	.w8(32'h3be8ae81),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b678347),
	.w1(32'hbae81f49),
	.w2(32'h3b978f2c),
	.w3(32'h3b0ce24c),
	.w4(32'hbae02a57),
	.w5(32'hbb44443e),
	.w6(32'hbb4031df),
	.w7(32'hb848dd55),
	.w8(32'h3a128c58),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9c46c),
	.w1(32'hba1fd9b8),
	.w2(32'hba3c97e6),
	.w3(32'hb9481c43),
	.w4(32'hbb26455c),
	.w5(32'h3aa4b962),
	.w6(32'h3b095ff7),
	.w7(32'hbaa7d779),
	.w8(32'hbb334a60),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0a9a3),
	.w1(32'hbb0bbf5f),
	.w2(32'h398e1d3a),
	.w3(32'hba7453d6),
	.w4(32'h3b69db5f),
	.w5(32'hbb2cb124),
	.w6(32'hbc04d19c),
	.w7(32'h3cb97c89),
	.w8(32'h3b1ff075),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6107e),
	.w1(32'h3aed0e05),
	.w2(32'hba06c9c8),
	.w3(32'hb7c4ab7c),
	.w4(32'hbaed4056),
	.w5(32'hbb4d9811),
	.w6(32'hba978291),
	.w7(32'hbae8a662),
	.w8(32'hbb356538),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49710f),
	.w1(32'h3b591109),
	.w2(32'h38fee7b3),
	.w3(32'h3c89946e),
	.w4(32'h3c44c0a0),
	.w5(32'h3c1039a0),
	.w6(32'h3ab9647e),
	.w7(32'h3a5eaefe),
	.w8(32'hbaf1d9cb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b5d2),
	.w1(32'hbc0720f6),
	.w2(32'h3c1a25bc),
	.w3(32'hb8a5ef69),
	.w4(32'hb98ccc41),
	.w5(32'h3bb75a73),
	.w6(32'hb98798ef),
	.w7(32'hba54c4d6),
	.w8(32'hbb7663a2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cc2d4),
	.w1(32'h3a1fa890),
	.w2(32'hba7d49b5),
	.w3(32'hbae5e02c),
	.w4(32'hb9a883c8),
	.w5(32'hbb5a9895),
	.w6(32'hbb4cd083),
	.w7(32'hbbba677c),
	.w8(32'h395d8077),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb221af8),
	.w1(32'hb53713a4),
	.w2(32'h3ab3dc47),
	.w3(32'h3b0221b6),
	.w4(32'h3b96927c),
	.w5(32'hb813b51b),
	.w6(32'hbbea0875),
	.w7(32'h38743e8c),
	.w8(32'h38915f38),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f49ef),
	.w1(32'h36f9efdf),
	.w2(32'hb9ba1fc8),
	.w3(32'hbacf6dfd),
	.w4(32'h3a0dfe57),
	.w5(32'h3c32acb6),
	.w6(32'h3a5179b5),
	.w7(32'hbaec4be8),
	.w8(32'hbb9c4eac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038442),
	.w1(32'h3b2c800f),
	.w2(32'hbb8ca44b),
	.w3(32'hbb6eea19),
	.w4(32'h3babda55),
	.w5(32'hbc143b8f),
	.w6(32'hbc04e4db),
	.w7(32'h3b61a935),
	.w8(32'hbaa2dafd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af731c6),
	.w1(32'hbb4f93bf),
	.w2(32'h3a97a497),
	.w3(32'h3ab1fb94),
	.w4(32'hbae699f3),
	.w5(32'h3abc9d56),
	.w6(32'h3a129795),
	.w7(32'hbb5269eb),
	.w8(32'h3c85e1cb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6c82b),
	.w1(32'hbaa23740),
	.w2(32'h3ca6d32a),
	.w3(32'hbacf1433),
	.w4(32'h3af9205f),
	.w5(32'h3aa1d408),
	.w6(32'hba8e98bd),
	.w7(32'h3b51dd59),
	.w8(32'hbb4321f2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae54fce),
	.w1(32'h3aaf6077),
	.w2(32'hba01156a),
	.w3(32'h3c41bcce),
	.w4(32'h3a9d7be8),
	.w5(32'hbb40b514),
	.w6(32'hba0825e1),
	.w7(32'hbc434d95),
	.w8(32'hba015d0d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb696574),
	.w1(32'h3be99d61),
	.w2(32'hb9ce4a15),
	.w3(32'hbbcc5500),
	.w4(32'hbb84d73e),
	.w5(32'h3b44d238),
	.w6(32'h3b45c54b),
	.w7(32'h39c0ecaa),
	.w8(32'h3b66e1c5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb401964),
	.w1(32'hbb0f0d48),
	.w2(32'h3a39f8ee),
	.w3(32'h3af3f04c),
	.w4(32'h3bd3d24c),
	.w5(32'hbaa01823),
	.w6(32'h3b202cd6),
	.w7(32'hba1f9be0),
	.w8(32'h3b3c5103),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a7e3),
	.w1(32'h3b7fbf62),
	.w2(32'h3b8bc697),
	.w3(32'h3ba22c41),
	.w4(32'h39ccebfb),
	.w5(32'h3b23c938),
	.w6(32'hbc017104),
	.w7(32'hbad18b51),
	.w8(32'h3b1fc14b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7af8f),
	.w1(32'hbb718cd8),
	.w2(32'hbb912a1b),
	.w3(32'hbbba0371),
	.w4(32'hbc62c6f9),
	.w5(32'hbb709d65),
	.w6(32'hbbc03996),
	.w7(32'hbaf1a23c),
	.w8(32'hbae14693),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a045b85),
	.w1(32'hba5a28ff),
	.w2(32'hbacd0f17),
	.w3(32'h3b1020a0),
	.w4(32'h3a42eb1b),
	.w5(32'hbb065a3b),
	.w6(32'h3adbb508),
	.w7(32'h399374e3),
	.w8(32'h3b62787b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370ce1bf),
	.w1(32'h39f4c73d),
	.w2(32'h3a699f58),
	.w3(32'h3980aed4),
	.w4(32'h3c3d803d),
	.w5(32'h3acde632),
	.w6(32'hba31efdf),
	.w7(32'hbc230a69),
	.w8(32'h3b7fde7b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3d62c),
	.w1(32'hba3255f3),
	.w2(32'h3a96f80e),
	.w3(32'hbbb3cf5b),
	.w4(32'hba89a372),
	.w5(32'h3b1d3029),
	.w6(32'hbb77631b),
	.w7(32'hbb6314dd),
	.w8(32'h3b45eac6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac072d8),
	.w1(32'hbab37cba),
	.w2(32'h39af9b4f),
	.w3(32'h39a18cf6),
	.w4(32'h3b59aa7d),
	.w5(32'h3b017996),
	.w6(32'hbace8445),
	.w7(32'h3ad27279),
	.w8(32'h39f9b82d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7ae8d),
	.w1(32'hba99cadb),
	.w2(32'hb84a14f4),
	.w3(32'h3a7942ad),
	.w4(32'hbab24f6a),
	.w5(32'hbac3c9d6),
	.w6(32'hbaf0268c),
	.w7(32'h3aa07f43),
	.w8(32'hbabd7318),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596a93),
	.w1(32'h3b85314a),
	.w2(32'h3963731b),
	.w3(32'h3ad19b0b),
	.w4(32'hbb18f9e9),
	.w5(32'hbb77db9f),
	.w6(32'h3a4a84bd),
	.w7(32'h388b3d7f),
	.w8(32'hbb1096f2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae428dd),
	.w1(32'h3cea1b30),
	.w2(32'hbaae5c71),
	.w3(32'h3c0ac18e),
	.w4(32'h3c047cb5),
	.w5(32'h3a452bdd),
	.w6(32'h3c0a5880),
	.w7(32'hbd39e33b),
	.w8(32'h3b0f8cdc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e05b),
	.w1(32'h3af1b116),
	.w2(32'hbb4d96ff),
	.w3(32'hba5ae565),
	.w4(32'h3d403c3a),
	.w5(32'h3b25e8e4),
	.w6(32'hbad53fad),
	.w7(32'hbbce55d8),
	.w8(32'h3b29cdc2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb682bf3),
	.w1(32'h3aade924),
	.w2(32'hba7e604f),
	.w3(32'hbb5a543e),
	.w4(32'h3b8b2d4f),
	.w5(32'hba55a4fd),
	.w6(32'h3d4c5348),
	.w7(32'h3b009c5a),
	.w8(32'hbb58b85f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8808e6),
	.w1(32'h3a931e10),
	.w2(32'h3cdf6fec),
	.w3(32'hbab7b825),
	.w4(32'hbc146fb1),
	.w5(32'hbafaeb30),
	.w6(32'h3b103dea),
	.w7(32'hbb04652a),
	.w8(32'h3ae4b441),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa9fdd),
	.w1(32'hbb559beb),
	.w2(32'h3b280eda),
	.w3(32'hba15155a),
	.w4(32'hbb0348fa),
	.w5(32'hba84e2a3),
	.w6(32'h3b19dbe1),
	.w7(32'hbbb2498a),
	.w8(32'hba1ab71e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8433688),
	.w1(32'hbb95ab47),
	.w2(32'h3b9d20cb),
	.w3(32'h3c2c3b34),
	.w4(32'h3ac35380),
	.w5(32'hbba62386),
	.w6(32'h3b052e57),
	.w7(32'hbbe8578e),
	.w8(32'hbb3c5049),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8418),
	.w1(32'hbc093543),
	.w2(32'h3ac0d842),
	.w3(32'h3a8250e2),
	.w4(32'h3b50bec2),
	.w5(32'h3b84a7b4),
	.w6(32'hbb536485),
	.w7(32'hbaee750b),
	.w8(32'hba880b8c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc64d1),
	.w1(32'hbb0ce270),
	.w2(32'hbc0f0c61),
	.w3(32'hbb697cae),
	.w4(32'h3a5aaaa8),
	.w5(32'h365b55a3),
	.w6(32'hba21b03f),
	.w7(32'h3b79c05b),
	.w8(32'hbb2d9a8a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79df25),
	.w1(32'hbb909eac),
	.w2(32'h3abfd73c),
	.w3(32'hba5f348b),
	.w4(32'hbaaa2d0c),
	.w5(32'hbbe45602),
	.w6(32'h3ba03dc8),
	.w7(32'hba4e7022),
	.w8(32'h3be06f95),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a01ee),
	.w1(32'h3a8eb853),
	.w2(32'h36e28901),
	.w3(32'hba92ebe5),
	.w4(32'h39ece5c1),
	.w5(32'hba781d3e),
	.w6(32'h3c7a698e),
	.w7(32'hbd108628),
	.w8(32'h3bac7505),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b552b),
	.w1(32'hba882df7),
	.w2(32'hb8b1b505),
	.w3(32'hba95a2d0),
	.w4(32'hbb2255d4),
	.w5(32'h3c7eab95),
	.w6(32'h3bdfcfc1),
	.w7(32'hbb1d45d5),
	.w8(32'h3ac4b8a7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e0ac),
	.w1(32'h390ce3e4),
	.w2(32'hbb8f3f86),
	.w3(32'hb9c4b7ef),
	.w4(32'h3a08efda),
	.w5(32'hbae81155),
	.w6(32'hbad276d3),
	.w7(32'hb9c91730),
	.w8(32'hbaac1960),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d482c2f),
	.w1(32'hba7d5aa5),
	.w2(32'h3c0e83dd),
	.w3(32'h396be5f7),
	.w4(32'h3a33f11e),
	.w5(32'hb8f67572),
	.w6(32'h3d1ed29b),
	.w7(32'hb9e824eb),
	.w8(32'h3b72f309),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960387d),
	.w1(32'hba95f7c5),
	.w2(32'hb88a151e),
	.w3(32'hbac4b377),
	.w4(32'hbbae177f),
	.w5(32'hbaaa0e8b),
	.w6(32'hbb10cdd2),
	.w7(32'hbb07d55b),
	.w8(32'hbb9fb0f7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35040),
	.w1(32'h3b64be0c),
	.w2(32'hbc2acebf),
	.w3(32'h3aeaea7e),
	.w4(32'hbc0d5ea3),
	.w5(32'hbd0e82be),
	.w6(32'hbd0cec6d),
	.w7(32'h3ad589fc),
	.w8(32'h39ead468),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae894ac),
	.w1(32'hba187fc4),
	.w2(32'h3ba6b62f),
	.w3(32'hbbdbd13b),
	.w4(32'h3b8a626d),
	.w5(32'h3bf5850b),
	.w6(32'h3a3363a5),
	.w7(32'h399f6e27),
	.w8(32'hb9a9753e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29cdd1),
	.w1(32'hbc165bd4),
	.w2(32'hb93baa9f),
	.w3(32'hbb018181),
	.w4(32'hbaab01d3),
	.w5(32'h3b2cf038),
	.w6(32'hbb2b0d77),
	.w7(32'h3a0da266),
	.w8(32'h3ad1715b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c1724a),
	.w1(32'h3ae261b9),
	.w2(32'hba15d569),
	.w3(32'hbcb06c59),
	.w4(32'hba84c6bb),
	.w5(32'hbae0cc74),
	.w6(32'hbb9fb253),
	.w7(32'hbd21ff74),
	.w8(32'h3b00e114),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8d372),
	.w1(32'h3ab9afa6),
	.w2(32'h3a7f2658),
	.w3(32'hbb310389),
	.w4(32'h3ad59cdf),
	.w5(32'h3c83693d),
	.w6(32'h3b2a2239),
	.w7(32'h3d0477d5),
	.w8(32'h3d022467),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3f93c),
	.w1(32'h3a1cd411),
	.w2(32'hbad43949),
	.w3(32'hba86aba2),
	.w4(32'hb9fe5af6),
	.w5(32'hbb9a6c79),
	.w6(32'hbb5a8303),
	.w7(32'h3ca7171c),
	.w8(32'hbc1a7cbe),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36db3a),
	.w1(32'hbb174bb0),
	.w2(32'h3a81b738),
	.w3(32'h3a831cc2),
	.w4(32'hbb0f1e68),
	.w5(32'h3a9d1365),
	.w6(32'h3cfbdeaf),
	.w7(32'hbbce79a3),
	.w8(32'hbb4224c0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b40c55),
	.w1(32'h3a44d19d),
	.w2(32'h3b505968),
	.w3(32'hbb66eeba),
	.w4(32'hbb02ddc5),
	.w5(32'h3ace68ca),
	.w6(32'h3ad81807),
	.w7(32'hbb84c847),
	.w8(32'hbba7e598),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f5101),
	.w1(32'hb96f5604),
	.w2(32'h3939bd44),
	.w3(32'h3bc84378),
	.w4(32'h39aa259b),
	.w5(32'h39cfd367),
	.w6(32'h3ba4ae45),
	.w7(32'hbb586fa4),
	.w8(32'hbb9d0136),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d419b),
	.w1(32'hbac48862),
	.w2(32'h3b1f559d),
	.w3(32'h3a14b381),
	.w4(32'hbb01de6e),
	.w5(32'h3a6fc2d9),
	.w6(32'hbb97b9dd),
	.w7(32'hba357a24),
	.w8(32'h3b9eb15b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bdeb7),
	.w1(32'hbbaeb312),
	.w2(32'hba3efd6f),
	.w3(32'hbba045fb),
	.w4(32'h38c0314f),
	.w5(32'h3b479003),
	.w6(32'h3aac90af),
	.w7(32'h3bb97c0e),
	.w8(32'h3bf8e87d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd8459),
	.w1(32'h3a92d1db),
	.w2(32'h3c97043c),
	.w3(32'hbaa5227e),
	.w4(32'h3aa0b8fc),
	.w5(32'hbb491130),
	.w6(32'h3b1e8a8e),
	.w7(32'hbbe8c6b3),
	.w8(32'h3a78cc9b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac21d4),
	.w1(32'hbb0d9854),
	.w2(32'h3c3a4fcd),
	.w3(32'h3bfa1084),
	.w4(32'hbb8a3f3a),
	.w5(32'h38a8425c),
	.w6(32'h3b2582cf),
	.w7(32'h3bc12e7e),
	.w8(32'hbb8edf7f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c6691),
	.w1(32'hbb5904d0),
	.w2(32'h39d4d170),
	.w3(32'hb949f1d0),
	.w4(32'hba196354),
	.w5(32'hbb6a1763),
	.w6(32'h3b2890a5),
	.w7(32'hbb98be83),
	.w8(32'hbbd5fe62),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a899fcf),
	.w1(32'h3a4646f4),
	.w2(32'hbad6f9a6),
	.w3(32'hbb32955c),
	.w4(32'h3ac46abb),
	.w5(32'h3ba8f765),
	.w6(32'hbc12aa04),
	.w7(32'hbaa31594),
	.w8(32'hbb4590e0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4df249),
	.w1(32'hb9d91b7f),
	.w2(32'h3b651f60),
	.w3(32'hbadfa2bf),
	.w4(32'hbb440520),
	.w5(32'hba510fad),
	.w6(32'hbad69311),
	.w7(32'hbc090c80),
	.w8(32'h3abaf60c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90baf5),
	.w1(32'hb97d5d4a),
	.w2(32'hbc3fa92a),
	.w3(32'h3b9009bc),
	.w4(32'hb955481d),
	.w5(32'hbc64230f),
	.w6(32'h3bc3ae7a),
	.w7(32'hbae823be),
	.w8(32'h3bc5bdbf),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fbbbc),
	.w1(32'hba6b07b3),
	.w2(32'hba0795c6),
	.w3(32'hbc10e8c1),
	.w4(32'hbb9d874e),
	.w5(32'hbb5a5a7c),
	.w6(32'hba18a270),
	.w7(32'hbbc913c2),
	.w8(32'h3b466002),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0596a9),
	.w1(32'h3b24f6a6),
	.w2(32'hbb1ecc25),
	.w3(32'hbb4188f1),
	.w4(32'hbb1bc1ca),
	.w5(32'h3d0852c0),
	.w6(32'h3b946bd0),
	.w7(32'h3a44c1cb),
	.w8(32'h3a000a32),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d845c),
	.w1(32'hbbc9cee9),
	.w2(32'hbbb523ca),
	.w3(32'h3b50324e),
	.w4(32'h3b5472c2),
	.w5(32'hbb58d29a),
	.w6(32'hbb2e1623),
	.w7(32'hbbd403bc),
	.w8(32'hbb925d7a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa777c),
	.w1(32'hbc0f7073),
	.w2(32'hba5733c4),
	.w3(32'h3bace357),
	.w4(32'hba582392),
	.w5(32'hbae36d3f),
	.w6(32'hbb2cf01a),
	.w7(32'hba5e6788),
	.w8(32'hba2ef3e2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba688d3f),
	.w1(32'h3837ed6d),
	.w2(32'h3be5c10a),
	.w3(32'h3a3c3b8f),
	.w4(32'h3aaf7de6),
	.w5(32'h3b5d046a),
	.w6(32'h3b9efab7),
	.w7(32'hbae42252),
	.w8(32'hbc02e601),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3d7f),
	.w1(32'hbb718622),
	.w2(32'hbc0f1fd2),
	.w3(32'hbb4c78ce),
	.w4(32'h3ab17fd6),
	.w5(32'h3b085e13),
	.w6(32'hbb4bb89c),
	.w7(32'h3bc90162),
	.w8(32'h3c2c9a12),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81855),
	.w1(32'h3c601af2),
	.w2(32'hba9a0e95),
	.w3(32'hbad52a91),
	.w4(32'h3b8ad904),
	.w5(32'h3ba6d24e),
	.w6(32'hbb43ff9d),
	.w7(32'h3c0d1562),
	.w8(32'hbb9c7905),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d5b0),
	.w1(32'h3b7a35b3),
	.w2(32'h3d1954d9),
	.w3(32'hbb399db9),
	.w4(32'hbbac8275),
	.w5(32'h3be280f5),
	.w6(32'h391d7d23),
	.w7(32'hb88a3634),
	.w8(32'h3aa7d766),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46166a),
	.w1(32'h3bd098dc),
	.w2(32'h3aa05f84),
	.w3(32'h3b83876d),
	.w4(32'hb7cec871),
	.w5(32'h3b82c0e0),
	.w6(32'hbb4171f5),
	.w7(32'hbbefb0aa),
	.w8(32'hbaf50846),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01abcf),
	.w1(32'h3b0f5aab),
	.w2(32'h3b46111b),
	.w3(32'hbbb84702),
	.w4(32'h3c35bc45),
	.w5(32'h3c186320),
	.w6(32'hbc317494),
	.w7(32'hba712b60),
	.w8(32'h3b35f89a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba634e9),
	.w1(32'h3cc3335a),
	.w2(32'h3ad78341),
	.w3(32'h3d0243a7),
	.w4(32'hb907d6f2),
	.w5(32'h3aaae793),
	.w6(32'h36e8bb06),
	.w7(32'hbb7ac673),
	.w8(32'hbba79882),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886d14),
	.w1(32'hbb2c1d74),
	.w2(32'h3ca1d666),
	.w3(32'h3b39a547),
	.w4(32'h3ae97c03),
	.w5(32'h3c81a1ff),
	.w6(32'h3c24465e),
	.w7(32'h3a5df8d6),
	.w8(32'hbbf034c4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1ac7b),
	.w1(32'h39a647b9),
	.w2(32'h3d536751),
	.w3(32'h3d24df16),
	.w4(32'hbad608fe),
	.w5(32'hbb3adfcc),
	.w6(32'h39a9b30e),
	.w7(32'h3c3b333a),
	.w8(32'hbc28295c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39956533),
	.w1(32'h3ab797c7),
	.w2(32'hbbdb6b6b),
	.w3(32'h3b14a92b),
	.w4(32'hbadd3b37),
	.w5(32'h3a609fda),
	.w6(32'h3bc1499e),
	.w7(32'hba62627d),
	.w8(32'hbc0b39ea),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafde632),
	.w1(32'hba86ab0e),
	.w2(32'hbb738155),
	.w3(32'hba8864b4),
	.w4(32'h3c26aaf6),
	.w5(32'hbaf35ca5),
	.w6(32'h3b366600),
	.w7(32'hbb822ad2),
	.w8(32'h3bc1caf0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf7167),
	.w1(32'hbb00af71),
	.w2(32'h3bcf6d30),
	.w3(32'hbb667471),
	.w4(32'hbc03bc2c),
	.w5(32'h3b105ed0),
	.w6(32'hbc1bd20a),
	.w7(32'hbb724e58),
	.w8(32'h3c048471),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02746c),
	.w1(32'h3c227fec),
	.w2(32'hbb56c30a),
	.w3(32'h3bd41bf8),
	.w4(32'h3ae5d6b8),
	.w5(32'hbaecb057),
	.w6(32'h3c019e12),
	.w7(32'hbab06539),
	.w8(32'h3b657839),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb82e8),
	.w1(32'hbb00f6d0),
	.w2(32'h3c469ac7),
	.w3(32'h3b56ce6b),
	.w4(32'h3cf6f6e5),
	.w5(32'hbb332d72),
	.w6(32'hbb0b853f),
	.w7(32'hbb95a9da),
	.w8(32'hba53e346),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c7efe3),
	.w1(32'h3c155ba4),
	.w2(32'h3b68eeb4),
	.w3(32'hba9f9a2b),
	.w4(32'h3b979b6f),
	.w5(32'h3b540212),
	.w6(32'hbaee67be),
	.w7(32'hbb8e0961),
	.w8(32'hbb58bd7d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c481539),
	.w1(32'h3bb37882),
	.w2(32'hbac6bae6),
	.w3(32'hbb820427),
	.w4(32'hbbf8807e),
	.w5(32'h3a4a8341),
	.w6(32'h3c240f0d),
	.w7(32'h3a08786e),
	.w8(32'hbadd0b37),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8304b3),
	.w1(32'h3bc57e6b),
	.w2(32'h3bc73d46),
	.w3(32'hb85765c4),
	.w4(32'h39b35fe8),
	.w5(32'h3b177eaa),
	.w6(32'hb914fabb),
	.w7(32'h3ae90cd7),
	.w8(32'h39d1cc69),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a33b5),
	.w1(32'hbc416700),
	.w2(32'hbab89cfb),
	.w3(32'hbb62663b),
	.w4(32'h3b5ffa5b),
	.w5(32'hbb2ff4eb),
	.w6(32'hbb4a3cf1),
	.w7(32'h3c4548e2),
	.w8(32'hbc005545),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c174053),
	.w1(32'hbbac9675),
	.w2(32'hbb56b1bb),
	.w3(32'hbb853b15),
	.w4(32'h3b848c33),
	.w5(32'hbb1771ca),
	.w6(32'h3c272c83),
	.w7(32'h3c349d64),
	.w8(32'h3a2c904a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107612),
	.w1(32'h3a7ae88b),
	.w2(32'hbc064e3a),
	.w3(32'h3bd81ef5),
	.w4(32'hbc3335c2),
	.w5(32'hbbb60db1),
	.w6(32'h3a9d54f1),
	.w7(32'hbbb7ed6b),
	.w8(32'hbb8a81cf),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4dded),
	.w1(32'hbc16391a),
	.w2(32'hbb8db45a),
	.w3(32'hbce186f1),
	.w4(32'hbb26e139),
	.w5(32'h3b49b914),
	.w6(32'hba4d408a),
	.w7(32'h3a950381),
	.w8(32'h3b8564e0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5706f),
	.w1(32'hbc41111f),
	.w2(32'h3bab7342),
	.w3(32'hbbd32ba4),
	.w4(32'hbaea3ca8),
	.w5(32'hbb92bd3f),
	.w6(32'hbaff63ce),
	.w7(32'hbb4c19fe),
	.w8(32'hbab5b69f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2b93a),
	.w1(32'hbaa987f6),
	.w2(32'hbc02a875),
	.w3(32'hb93c213e),
	.w4(32'h3b12b76b),
	.w5(32'hbb99de36),
	.w6(32'hbc2253fc),
	.w7(32'h3b0cc70d),
	.w8(32'hb9c055bb),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f3da3),
	.w1(32'h3b888ab1),
	.w2(32'h39a216b0),
	.w3(32'hbb479b6c),
	.w4(32'h3be634ce),
	.w5(32'h3be5a664),
	.w6(32'hbb36ce89),
	.w7(32'h39f650f4),
	.w8(32'hbaf4e921),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28d1a7),
	.w1(32'hbb0ed43f),
	.w2(32'h3b69963d),
	.w3(32'h3c2a047e),
	.w4(32'hbac99db3),
	.w5(32'hba33fb12),
	.w6(32'h3b7bfbab),
	.w7(32'h3b9e60c0),
	.w8(32'hbb86ab83),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb77169),
	.w1(32'hbd30bc1d),
	.w2(32'hbb4c3f2f),
	.w3(32'h3b59a1dc),
	.w4(32'hbb8b316f),
	.w5(32'hbc6c69c9),
	.w6(32'h3a400fd3),
	.w7(32'h3ac1b307),
	.w8(32'h3b682505),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab16c),
	.w1(32'hbae1f7d2),
	.w2(32'h3b0d61fc),
	.w3(32'hbbc85e7b),
	.w4(32'hb9cc01c5),
	.w5(32'hbb5a7166),
	.w6(32'hbd1d1974),
	.w7(32'hbc46bcc2),
	.w8(32'h3aa9d3a5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34d212),
	.w1(32'hb78495c0),
	.w2(32'h3b221bf5),
	.w3(32'h3bfec9ab),
	.w4(32'h3ae0784a),
	.w5(32'hbb885a76),
	.w6(32'h3a6c302a),
	.w7(32'hbb379063),
	.w8(32'h394b4e54),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca5360),
	.w1(32'hbb1d337a),
	.w2(32'hbb0c0175),
	.w3(32'h3bd2a0a2),
	.w4(32'hba51fc52),
	.w5(32'hba2b04ee),
	.w6(32'hb9ac1dec),
	.w7(32'hbba022a3),
	.w8(32'h3bd60ddb),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ad1b),
	.w1(32'hbab75d41),
	.w2(32'h3add2dc9),
	.w3(32'hbb183cb7),
	.w4(32'hbc044b70),
	.w5(32'h3ba7e644),
	.w6(32'hbb839681),
	.w7(32'h3bc01ea1),
	.w8(32'h3c2cb29e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65f513),
	.w1(32'hbc4b1c65),
	.w2(32'hba5c3819),
	.w3(32'h3c619f6d),
	.w4(32'hbb4a1cf3),
	.w5(32'hbad6ebbd),
	.w6(32'h3bb9a4e0),
	.w7(32'h3bbb762d),
	.w8(32'hbb5c3ed7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043272),
	.w1(32'h3a639c07),
	.w2(32'hbbe789f9),
	.w3(32'hbae7e7da),
	.w4(32'hbaf4e78d),
	.w5(32'hbadf9d81),
	.w6(32'hbc7c01f1),
	.w7(32'hbc0d3c00),
	.w8(32'h3c19f400),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba421e20),
	.w1(32'hba82a983),
	.w2(32'h3ab2d2de),
	.w3(32'h3d5d2555),
	.w4(32'hba36df3f),
	.w5(32'hbc2d9712),
	.w6(32'h3a946f11),
	.w7(32'h39c92ee8),
	.w8(32'h3ba700d2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b5ef0),
	.w1(32'h3a5f1920),
	.w2(32'h38843662),
	.w3(32'hbaaf4703),
	.w4(32'h397f6ca9),
	.w5(32'hbb7135b3),
	.w6(32'hbbee0413),
	.w7(32'h3bf9020f),
	.w8(32'h3a3844dd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4095),
	.w1(32'h3b29b405),
	.w2(32'h38a8f74d),
	.w3(32'hbac1dfa5),
	.w4(32'h3c2dcb7a),
	.w5(32'h3d47b48a),
	.w6(32'hbb3a6376),
	.w7(32'h3d1c534f),
	.w8(32'h37dc1479),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4b9ec),
	.w1(32'h3bb9e701),
	.w2(32'h3b35780c),
	.w3(32'h3bc9ae1a),
	.w4(32'hbadec978),
	.w5(32'hbb7670aa),
	.w6(32'hbb341f19),
	.w7(32'h3b526260),
	.w8(32'hbb8c327c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978d39b),
	.w1(32'hbc3e1205),
	.w2(32'h3c2babd0),
	.w3(32'hbb45ff02),
	.w4(32'h3ce9a889),
	.w5(32'h3987de96),
	.w6(32'hbc2d1bac),
	.w7(32'hbd8ba342),
	.w8(32'h3b6dcdf8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d227d),
	.w1(32'hba66920b),
	.w2(32'hb9422b1f),
	.w3(32'hbcbabf57),
	.w4(32'hba3b5b7e),
	.w5(32'h39948ca6),
	.w6(32'hba50a539),
	.w7(32'hbba1efb9),
	.w8(32'hbb2df011),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb231858),
	.w1(32'h3a16ec90),
	.w2(32'h3a2a6e44),
	.w3(32'hba514021),
	.w4(32'h39dbeda4),
	.w5(32'hbb86f092),
	.w6(32'hbb23b22f),
	.w7(32'hba87ba8a),
	.w8(32'hbbc6c889),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b12b),
	.w1(32'h3649548d),
	.w2(32'hbc02e102),
	.w3(32'h3ae89095),
	.w4(32'h3c2d6c78),
	.w5(32'hb9fb6b30),
	.w6(32'hbb91dfa3),
	.w7(32'hb8d90d0f),
	.w8(32'hbb7d3cc1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e5db),
	.w1(32'hbbc1b236),
	.w2(32'h3b567ff9),
	.w3(32'hbb56389a),
	.w4(32'h38d68f89),
	.w5(32'h3a4a76d6),
	.w6(32'h3ac73cc5),
	.w7(32'hbbd478e1),
	.w8(32'hb88f6c20),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a4ac9),
	.w1(32'h3a81ca1a),
	.w2(32'h3b44f713),
	.w3(32'hb9412f95),
	.w4(32'hbccd5cdf),
	.w5(32'hbba7fbee),
	.w6(32'hbb452d04),
	.w7(32'hbc2bd773),
	.w8(32'hbceefd1b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2d350),
	.w1(32'hbba94041),
	.w2(32'hbbe5218c),
	.w3(32'hbc023b21),
	.w4(32'hbc85f0a3),
	.w5(32'hbc45c750),
	.w6(32'hbbde6b3d),
	.w7(32'h395a7a67),
	.w8(32'h3b9bf14d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac457c),
	.w1(32'hbbea7dc1),
	.w2(32'hbba625e6),
	.w3(32'hbc320ce0),
	.w4(32'hbbdae02c),
	.w5(32'hbc81e1bc),
	.w6(32'hbb7514d3),
	.w7(32'hbb31787d),
	.w8(32'h3a4e78b7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfa7d2),
	.w1(32'hbb9ddb4a),
	.w2(32'h39a7049d),
	.w3(32'hbba254ea),
	.w4(32'hbbde1924),
	.w5(32'hbae04bd9),
	.w6(32'h3a8165bd),
	.w7(32'h397dfe1c),
	.w8(32'hba212d84),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58a6bb),
	.w1(32'hba172970),
	.w2(32'h3afedef7),
	.w3(32'hba1912c4),
	.w4(32'h3a928676),
	.w5(32'hbc6ba563),
	.w6(32'h3b85a6f8),
	.w7(32'hbba58f6b),
	.w8(32'h3c42b8d9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe84ec6),
	.w1(32'hb914950f),
	.w2(32'hbc8c18ee),
	.w3(32'hbabaefeb),
	.w4(32'hbadb1c8e),
	.w5(32'h3c006d09),
	.w6(32'h3b475be7),
	.w7(32'h3b3129ca),
	.w8(32'hbbf637a3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f1f80),
	.w1(32'h3aada251),
	.w2(32'hbb1a5853),
	.w3(32'h39d37b96),
	.w4(32'hbb10d5ce),
	.w5(32'h3b017636),
	.w6(32'h3b008b42),
	.w7(32'hbc26be71),
	.w8(32'hbb61099f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a969c8b),
	.w1(32'h3bac2505),
	.w2(32'h3af5e4a6),
	.w3(32'hbbe3b225),
	.w4(32'h3b506731),
	.w5(32'hbbe368cb),
	.w6(32'hbb424d6d),
	.w7(32'h3b57d800),
	.w8(32'hbbbb2d8a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c4b4e),
	.w1(32'hbbae2b58),
	.w2(32'hba4afa84),
	.w3(32'h3ba3e336),
	.w4(32'h3b2d0375),
	.w5(32'hbb616cdc),
	.w6(32'h3c3e3e30),
	.w7(32'hb9b2ce53),
	.w8(32'h3a990eaf),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d567),
	.w1(32'hb992a376),
	.w2(32'h3c02a4f2),
	.w3(32'hbb8af452),
	.w4(32'hb9911c44),
	.w5(32'hbb3570a7),
	.w6(32'h3b808e31),
	.w7(32'hbac8a1f3),
	.w8(32'h3c1fe947),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f24278),
	.w1(32'hbb912232),
	.w2(32'hba359e8b),
	.w3(32'h3b1deabd),
	.w4(32'hbb343e0c),
	.w5(32'h3a5bf29f),
	.w6(32'hb9c7d0b2),
	.w7(32'hbb1e1429),
	.w8(32'hbb6ee7f8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf858ab),
	.w1(32'hbbcdf1d2),
	.w2(32'hbb081e19),
	.w3(32'h3ba11d27),
	.w4(32'hba123eda),
	.w5(32'hbaade20c),
	.w6(32'h3b6f7543),
	.w7(32'hbc01323d),
	.w8(32'h3b32cbef),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf087),
	.w1(32'h3b083374),
	.w2(32'h3a23ab8d),
	.w3(32'h38bbf2c1),
	.w4(32'h3b011032),
	.w5(32'h3b5ee56d),
	.w6(32'h39bd292f),
	.w7(32'h393659e9),
	.w8(32'h3bc2841e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69e83a),
	.w1(32'hbb86533f),
	.w2(32'h3bb1c02e),
	.w3(32'hbb8debc9),
	.w4(32'hbb43a059),
	.w5(32'hbb598cd3),
	.w6(32'hb9836053),
	.w7(32'hbba4c1d2),
	.w8(32'h3c1bc091),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02dcbe),
	.w1(32'h3b0255fa),
	.w2(32'hba9e30d2),
	.w3(32'h3b0c62ad),
	.w4(32'hbae78cd1),
	.w5(32'hb9a0f901),
	.w6(32'h3b07f829),
	.w7(32'h3b2f7bcc),
	.w8(32'hbac53310),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa260c8),
	.w1(32'hb985b567),
	.w2(32'h3a8e254c),
	.w3(32'h3a9a0837),
	.w4(32'hb96a7fdd),
	.w5(32'h3b8ae76b),
	.w6(32'h3b3b9621),
	.w7(32'hbba9f4ee),
	.w8(32'hba300ae6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f5fdd),
	.w1(32'h3a0aad69),
	.w2(32'hbad4e9b8),
	.w3(32'hba993b7e),
	.w4(32'hbab78614),
	.w5(32'hbbb5b685),
	.w6(32'h3a886e49),
	.w7(32'h3b1467a7),
	.w8(32'hbb8b6a1f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d666a8),
	.w1(32'h3b0019d2),
	.w2(32'hbc0db492),
	.w3(32'h3a01f8b2),
	.w4(32'h3cb69a2d),
	.w5(32'h3bbdd690),
	.w6(32'hba76f1a5),
	.w7(32'hbbab3b86),
	.w8(32'h399c7a5e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34d766),
	.w1(32'h3ae6f060),
	.w2(32'hbb16d6d6),
	.w3(32'hbb6f3be6),
	.w4(32'h3bb6a3c0),
	.w5(32'hbb344f35),
	.w6(32'h3b8cc6f3),
	.w7(32'hbb2de707),
	.w8(32'h3ba78c53),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3034eb),
	.w1(32'h39da0a69),
	.w2(32'h3b385fc2),
	.w3(32'hbab0e18a),
	.w4(32'h3692a37e),
	.w5(32'h3c0e27e7),
	.w6(32'h3b471a79),
	.w7(32'hbc862b4b),
	.w8(32'h3842b204),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390de67c),
	.w1(32'h3b35a2c0),
	.w2(32'h39d4fa26),
	.w3(32'hbbb50e3e),
	.w4(32'hb909f5fe),
	.w5(32'h3b1caf4a),
	.w6(32'h3b87925c),
	.w7(32'hbb7563ef),
	.w8(32'h39e0fb10),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63d7a5),
	.w1(32'hbbeb0617),
	.w2(32'hbb13fb82),
	.w3(32'hbab15fc1),
	.w4(32'hbb0d512f),
	.w5(32'hb986bd72),
	.w6(32'hb83cc5ca),
	.w7(32'hb824ebbf),
	.w8(32'hbb0b63c6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d4775),
	.w1(32'hb95db466),
	.w2(32'hb90a164a),
	.w3(32'h39fe7e99),
	.w4(32'h3b0d2c54),
	.w5(32'hbc0542b5),
	.w6(32'hbc182596),
	.w7(32'hba7e86b1),
	.w8(32'h3a8d4424),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ccdc5),
	.w1(32'hb945bbe0),
	.w2(32'hbb100539),
	.w3(32'h3a745985),
	.w4(32'h3a0278f1),
	.w5(32'hbb85cd0d),
	.w6(32'hbaffc03c),
	.w7(32'h3c8ae463),
	.w8(32'hbba94fdd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c960d46),
	.w1(32'hbaed6b8a),
	.w2(32'hbae4e2fa),
	.w3(32'h3b8f03ce),
	.w4(32'hbaf7a941),
	.w5(32'hba8964d6),
	.w6(32'hbbd63026),
	.w7(32'h3b560601),
	.w8(32'hbac9d442),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825e8b),
	.w1(32'h3a366476),
	.w2(32'h3b08c543),
	.w3(32'h39bcefaf),
	.w4(32'hbaa3a5fa),
	.w5(32'hb9f053fa),
	.w6(32'hb8fbe862),
	.w7(32'hbba07cb6),
	.w8(32'h3b070c7d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf032ad),
	.w1(32'hbb258e23),
	.w2(32'hba6a44cc),
	.w3(32'hb9a12813),
	.w4(32'h3c17e3b9),
	.w5(32'hbb1629b6),
	.w6(32'h3ad3cc39),
	.w7(32'h391dd566),
	.w8(32'h3bcad174),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6722af7),
	.w1(32'hbac85bce),
	.w2(32'h3a4b4356),
	.w3(32'h39f1a063),
	.w4(32'hb9f158fa),
	.w5(32'h3bb55143),
	.w6(32'hbb973ac2),
	.w7(32'hba3efd9f),
	.w8(32'hbbcb44d3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27859e),
	.w1(32'h398855e3),
	.w2(32'h3b3e38ca),
	.w3(32'hbc6c7fb4),
	.w4(32'h3b736984),
	.w5(32'hbb495c1f),
	.w6(32'h3a01d34f),
	.w7(32'h3b56a431),
	.w8(32'hbb2e484e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb684115),
	.w1(32'hbb2ddec0),
	.w2(32'hb9d27ee3),
	.w3(32'h38bab7fd),
	.w4(32'h3ac7145e),
	.w5(32'h3a9712e1),
	.w6(32'hbbb55307),
	.w7(32'h3abb043f),
	.w8(32'h3aa8c559),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4b0f6),
	.w1(32'hba287d45),
	.w2(32'h3a1f7b37),
	.w3(32'hbb07a736),
	.w4(32'hbacb52ad),
	.w5(32'hba23158e),
	.w6(32'h3a2c5ca2),
	.w7(32'hbb107101),
	.w8(32'h3a7add9b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b551508),
	.w1(32'h3b29910a),
	.w2(32'hba092a0b),
	.w3(32'h3b198648),
	.w4(32'hb9b6810e),
	.w5(32'h39881e81),
	.w6(32'h3af32acf),
	.w7(32'hb9500b77),
	.w8(32'hb9d90c39),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbef87),
	.w1(32'h3b14ab6e),
	.w2(32'hbb036b2e),
	.w3(32'hb9306273),
	.w4(32'hba741133),
	.w5(32'hb9dbecae),
	.w6(32'hbb0b7d02),
	.w7(32'h3b32daaa),
	.w8(32'h39ef5c26),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39879b46),
	.w1(32'hbc5482ee),
	.w2(32'h3b96fe0f),
	.w3(32'h3aa989c4),
	.w4(32'h3bb9c749),
	.w5(32'h3a311339),
	.w6(32'hbb71f097),
	.w7(32'h3a93f36b),
	.w8(32'h3ba0bafc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51bd78),
	.w1(32'hbaedd486),
	.w2(32'hbb08ed09),
	.w3(32'hb9b1e21c),
	.w4(32'h39c1fdef),
	.w5(32'h3af301c2),
	.w6(32'h3ae59863),
	.w7(32'h3b292a61),
	.w8(32'h3b93fbc6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55e835),
	.w1(32'h3b47a06e),
	.w2(32'h39859d9f),
	.w3(32'hbb7cf19e),
	.w4(32'h3b66cc18),
	.w5(32'hba5cdb30),
	.w6(32'h3a4846da),
	.w7(32'h3b8097ac),
	.w8(32'hb93d01fe),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e07f),
	.w1(32'hbb730356),
	.w2(32'hbae0cc39),
	.w3(32'hbb10dda8),
	.w4(32'h3ab6d436),
	.w5(32'h3bab77ed),
	.w6(32'hbbb09bb2),
	.w7(32'h3b10dadb),
	.w8(32'h3af15a1d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f83d),
	.w1(32'hbaee2339),
	.w2(32'h3b7496ca),
	.w3(32'hbaefaa16),
	.w4(32'h3a867aa5),
	.w5(32'h3ab749f2),
	.w6(32'h3b3c2719),
	.w7(32'hbb951499),
	.w8(32'hbc17273f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba42ce1),
	.w1(32'h3d07ed97),
	.w2(32'hbb9ee4a8),
	.w3(32'h3d4d50d0),
	.w4(32'h3abfa6fa),
	.w5(32'h3addeefc),
	.w6(32'hbaff4a4b),
	.w7(32'hbb3cc0b8),
	.w8(32'h3ae4fa9e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule