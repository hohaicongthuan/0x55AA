module layer_10_featuremap_17(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e0c8),
	.w1(32'hbbc49465),
	.w2(32'h3b21b2b8),
	.w3(32'h3b11629f),
	.w4(32'hba0863c2),
	.w5(32'hba4619b2),
	.w6(32'h3a4ded5f),
	.w7(32'hbafb6c09),
	.w8(32'hbb69f410),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b567db4),
	.w1(32'h3c1b50bc),
	.w2(32'hbb0f9c5f),
	.w3(32'h3b0122ff),
	.w4(32'h3bf6aff1),
	.w5(32'hbbbcc7cb),
	.w6(32'hbb190cad),
	.w7(32'hbb85eb97),
	.w8(32'hbb4769c4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba23e6b),
	.w1(32'hbb66e589),
	.w2(32'hbb5e4002),
	.w3(32'hbb266141),
	.w4(32'hbb107af3),
	.w5(32'hbbc843ac),
	.w6(32'hbb7d8eb7),
	.w7(32'h39a4fe68),
	.w8(32'h3b1baae0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2014bc),
	.w1(32'hbb8493dd),
	.w2(32'h3b78eb83),
	.w3(32'h3b640d93),
	.w4(32'hb96eb4d2),
	.w5(32'hbb83dc10),
	.w6(32'hbab9c4cf),
	.w7(32'h3b105cc5),
	.w8(32'h38c4b3f0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1b897),
	.w1(32'hbae1718f),
	.w2(32'h3a9f9fd6),
	.w3(32'hbb92ed39),
	.w4(32'h3bab8fcc),
	.w5(32'hbbb3611c),
	.w6(32'h3bfb95b2),
	.w7(32'h3c29aca4),
	.w8(32'hbb4bbcd4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2376f5),
	.w1(32'h3acad761),
	.w2(32'hbce024f4),
	.w3(32'hbb0290a8),
	.w4(32'hbb20d5da),
	.w5(32'h3c47e32c),
	.w6(32'h39d64c79),
	.w7(32'h3b875e05),
	.w8(32'h3ce19cb1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f60c),
	.w1(32'hbc6cd8dc),
	.w2(32'hbb28fdab),
	.w3(32'h3db94ce2),
	.w4(32'h3d770c42),
	.w5(32'hbc007050),
	.w6(32'h3dd908b7),
	.w7(32'h3d83a1de),
	.w8(32'h3b0b2948),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dfcab),
	.w1(32'hbc20f83e),
	.w2(32'h3897deef),
	.w3(32'hbba5a914),
	.w4(32'hbc73192e),
	.w5(32'hba888b95),
	.w6(32'h3c1ead34),
	.w7(32'h3b7c8ff7),
	.w8(32'h3b8c596f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2570be),
	.w1(32'hbbc5c2d2),
	.w2(32'hbad3a6e0),
	.w3(32'h3aa375e5),
	.w4(32'hbb2fa108),
	.w5(32'hbb36a439),
	.w6(32'h3b5e830b),
	.w7(32'hb83e0539),
	.w8(32'h3aeaa299),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136b7e),
	.w1(32'hbba07547),
	.w2(32'hbc2f3499),
	.w3(32'h3a502373),
	.w4(32'h3a45d49c),
	.w5(32'hba55579e),
	.w6(32'h3b4ea79e),
	.w7(32'hbbb4669c),
	.w8(32'h3c52e31a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f66f),
	.w1(32'hbb1e125d),
	.w2(32'hb995a39f),
	.w3(32'h3cc9931d),
	.w4(32'h3ccbc928),
	.w5(32'hbb4f4d82),
	.w6(32'h3d1d31ac),
	.w7(32'h3d1231c9),
	.w8(32'h3a7ba061),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d693),
	.w1(32'hbb5d6be5),
	.w2(32'h382f91b6),
	.w3(32'h3bd079d2),
	.w4(32'h3b5dad15),
	.w5(32'hbbc88bde),
	.w6(32'h3c591e7c),
	.w7(32'hbaeaf616),
	.w8(32'hbc33efec),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc158c82),
	.w1(32'hbc1a4ee6),
	.w2(32'hbb1b342c),
	.w3(32'hbc7fd191),
	.w4(32'hbc6cb6f8),
	.w5(32'hbab61717),
	.w6(32'hbc81819f),
	.w7(32'hbc9ee0ca),
	.w8(32'hbbe250fe),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb28c),
	.w1(32'hb9553675),
	.w2(32'h3c276687),
	.w3(32'hbb7349da),
	.w4(32'hbb03cca4),
	.w5(32'h3b7edc55),
	.w6(32'hbc16b9a0),
	.w7(32'hbbd79dde),
	.w8(32'hbac36601),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ba1a9),
	.w1(32'h3bea3319),
	.w2(32'hb9ac7218),
	.w3(32'h3b6c0a51),
	.w4(32'h3b497386),
	.w5(32'h3a44214f),
	.w6(32'hbbc0c75a),
	.w7(32'hbb9ee565),
	.w8(32'hb9c76d12),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb634ac7),
	.w1(32'h3bb6a96f),
	.w2(32'hbc7aec8f),
	.w3(32'hbc0cba7b),
	.w4(32'h3b441a30),
	.w5(32'h3c2fc73a),
	.w6(32'hbb788e51),
	.w7(32'hb8c86ba8),
	.w8(32'h3cf1551c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd23cab),
	.w1(32'hba16573d),
	.w2(32'h39485cd2),
	.w3(32'h3d5ace6d),
	.w4(32'h3d46e077),
	.w5(32'hbae4aa9c),
	.w6(32'h3d986cb6),
	.w7(32'h3d7e7505),
	.w8(32'h3bbb1099),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946765),
	.w1(32'hbb34e53c),
	.w2(32'h3b30ba35),
	.w3(32'hbb6423ed),
	.w4(32'hbbdd5d3b),
	.w5(32'hbbea3901),
	.w6(32'h3be45817),
	.w7(32'hba61b828),
	.w8(32'h3b01b879),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadbd62),
	.w1(32'hbb8cb31b),
	.w2(32'h3adcaa88),
	.w3(32'hbbbac194),
	.w4(32'hbb8935e4),
	.w5(32'h3b486712),
	.w6(32'hbb86a5af),
	.w7(32'hbb9993af),
	.w8(32'h3b5456c5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2187c3),
	.w1(32'h3bbd8a9a),
	.w2(32'hbb918207),
	.w3(32'h3c4217e6),
	.w4(32'h3bc44a7b),
	.w5(32'h3a352048),
	.w6(32'h3af0ac11),
	.w7(32'h3b789e1a),
	.w8(32'hb9c0c9e0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac52c1b),
	.w1(32'h39f99cb2),
	.w2(32'h3ba77c52),
	.w3(32'h3920affe),
	.w4(32'hbb0005f9),
	.w5(32'hbb8bf692),
	.w6(32'h38a5453a),
	.w7(32'h3a9ce8ea),
	.w8(32'h3afdbade),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae11357),
	.w1(32'h3b71a549),
	.w2(32'h3b5b7639),
	.w3(32'h39510fd6),
	.w4(32'h3a12e0c2),
	.w5(32'hba29f8b3),
	.w6(32'hba13e32e),
	.w7(32'h3b112070),
	.w8(32'hbb12a123),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dcd3e),
	.w1(32'hbb27ad9c),
	.w2(32'h3c894758),
	.w3(32'h3b256804),
	.w4(32'hbba6eca0),
	.w5(32'hbacc9903),
	.w6(32'hbbfdfbe7),
	.w7(32'hbb9e8308),
	.w8(32'hbb8147be),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092265),
	.w1(32'h3c374937),
	.w2(32'h3a4d27aa),
	.w3(32'hbc933629),
	.w4(32'hbbc7616e),
	.w5(32'hba062c24),
	.w6(32'hbc91eca1),
	.w7(32'hbc28d4de),
	.w8(32'hbbe84eca),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1af6),
	.w1(32'hbb1b1568),
	.w2(32'hbb9bf854),
	.w3(32'h3a7bfabe),
	.w4(32'hbb113c54),
	.w5(32'hbaf10883),
	.w6(32'hbc3421cd),
	.w7(32'hbbc810b6),
	.w8(32'h3be58f77),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86fbf9),
	.w1(32'hbb2c588f),
	.w2(32'hbb048ad7),
	.w3(32'h3bac24cb),
	.w4(32'h3b8b4b81),
	.w5(32'hbbb8f5b2),
	.w6(32'h3c407432),
	.w7(32'hbb294ccb),
	.w8(32'h3a85cef3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b970389),
	.w1(32'h3b66766c),
	.w2(32'h39eab68a),
	.w3(32'hba2ae803),
	.w4(32'h3a5ad30a),
	.w5(32'hb9eedab3),
	.w6(32'h3a69b978),
	.w7(32'h3bef2c52),
	.w8(32'h39f7495f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca9585),
	.w1(32'h3bc73869),
	.w2(32'hbc156689),
	.w3(32'hbbb49fca),
	.w4(32'h3bff8d64),
	.w5(32'h3a65d752),
	.w6(32'hbbf7fe2a),
	.w7(32'h3a3ee4d8),
	.w8(32'h3b6fdf65),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0da66d),
	.w1(32'h3a48bead),
	.w2(32'h3b5d7e10),
	.w3(32'h3c39515b),
	.w4(32'h3c5133d2),
	.w5(32'hbb285852),
	.w6(32'h3b5bf584),
	.w7(32'h3b861be9),
	.w8(32'hbbc19528),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c255567),
	.w1(32'h3c053400),
	.w2(32'hb9ac70ac),
	.w3(32'h3b3eef74),
	.w4(32'hb8a088b8),
	.w5(32'hbb53d7a6),
	.w6(32'hbad88461),
	.w7(32'hbc14a569),
	.w8(32'hbaab16e5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9eae),
	.w1(32'hbaaa2cd1),
	.w2(32'h3b27b0b0),
	.w3(32'hbbff5516),
	.w4(32'hbb45cdb9),
	.w5(32'h3c355dd6),
	.w6(32'hbb3eebc7),
	.w7(32'hb8a4e531),
	.w8(32'h3c9774c6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a534813),
	.w1(32'h3b77cde3),
	.w2(32'hbc3b298c),
	.w3(32'h3c1e015d),
	.w4(32'h3b4211c8),
	.w5(32'h3b598b9e),
	.w6(32'h3ca26ffa),
	.w7(32'h3c5faf11),
	.w8(32'h3c6934f9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa1b1e),
	.w1(32'hbb0c861a),
	.w2(32'h3ba68427),
	.w3(32'h3cc5ff4b),
	.w4(32'h3ca9364d),
	.w5(32'h3c1544ca),
	.w6(32'h3ca85d3d),
	.w7(32'h3c0b310e),
	.w8(32'h3b5a449c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d8728),
	.w1(32'h3b7d8419),
	.w2(32'hbb495871),
	.w3(32'h3be484e6),
	.w4(32'h3b91f657),
	.w5(32'hbc5c5f3a),
	.w6(32'hbb6b3e9d),
	.w7(32'hba492051),
	.w8(32'hbca74bed),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aa36e),
	.w1(32'hbbc45684),
	.w2(32'h3a96e261),
	.w3(32'hbce3b0a6),
	.w4(32'hbc1234e5),
	.w5(32'h3ab6ef2a),
	.w6(32'hbc5eb3cc),
	.w7(32'h3c0fbd5b),
	.w8(32'hbbad8326),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2bc71),
	.w1(32'hb94c4c22),
	.w2(32'hbc1fead2),
	.w3(32'h3b5c7726),
	.w4(32'hbbb973c4),
	.w5(32'hbc0b9d35),
	.w6(32'hbb99a4e3),
	.w7(32'hbbea15f8),
	.w8(32'h3aa8353c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1e880),
	.w1(32'hbc3d6a0b),
	.w2(32'h39f24bc0),
	.w3(32'h3bc2a873),
	.w4(32'hbc21bf4d),
	.w5(32'h3ac5dc90),
	.w6(32'h3b922b6f),
	.w7(32'hbbca771e),
	.w8(32'hbbe52de9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc931ea),
	.w1(32'hbbaa8719),
	.w2(32'h3b9841f8),
	.w3(32'hba99589d),
	.w4(32'h3a925ea8),
	.w5(32'h3bad13b6),
	.w6(32'hbcaefd72),
	.w7(32'hbc35c157),
	.w8(32'h3c20e989),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d606d),
	.w1(32'h3bbb1ffa),
	.w2(32'hba943d64),
	.w3(32'h3c35cebf),
	.w4(32'h3c024851),
	.w5(32'h3a475a2f),
	.w6(32'hb99d3058),
	.w7(32'hbb921947),
	.w8(32'hbc3cee8e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd3d8),
	.w1(32'h39d60674),
	.w2(32'h3ba59b7f),
	.w3(32'h3b06f949),
	.w4(32'hbbbcb70e),
	.w5(32'h3b83f51e),
	.w6(32'hbc692882),
	.w7(32'hbc756b18),
	.w8(32'h3a9e7b03),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5f03),
	.w1(32'h3ba26431),
	.w2(32'hbb8a3fde),
	.w3(32'h3ba3a789),
	.w4(32'h3bacdfcf),
	.w5(32'h3c4e2a56),
	.w6(32'h3b9755f6),
	.w7(32'h3bcb94d2),
	.w8(32'h3cfe5293),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e1380),
	.w1(32'h3b0bac3c),
	.w2(32'hbc14afae),
	.w3(32'h3cb1f916),
	.w4(32'h3cd1ba47),
	.w5(32'hbc54957c),
	.w6(32'h3d0b64ed),
	.w7(32'h3cd066e9),
	.w8(32'hbc07e644),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeddce2),
	.w1(32'hbc3a272a),
	.w2(32'h3aead504),
	.w3(32'hbc748acf),
	.w4(32'hbc47ff69),
	.w5(32'h3b7209b8),
	.w6(32'hbc6d66ce),
	.w7(32'hbc6e8de9),
	.w8(32'h3ac01d65),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8e980),
	.w1(32'h3a999a18),
	.w2(32'hbc01eb33),
	.w3(32'hbbba06e8),
	.w4(32'h3accb4be),
	.w5(32'h3b4643e0),
	.w6(32'hbb95b66a),
	.w7(32'hbb00b932),
	.w8(32'h3b3eaf23),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba71fb7),
	.w1(32'hbc73542b),
	.w2(32'h3bc87e18),
	.w3(32'h3b95b990),
	.w4(32'h3ab54e87),
	.w5(32'h3c79989a),
	.w6(32'h3c1d66ca),
	.w7(32'hba9dd897),
	.w8(32'h3bd35e4b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3f25f),
	.w1(32'hbb66e1f0),
	.w2(32'hbb1a75df),
	.w3(32'h3c27d6bb),
	.w4(32'h3c09e909),
	.w5(32'h3aa543f8),
	.w6(32'h3b40d19b),
	.w7(32'hbba53898),
	.w8(32'h3a13ffb1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1ea53),
	.w1(32'hbbc55ee7),
	.w2(32'hbb197dd2),
	.w3(32'hbb04ee41),
	.w4(32'hbb027ad0),
	.w5(32'hbc0c749e),
	.w6(32'hbb196ea5),
	.w7(32'hba58fc99),
	.w8(32'h3a97c81a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0857d9),
	.w1(32'hbb844069),
	.w2(32'hbb61117b),
	.w3(32'hbc58687a),
	.w4(32'hbbac0e49),
	.w5(32'hbb8f1716),
	.w6(32'h3c057623),
	.w7(32'hba865c19),
	.w8(32'hbb12e0d1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f5b3),
	.w1(32'h3a2cb617),
	.w2(32'hb8f0b2f9),
	.w3(32'h3adcee85),
	.w4(32'h3a386714),
	.w5(32'hbc10d0f9),
	.w6(32'hba0495c6),
	.w7(32'hbadcd514),
	.w8(32'hbc81f964),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5a6e9),
	.w1(32'hbac60fa0),
	.w2(32'h39ecf64b),
	.w3(32'hbc1d3106),
	.w4(32'hbc56619d),
	.w5(32'hbb23eec0),
	.w6(32'hbc557d23),
	.w7(32'hbb57ebb0),
	.w8(32'hbb9debb7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc454581),
	.w1(32'hbb50f56a),
	.w2(32'hbc339037),
	.w3(32'hbc1426dd),
	.w4(32'hbbf6449a),
	.w5(32'hbb09c31a),
	.w6(32'hbb8de62a),
	.w7(32'hbafe0c22),
	.w8(32'h3c4e877e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5476f),
	.w1(32'hbc0a9e1e),
	.w2(32'h3a77e18c),
	.w3(32'h3baf424f),
	.w4(32'h3c6f31e9),
	.w5(32'h3aec4945),
	.w6(32'h3c93ad83),
	.w7(32'h3c8d4f8a),
	.w8(32'hbbb65d75),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93cd32),
	.w1(32'hbbaed874),
	.w2(32'hbbc2836c),
	.w3(32'hbba3cee7),
	.w4(32'h3ac94429),
	.w5(32'hbb606bb7),
	.w6(32'h39679268),
	.w7(32'h3afe41df),
	.w8(32'h3c07142f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba286e3),
	.w1(32'hbb9d4f10),
	.w2(32'h3c27c5cc),
	.w3(32'hbbe8ad26),
	.w4(32'hbbbc6f09),
	.w5(32'hbc04f891),
	.w6(32'h3c069345),
	.w7(32'h3a5eee55),
	.w8(32'h3ba02987),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56093),
	.w1(32'hbb868d91),
	.w2(32'h3b81acf7),
	.w3(32'hbc2e95b9),
	.w4(32'hbbc92412),
	.w5(32'hbb140e93),
	.w6(32'hbb2c3fa4),
	.w7(32'h3bfdbaf5),
	.w8(32'hbc723116),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7d2b5),
	.w1(32'hbafc8a29),
	.w2(32'hbc75405a),
	.w3(32'hbc5a163c),
	.w4(32'hbc655ba7),
	.w5(32'hbbebbe65),
	.w6(32'hbc9ccc52),
	.w7(32'hbca69186),
	.w8(32'h3b954858),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e394),
	.w1(32'hbbf8391d),
	.w2(32'hbba4c261),
	.w3(32'hbbba1d49),
	.w4(32'hbb76b5bd),
	.w5(32'h3b4aaab5),
	.w6(32'h3abde710),
	.w7(32'h3b5f7fce),
	.w8(32'h3b880c24),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ef7a6),
	.w1(32'h3a92ea64),
	.w2(32'hb98cdf1c),
	.w3(32'h3ba1c119),
	.w4(32'h3b42d81d),
	.w5(32'h3a9bf381),
	.w6(32'h3ba3ab4b),
	.w7(32'hb9f1db20),
	.w8(32'hb99e7788),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16d0a7),
	.w1(32'h3b2eff70),
	.w2(32'hbb0352fd),
	.w3(32'h3b880b5c),
	.w4(32'h3b98933d),
	.w5(32'h3c7b6c13),
	.w6(32'hbbaa8f33),
	.w7(32'hbadda825),
	.w8(32'h3cce54c1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8a13),
	.w1(32'h3bd50f6c),
	.w2(32'hbc74c1ea),
	.w3(32'h3cfb63ee),
	.w4(32'h3cac00e6),
	.w5(32'hbcf51066),
	.w6(32'h3ce6993f),
	.w7(32'h3caf8498),
	.w8(32'hbc2d9522),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd81234),
	.w1(32'hbcbe54c7),
	.w2(32'h3b83d04b),
	.w3(32'hbcefd203),
	.w4(32'hbc3cee17),
	.w5(32'h3b351e65),
	.w6(32'h3bb08a3b),
	.w7(32'h3bacd942),
	.w8(32'h3bb3c902),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849dc5),
	.w1(32'h3c030c72),
	.w2(32'h396a695f),
	.w3(32'hbb4080fd),
	.w4(32'h3c246148),
	.w5(32'h3b413f00),
	.w6(32'hbbf1bf8f),
	.w7(32'h3b0a3d27),
	.w8(32'h3b8ed537),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22bf2b),
	.w1(32'h3b2ed9b7),
	.w2(32'hbb4500cc),
	.w3(32'h3b8b4460),
	.w4(32'h3b3f2d05),
	.w5(32'h3bf6d3b1),
	.w6(32'h3b02c574),
	.w7(32'hbad459eb),
	.w8(32'hba82c1c3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90dd293),
	.w1(32'hbb59a38c),
	.w2(32'hb993ae8e),
	.w3(32'h3c809b1d),
	.w4(32'h3c277506),
	.w5(32'hba178df5),
	.w6(32'h3b5628d1),
	.w7(32'h3bde1c6a),
	.w8(32'hbab579d7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8159d1),
	.w1(32'h3bdf5d35),
	.w2(32'hbb38b95d),
	.w3(32'hbbdc444c),
	.w4(32'h3b7c659c),
	.w5(32'hbbcbdb2b),
	.w6(32'h3bd10e25),
	.w7(32'h3bd3d2b4),
	.w8(32'hbbb44a0a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8774d),
	.w1(32'hbb2d4d52),
	.w2(32'hbad1296d),
	.w3(32'hbbcd286e),
	.w4(32'hbba23ca8),
	.w5(32'h3bcdc743),
	.w6(32'hbbbc9ad2),
	.w7(32'hbb86cc20),
	.w8(32'h3b564e0b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31eb6a),
	.w1(32'h3c2761fa),
	.w2(32'h3c4b1516),
	.w3(32'h3b2b78f9),
	.w4(32'h3c5c0839),
	.w5(32'h3c626408),
	.w6(32'hbbfb834a),
	.w7(32'hbaa69eca),
	.w8(32'h3b5e0887),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25408a),
	.w1(32'hbb52a12b),
	.w2(32'h3c57604a),
	.w3(32'h3b9fed99),
	.w4(32'hbb7ec765),
	.w5(32'h3bb4dfc1),
	.w6(32'h3a758ff4),
	.w7(32'h3bc3a7ce),
	.w8(32'h3be27f7c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bd1b3),
	.w1(32'h3bfcbc69),
	.w2(32'hbb617ffd),
	.w3(32'h3c29b94d),
	.w4(32'h3c08b7d4),
	.w5(32'hbb6a6309),
	.w6(32'h3b703407),
	.w7(32'h3bdc094c),
	.w8(32'h3a6463ba),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae8405),
	.w1(32'h3a8adecb),
	.w2(32'hbb8e225c),
	.w3(32'h3b6533e4),
	.w4(32'h3b9dfb51),
	.w5(32'hbbbd9c20),
	.w6(32'h3a9a4ad4),
	.w7(32'hb9bb9bcb),
	.w8(32'hbc0f7676),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98600a),
	.w1(32'h397bb4d6),
	.w2(32'h3a430cdf),
	.w3(32'hbae51d8c),
	.w4(32'h39a9c72a),
	.w5(32'hbbccbd71),
	.w6(32'hbb384593),
	.w7(32'hb9ae35c7),
	.w8(32'hbbeb8d11),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9164ec),
	.w1(32'hbbaf2011),
	.w2(32'h3bba7b2b),
	.w3(32'hbc12a970),
	.w4(32'hbc1cee92),
	.w5(32'h3c6d8d82),
	.w6(32'hbc20e0d5),
	.w7(32'hbbc63e37),
	.w8(32'h3c1ea1a7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c193d60),
	.w1(32'h3c27c351),
	.w2(32'h3905e2ef),
	.w3(32'h3c3b0265),
	.w4(32'h3c3e7732),
	.w5(32'hbb5d8e14),
	.w6(32'h3c0fb1d5),
	.w7(32'h3c0f94e7),
	.w8(32'hbbee283a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b5d70),
	.w1(32'hbb73c3c9),
	.w2(32'h3bd90170),
	.w3(32'h3ab613c4),
	.w4(32'hbab27572),
	.w5(32'h39cee821),
	.w6(32'hbc0be355),
	.w7(32'hbba7e10e),
	.w8(32'h3ba88fcc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b527c6),
	.w1(32'h3b4e31f0),
	.w2(32'h3b6771c7),
	.w3(32'hbc0c9a35),
	.w4(32'hbbbe9885),
	.w5(32'h3a723b4e),
	.w6(32'hbb8247ae),
	.w7(32'hbb011473),
	.w8(32'hbb9b7e60),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af32f53),
	.w1(32'hb904e96e),
	.w2(32'hbb0d9a25),
	.w3(32'hbb94dcaa),
	.w4(32'hbbc6fadd),
	.w5(32'h3a80a08c),
	.w6(32'hbc11b317),
	.w7(32'hbc1681a4),
	.w8(32'hb90b72a9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514604),
	.w1(32'h3b827570),
	.w2(32'h3b9991f9),
	.w3(32'h3c70a2ce),
	.w4(32'hba541a31),
	.w5(32'hbb1c4079),
	.w6(32'h3b9c264a),
	.w7(32'h3bd1607c),
	.w8(32'hbb43d8f2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8c8e),
	.w1(32'hbb56a9d3),
	.w2(32'hbc396117),
	.w3(32'h3b910061),
	.w4(32'hbae19bce),
	.w5(32'hbb41ce40),
	.w6(32'h3aa6ffd1),
	.w7(32'h3b8aefa1),
	.w8(32'hbb88bbd8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65ec99),
	.w1(32'hbb91c095),
	.w2(32'h3ac5d7b1),
	.w3(32'hbc1e0b06),
	.w4(32'hba1f9294),
	.w5(32'h39f6a442),
	.w6(32'h3b938cad),
	.w7(32'h3b27469b),
	.w8(32'h3a9a31dc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55aaf4),
	.w1(32'h3b3c00a5),
	.w2(32'hbbc816db),
	.w3(32'hbb7c7aed),
	.w4(32'h3a15c4cc),
	.w5(32'hbbca1a6c),
	.w6(32'hbabd2941),
	.w7(32'hbb0bff08),
	.w8(32'hbb38815f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc424900),
	.w1(32'hba0a772c),
	.w2(32'hbb4ccdd8),
	.w3(32'hbbc8004b),
	.w4(32'hbb925229),
	.w5(32'hbb5b7d66),
	.w6(32'hbc1004d4),
	.w7(32'hbc04a96a),
	.w8(32'hb8e8a51a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178d7f),
	.w1(32'hbc15519d),
	.w2(32'hbb00fbf4),
	.w3(32'hbc2deb50),
	.w4(32'hbbfaeb49),
	.w5(32'hb962478e),
	.w6(32'hbbccb506),
	.w7(32'hbb579952),
	.w8(32'h3b918ffd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a337812),
	.w1(32'hb982fb7f),
	.w2(32'h3bb3ca24),
	.w3(32'h3b538ac3),
	.w4(32'h3b2a704a),
	.w5(32'hbc0cef7c),
	.w6(32'h3bbdb4b5),
	.w7(32'h3c15a086),
	.w8(32'hbbcf49b3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7de143),
	.w1(32'h3b702da5),
	.w2(32'h39ee35e0),
	.w3(32'hbc0f148f),
	.w4(32'hbc1a712c),
	.w5(32'h3bd7538b),
	.w6(32'hbc605932),
	.w7(32'hbc3c0583),
	.w8(32'h3ba39849),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a08dc),
	.w1(32'h3b478b2e),
	.w2(32'h3add38ed),
	.w3(32'h3b838645),
	.w4(32'h3b801f70),
	.w5(32'hbba3b494),
	.w6(32'h3b07da45),
	.w7(32'h3b0af1f9),
	.w8(32'hba105bb6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca749),
	.w1(32'hbab65942),
	.w2(32'h3b380fad),
	.w3(32'hbc2a8b0d),
	.w4(32'h3afa679c),
	.w5(32'h3b88204f),
	.w6(32'h39f74daa),
	.w7(32'h3c1c2a14),
	.w8(32'h3b3ec4b3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24492a),
	.w1(32'h3bf25406),
	.w2(32'hba6a489b),
	.w3(32'h3bad8e9c),
	.w4(32'h3bfb1b10),
	.w5(32'hb9a74403),
	.w6(32'hbb8e7b78),
	.w7(32'h3b3bd877),
	.w8(32'hbb76108f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb877c0f6),
	.w1(32'h3b07774a),
	.w2(32'h3aca8747),
	.w3(32'hbabaf847),
	.w4(32'hba4b7f87),
	.w5(32'hbae78a45),
	.w6(32'hbaca9b6d),
	.w7(32'hbb0607aa),
	.w8(32'h3b1592bd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3776b8),
	.w1(32'h3a5cc404),
	.w2(32'h3c53a365),
	.w3(32'hb9a2dbdc),
	.w4(32'h3a89a992),
	.w5(32'hbcf3948b),
	.w6(32'hbb173987),
	.w7(32'h3aa73cc4),
	.w8(32'hbd1ed147),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a005),
	.w1(32'hbc10a944),
	.w2(32'h3b5b9a3d),
	.w3(32'hbd4b87fb),
	.w4(32'hbd1b2fdb),
	.w5(32'hbbaa27f0),
	.w6(32'hbd05f999),
	.w7(32'hbc9291f3),
	.w8(32'hbbb8d5be),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04da2e),
	.w1(32'hbbd38f7f),
	.w2(32'hbc2921ae),
	.w3(32'hbc4d862f),
	.w4(32'hbc10cdff),
	.w5(32'h3b3c4f0b),
	.w6(32'hbc479a8c),
	.w7(32'hbbf97c35),
	.w8(32'h3b94e365),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98dc49),
	.w1(32'hbbbbedb9),
	.w2(32'h3bfda173),
	.w3(32'h3ca1e9d6),
	.w4(32'h3c153ddf),
	.w5(32'h3bbed860),
	.w6(32'h3c2689d3),
	.w7(32'h3a0c7335),
	.w8(32'hbb8d4214),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62b22c),
	.w1(32'h3aed375a),
	.w2(32'hbbdc901f),
	.w3(32'h3ad01754),
	.w4(32'h3af56856),
	.w5(32'hbb99c46e),
	.w6(32'hbb30a595),
	.w7(32'h3a01d451),
	.w8(32'hba0e26da),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc357a71),
	.w1(32'hbab61061),
	.w2(32'h3c0ca483),
	.w3(32'hbbea3f11),
	.w4(32'h38b643de),
	.w5(32'h3c8c312d),
	.w6(32'hba726607),
	.w7(32'hba3a4797),
	.w8(32'h3ba01a01),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e95f),
	.w1(32'h3c57f5d8),
	.w2(32'h3bb0c6bb),
	.w3(32'h3c1ccf74),
	.w4(32'h3c32c93c),
	.w5(32'h3c0a8e90),
	.w6(32'h3b90b831),
	.w7(32'h38ac70f7),
	.w8(32'h3b616209),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0da95),
	.w1(32'h3bfb05fb),
	.w2(32'h3b837969),
	.w3(32'h3c0020ee),
	.w4(32'h3c0fe97d),
	.w5(32'hbb5fe559),
	.w6(32'h3be0e9a3),
	.w7(32'h3b9fe09a),
	.w8(32'hbc41fafc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7518fd),
	.w1(32'h3b306855),
	.w2(32'h3bc8d48f),
	.w3(32'hbc64f332),
	.w4(32'hbc3d9dd3),
	.w5(32'h3b382404),
	.w6(32'hbc731c33),
	.w7(32'hbc562d25),
	.w8(32'h3bdf33cd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59ba36),
	.w1(32'h3b9a545e),
	.w2(32'hbc4e6d7a),
	.w3(32'h3b59616f),
	.w4(32'h397f32e3),
	.w5(32'h3b17cb1c),
	.w6(32'h3b8bb962),
	.w7(32'hba0f838d),
	.w8(32'h3c55ffc3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8b64),
	.w1(32'hbbb0d8e2),
	.w2(32'hb9a26f60),
	.w3(32'h3bcd0915),
	.w4(32'h3c12863c),
	.w5(32'h3c21b5de),
	.w6(32'h3c5b6f07),
	.w7(32'h3b68427e),
	.w8(32'h3b5a9754),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3640f2),
	.w1(32'hbc82b224),
	.w2(32'hbb6cc692),
	.w3(32'h3b8840ec),
	.w4(32'hbc3b2bbf),
	.w5(32'hbc122c81),
	.w6(32'hbc1ad445),
	.w7(32'hbbdf0a7f),
	.w8(32'hb9a926c2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877aca),
	.w1(32'h3b8c7d2c),
	.w2(32'h3bddd1b1),
	.w3(32'h3ab51c93),
	.w4(32'hbb70b3c9),
	.w5(32'h3c1a4d79),
	.w6(32'hbc08b74a),
	.w7(32'hbac761f5),
	.w8(32'hbb802ed8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696b04),
	.w1(32'hbaf0af3d),
	.w2(32'hbc29d77f),
	.w3(32'hba27b155),
	.w4(32'h39b082b6),
	.w5(32'hbc1a540d),
	.w6(32'hbb39d3b8),
	.w7(32'h3ab0dade),
	.w8(32'hbb0cebdc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817039),
	.w1(32'hbb9afc0f),
	.w2(32'h3a8801e9),
	.w3(32'h3bf4d5cb),
	.w4(32'hbbd2b943),
	.w5(32'hbc1336e4),
	.w6(32'hba9aba8b),
	.w7(32'hba2cb8fa),
	.w8(32'hbabebb98),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb329af1),
	.w1(32'h3a0f84e4),
	.w2(32'hbbde215a),
	.w3(32'hbc8f7ca5),
	.w4(32'hbc858670),
	.w5(32'hbb4cfbcd),
	.w6(32'hbc49144a),
	.w7(32'hbbc6fbba),
	.w8(32'hbb19844f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59eb03),
	.w1(32'hbca32351),
	.w2(32'hbb42bff0),
	.w3(32'hbbdc5738),
	.w4(32'hbc4513fd),
	.w5(32'h3b71ba32),
	.w6(32'h3b19e098),
	.w7(32'h3b89236a),
	.w8(32'hba7496a5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea88a2),
	.w1(32'hba9131c3),
	.w2(32'hbc0f0190),
	.w3(32'h3c277599),
	.w4(32'h3b12b8f5),
	.w5(32'hbbc2717b),
	.w6(32'h3ba6f632),
	.w7(32'h3b8b076a),
	.w8(32'hbb17a5b9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9b22d),
	.w1(32'h3c0683a6),
	.w2(32'hbbed214d),
	.w3(32'h3b4ddbb4),
	.w4(32'h3bed5005),
	.w5(32'hbba19941),
	.w6(32'hbb18206c),
	.w7(32'h3ad498bd),
	.w8(32'h3bcad122),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886f5c),
	.w1(32'h3b5e0cbf),
	.w2(32'hbacabfb1),
	.w3(32'h3bb82ed8),
	.w4(32'h3c52e525),
	.w5(32'h3bef6e93),
	.w6(32'h3acf3047),
	.w7(32'h3bca9f34),
	.w8(32'hba0df065),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398a5b),
	.w1(32'hbb738932),
	.w2(32'hbb308d40),
	.w3(32'h3b8b4292),
	.w4(32'hbbfdaeef),
	.w5(32'hba2cb537),
	.w6(32'h3baf4869),
	.w7(32'hbbba6f9b),
	.w8(32'hbbe65ba9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea369a),
	.w1(32'hbba1e391),
	.w2(32'h3bcb3f8a),
	.w3(32'h3c0a782c),
	.w4(32'h3ad86a5b),
	.w5(32'hbb805268),
	.w6(32'hbb0c915e),
	.w7(32'hba7c422b),
	.w8(32'hbba4f95b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be40758),
	.w1(32'h3b2f0d74),
	.w2(32'hbb14b744),
	.w3(32'h3b1b6eea),
	.w4(32'h3b6c1d2c),
	.w5(32'hbbf7c6f1),
	.w6(32'hbba7b986),
	.w7(32'hbc1cd213),
	.w8(32'hbc642c49),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc210d),
	.w1(32'h3b5ee0b5),
	.w2(32'h3aefe34e),
	.w3(32'hbc967396),
	.w4(32'hbba35ec4),
	.w5(32'h3c2bbc90),
	.w6(32'hbb37e917),
	.w7(32'hbb1f261f),
	.w8(32'h3c4a83c9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33b2d4),
	.w1(32'hbacb70d6),
	.w2(32'h3b0cc9ed),
	.w3(32'h3cb5d8a0),
	.w4(32'h3c302073),
	.w5(32'hbc49a14d),
	.w6(32'h3cd01bbd),
	.w7(32'h3c6c2167),
	.w8(32'hbba428c2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a24ee),
	.w1(32'hbbe181ad),
	.w2(32'hbc7c7b21),
	.w3(32'hbc21e1bd),
	.w4(32'hbc870831),
	.w5(32'hbb0c98af),
	.w6(32'hbc1220eb),
	.w7(32'hbbf57978),
	.w8(32'hba9315a7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f2999),
	.w1(32'hbc6870e2),
	.w2(32'hbb58517f),
	.w3(32'hba761d6e),
	.w4(32'hba754268),
	.w5(32'h3b982ea4),
	.w6(32'h3b492dcb),
	.w7(32'h39976601),
	.w8(32'h3c11fa7c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81ecd1),
	.w1(32'h3b1d23b7),
	.w2(32'hbb2ecc65),
	.w3(32'h3c31b51a),
	.w4(32'h3bdb3171),
	.w5(32'hbc990011),
	.w6(32'h3c510dc4),
	.w7(32'h3bbc73ae),
	.w8(32'hbcc34d91),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dd81a),
	.w1(32'hbc65b1b1),
	.w2(32'hbb7e2b57),
	.w3(32'hbce295f2),
	.w4(32'hbcaedc6a),
	.w5(32'h3bd3591c),
	.w6(32'hbcd2fbf0),
	.w7(32'hbcc57578),
	.w8(32'h3c128a3d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e1310f),
	.w1(32'h3b538533),
	.w2(32'h3bc5a67f),
	.w3(32'h3c6cec55),
	.w4(32'h3c7e945b),
	.w5(32'h3c9a8176),
	.w6(32'h3c43885e),
	.w7(32'h3c37b22a),
	.w8(32'h3c48ee86),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab6e7),
	.w1(32'h3bf4303a),
	.w2(32'hbabc8038),
	.w3(32'h3d06638d),
	.w4(32'h3cdf610b),
	.w5(32'hbbbf8d44),
	.w6(32'h3c456beb),
	.w7(32'h3bead53b),
	.w8(32'h3b15605c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74d9cf),
	.w1(32'hbb5e58b5),
	.w2(32'hba8815e1),
	.w3(32'hbbf1ed83),
	.w4(32'hbb3341eb),
	.w5(32'h3bbf2b71),
	.w6(32'hb9499a95),
	.w7(32'h3bec9362),
	.w8(32'h3a6e23a1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab57e3d),
	.w1(32'h39820f4f),
	.w2(32'h394dae23),
	.w3(32'hbb82cd4b),
	.w4(32'hba9ab938),
	.w5(32'hbb0f0cfc),
	.w6(32'h3a6ff84d),
	.w7(32'hb9f7d70f),
	.w8(32'hbabd227f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb898b99),
	.w1(32'hbb7b61e9),
	.w2(32'hbafd6aaa),
	.w3(32'hbb8a6583),
	.w4(32'hbbbe9e25),
	.w5(32'hbb854ff6),
	.w6(32'hbb574d5a),
	.w7(32'hbbd8cd46),
	.w8(32'hbb6e1969),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886900),
	.w1(32'h3b4c6b1a),
	.w2(32'h3ba4a146),
	.w3(32'hbc1e8b95),
	.w4(32'hbb234d80),
	.w5(32'h3c09d8da),
	.w6(32'hbc2baa5b),
	.w7(32'hbc1dc50c),
	.w8(32'hbbd3aff0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d61d5),
	.w1(32'h3bb372ab),
	.w2(32'hbbb9f429),
	.w3(32'h3c3a96a1),
	.w4(32'h3aff3bd9),
	.w5(32'h38092972),
	.w6(32'hbc45f62b),
	.w7(32'hbbcae12c),
	.w8(32'h3bb27459),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b107251),
	.w1(32'h3aff8fb7),
	.w2(32'hbc11eb6a),
	.w3(32'h3c081175),
	.w4(32'h3be066ab),
	.w5(32'h398697e7),
	.w6(32'h3c14b7dd),
	.w7(32'h3bc4039c),
	.w8(32'h3bd5d651),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85058b),
	.w1(32'hbbb59327),
	.w2(32'h3b807cbe),
	.w3(32'h3c567c9b),
	.w4(32'h3a232ad3),
	.w5(32'h3bf94657),
	.w6(32'hbae2632d),
	.w7(32'hbb81c896),
	.w8(32'h3c24545e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b271f38),
	.w1(32'hbb35dbeb),
	.w2(32'h3c384c04),
	.w3(32'h3b214ba4),
	.w4(32'h3ba862ea),
	.w5(32'h3c28ceb2),
	.w6(32'h3c39f4a9),
	.w7(32'h3c4dbf32),
	.w8(32'h3b9faec9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c916eee),
	.w1(32'h3bf7d8b8),
	.w2(32'hbbdda738),
	.w3(32'h3c63ba13),
	.w4(32'h3c06f6db),
	.w5(32'hbc347568),
	.w6(32'h3c048a41),
	.w7(32'h3bb66716),
	.w8(32'h3b6400d6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4ae0c),
	.w1(32'h3aea99e4),
	.w2(32'h3af32c5f),
	.w3(32'hbc1b338d),
	.w4(32'hbacf373e),
	.w5(32'h3baf5c03),
	.w6(32'h3b994609),
	.w7(32'h3b521842),
	.w8(32'h3c0a6abd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878bc9),
	.w1(32'h3c0f4cd5),
	.w2(32'hbb950cdc),
	.w3(32'h3a6ea83e),
	.w4(32'h39e3eba1),
	.w5(32'hbbcdb32f),
	.w6(32'h3bc21f55),
	.w7(32'h3b91d67c),
	.w8(32'h3c4cdb0e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec25f4),
	.w1(32'h3b45b087),
	.w2(32'h3a68cf61),
	.w3(32'h3bf0f0de),
	.w4(32'h3b503abe),
	.w5(32'h3bb151dd),
	.w6(32'h3ca48110),
	.w7(32'h3c99761c),
	.w8(32'h3b341804),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b313f53),
	.w1(32'hbb3a4e07),
	.w2(32'h3bdf07e6),
	.w3(32'h3be5e4bb),
	.w4(32'h3b61c03f),
	.w5(32'hbcbb236d),
	.w6(32'h3b967297),
	.w7(32'h3a198744),
	.w8(32'hbcd9d53f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7bddd),
	.w1(32'hbbdd2983),
	.w2(32'h3c5ff9fc),
	.w3(32'hbd068c4e),
	.w4(32'hbccec25b),
	.w5(32'h3c2ca4e3),
	.w6(32'hbc95420f),
	.w7(32'hbbfe7104),
	.w8(32'h3b66362b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6bddf),
	.w1(32'h3c34e1b4),
	.w2(32'h3af94a30),
	.w3(32'h3bffb4de),
	.w4(32'h3bed0879),
	.w5(32'hbb4b4c7c),
	.w6(32'hb95a0e5e),
	.w7(32'h3c0b690f),
	.w8(32'hb96cd6d4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb468b5e),
	.w1(32'hbbb0afd4),
	.w2(32'hbb851cd0),
	.w3(32'hbc676752),
	.w4(32'hbc302ef4),
	.w5(32'hba75416f),
	.w6(32'hbbd30a10),
	.w7(32'hbbb4d8d0),
	.w8(32'h3c0642b6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab56c),
	.w1(32'h3ac2a403),
	.w2(32'h3a9f8dd6),
	.w3(32'h3bf43be1),
	.w4(32'h3b809c3f),
	.w5(32'hbc644286),
	.w6(32'h3c1f7283),
	.w7(32'h3bdd7abc),
	.w8(32'hbc828a76),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbfc87),
	.w1(32'hbbe03020),
	.w2(32'h3c02164e),
	.w3(32'hbcb2760d),
	.w4(32'hbc4de596),
	.w5(32'h3c1396f7),
	.w6(32'hbc98b429),
	.w7(32'hbc2bacff),
	.w8(32'h3bf0f122),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b828a60),
	.w1(32'h3b2ba070),
	.w2(32'h39dbf4cf),
	.w3(32'h3bac18cf),
	.w4(32'hbb14673a),
	.w5(32'hb95669e2),
	.w6(32'h3b8185ec),
	.w7(32'hbba9d6aa),
	.w8(32'h3af2d7e5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6efc66),
	.w1(32'hbb3aec56),
	.w2(32'h3bbce385),
	.w3(32'hba879778),
	.w4(32'h3b1092b8),
	.w5(32'h3a060714),
	.w6(32'h3a144b01),
	.w7(32'h3b54a495),
	.w8(32'h3a3663a8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5dc3e),
	.w1(32'h3bb511a3),
	.w2(32'hbb1b91ee),
	.w3(32'h3a85c9ff),
	.w4(32'hbb3b6284),
	.w5(32'hbae99b73),
	.w6(32'h3b49966b),
	.w7(32'hbb66eb66),
	.w8(32'hbbb2cf7d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08ba30),
	.w1(32'hbb8ce200),
	.w2(32'h3c0d5a4d),
	.w3(32'hbbdf9b94),
	.w4(32'hbb8715fa),
	.w5(32'hb9271b2c),
	.w6(32'hbb300735),
	.w7(32'hbbaa95b7),
	.w8(32'h3c1b81b9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be602cd),
	.w1(32'h3b8ac94d),
	.w2(32'h3aa98eb4),
	.w3(32'h3c1db5ab),
	.w4(32'hbb6f469b),
	.w5(32'h39da7386),
	.w6(32'h3c1adda3),
	.w7(32'h3b7a06eb),
	.w8(32'hba138716),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01ebab),
	.w1(32'h3ae1ff66),
	.w2(32'hb7be1d01),
	.w3(32'hb96530a0),
	.w4(32'h3ba8689d),
	.w5(32'h3c1d2374),
	.w6(32'h3a27bec9),
	.w7(32'h3aa8f060),
	.w8(32'h3c13edd6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ddaf),
	.w1(32'h3b27e09b),
	.w2(32'hbb0b7d3f),
	.w3(32'h3c80a063),
	.w4(32'h3c3117e8),
	.w5(32'hb9e6e9f7),
	.w6(32'h3c2321cd),
	.w7(32'h3bf70dcf),
	.w8(32'h3b382750),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ebe6),
	.w1(32'hbb6bdfde),
	.w2(32'hbbd0dded),
	.w3(32'hba9bccea),
	.w4(32'h3ad93953),
	.w5(32'hbbaa0f2b),
	.w6(32'h3b875316),
	.w7(32'h3ba48378),
	.w8(32'hbb8e114a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9a0be),
	.w1(32'hbb437817),
	.w2(32'h3ac6cd78),
	.w3(32'hbbba3ad5),
	.w4(32'hbbb4fb67),
	.w5(32'h39864f35),
	.w6(32'hbbb17f8a),
	.w7(32'hbb9a9bb3),
	.w8(32'h3b9150e5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a662419),
	.w1(32'h3b81c23e),
	.w2(32'hbb66f9fe),
	.w3(32'h3bb599ee),
	.w4(32'h3a42ce30),
	.w5(32'hbb8fffed),
	.w6(32'h3b09c5b0),
	.w7(32'hba06fa6f),
	.w8(32'h3bf2740c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222ae8),
	.w1(32'hbbe5af48),
	.w2(32'hbbe73585),
	.w3(32'hba89391d),
	.w4(32'h3a4687a0),
	.w5(32'hbb78f3d1),
	.w6(32'h3b83a5bf),
	.w7(32'hbb0578f2),
	.w8(32'h3b0c43d2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b0e08),
	.w1(32'h3a7bb090),
	.w2(32'h3b774656),
	.w3(32'hbb63f8da),
	.w4(32'hbbbf59cd),
	.w5(32'h3983d834),
	.w6(32'hbba5d04c),
	.w7(32'hbbe5e980),
	.w8(32'h3b7cbb54),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abef8b8),
	.w1(32'h3a027188),
	.w2(32'h3b420575),
	.w3(32'h3ae56694),
	.w4(32'hb94d0a6d),
	.w5(32'hbc0ffdad),
	.w6(32'h3ad1184b),
	.w7(32'hbb85a284),
	.w8(32'hbc901353),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c40ca),
	.w1(32'hbb67ef6e),
	.w2(32'hbaefda1d),
	.w3(32'hbc274aca),
	.w4(32'hbc12ddb1),
	.w5(32'hbb41916e),
	.w6(32'hbc113582),
	.w7(32'hbc014347),
	.w8(32'hbb65725b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde86a8),
	.w1(32'hbae860a8),
	.w2(32'h3b97af54),
	.w3(32'hbbb50bea),
	.w4(32'hbb97b084),
	.w5(32'h3ada5d5d),
	.w6(32'hbaea3111),
	.w7(32'hbb774aa0),
	.w8(32'h3be4feb3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f785),
	.w1(32'h3c1abc34),
	.w2(32'hbc2059b4),
	.w3(32'h3c2fd836),
	.w4(32'h3c1a90d4),
	.w5(32'hbbfda932),
	.w6(32'h3b05ca9c),
	.w7(32'h3b77f797),
	.w8(32'hbc131a38),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b9b9),
	.w1(32'h3a0c9bab),
	.w2(32'hbb1d1d88),
	.w3(32'h3a38f8a5),
	.w4(32'hbb2473fb),
	.w5(32'h3c1ccd65),
	.w6(32'hbbc43d52),
	.w7(32'hbc0a3e81),
	.w8(32'h3bd174e7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e1577),
	.w1(32'h3bc9553e),
	.w2(32'hba691e2e),
	.w3(32'h3c33803f),
	.w4(32'h3bec8eb7),
	.w5(32'hbafc988a),
	.w6(32'h3c2a2d5a),
	.w7(32'h39d91c64),
	.w8(32'hb96214be),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90d0c),
	.w1(32'h3b4b550d),
	.w2(32'h3c63b847),
	.w3(32'hbbd5130a),
	.w4(32'h3b98023d),
	.w5(32'h3c0e3e3a),
	.w6(32'hbb277a4b),
	.w7(32'h3ba4dae4),
	.w8(32'h3bd496fa),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7304ca),
	.w1(32'h3c2c3c96),
	.w2(32'h3c3c1761),
	.w3(32'hbc6bd96a),
	.w4(32'h3bcd5b32),
	.w5(32'h3c5acd5b),
	.w6(32'hbc7491cb),
	.w7(32'h3c2c3625),
	.w8(32'h3b46c8a4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d28ff),
	.w1(32'h3c2522b1),
	.w2(32'hbc45567b),
	.w3(32'h3c2d0022),
	.w4(32'h3c3a5010),
	.w5(32'hbc3d4e27),
	.w6(32'h3c5529b0),
	.w7(32'h3c1a2a82),
	.w8(32'hbb1573db),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a8442),
	.w1(32'hbb05712c),
	.w2(32'h3b027cc3),
	.w3(32'hbbb9b0fa),
	.w4(32'h3ba2b7f4),
	.w5(32'hbc0a1ee4),
	.w6(32'h3b5828d4),
	.w7(32'h3c0fc23d),
	.w8(32'hba93b487),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3573d),
	.w1(32'h3949e7d3),
	.w2(32'hb9b90541),
	.w3(32'hbb6611af),
	.w4(32'h39b39f3c),
	.w5(32'hbc173bee),
	.w6(32'hbbab50fe),
	.w7(32'hbc1fba21),
	.w8(32'hbba38b76),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc91ae0),
	.w1(32'hbae41b15),
	.w2(32'hbca69587),
	.w3(32'h3b10f9fd),
	.w4(32'h3b37fb76),
	.w5(32'hbc5421ec),
	.w6(32'h3b28c19e),
	.w7(32'h3b5a453b),
	.w8(32'hba100766),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43f661),
	.w1(32'h3aa88e0a),
	.w2(32'h3ba30c8e),
	.w3(32'h3bad6d68),
	.w4(32'h3cc8f4e8),
	.w5(32'hbaa99834),
	.w6(32'h3ca59da6),
	.w7(32'h3d08136e),
	.w8(32'hbbfc8957),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba676ae),
	.w1(32'h3afef69a),
	.w2(32'hbbaceef9),
	.w3(32'hbc37d02f),
	.w4(32'hbac82fa2),
	.w5(32'hb9e28f8a),
	.w6(32'hbbdf3677),
	.w7(32'hbbe449d0),
	.w8(32'h3930db6a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb687b),
	.w1(32'hbb5e76e0),
	.w2(32'h3c819dae),
	.w3(32'hba88f402),
	.w4(32'h3bc38cd2),
	.w5(32'h3c598662),
	.w6(32'h3ad4eb3e),
	.w7(32'h3ba9fad9),
	.w8(32'h3c466fb9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50f54d),
	.w1(32'h3bde602b),
	.w2(32'hbd00f876),
	.w3(32'h3c01d59d),
	.w4(32'h3bf61f0b),
	.w5(32'hbcf187bf),
	.w6(32'h3c367b87),
	.w7(32'h3c0f4fbf),
	.w8(32'hbbdad6e0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbf2fc),
	.w1(32'hbb3cd425),
	.w2(32'h3c5f51eb),
	.w3(32'hbc126093),
	.w4(32'h3cc73e8d),
	.w5(32'h3c8c795a),
	.w6(32'h3cb5d692),
	.w7(32'h3d415230),
	.w8(32'h3bf16271),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b5dea),
	.w1(32'h3b2e6d9f),
	.w2(32'hbb83a23d),
	.w3(32'h3bd3fdfc),
	.w4(32'hba3a226d),
	.w5(32'hbb52ff76),
	.w6(32'hbaeae94c),
	.w7(32'hb97a910e),
	.w8(32'h3b5b5b67),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fafa9),
	.w1(32'h3a641272),
	.w2(32'h3bbd5ee3),
	.w3(32'h3b0979c6),
	.w4(32'hbbbfde55),
	.w5(32'h3add1431),
	.w6(32'h3c1da144),
	.w7(32'hbbc9b792),
	.w8(32'h3b84b2ef),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbb2f7),
	.w1(32'h3b6b52fb),
	.w2(32'hbadebe45),
	.w3(32'h3b87bd14),
	.w4(32'hbc395609),
	.w5(32'hbc73b3d0),
	.w6(32'hbc1e0e5c),
	.w7(32'hbc5c3d8c),
	.w8(32'hbbc6d1f1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad95d71),
	.w1(32'h3bad64cc),
	.w2(32'hb8243a91),
	.w3(32'hbbf173c6),
	.w4(32'hbb979610),
	.w5(32'h3c7c31c7),
	.w6(32'hbc3bd37f),
	.w7(32'hbb2cb41e),
	.w8(32'h3bdecc60),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25e456),
	.w1(32'h3c2dfb37),
	.w2(32'hbb65b053),
	.w3(32'h3c4e67c9),
	.w4(32'h3c09e192),
	.w5(32'h3abd04dd),
	.w6(32'h3c5306e5),
	.w7(32'h3be5b8ea),
	.w8(32'h3a9e3118),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4856ba),
	.w1(32'h3c12c74d),
	.w2(32'hb9a4ff1c),
	.w3(32'h3b1ecfc5),
	.w4(32'h3c826b83),
	.w5(32'h3ac509d3),
	.w6(32'h3c0bb1c7),
	.w7(32'h3c9c6700),
	.w8(32'hbb974411),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4789f),
	.w1(32'h3adb2d69),
	.w2(32'hbc32d152),
	.w3(32'hbc163178),
	.w4(32'h3b591c46),
	.w5(32'hbbd2f4b3),
	.w6(32'hbb42fc28),
	.w7(32'hba314af8),
	.w8(32'h3ae71c86),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44c5a5),
	.w1(32'hba84c5fc),
	.w2(32'h3c1458b9),
	.w3(32'hbc10b4a1),
	.w4(32'hbb93f3bf),
	.w5(32'h3c381767),
	.w6(32'hbc44b4ef),
	.w7(32'h39a25e68),
	.w8(32'h3b045ced),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be49c19),
	.w1(32'hbb507094),
	.w2(32'hbbdf9705),
	.w3(32'h3ad6e7e7),
	.w4(32'hbbf5d5bc),
	.w5(32'hbb831ccb),
	.w6(32'h3b1addf5),
	.w7(32'hbb924c07),
	.w8(32'h3af31ee8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8d9f),
	.w1(32'hb88df7c5),
	.w2(32'hbb19704a),
	.w3(32'h3bda7614),
	.w4(32'h3bb62a75),
	.w5(32'hb9228c5b),
	.w6(32'h3c3a3b56),
	.w7(32'h3c30843d),
	.w8(32'h39ec480f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b855),
	.w1(32'h3a2d0e26),
	.w2(32'hbac00163),
	.w3(32'hbb243eaa),
	.w4(32'h3a82558e),
	.w5(32'hbc4b524b),
	.w6(32'h3a3b4c4b),
	.w7(32'h3b946588),
	.w8(32'hbc4170ab),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79586a),
	.w1(32'hbc1d5350),
	.w2(32'h3c11a239),
	.w3(32'hbce7dcde),
	.w4(32'hbcb1f4c7),
	.w5(32'h3c4ac39e),
	.w6(32'hbcfbf21d),
	.w7(32'hbcd5f9db),
	.w8(32'h3ba220d5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2382c),
	.w1(32'h3c27f7b9),
	.w2(32'h3ad63a5d),
	.w3(32'h3c56b89f),
	.w4(32'h3bc02044),
	.w5(32'h3b88252a),
	.w6(32'h3bf30c9a),
	.w7(32'h3b87d1b8),
	.w8(32'h3c24e16c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b135374),
	.w1(32'h3c01ff4d),
	.w2(32'h3c22b605),
	.w3(32'h3c9999e2),
	.w4(32'h3c85a3a5),
	.w5(32'h3c571f72),
	.w6(32'h3cb687b8),
	.w7(32'h3b50c726),
	.w8(32'h3a4ddbef),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae299af),
	.w1(32'h3bc51356),
	.w2(32'hbbaaf2a6),
	.w3(32'hbc129f57),
	.w4(32'hbb8784ec),
	.w5(32'hbb34748b),
	.w6(32'hbbdce301),
	.w7(32'h3b339504),
	.w8(32'h3bab2f3a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c434a1d),
	.w1(32'h3c8e4094),
	.w2(32'hbc51ce1b),
	.w3(32'h3c8e0bf8),
	.w4(32'h3cc430d8),
	.w5(32'hbc378303),
	.w6(32'h3bacca04),
	.w7(32'hbb4a9cbd),
	.w8(32'hbc7e1ccb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ac627),
	.w1(32'h3ab4f782),
	.w2(32'hbb12e33e),
	.w3(32'hbcad97aa),
	.w4(32'hbbe53b4d),
	.w5(32'hbbddc15f),
	.w6(32'hb987d2b6),
	.w7(32'hbc145434),
	.w8(32'hbb937727),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031444),
	.w1(32'h3b390206),
	.w2(32'h3a6d3e2f),
	.w3(32'hbbd0d195),
	.w4(32'h3b700bab),
	.w5(32'hbba1cf39),
	.w6(32'hbc18fc88),
	.w7(32'hbb8c7ae8),
	.w8(32'h3b4c306a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b212135),
	.w1(32'hbbc360dd),
	.w2(32'hbcf3a140),
	.w3(32'hbc45c14f),
	.w4(32'hbbc470f1),
	.w5(32'hbd592519),
	.w6(32'h3a019f68),
	.w7(32'hbb9f7fff),
	.w8(32'hbd6a0673),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd70ec61),
	.w1(32'hbd29773c),
	.w2(32'hbb954039),
	.w3(32'hbdae3f49),
	.w4(32'hbd544956),
	.w5(32'hbbdf19fc),
	.w6(32'hbda62ae1),
	.w7(32'hbd007962),
	.w8(32'h3c1e1d50),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd571e0),
	.w1(32'h3bc4b28e),
	.w2(32'hbc658c52),
	.w3(32'hbb61cbc6),
	.w4(32'h3c3db334),
	.w5(32'hbd02fdcf),
	.w6(32'h3c7b810a),
	.w7(32'h3ced64ed),
	.w8(32'hbcfd70c6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05d6ca),
	.w1(32'hbce8e135),
	.w2(32'h3aa439ad),
	.w3(32'hbd511576),
	.w4(32'hbd359708),
	.w5(32'h3ac9cf8f),
	.w6(32'hbcd3c098),
	.w7(32'hbc1faf70),
	.w8(32'h3c8cd59e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dcd38),
	.w1(32'h3cbbd41d),
	.w2(32'h3b7e5aea),
	.w3(32'hbb77eb53),
	.w4(32'h3c3cb783),
	.w5(32'h3c8a28fb),
	.w6(32'hbc4910fe),
	.w7(32'h39bf761e),
	.w8(32'h3becc851),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47656b),
	.w1(32'h3a8424cb),
	.w2(32'h3a61d8a0),
	.w3(32'h3c41401a),
	.w4(32'hbbb1f016),
	.w5(32'hbb2abfaf),
	.w6(32'h3ba93a65),
	.w7(32'hbb787326),
	.w8(32'hbac08171),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57ba84),
	.w1(32'h3b1aa684),
	.w2(32'h3b19be6c),
	.w3(32'hbaf5eda1),
	.w4(32'hbc2aece7),
	.w5(32'h3ba6b6c2),
	.w6(32'hbb3b7ae4),
	.w7(32'hbbb36c66),
	.w8(32'h3bb775eb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027f7e),
	.w1(32'h3b74c775),
	.w2(32'hbbda8eb7),
	.w3(32'hbaa85bcd),
	.w4(32'h39607c6c),
	.w5(32'hbb94c43b),
	.w6(32'hbc57ce48),
	.w7(32'hbcb74aaf),
	.w8(32'hbb445a1b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c7d5),
	.w1(32'hbae32018),
	.w2(32'hbae7cb47),
	.w3(32'hbad06efb),
	.w4(32'h390bbbd8),
	.w5(32'hbbfbb0e3),
	.w6(32'hbba4973b),
	.w7(32'hbb0421db),
	.w8(32'hbbbfd0e8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25b168),
	.w1(32'h3b1c0914),
	.w2(32'h3b326cac),
	.w3(32'hbbfc271c),
	.w4(32'hba9a3873),
	.w5(32'h3b85602b),
	.w6(32'hbc1ddd60),
	.w7(32'hbbddb158),
	.w8(32'h3b855cfa),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d4d15),
	.w1(32'h3b949903),
	.w2(32'h3b88f151),
	.w3(32'h3c0dca14),
	.w4(32'h3c768739),
	.w5(32'hbad85dba),
	.w6(32'h3c53bbbc),
	.w7(32'h3c8c6c3c),
	.w8(32'hbb8bbfef),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2f8be),
	.w1(32'h3bc64204),
	.w2(32'hbbc5f149),
	.w3(32'hbc3c061c),
	.w4(32'h3a83f546),
	.w5(32'hbba27126),
	.w6(32'hbba36902),
	.w7(32'hba5942c4),
	.w8(32'hbb54cf4c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abab245),
	.w1(32'h3ba82691),
	.w2(32'h3b8f262f),
	.w3(32'h3bb9c192),
	.w4(32'h3bacfa26),
	.w5(32'h3ad0908a),
	.w6(32'hbb190360),
	.w7(32'h3a851662),
	.w8(32'hbb675fce),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42df3),
	.w1(32'hbb9ba537),
	.w2(32'h3c60b006),
	.w3(32'hbc06b982),
	.w4(32'hbbee9420),
	.w5(32'h3d177cf5),
	.w6(32'hbc43c649),
	.w7(32'hbc4b2d52),
	.w8(32'h3d491e32),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51dc14),
	.w1(32'h3be29c53),
	.w2(32'hbc2c32f3),
	.w3(32'h3d2dfe76),
	.w4(32'h3c213e36),
	.w5(32'hbc38c775),
	.w6(32'h3d16d4f3),
	.w7(32'hb968f0d5),
	.w8(32'hbb44f1c7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc471332),
	.w1(32'h3b2d94ce),
	.w2(32'h39fc8380),
	.w3(32'hbc5e3e57),
	.w4(32'hbaedbe6a),
	.w5(32'h3adc20e6),
	.w6(32'hbc18c2aa),
	.w7(32'h3a88e00a),
	.w8(32'h392dbd7c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a83cb),
	.w1(32'h3a8fd221),
	.w2(32'h3b678781),
	.w3(32'hb9149744),
	.w4(32'h392fec78),
	.w5(32'hbbaade91),
	.w6(32'h3bac05f6),
	.w7(32'hbb15a3b0),
	.w8(32'h3c2826d8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9316e9),
	.w1(32'h3b57e57c),
	.w2(32'hb9925e8b),
	.w3(32'h3b3bd142),
	.w4(32'h3be4bee9),
	.w5(32'hb9ce0cc0),
	.w6(32'h3c36dde8),
	.w7(32'h3c0badf3),
	.w8(32'h3bc3e3c7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e4d45),
	.w1(32'h3c2c9776),
	.w2(32'hbcd1ec69),
	.w3(32'hbbb79c09),
	.w4(32'h3c1f765e),
	.w5(32'hbc9f02cd),
	.w6(32'h3b650ead),
	.w7(32'h3c6c2ae1),
	.w8(32'hbc0cb4af),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7e8b3),
	.w1(32'h3a5617bb),
	.w2(32'hb98925d7),
	.w3(32'hbbc66773),
	.w4(32'h3ca74aa8),
	.w5(32'hbb940a4d),
	.w6(32'h3a0c9c71),
	.w7(32'h3ce3741c),
	.w8(32'h3b3799fe),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb789bb9c),
	.w1(32'h3b5ec430),
	.w2(32'h3978245e),
	.w3(32'hbb27f8ad),
	.w4(32'hbba240a8),
	.w5(32'h39012302),
	.w6(32'hbb53d978),
	.w7(32'hbb8e8e9d),
	.w8(32'h3bc073c7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe3e71),
	.w1(32'h3b280d56),
	.w2(32'hbc264dff),
	.w3(32'h3abd8008),
	.w4(32'h3bd5ee05),
	.w5(32'hbc3784c2),
	.w6(32'h3a7bf376),
	.w7(32'hba3b1fcc),
	.w8(32'hbbffc6b2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910873),
	.w1(32'hb997b6a5),
	.w2(32'hbb347954),
	.w3(32'hbc201de1),
	.w4(32'hbb9858c0),
	.w5(32'hbb9475c6),
	.w6(32'hbc8ad032),
	.w7(32'hbbc1fe09),
	.w8(32'hb9b9ca9d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0700a),
	.w1(32'h3adfbe67),
	.w2(32'hbc1ffa3a),
	.w3(32'hbc44658d),
	.w4(32'hb9e5a307),
	.w5(32'h39810d7f),
	.w6(32'hbba49de1),
	.w7(32'h3b46dbd6),
	.w8(32'h3b736623),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61a4c2),
	.w1(32'hbc1dcd30),
	.w2(32'hbc71ebfc),
	.w3(32'h3a21bc99),
	.w4(32'hb76dc7d4),
	.w5(32'hbc587e19),
	.w6(32'h3bceb23d),
	.w7(32'hbbcafbe2),
	.w8(32'hbb0e0bc8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc154a3d),
	.w1(32'h3b991638),
	.w2(32'hba438dd7),
	.w3(32'hbb91668d),
	.w4(32'h3c4c0aa6),
	.w5(32'h3ac77a0d),
	.w6(32'h3b19b5b8),
	.w7(32'h3c8ad5b5),
	.w8(32'h3a10706e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03be91),
	.w1(32'hbbd46d1b),
	.w2(32'h3c4ad407),
	.w3(32'hbc011bdd),
	.w4(32'hbbce03cd),
	.w5(32'h3bcde1b3),
	.w6(32'hbbecd4e0),
	.w7(32'hbbe0d306),
	.w8(32'h3b1abd9c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f352b),
	.w1(32'h3c05ccf8),
	.w2(32'h3ae267fd),
	.w3(32'h3c586d78),
	.w4(32'h3b8f67ca),
	.w5(32'h3ab6de06),
	.w6(32'h3b493a73),
	.w7(32'h3a08b791),
	.w8(32'h3bd6691c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6f76a),
	.w1(32'hba7cea54),
	.w2(32'h3c870197),
	.w3(32'h3c16dbdd),
	.w4(32'h3b3af715),
	.w5(32'h3c957571),
	.w6(32'h3bbf7b6c),
	.w7(32'h3b2e6ad9),
	.w8(32'h3c407709),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a7775),
	.w1(32'h3c0bf9ee),
	.w2(32'hbc7814b6),
	.w3(32'h3bb840de),
	.w4(32'h3b03de47),
	.w5(32'hbcc0afb2),
	.w6(32'hbb819af6),
	.w7(32'hbb3de707),
	.w8(32'hbc9c8799),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd613e),
	.w1(32'hbb8aa142),
	.w2(32'hbbaac1b2),
	.w3(32'hbd10f553),
	.w4(32'hbc66366a),
	.w5(32'hbbf43a54),
	.w6(32'hbcf52b30),
	.w7(32'hbc9b542d),
	.w8(32'hbc4901ed),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b58c9),
	.w1(32'hbbd185d5),
	.w2(32'h3bc61d4f),
	.w3(32'hbc4d9940),
	.w4(32'hbc1710b9),
	.w5(32'hbae95323),
	.w6(32'hbc53005c),
	.w7(32'hbc3720b9),
	.w8(32'hbb8e93ab),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af417c7),
	.w1(32'hba265a63),
	.w2(32'h3ae38b25),
	.w3(32'hbb97f786),
	.w4(32'h3be66597),
	.w5(32'hb9d39bde),
	.w6(32'hbb6736fd),
	.w7(32'h3b87f607),
	.w8(32'hb8e0bd5e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06fdf8),
	.w1(32'hbbb925b9),
	.w2(32'h3a25b7d2),
	.w3(32'h3c314b6f),
	.w4(32'h3b740210),
	.w5(32'hbbf59d08),
	.w6(32'h3c5d6729),
	.w7(32'h3c4bd851),
	.w8(32'hbc325e40),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1565b9),
	.w1(32'hbaeb9404),
	.w2(32'h3d515da2),
	.w3(32'h3aca198f),
	.w4(32'h3c843a9e),
	.w5(32'h3d3ae355),
	.w6(32'h3c88cc92),
	.w7(32'h3c97978a),
	.w8(32'h3d03ecab),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d24f3b5),
	.w1(32'h3c5eeae3),
	.w2(32'hbc3e8f8e),
	.w3(32'h3cde760a),
	.w4(32'hbc1ca8b3),
	.w5(32'hbc3b5218),
	.w6(32'h39fb105e),
	.w7(32'hbccde5cd),
	.w8(32'hbc0b6f90),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194fb7),
	.w1(32'hbb860893),
	.w2(32'hbaa2337d),
	.w3(32'hbb40cb21),
	.w4(32'h3a221cf1),
	.w5(32'h3a150407),
	.w6(32'hbb9d4496),
	.w7(32'hbb2d35cf),
	.w8(32'hbbca73ca),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de3c89),
	.w1(32'hbb789e07),
	.w2(32'hbb456b76),
	.w3(32'hbb9a23af),
	.w4(32'hbc3159b3),
	.w5(32'hba8d409b),
	.w6(32'hbc73c52c),
	.w7(32'hbc920f9e),
	.w8(32'hbb4b01d8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01e8a1),
	.w1(32'h3b2b06e3),
	.w2(32'h3b8ea8e8),
	.w3(32'hba253011),
	.w4(32'h374a9301),
	.w5(32'h3c2ac546),
	.w6(32'hbb29fa69),
	.w7(32'h3b65d1f5),
	.w8(32'h3afc7bbb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb334d19),
	.w1(32'h3a3a4443),
	.w2(32'hbc8653bd),
	.w3(32'h3bb6c41a),
	.w4(32'h3bbd8d27),
	.w5(32'hbcf7037a),
	.w6(32'hbb391af9),
	.w7(32'h3be65c79),
	.w8(32'hbbbea1b8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbc312),
	.w1(32'hbc2a035b),
	.w2(32'h3c0d49bb),
	.w3(32'hbcf6be4d),
	.w4(32'hbb9799b3),
	.w5(32'h3b6f7ac2),
	.w6(32'hbb6c12c2),
	.w7(32'h3c875330),
	.w8(32'h3ae9b994),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301478),
	.w1(32'h3b987c4e),
	.w2(32'hbc2ad9be),
	.w3(32'h3b406030),
	.w4(32'h3b46b93c),
	.w5(32'hbc7e6a10),
	.w6(32'h3bee213e),
	.w7(32'h3c15f35b),
	.w8(32'hbc66ae69),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc619176),
	.w1(32'hbbbbafa6),
	.w2(32'hbc5daeee),
	.w3(32'hbc8f1fa9),
	.w4(32'hbc38437f),
	.w5(32'hbb8b18fa),
	.w6(32'hbc7d09b9),
	.w7(32'hb8d2d442),
	.w8(32'h39c9cb45),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30cd9c),
	.w1(32'hbc1a17b6),
	.w2(32'h3b809a0d),
	.w3(32'hb95388bc),
	.w4(32'h3ae823bb),
	.w5(32'hbb75b7cd),
	.w6(32'h3c91801c),
	.w7(32'h3c0e3f67),
	.w8(32'hbba8449f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac61375),
	.w1(32'h3ae22b57),
	.w2(32'hbb7630b4),
	.w3(32'h3a24f301),
	.w4(32'h3b7d8959),
	.w5(32'hbae41219),
	.w6(32'hbba65190),
	.w7(32'hbb229903),
	.w8(32'hbac69bdc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8243e),
	.w1(32'h3b249a7f),
	.w2(32'hbbfddd6b),
	.w3(32'hbb8a7be6),
	.w4(32'hbb0a952d),
	.w5(32'hbc5f47b6),
	.w6(32'hb92ccfb6),
	.w7(32'h3b4f2638),
	.w8(32'hbc17c19d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd14404),
	.w1(32'hbbf84a2c),
	.w2(32'h3a7f6010),
	.w3(32'hbcd62e68),
	.w4(32'hbcc66c2a),
	.w5(32'h3c67d3bf),
	.w6(32'hbca0e2da),
	.w7(32'hbc8b13cb),
	.w8(32'h3c636368),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c86a5),
	.w1(32'h3c1a0dd3),
	.w2(32'h3b968d5e),
	.w3(32'h3cc9dbfe),
	.w4(32'h3c6af9d4),
	.w5(32'hbb897cf9),
	.w6(32'h3c7f7752),
	.w7(32'h3b40581c),
	.w8(32'h3b311180),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c26e),
	.w1(32'h3b36ab37),
	.w2(32'hbc0b5b30),
	.w3(32'hbbddfd29),
	.w4(32'h3a8f9ed9),
	.w5(32'hbc7423f7),
	.w6(32'h3b6edf62),
	.w7(32'h3c0185b7),
	.w8(32'hbc5dcbd2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca95923),
	.w1(32'hbc0824fb),
	.w2(32'hbcbcfee5),
	.w3(32'hbceacd81),
	.w4(32'hbc6d1878),
	.w5(32'hbcbfd1e6),
	.w6(32'hbce4fd4e),
	.w7(32'hbc9220a5),
	.w8(32'hbc9e0c7a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7aea0),
	.w1(32'hbc329eb7),
	.w2(32'hbbc64aaa),
	.w3(32'hbcea5e84),
	.w4(32'hbb5f86e9),
	.w5(32'hbbd4ae10),
	.w6(32'hbce8b4e2),
	.w7(32'hbb9aa24d),
	.w8(32'h3b1fff88),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a508a),
	.w1(32'hbba54a23),
	.w2(32'h3bbd9c56),
	.w3(32'hbc4ec0ab),
	.w4(32'hbc5d831c),
	.w5(32'h3b756455),
	.w6(32'h3b13204c),
	.w7(32'hba7fd896),
	.w8(32'hbac5cd00),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afabe45),
	.w1(32'h3aa69556),
	.w2(32'h3ad1fe3a),
	.w3(32'hba9eea16),
	.w4(32'h39360691),
	.w5(32'hbbd1f006),
	.w6(32'h3b625d2b),
	.w7(32'hba94c4bc),
	.w8(32'hbba03031),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb203985),
	.w1(32'h3ba9f9fe),
	.w2(32'h3ba356f7),
	.w3(32'hbc1e0699),
	.w4(32'hbc008f0f),
	.w5(32'h3b0ed8e2),
	.w6(32'hbc7684c8),
	.w7(32'hbc2dbc6e),
	.w8(32'h3b264ee0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cd7a2),
	.w1(32'h3a83e695),
	.w2(32'hbbb1af10),
	.w3(32'h3beb5716),
	.w4(32'hb855f796),
	.w5(32'hbbe43d79),
	.w6(32'h3b8876be),
	.w7(32'h3bcf3413),
	.w8(32'hba5a8dd3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb14d7d),
	.w1(32'h376244ac),
	.w2(32'hbb568cd7),
	.w3(32'h3a94a162),
	.w4(32'h3b82faca),
	.w5(32'h3b3a9ce6),
	.w6(32'h3ae0367e),
	.w7(32'h3af03645),
	.w8(32'h3ac51e25),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc198e1f),
	.w1(32'hba0ceedd),
	.w2(32'h3b34a6af),
	.w3(32'hbc70c1b6),
	.w4(32'hbaec5090),
	.w5(32'h3becb897),
	.w6(32'hbbe1fdbf),
	.w7(32'hbc8fd638),
	.w8(32'h3b77cf29),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d5686),
	.w1(32'h3b8f9e7c),
	.w2(32'hbc5a291f),
	.w3(32'hbbc28ead),
	.w4(32'h3acf5d41),
	.w5(32'hbc6cc6b6),
	.w6(32'hbb8bc24c),
	.w7(32'h3bc699f5),
	.w8(32'hbc0180a4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ce04b),
	.w1(32'hbbfb8d37),
	.w2(32'hbc0312c4),
	.w3(32'hbc50faef),
	.w4(32'hbc07f72b),
	.w5(32'hbc2cd378),
	.w6(32'hbc72858b),
	.w7(32'hbb906284),
	.w8(32'hbb35b9e3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b1a84),
	.w1(32'hbc5c5dd0),
	.w2(32'h3bf9eb95),
	.w3(32'hbcd88b9c),
	.w4(32'hbcda45db),
	.w5(32'h3c8b50bd),
	.w6(32'hbc5d3a1b),
	.w7(32'hbc6a23d8),
	.w8(32'h3c91e2b2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8d708),
	.w1(32'h3cdda059),
	.w2(32'hbc31c65b),
	.w3(32'h3d09e681),
	.w4(32'h3ce112ae),
	.w5(32'hbcb6b033),
	.w6(32'h3c0a1047),
	.w7(32'hbc4637ed),
	.w8(32'hbc21819a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5122e2),
	.w1(32'hbc0a6ea5),
	.w2(32'hba9f391a),
	.w3(32'hbd03e2bc),
	.w4(32'hbcd17373),
	.w5(32'h3c1db1ca),
	.w6(32'hbcc34769),
	.w7(32'hbcb35e63),
	.w8(32'h3bc16af9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe4c58),
	.w1(32'h3c031dec),
	.w2(32'hba611d39),
	.w3(32'h390c7c25),
	.w4(32'hba5c7aa7),
	.w5(32'hbbe60906),
	.w6(32'h393c3c68),
	.w7(32'hbbe9d663),
	.w8(32'hbc02b71d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f53f7),
	.w1(32'hbb0b1f84),
	.w2(32'hbc2bb96d),
	.w3(32'hbbce0bf8),
	.w4(32'h3ab51165),
	.w5(32'hbc051375),
	.w6(32'hbbf00d7c),
	.w7(32'hba4eba0e),
	.w8(32'hbbc68d8c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b658),
	.w1(32'h3abef04e),
	.w2(32'hb907feca),
	.w3(32'h3ab589d6),
	.w4(32'h3a594976),
	.w5(32'hbb24cb81),
	.w6(32'h3b2e8538),
	.w7(32'h3b61b3df),
	.w8(32'hbac4241b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b28a3),
	.w1(32'h3a1f80b1),
	.w2(32'hbbc7461e),
	.w3(32'hbb33096d),
	.w4(32'hbaa5f8e1),
	.w5(32'hbc05eb00),
	.w6(32'hbb828d0d),
	.w7(32'hbb0fb3db),
	.w8(32'hbb281e44),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffc7e7),
	.w1(32'hbb177d76),
	.w2(32'hbc9f2aca),
	.w3(32'hbbb43610),
	.w4(32'hbae5f395),
	.w5(32'hbc8e7e08),
	.w6(32'hbb8b5520),
	.w7(32'hbb41e3ad),
	.w8(32'hbc657d21),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc959b79),
	.w1(32'hbb7fc972),
	.w2(32'hbb9a7b83),
	.w3(32'hbcdd182f),
	.w4(32'hbc7ae442),
	.w5(32'hbca694a2),
	.w6(32'hbc561cf8),
	.w7(32'hbc7793ce),
	.w8(32'hbc8d338b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60d82f),
	.w1(32'hbc0a4b69),
	.w2(32'h3ad5a8e4),
	.w3(32'hbd13b95c),
	.w4(32'hbccbce3f),
	.w5(32'hbb203080),
	.w6(32'hbd0d50b0),
	.w7(32'hbca48fcd),
	.w8(32'hbb840f30),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93045e),
	.w1(32'h3c7544e2),
	.w2(32'h3c506e75),
	.w3(32'hbca79ce4),
	.w4(32'hbb26f395),
	.w5(32'h3c28237e),
	.w6(32'hbcaa1495),
	.w7(32'hbc86e250),
	.w8(32'h3bbcf11d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b240f),
	.w1(32'h3b138f16),
	.w2(32'hbad3cadf),
	.w3(32'h3afc0db4),
	.w4(32'h3c067c25),
	.w5(32'hbbc34ffd),
	.w6(32'hbc1056b9),
	.w7(32'h3b34fec7),
	.w8(32'hbbbdec52),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc148efb),
	.w1(32'h3bd86e9a),
	.w2(32'h3c2189f0),
	.w3(32'h3aa8b56d),
	.w4(32'h3c4061b0),
	.w5(32'h3c72de39),
	.w6(32'h3b0fe97f),
	.w7(32'h3c331c78),
	.w8(32'h3c5b2cef),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule