module layer_10_featuremap_58(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee9ee6),
	.w1(32'h3a5e0cdb),
	.w2(32'h3c961921),
	.w3(32'h3bbf0970),
	.w4(32'h3b905725),
	.w5(32'h3d0b5cd3),
	.w6(32'h3bd0cbcd),
	.w7(32'h3b948d91),
	.w8(32'h3cf3467f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fcd22),
	.w1(32'hbc419311),
	.w2(32'hbc06d403),
	.w3(32'h3beed5a2),
	.w4(32'hbba76e2b),
	.w5(32'hbc187b29),
	.w6(32'h3bd00921),
	.w7(32'hbaf6db86),
	.w8(32'hbc1979a2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd55b6),
	.w1(32'hbb30f39e),
	.w2(32'hbc37e325),
	.w3(32'h3b5d581b),
	.w4(32'hb93eb8c7),
	.w5(32'hbcaa9bf2),
	.w6(32'h38d25c68),
	.w7(32'hbb172504),
	.w8(32'hbc826d9c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69f127),
	.w1(32'hbbf65403),
	.w2(32'h3b225737),
	.w3(32'hbcd403d0),
	.w4(32'hbc97b5c3),
	.w5(32'hbb6e53e7),
	.w6(32'hbc965479),
	.w7(32'hbc1577e4),
	.w8(32'h3bd2aedc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e4c7),
	.w1(32'hbc0fee8f),
	.w2(32'h3bf7552f),
	.w3(32'hbbae93a9),
	.w4(32'hbc523f97),
	.w5(32'h3b6990cf),
	.w6(32'hbba888a5),
	.w7(32'hbc46c2a9),
	.w8(32'hbb4c65a4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d754),
	.w1(32'h3c181f05),
	.w2(32'h3a395fa9),
	.w3(32'h3aab08a3),
	.w4(32'h3bc35197),
	.w5(32'h3ad4cb30),
	.w6(32'hbb5aa3ba),
	.w7(32'hbaebae7f),
	.w8(32'h3afa2fc5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43aa1),
	.w1(32'hbb3198c8),
	.w2(32'h3a8e63c5),
	.w3(32'h3b426873),
	.w4(32'h3b1e6b93),
	.w5(32'hb71b03d6),
	.w6(32'h3b3a3471),
	.w7(32'h39dda0a9),
	.w8(32'hba90b144),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fd9b3),
	.w1(32'hba88080d),
	.w2(32'h3aa3012a),
	.w3(32'h3ba9a186),
	.w4(32'h3ab48d91),
	.w5(32'hba7cfb83),
	.w6(32'hba7a5b38),
	.w7(32'hbbb9a5b1),
	.w8(32'hbb4ec99f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2de7be),
	.w1(32'hbb2e8ac2),
	.w2(32'h3bc1ccd6),
	.w3(32'hb9f355bf),
	.w4(32'hbc02ff3a),
	.w5(32'h3bd029f0),
	.w6(32'hba118baf),
	.w7(32'hbb8fd8c9),
	.w8(32'h3c05be7b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf19876),
	.w1(32'h3bb2e4e0),
	.w2(32'hb9599536),
	.w3(32'h3ba35ce3),
	.w4(32'h3856c441),
	.w5(32'hbac39242),
	.w6(32'hbab09441),
	.w7(32'hba900c48),
	.w8(32'hb9d3b39f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55db5e),
	.w1(32'hba9555f7),
	.w2(32'hbbfc89b9),
	.w3(32'hbacdcb0c),
	.w4(32'hbb3f279e),
	.w5(32'hbc7a3189),
	.w6(32'hbab5f723),
	.w7(32'hbb40799f),
	.w8(32'hbc7b7290),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f64c),
	.w1(32'hbbc17742),
	.w2(32'h3a44d781),
	.w3(32'hbca2ce80),
	.w4(32'hbb97a203),
	.w5(32'h3b72dfa6),
	.w6(32'hbc786baa),
	.w7(32'hbc1368cf),
	.w8(32'h3ad63045),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f8abf),
	.w1(32'h3a881a0f),
	.w2(32'h3b790d65),
	.w3(32'h3b92f8fc),
	.w4(32'h3b7f0652),
	.w5(32'h3b1832e4),
	.w6(32'h3b5a9148),
	.w7(32'h3b905880),
	.w8(32'h39fee66c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f8895),
	.w1(32'hbc0d6055),
	.w2(32'hbb2f5c9a),
	.w3(32'h3cda031d),
	.w4(32'hbc0ba44d),
	.w5(32'hbbaf1989),
	.w6(32'h3cc82ee6),
	.w7(32'hbc3e8998),
	.w8(32'hb80ceaa6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02137b),
	.w1(32'hbaffd4f1),
	.w2(32'h3a523121),
	.w3(32'h3b670ae6),
	.w4(32'hbbe1d297),
	.w5(32'h3ab9ed58),
	.w6(32'hbba20311),
	.w7(32'hbbc1fa56),
	.w8(32'hbb02584a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c4799),
	.w1(32'hbb9469aa),
	.w2(32'hb8ba23da),
	.w3(32'h3b42e1b1),
	.w4(32'hb9c31633),
	.w5(32'hb92a3a1a),
	.w6(32'hb9eacaa6),
	.w7(32'hbbc3e84a),
	.w8(32'h384c64b5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf9cc7),
	.w1(32'hba31bed9),
	.w2(32'hbb1351b4),
	.w3(32'h3a60bb8c),
	.w4(32'hba93a1d1),
	.w5(32'hbbb03913),
	.w6(32'hb8776a68),
	.w7(32'hbaa9e0ee),
	.w8(32'hbafa38f9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b178),
	.w1(32'hbb7467dc),
	.w2(32'hbb0e75ad),
	.w3(32'hbb96a3ec),
	.w4(32'hbb9ffd78),
	.w5(32'hba7868c2),
	.w6(32'h3a518874),
	.w7(32'h392bf826),
	.w8(32'hba70f832),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46e6de),
	.w1(32'hbbb22697),
	.w2(32'hbbf184c5),
	.w3(32'h3c1f5b63),
	.w4(32'hbbfb25fe),
	.w5(32'hbb046362),
	.w6(32'h3bccedfc),
	.w7(32'hbb3066c4),
	.w8(32'hbc0a6d75),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fdddd),
	.w1(32'hbbef4040),
	.w2(32'hb84af8c8),
	.w3(32'hbbd67464),
	.w4(32'hbb380a7b),
	.w5(32'hbaf83d2e),
	.w6(32'hbc7f57b5),
	.w7(32'hbc207abb),
	.w8(32'hbb167ea3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad860f3),
	.w1(32'hbab4fd3d),
	.w2(32'hbc16794e),
	.w3(32'hbb45d2b5),
	.w4(32'hbaf1db2e),
	.w5(32'hbc9642b9),
	.w6(32'hbb70a26f),
	.w7(32'hbae9c290),
	.w8(32'hbc3e6173),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bfdbd),
	.w1(32'hbb46d985),
	.w2(32'hbb8cdb5c),
	.w3(32'hbcdd6f19),
	.w4(32'hbc23b592),
	.w5(32'hbbeed947),
	.w6(32'hbc6d2f07),
	.w7(32'hba37d49e),
	.w8(32'hbc0a5887),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28171),
	.w1(32'hbb0abdfb),
	.w2(32'h3a7451e3),
	.w3(32'h39c691ca),
	.w4(32'h3b5cf39d),
	.w5(32'h3a7cf3d4),
	.w6(32'hbb6c7aaa),
	.w7(32'h3a8a66d9),
	.w8(32'h3a85cb98),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91ab42),
	.w1(32'h3a8e9371),
	.w2(32'h3b9e9bb3),
	.w3(32'hb9c4cea5),
	.w4(32'h3a94df8a),
	.w5(32'h3c1dd40e),
	.w6(32'hba4bddef),
	.w7(32'h3a21aa4a),
	.w8(32'h3b83e771),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca84771),
	.w1(32'hbc01c1dd),
	.w2(32'hba636783),
	.w3(32'h3cc516c0),
	.w4(32'hbb578412),
	.w5(32'h3c0a3052),
	.w6(32'h3c7760c6),
	.w7(32'hbbc02247),
	.w8(32'h3c1d3d44),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be9a8),
	.w1(32'hbc132a3d),
	.w2(32'h3b991f75),
	.w3(32'h3b097964),
	.w4(32'hb9443192),
	.w5(32'h3bea4b97),
	.w6(32'hbb8fc3e2),
	.w7(32'hbbff44db),
	.w8(32'h3bd24c5d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c534f37),
	.w1(32'h3b27360d),
	.w2(32'hb99f0138),
	.w3(32'h3c57f9d1),
	.w4(32'h3b8ef9cb),
	.w5(32'hb7dd49b3),
	.w6(32'h3c60dc16),
	.w7(32'h3beac73c),
	.w8(32'hba2a5cc7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f541e),
	.w1(32'hb98acca5),
	.w2(32'h3a891e55),
	.w3(32'h3a55e216),
	.w4(32'hb8eac37a),
	.w5(32'h3a8adbbe),
	.w6(32'h39bdb814),
	.w7(32'hb9ef2984),
	.w8(32'hb91f6605),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a224d),
	.w1(32'hbb93723a),
	.w2(32'hbb757248),
	.w3(32'h39256b57),
	.w4(32'hbba13cb3),
	.w5(32'hbbcb2d42),
	.w6(32'h3b4abd98),
	.w7(32'hbadf8d32),
	.w8(32'hbc1a2eb1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806ba4),
	.w1(32'h3ba3ca1b),
	.w2(32'h3b132896),
	.w3(32'hbb95dbb4),
	.w4(32'h3b6b82b4),
	.w5(32'h3b0a2080),
	.w6(32'hbc2cf0e5),
	.w7(32'hbb96fbf7),
	.w8(32'h3aec28f8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50268c),
	.w1(32'h3b18917b),
	.w2(32'h394be9f3),
	.w3(32'h3b5c6989),
	.w4(32'h3b33b6e4),
	.w5(32'hbbb5c9e7),
	.w6(32'h3b231f79),
	.w7(32'h3ad0aea6),
	.w8(32'hbb307dab),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8852c3),
	.w1(32'hbae3e3c1),
	.w2(32'h3a47ba87),
	.w3(32'hbbd3e923),
	.w4(32'hb837a05c),
	.w5(32'hbb7265b3),
	.w6(32'hbb9e438f),
	.w7(32'hbb0d4ca2),
	.w8(32'hbb96f7cd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227d9c),
	.w1(32'h3aadde2a),
	.w2(32'hbb6f4c56),
	.w3(32'hbaee7274),
	.w4(32'hbb32ee8a),
	.w5(32'hbadb6d23),
	.w6(32'hbaf06ef9),
	.w7(32'hb6964de6),
	.w8(32'hbabce736),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3cd99),
	.w1(32'hbaa789dc),
	.w2(32'h3ba92e74),
	.w3(32'h39c3968c),
	.w4(32'hbad19205),
	.w5(32'h3b976a82),
	.w6(32'hb7cda9be),
	.w7(32'hbb0cc8e5),
	.w8(32'h3bfbab10),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86cb7a),
	.w1(32'h3af78bc8),
	.w2(32'hba0460f3),
	.w3(32'h3bca3179),
	.w4(32'h3b780ebc),
	.w5(32'hb8cfbeab),
	.w6(32'h3b9d2894),
	.w7(32'h3ad4f09a),
	.w8(32'hb9c7cada),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba253a59),
	.w1(32'hb9bfc77d),
	.w2(32'hb9c97d1a),
	.w3(32'hba0e3591),
	.w4(32'hbafefeda),
	.w5(32'hbb6eb8ed),
	.w6(32'hb9ef160f),
	.w7(32'hbaa36e31),
	.w8(32'hbb923258),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3cc88),
	.w1(32'h3982c7f0),
	.w2(32'hbc0a4183),
	.w3(32'hbb15e6bb),
	.w4(32'hb9b0692e),
	.w5(32'hbbb2a615),
	.w6(32'h3a599b71),
	.w7(32'h3b114013),
	.w8(32'hbb91205e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf84bf1),
	.w1(32'hbc0728c8),
	.w2(32'hbb6a18f0),
	.w3(32'hbba38cd8),
	.w4(32'hbbf73ec8),
	.w5(32'hbb12d4c2),
	.w6(32'hbb6ca0a0),
	.w7(32'hbbde3384),
	.w8(32'h3b88f06f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae91b3e),
	.w1(32'h3a0288d6),
	.w2(32'h3b689ced),
	.w3(32'hb9962214),
	.w4(32'hba5368d1),
	.w5(32'hba1ad41f),
	.w6(32'hbaf70a41),
	.w7(32'h3b43f254),
	.w8(32'hbab83f92),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb222c2),
	.w1(32'h3b5f88a7),
	.w2(32'h3b3d35c0),
	.w3(32'h397324bc),
	.w4(32'hba4ad220),
	.w5(32'h3a8eef0f),
	.w6(32'h3be80a0a),
	.w7(32'h3b456256),
	.w8(32'h3960d619),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84fe57),
	.w1(32'h3c056fb7),
	.w2(32'hbad652fd),
	.w3(32'h3ba27b12),
	.w4(32'h3bd9713c),
	.w5(32'h37e48fb6),
	.w6(32'h3b2ee02b),
	.w7(32'h3b9d8e33),
	.w8(32'h3b6a5f94),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d9343),
	.w1(32'hbae4eed7),
	.w2(32'hbbea989e),
	.w3(32'h393d449b),
	.w4(32'hbb28d35b),
	.w5(32'hbc2ac3e3),
	.w6(32'hbaa5dc08),
	.w7(32'hbb67da51),
	.w8(32'hbc061079),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfc0c7),
	.w1(32'h3a57d71b),
	.w2(32'h39e4e8eb),
	.w3(32'hbc5ad1fd),
	.w4(32'hbbd418b9),
	.w5(32'h3a30ddb6),
	.w6(32'hbc40b4ea),
	.w7(32'hbbc591e5),
	.w8(32'h3a19953d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82ab73),
	.w1(32'hb9bdbda1),
	.w2(32'hbc0f5f3c),
	.w3(32'hba9e98fb),
	.w4(32'hb9b56718),
	.w5(32'hbc000dc6),
	.w6(32'hb9ba9e48),
	.w7(32'h3aad199a),
	.w8(32'hbbe8784a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4e64f),
	.w1(32'hbafde416),
	.w2(32'hbbdd84bd),
	.w3(32'hbbded999),
	.w4(32'hbbac9051),
	.w5(32'hbbaf7a09),
	.w6(32'hbc0a4597),
	.w7(32'hbc13ba5d),
	.w8(32'hbb9c0974),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2aad9),
	.w1(32'h3b42a2b4),
	.w2(32'hb9dda264),
	.w3(32'h392e821e),
	.w4(32'h3b014484),
	.w5(32'hba238c33),
	.w6(32'hbb6ad3c1),
	.w7(32'h3ba29a5a),
	.w8(32'hbb5432fb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b0c3),
	.w1(32'hbb6f4f19),
	.w2(32'hba9c0ac5),
	.w3(32'hbbfa186d),
	.w4(32'hbb59187b),
	.w5(32'hba3fffc7),
	.w6(32'hbbc58449),
	.w7(32'hba01509d),
	.w8(32'h3bcaa587),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe495d2),
	.w1(32'hbbdbe96c),
	.w2(32'h3a8bc47a),
	.w3(32'hbb70b381),
	.w4(32'hbb8cdca3),
	.w5(32'h38dbaad6),
	.w6(32'hbb3ee374),
	.w7(32'hbac798b8),
	.w8(32'hb9d49b78),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc7184),
	.w1(32'hba6a2549),
	.w2(32'h3a3b1cec),
	.w3(32'hbafda07b),
	.w4(32'hba6ba7da),
	.w5(32'h3bcd0fb5),
	.w6(32'hbaf2ca86),
	.w7(32'hb914a340),
	.w8(32'h3ba2dd9c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba438e2),
	.w1(32'hba4031a9),
	.w2(32'hbbf25245),
	.w3(32'h3a79ffaa),
	.w4(32'hbaf1adee),
	.w5(32'h39b77e8a),
	.w6(32'h3a5c74d3),
	.w7(32'h3b6064c9),
	.w8(32'hbb8cfd2a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb36dd8),
	.w1(32'hbbbce51f),
	.w2(32'h3b881a36),
	.w3(32'hba1ee90e),
	.w4(32'hbb223edc),
	.w5(32'hbb2c8fa0),
	.w6(32'hbb95b492),
	.w7(32'hbae8a624),
	.w8(32'hbb64bb26),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b883ab),
	.w1(32'h3b2eb6f1),
	.w2(32'hbb513385),
	.w3(32'h3b80d359),
	.w4(32'h3be3a5d8),
	.w5(32'hbbb8edf1),
	.w6(32'h39a6e90b),
	.w7(32'h3bb9d45c),
	.w8(32'hbaab28c2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe83df),
	.w1(32'hbb55a911),
	.w2(32'h38dd227d),
	.w3(32'h39f6904c),
	.w4(32'h3b29dbf1),
	.w5(32'hb9d61e70),
	.w6(32'hbb072cba),
	.w7(32'h3b8abe59),
	.w8(32'hb9957e5d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eb00d),
	.w1(32'hb99053c8),
	.w2(32'h3aa0dac5),
	.w3(32'h3b061d42),
	.w4(32'h3b468f3f),
	.w5(32'hbbc22331),
	.w6(32'hb9b72575),
	.w7(32'hbb1cad9d),
	.w8(32'hbb885628),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0c83),
	.w1(32'hba608763),
	.w2(32'h3bbb0b2f),
	.w3(32'hbb1de2dd),
	.w4(32'h3a627da5),
	.w5(32'h3a9fb378),
	.w6(32'hbbf7b71f),
	.w7(32'hbbc93ee9),
	.w8(32'h3b0dacd5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c228694),
	.w1(32'h3c07a029),
	.w2(32'h3b43d175),
	.w3(32'h3b30a97b),
	.w4(32'h3ae65311),
	.w5(32'h3a73c803),
	.w6(32'h3c1a9a1d),
	.w7(32'h3bb78b32),
	.w8(32'h3adb5669),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafbe08),
	.w1(32'hbb856b0f),
	.w2(32'h3b9e00b2),
	.w3(32'hbb3e2e3c),
	.w4(32'hbb56af65),
	.w5(32'h3acd4c00),
	.w6(32'hbb4404e2),
	.w7(32'hbae9bce8),
	.w8(32'h3a11e16c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c4808),
	.w1(32'h3913d9cc),
	.w2(32'hb97b4b5e),
	.w3(32'hba08e4c3),
	.w4(32'hbb22eae9),
	.w5(32'hb9493ced),
	.w6(32'hbb5adf20),
	.w7(32'hbb5641fe),
	.w8(32'hbaa3c06e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3be29b),
	.w1(32'hb8e8cf42),
	.w2(32'h3a0611d0),
	.w3(32'hb99066ac),
	.w4(32'hbaf98da1),
	.w5(32'hbb7c812d),
	.w6(32'hba8507a6),
	.w7(32'hbb1c9ad1),
	.w8(32'hba9ad450),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b899a),
	.w1(32'hba5ec1b3),
	.w2(32'h3b073d50),
	.w3(32'hbb6bac25),
	.w4(32'hbab316b0),
	.w5(32'h3bae00c9),
	.w6(32'hbb5c9f27),
	.w7(32'hbb4313c1),
	.w8(32'h3b2e336e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96ea79),
	.w1(32'h3bab9539),
	.w2(32'hbb22c99f),
	.w3(32'h3b61319d),
	.w4(32'h3b60df76),
	.w5(32'hbb8bc08a),
	.w6(32'hbae9a99b),
	.w7(32'h3a8b7ac6),
	.w8(32'hbbcaf4c7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab51dd7),
	.w1(32'h3b95802d),
	.w2(32'hbb8edaef),
	.w3(32'hbb0303c8),
	.w4(32'h3b790c4d),
	.w5(32'hbbda5a20),
	.w6(32'h3a7a0289),
	.w7(32'h3c14d189),
	.w8(32'hb94a7117),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fabb4),
	.w1(32'hbb04df60),
	.w2(32'hb7dcf3b8),
	.w3(32'hbbb81e81),
	.w4(32'hbbada518),
	.w5(32'h399cc60b),
	.w6(32'h3a882c8f),
	.w7(32'hba7fbe11),
	.w8(32'h3abe64e4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a8648),
	.w1(32'h3abf1dc6),
	.w2(32'h3b5e8d25),
	.w3(32'hb92d4ef9),
	.w4(32'h3af5933e),
	.w5(32'h3b02e38e),
	.w6(32'h3a9a96f5),
	.w7(32'h3aafca44),
	.w8(32'h3bacb2ca),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2afcc4),
	.w1(32'h3a1d3d04),
	.w2(32'h3a17c8f0),
	.w3(32'h3b7e9d30),
	.w4(32'hba8d7fd2),
	.w5(32'h3a895d7e),
	.w6(32'h3b31b1ab),
	.w7(32'h3addb61f),
	.w8(32'h399ef470),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba563505),
	.w1(32'hbb0a0c91),
	.w2(32'h39622527),
	.w3(32'h3b042dbf),
	.w4(32'h393c84ea),
	.w5(32'h39ac12c5),
	.w6(32'h3a7a6359),
	.w7(32'hba8416ba),
	.w8(32'h3a0b5434),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75487a),
	.w1(32'h3ab5aafd),
	.w2(32'hba74cf19),
	.w3(32'h3a6a2f31),
	.w4(32'h39cf5591),
	.w5(32'h3aba7531),
	.w6(32'h3a53c690),
	.w7(32'h3a7dff53),
	.w8(32'hbaa28e26),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad106ad),
	.w1(32'h3b3d0770),
	.w2(32'hba14ad46),
	.w3(32'h3b2b79e9),
	.w4(32'h3b1135f7),
	.w5(32'hba852b4c),
	.w6(32'hb896a0fc),
	.w7(32'h3b501e5e),
	.w8(32'hba8651c0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b372548),
	.w1(32'h38cb237a),
	.w2(32'hb9c3a8c1),
	.w3(32'h3ae147df),
	.w4(32'hb968e3ca),
	.w5(32'hba56ae0f),
	.w6(32'h3b61e733),
	.w7(32'hbab078f0),
	.w8(32'hba7038f5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01d755),
	.w1(32'hba10eade),
	.w2(32'hbac16516),
	.w3(32'hbadd3bb2),
	.w4(32'hba316f73),
	.w5(32'hbb4312c6),
	.w6(32'hba9eee01),
	.w7(32'hb9c717f6),
	.w8(32'hba3352fb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02815e),
	.w1(32'h3b43286d),
	.w2(32'h3aa330a6),
	.w3(32'hba9c5cf1),
	.w4(32'h3b3f17ac),
	.w5(32'hbb3ad8e1),
	.w6(32'h3aba4b49),
	.w7(32'h3b578299),
	.w8(32'hbb763ce5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c040f),
	.w1(32'hba9900e0),
	.w2(32'h3b6ab527),
	.w3(32'hba3448a7),
	.w4(32'h3989a955),
	.w5(32'h3ae4fb70),
	.w6(32'hbabb9247),
	.w7(32'hb9ac433e),
	.w8(32'hbb1b35de),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf39f07),
	.w1(32'h3b4e0d47),
	.w2(32'hbc262276),
	.w3(32'hbb59fbb9),
	.w4(32'hbb283d46),
	.w5(32'hbc5a77e9),
	.w6(32'hbbd42577),
	.w7(32'hbad01d3c),
	.w8(32'hbbb4fc82),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb5b9f),
	.w1(32'hbb2a58ab),
	.w2(32'h3af4da24),
	.w3(32'hbc076630),
	.w4(32'h3a8e4eaa),
	.w5(32'h3af04f47),
	.w6(32'hbb4d954b),
	.w7(32'h3b3b2d8b),
	.w8(32'h3b0571b8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b5c1b5),
	.w1(32'h39e5090b),
	.w2(32'h3aa8b0fa),
	.w3(32'h3a13452d),
	.w4(32'h3ae31ccb),
	.w5(32'h3af35868),
	.w6(32'h3a9967df),
	.w7(32'h3acacfd4),
	.w8(32'h3aa92133),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b189c72),
	.w1(32'h3adffe79),
	.w2(32'h3afb7a81),
	.w3(32'h3ab939e5),
	.w4(32'h3a13a9e8),
	.w5(32'hb9efef6c),
	.w6(32'hb99cf113),
	.w7(32'h3aafbe84),
	.w8(32'hba3273d8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e9383),
	.w1(32'hbb5b6f6a),
	.w2(32'h3b54eff9),
	.w3(32'h3ae9f6d9),
	.w4(32'h3af2579e),
	.w5(32'h3a441c8c),
	.w6(32'hba890202),
	.w7(32'h3ac40d32),
	.w8(32'h3b02e27d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab51402),
	.w1(32'hbbabf179),
	.w2(32'h3bdc1dcc),
	.w3(32'hba9cd801),
	.w4(32'hba913bf3),
	.w5(32'h39a289f6),
	.w6(32'hbb90b58b),
	.w7(32'hbb9507f0),
	.w8(32'h3b14420f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92aaf9f),
	.w1(32'hba63cf7d),
	.w2(32'hb804dfdc),
	.w3(32'hbb84b577),
	.w4(32'hbb7b205c),
	.w5(32'h3a785ac3),
	.w6(32'hba04c349),
	.w7(32'hbac31ab5),
	.w8(32'h399b3bba),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c77e3),
	.w1(32'h3a675d72),
	.w2(32'h3a981fcf),
	.w3(32'h3979e6ed),
	.w4(32'h3a7a086a),
	.w5(32'h3ad7f6ce),
	.w6(32'h39613c77),
	.w7(32'h3a54cb48),
	.w8(32'h3a4af4f1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b6fd5),
	.w1(32'hba851911),
	.w2(32'hbb3dec45),
	.w3(32'hb93a11dd),
	.w4(32'h3ad5fdca),
	.w5(32'hbb208f36),
	.w6(32'hba2c9073),
	.w7(32'h3a1a3b01),
	.w8(32'hbb3fcf7b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae897d9),
	.w1(32'hbb0f8c85),
	.w2(32'h3b353748),
	.w3(32'hba486d24),
	.w4(32'hbaf38499),
	.w5(32'h3abd949a),
	.w6(32'hbab9223f),
	.w7(32'hbb2f2526),
	.w8(32'hbad922ea),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf45a8),
	.w1(32'hbb0816be),
	.w2(32'hbc215027),
	.w3(32'h39162438),
	.w4(32'hbb19a20b),
	.w5(32'hbc39b621),
	.w6(32'hbb4d0a51),
	.w7(32'h3b04f6ee),
	.w8(32'hbc2cb43b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862ce8),
	.w1(32'hb9a9fb8a),
	.w2(32'h3aed60be),
	.w3(32'hbbba44a7),
	.w4(32'hbb7169d5),
	.w5(32'hbb3a4478),
	.w6(32'hbb96c43d),
	.w7(32'h3b44bac3),
	.w8(32'h3aa2dc27),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d8a99),
	.w1(32'h3aac5971),
	.w2(32'h3b695364),
	.w3(32'hbc049a9d),
	.w4(32'hbb5a223c),
	.w5(32'h3bd40fd6),
	.w6(32'hbae2a5bc),
	.w7(32'hbac682b4),
	.w8(32'h3b0cfcd2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ea852),
	.w1(32'h3b821f97),
	.w2(32'h3b1dc1c5),
	.w3(32'h3b1e8ffe),
	.w4(32'h3bcbd343),
	.w5(32'h3aa2be84),
	.w6(32'h39904913),
	.w7(32'h3b803273),
	.w8(32'h3a3325ff),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22197b),
	.w1(32'h3a82ccde),
	.w2(32'h3b22008a),
	.w3(32'hbaae40b9),
	.w4(32'h3b37c613),
	.w5(32'h3afc7037),
	.w6(32'hb9fac541),
	.w7(32'h3b7b6702),
	.w8(32'h3afd5d38),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cc0df),
	.w1(32'h3b95548c),
	.w2(32'hba9a2242),
	.w3(32'h3b4b5d1c),
	.w4(32'h3b45c0bc),
	.w5(32'h38d3d744),
	.w6(32'h3b06fd3d),
	.w7(32'h3b687497),
	.w8(32'h39c93490),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67229),
	.w1(32'hba0a9f9a),
	.w2(32'h3900127c),
	.w3(32'hbbb8a900),
	.w4(32'h3ac006e2),
	.w5(32'h39da1f73),
	.w6(32'hbb803d8c),
	.w7(32'h38a30757),
	.w8(32'hb9f0dc17),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e89cc),
	.w1(32'h394752ef),
	.w2(32'h3afe1509),
	.w3(32'h3ab2cfcd),
	.w4(32'h3b64039b),
	.w5(32'h3c0c6e21),
	.w6(32'hba1b4a95),
	.w7(32'hbb671f1c),
	.w8(32'h3bafb742),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b492e0a),
	.w1(32'hbaf2620f),
	.w2(32'h3a86bf2e),
	.w3(32'h3c0c5de3),
	.w4(32'h3ae9d9ae),
	.w5(32'h3a1f000a),
	.w6(32'h3bd5c1d8),
	.w7(32'hbae4c90a),
	.w8(32'h3aa00491),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae29651),
	.w1(32'h3b1bf93f),
	.w2(32'h3ac2cad7),
	.w3(32'h3b3b8f6e),
	.w4(32'hba807be9),
	.w5(32'h3a96b23d),
	.w6(32'h3b905084),
	.w7(32'hbafff48b),
	.w8(32'h3a87015d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91c9dd),
	.w1(32'h3b69ba3e),
	.w2(32'h3ba90d01),
	.w3(32'h3b752f9c),
	.w4(32'h3b59e232),
	.w5(32'h3b5de24a),
	.w6(32'h3b84b2ef),
	.w7(32'h3b9414e8),
	.w8(32'h3b4fbf2f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b859eeb),
	.w1(32'h3b6194f9),
	.w2(32'h3a815341),
	.w3(32'h3b4cddff),
	.w4(32'h3b21ca50),
	.w5(32'h39e59b32),
	.w6(32'h3b39fe8c),
	.w7(32'h3b4af598),
	.w8(32'h3ba50777),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f108),
	.w1(32'hbae846bb),
	.w2(32'hbae8f2b6),
	.w3(32'h3b16124b),
	.w4(32'hba611e83),
	.w5(32'h3b5a5d86),
	.w6(32'h3b1f94f4),
	.w7(32'h3a379b2d),
	.w8(32'h3b495e2a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9357d),
	.w1(32'hb97fa106),
	.w2(32'h3b47192d),
	.w3(32'h3bbbdf3c),
	.w4(32'h3af60c04),
	.w5(32'h3b9720cb),
	.w6(32'hbad1b5f9),
	.w7(32'hbbd960f8),
	.w8(32'h3b038db7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3259a1),
	.w1(32'hbae23aa1),
	.w2(32'hbabe55bd),
	.w3(32'h3b1445f5),
	.w4(32'hba93732a),
	.w5(32'hbbdd8fa9),
	.w6(32'hbaa7d65f),
	.w7(32'hba7cc02b),
	.w8(32'hba97b57f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde7325),
	.w1(32'hba6f42c5),
	.w2(32'hbb03fb41),
	.w3(32'hbc3156f5),
	.w4(32'hbbc60103),
	.w5(32'hbaf93c7d),
	.w6(32'hbb83ecd6),
	.w7(32'h3ae47c9d),
	.w8(32'h3a8e0a09),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc3c40),
	.w1(32'hbacf902b),
	.w2(32'hbb904193),
	.w3(32'hb844155e),
	.w4(32'h39ab7b17),
	.w5(32'hbada71df),
	.w6(32'h3b617065),
	.w7(32'hba3caee3),
	.w8(32'hb828c97d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0afa),
	.w1(32'h3b59c93f),
	.w2(32'hbb2cf2a1),
	.w3(32'hbb92a520),
	.w4(32'h3b1c0a8a),
	.w5(32'hbbff529b),
	.w6(32'hbb758865),
	.w7(32'h3b420f10),
	.w8(32'hbbf033a1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d6f8f),
	.w1(32'h39c2fef2),
	.w2(32'hba38510f),
	.w3(32'hbbbe445e),
	.w4(32'h3b21844c),
	.w5(32'hbb82e782),
	.w6(32'hbc2bae82),
	.w7(32'hbc080a51),
	.w8(32'hbb2b0376),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ac3c3),
	.w1(32'h3afd4f98),
	.w2(32'hba8c0780),
	.w3(32'h3b517730),
	.w4(32'h3b20aa2f),
	.w5(32'h3a3cc210),
	.w6(32'hbb212042),
	.w7(32'hbc23ad74),
	.w8(32'h39c802a5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa77a9b),
	.w1(32'hbabfbe52),
	.w2(32'hbaa28ea7),
	.w3(32'hba963b7f),
	.w4(32'h3b28637f),
	.w5(32'h3ab2add6),
	.w6(32'hba86f1b2),
	.w7(32'h3a7178be),
	.w8(32'h3a853a7b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3637d6),
	.w1(32'h3b6d1174),
	.w2(32'h3a79f3f6),
	.w3(32'h3abb4dbd),
	.w4(32'h3bc1dd2b),
	.w5(32'hba8f1109),
	.w6(32'h3a44a6d5),
	.w7(32'h3ba3c9f2),
	.w8(32'hbb1ca28d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4ab3e),
	.w1(32'h39094e56),
	.w2(32'h3b48b87c),
	.w3(32'hb9504148),
	.w4(32'hbb779f4b),
	.w5(32'h3aa3a82b),
	.w6(32'h3ae928dc),
	.w7(32'hbb59db87),
	.w8(32'hb99c4275),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9520e7),
	.w1(32'h3af1050f),
	.w2(32'h39eadeff),
	.w3(32'h3a1aec36),
	.w4(32'h3b9c249c),
	.w5(32'hba5e4b8d),
	.w6(32'h3b0d13da),
	.w7(32'h3b912204),
	.w8(32'hbae529aa),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a5f2),
	.w1(32'h3ae2862a),
	.w2(32'hbb9cfb43),
	.w3(32'hba5fe822),
	.w4(32'h3b286e60),
	.w5(32'hbbfe62d7),
	.w6(32'h39a982ee),
	.w7(32'h3b4b7688),
	.w8(32'hbba6db99),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ffd23),
	.w1(32'hbb59d8f4),
	.w2(32'hbb75625c),
	.w3(32'hbc12a0f4),
	.w4(32'hbb113f46),
	.w5(32'hbbe66202),
	.w6(32'hbbec0f4f),
	.w7(32'hba9c9c08),
	.w8(32'hbbe0f2ee),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb149032),
	.w1(32'hbad43f80),
	.w2(32'hba7935d9),
	.w3(32'hbbb90224),
	.w4(32'hbac17d3d),
	.w5(32'hbb2919fc),
	.w6(32'hbb0ec5fb),
	.w7(32'hbb3beb3d),
	.w8(32'hbac03413),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b146a87),
	.w1(32'h3b48f4ac),
	.w2(32'hbbad71db),
	.w3(32'hbb5ce8b6),
	.w4(32'h3b1d835e),
	.w5(32'hbc1566b7),
	.w6(32'hbbb9d83e),
	.w7(32'hbb04def8),
	.w8(32'hbbcf4b7e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae6f8b),
	.w1(32'h3994339a),
	.w2(32'hbab020ca),
	.w3(32'hbc4bc012),
	.w4(32'hbbdf18d0),
	.w5(32'h3a6bc470),
	.w6(32'hbbc94ae8),
	.w7(32'hb987506d),
	.w8(32'hb84a8b27),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ec764),
	.w1(32'h3adefc5b),
	.w2(32'hbabc644a),
	.w3(32'h3af4e9b2),
	.w4(32'h3bb69a37),
	.w5(32'h3b68e882),
	.w6(32'h3b9a6cbb),
	.w7(32'h3c041c0c),
	.w8(32'h3ac2aa12),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9458ff),
	.w1(32'h3b7a9b32),
	.w2(32'hbaefa880),
	.w3(32'h3b94d4eb),
	.w4(32'h3b439875),
	.w5(32'hbc46c37f),
	.w6(32'h3bf6d16a),
	.w7(32'h3bce015e),
	.w8(32'hbc1690d7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1db813),
	.w1(32'h3b8c419f),
	.w2(32'hbaa951fa),
	.w3(32'hbc0d1162),
	.w4(32'hbb1c4c7f),
	.w5(32'hbafea6e5),
	.w6(32'hbc0971f3),
	.w7(32'hb9de4df6),
	.w8(32'h3a34268a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14f41e),
	.w1(32'h37e3ebff),
	.w2(32'hbbd51a02),
	.w3(32'hb7e0a5c3),
	.w4(32'hbaa7ff11),
	.w5(32'hbba2bf5d),
	.w6(32'h3a7d307b),
	.w7(32'hba9cdebc),
	.w8(32'hbabe0901),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba779f1),
	.w1(32'hbb5505c6),
	.w2(32'h3b0801cf),
	.w3(32'hbb4c3dfa),
	.w4(32'hbaca5b6e),
	.w5(32'h3ae40ef3),
	.w6(32'hba95df45),
	.w7(32'hb9b53ba4),
	.w8(32'h396ff91c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b532fe3),
	.w1(32'h3b9fc530),
	.w2(32'hbb2c01b2),
	.w3(32'h3b8f9c5f),
	.w4(32'h3bc74e05),
	.w5(32'hbb067db3),
	.w6(32'h3afc15e8),
	.w7(32'h3b2f0303),
	.w8(32'h39f22cc1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1894),
	.w1(32'hbb572854),
	.w2(32'h39505492),
	.w3(32'hbb42effa),
	.w4(32'hbb45b3c6),
	.w5(32'hb969e1ad),
	.w6(32'hba9f2b47),
	.w7(32'hbb4bdb8a),
	.w8(32'hb9a43964),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39880b67),
	.w1(32'hbba45921),
	.w2(32'hbb43e666),
	.w3(32'hbadddd45),
	.w4(32'h3b4a33bf),
	.w5(32'hbb8bd1d1),
	.w6(32'hba01b6a7),
	.w7(32'hb973d7ee),
	.w8(32'hbb992364),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaa0d7),
	.w1(32'h3a90074c),
	.w2(32'hbb05dad0),
	.w3(32'h3a35ec27),
	.w4(32'h3b5124aa),
	.w5(32'hbad15f4a),
	.w6(32'hbb6e7a4e),
	.w7(32'hbbc17987),
	.w8(32'h3910e853),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb345c42),
	.w1(32'h3a8bac95),
	.w2(32'h3b34ee57),
	.w3(32'hbbf70146),
	.w4(32'hbbb972d2),
	.w5(32'h3b0d4aa9),
	.w6(32'hbac25d60),
	.w7(32'h3b64d506),
	.w8(32'h3b0e6e6e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52f408),
	.w1(32'h3b47308a),
	.w2(32'h3aabac69),
	.w3(32'h3b4a11e8),
	.w4(32'h3b613862),
	.w5(32'h3aae01f5),
	.w6(32'h3b3eef23),
	.w7(32'h3b566527),
	.w8(32'h3a253a63),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac17ae8),
	.w1(32'h3a8aab9b),
	.w2(32'hbb4b5f58),
	.w3(32'h3b056799),
	.w4(32'h3acc4cfc),
	.w5(32'hbb27bc8d),
	.w6(32'hb9c0e11a),
	.w7(32'hb94cc80e),
	.w8(32'h3a9a08d8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9017e1),
	.w1(32'hbb60733e),
	.w2(32'hba530673),
	.w3(32'hbaf63f15),
	.w4(32'hbaee0fc2),
	.w5(32'hbae128cb),
	.w6(32'hba7a103f),
	.w7(32'h3b87b9e3),
	.w8(32'hbaad725b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2f49),
	.w1(32'hb9dffeef),
	.w2(32'h3b0a1186),
	.w3(32'hbb5fb17c),
	.w4(32'hbabe62a5),
	.w5(32'h3b18ca9c),
	.w6(32'hbae70cd7),
	.w7(32'hba0f46e0),
	.w8(32'hbb040ab1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4f510),
	.w1(32'h3a147b4a),
	.w2(32'hbab76a19),
	.w3(32'hbaddb402),
	.w4(32'h3ac8dc97),
	.w5(32'h3b9b7d4d),
	.w6(32'hba314034),
	.w7(32'h3b6e45b1),
	.w8(32'h37f8712b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b89fe),
	.w1(32'h3bb83b4b),
	.w2(32'h3b5bfabd),
	.w3(32'hbaf24a4e),
	.w4(32'h3bb4bac9),
	.w5(32'h3b7fc6a7),
	.w6(32'hbb8b1abf),
	.w7(32'h3b8ab430),
	.w8(32'h3ae758b3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20aa05),
	.w1(32'h3b2c74b3),
	.w2(32'h3abbb977),
	.w3(32'hbb0ac7e9),
	.w4(32'h3a007385),
	.w5(32'hba43913e),
	.w6(32'hbbf3835d),
	.w7(32'hbb177272),
	.w8(32'hbbf2d56b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6d23),
	.w1(32'h3bfbd16c),
	.w2(32'h3ab1c752),
	.w3(32'hbaa0c698),
	.w4(32'h3ba44127),
	.w5(32'hba8d8e97),
	.w6(32'hbb28ae06),
	.w7(32'h3b94fae2),
	.w8(32'h3b4240bb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9f89a),
	.w1(32'hbc037ab0),
	.w2(32'h3a51d58e),
	.w3(32'hbb845f25),
	.w4(32'hbb979c10),
	.w5(32'hbb4c3889),
	.w6(32'h3b739417),
	.w7(32'h3b79e1a9),
	.w8(32'h3ac0070a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ee53a),
	.w1(32'h3b5cb872),
	.w2(32'hbbb412b3),
	.w3(32'hb9739055),
	.w4(32'hbb24b3d3),
	.w5(32'hbc2ca94a),
	.w6(32'h3bc9645c),
	.w7(32'h3b248764),
	.w8(32'hbc027a7d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2563c7),
	.w1(32'h386c0742),
	.w2(32'hba167bad),
	.w3(32'hbc333ad4),
	.w4(32'hbbad8e83),
	.w5(32'h398ecccf),
	.w6(32'hbbd6b510),
	.w7(32'hbb9501d2),
	.w8(32'hbbd087ee),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37be2a),
	.w1(32'hbbd1a9b0),
	.w2(32'hbb890e49),
	.w3(32'hbb041c2f),
	.w4(32'hbb63e77e),
	.w5(32'hbba3fa61),
	.w6(32'hbbcc3d10),
	.w7(32'hbb817112),
	.w8(32'hbbc35a3e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b0c02),
	.w1(32'h3a5acbcb),
	.w2(32'hb7fcc33f),
	.w3(32'hbb930b4b),
	.w4(32'h3ae136a0),
	.w5(32'hba937076),
	.w6(32'hbb0c4e07),
	.w7(32'h3b668d19),
	.w8(32'hba62cdfa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49c8a5),
	.w1(32'hba86d4e5),
	.w2(32'hbb8afa20),
	.w3(32'hbb19f02c),
	.w4(32'hbaefe69a),
	.w5(32'hbb80cea8),
	.w6(32'hbad5d067),
	.w7(32'hbad0d6a6),
	.w8(32'h39dca2f1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92d8eb),
	.w1(32'hbb58a8ac),
	.w2(32'hbaaccef2),
	.w3(32'hbb2a3430),
	.w4(32'hbb2682b2),
	.w5(32'hbb39ee30),
	.w6(32'hbb301b3b),
	.w7(32'hbbb7be67),
	.w8(32'hbb4980d7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7fb0f),
	.w1(32'hbb215475),
	.w2(32'hbb373c32),
	.w3(32'h370a9134),
	.w4(32'h3af0f999),
	.w5(32'h39c4cba3),
	.w6(32'hba98da12),
	.w7(32'hbaa20654),
	.w8(32'h39c93975),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab563ac),
	.w1(32'hba97e957),
	.w2(32'h3a8bc644),
	.w3(32'h3b3e2ab4),
	.w4(32'hbb35dff5),
	.w5(32'h3abaa440),
	.w6(32'h3afea741),
	.w7(32'hbb00da62),
	.w8(32'h3adfc79a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b088896),
	.w1(32'h3b1516a3),
	.w2(32'hba2da7b6),
	.w3(32'h3b3ed07c),
	.w4(32'h3ae8bbf9),
	.w5(32'hbc10559d),
	.w6(32'h3b127225),
	.w7(32'h3a5b1a84),
	.w8(32'hbbd2f257),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4faf6),
	.w1(32'h3b3fd942),
	.w2(32'h3aeb8ee1),
	.w3(32'hbc13c75a),
	.w4(32'hbb3f99ed),
	.w5(32'h39d88f9a),
	.w6(32'hbc2cebb8),
	.w7(32'hbad2b497),
	.w8(32'hb99cf497),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ec1bb),
	.w1(32'h3a966f7d),
	.w2(32'hbbde4882),
	.w3(32'h38866684),
	.w4(32'h39f891e2),
	.w5(32'hbb3688ac),
	.w6(32'h38806ac1),
	.w7(32'h3aad8c48),
	.w8(32'hbba87001),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba049ab),
	.w1(32'hbb64dca4),
	.w2(32'hbb0c07b3),
	.w3(32'hbbbc51d8),
	.w4(32'hbb0950e3),
	.w5(32'hb9a4ac39),
	.w6(32'hbb91afc4),
	.w7(32'hbb7ba38a),
	.w8(32'hbb264b0b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d36293),
	.w1(32'hba72e7b1),
	.w2(32'hbb62996b),
	.w3(32'h3ac7a96b),
	.w4(32'hbb7003fb),
	.w5(32'hbb96bb1b),
	.w6(32'hbb3fca67),
	.w7(32'hbbb6d9bc),
	.w8(32'hbae322d6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5260f5),
	.w1(32'hbb7b6aee),
	.w2(32'h3b01ba11),
	.w3(32'hbba57c5c),
	.w4(32'hbba9546e),
	.w5(32'h3ad696eb),
	.w6(32'hbb627d0b),
	.w7(32'hbbaadb57),
	.w8(32'h3ab771fe),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad5c6),
	.w1(32'h3ab6b29e),
	.w2(32'hb89fe176),
	.w3(32'h3b0af353),
	.w4(32'h3a6c5b72),
	.w5(32'h38577e60),
	.w6(32'h3ae9b01a),
	.w7(32'h3a319c7c),
	.w8(32'hba8cb228),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff17ef),
	.w1(32'hbb58f5c7),
	.w2(32'hbbdf78da),
	.w3(32'hba948ab6),
	.w4(32'hbb39ae97),
	.w5(32'hbb9a39af),
	.w6(32'hbadca3d1),
	.w7(32'hbb7e9418),
	.w8(32'hbb3ca9d0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f46a3),
	.w1(32'hbbae3994),
	.w2(32'hbab1573e),
	.w3(32'hbba598d8),
	.w4(32'hbb7eb676),
	.w5(32'hbc390365),
	.w6(32'hbb4d231b),
	.w7(32'hbb0a91d9),
	.w8(32'hbb717923),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78425a),
	.w1(32'h3b1e2c20),
	.w2(32'h3959152f),
	.w3(32'hbc25cdf6),
	.w4(32'hbb107eda),
	.w5(32'hb8fcda66),
	.w6(32'hbbca856d),
	.w7(32'hbb68965f),
	.w8(32'h39e9cd03),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98a52f),
	.w1(32'h3a6128e7),
	.w2(32'hba494af5),
	.w3(32'hbaa82bf8),
	.w4(32'h3b39e838),
	.w5(32'hbb25dd45),
	.w6(32'hba62bd56),
	.w7(32'h3ac3f4fb),
	.w8(32'hbb4da2eb),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba172c7e),
	.w1(32'hba22cf91),
	.w2(32'h3ae8fcf1),
	.w3(32'hbba24b65),
	.w4(32'hbb8f91a1),
	.w5(32'hb981f88b),
	.w6(32'hbae27b03),
	.w7(32'hbb0f4d7e),
	.w8(32'h3ab88008),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c726d3),
	.w1(32'h3b991462),
	.w2(32'h3b1698a9),
	.w3(32'h3a9814f3),
	.w4(32'h3c0f5bee),
	.w5(32'h3b07aacc),
	.w6(32'hb907cee4),
	.w7(32'h3c01b26e),
	.w8(32'h3b02f46e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ad27),
	.w1(32'h3b335c1e),
	.w2(32'hbbfadfeb),
	.w3(32'h3b7682cd),
	.w4(32'h3b805cf7),
	.w5(32'hbba23749),
	.w6(32'h3b24d010),
	.w7(32'h3b3b0fb9),
	.w8(32'hb821df38),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f614),
	.w1(32'hbbb6b56a),
	.w2(32'hbc479af7),
	.w3(32'hbb14634a),
	.w4(32'hbb608651),
	.w5(32'hbc09d6fb),
	.w6(32'hbb6b3de5),
	.w7(32'hbb0cd313),
	.w8(32'hbc105d20),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d1845),
	.w1(32'hbbe53068),
	.w2(32'hba09eb97),
	.w3(32'hbc45f6af),
	.w4(32'hbc0f369b),
	.w5(32'hba1583fd),
	.w6(32'hbc1416d0),
	.w7(32'hbbaba1b0),
	.w8(32'h3b011d86),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fd6b0),
	.w1(32'hbb343f3d),
	.w2(32'h39269fe4),
	.w3(32'h3b809cd5),
	.w4(32'hbb3cf8b1),
	.w5(32'hb84cec32),
	.w6(32'h3b3854c2),
	.w7(32'hbb9531bb),
	.w8(32'h390881a5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397345f3),
	.w1(32'h39697dba),
	.w2(32'h39e93fba),
	.w3(32'h38280255),
	.w4(32'h3911605a),
	.w5(32'hb9368f6d),
	.w6(32'h391628d2),
	.w7(32'h39afa7de),
	.w8(32'hbac0d8be),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabf220),
	.w1(32'hbad43e50),
	.w2(32'h3a2b9735),
	.w3(32'hb9c6801a),
	.w4(32'hbb8e039f),
	.w5(32'h3ad635d6),
	.w6(32'hbb0ce980),
	.w7(32'hbb9d7ecb),
	.w8(32'h3b237cba),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d0ea2),
	.w1(32'h3a7ecbc9),
	.w2(32'h38df685a),
	.w3(32'hba166ec0),
	.w4(32'hba290e0b),
	.w5(32'h3a63f646),
	.w6(32'h3834ea5f),
	.w7(32'hb9bbb426),
	.w8(32'h3a5ff92c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3be852),
	.w1(32'h3a3ef20d),
	.w2(32'h38d6f96c),
	.w3(32'h3ab551d6),
	.w4(32'h3ad94dc8),
	.w5(32'h3b62098b),
	.w6(32'h3ab6f642),
	.w7(32'h3addaae4),
	.w8(32'h3a8a2bfe),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ef306),
	.w1(32'h388f3d70),
	.w2(32'hbb5d7b84),
	.w3(32'h3b7983d4),
	.w4(32'h3b5d1add),
	.w5(32'hbabcc3b8),
	.w6(32'h3a87299c),
	.w7(32'h399b11c2),
	.w8(32'h3b752a02),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa7bc),
	.w1(32'hbb6de93f),
	.w2(32'hb9109673),
	.w3(32'hbb040db5),
	.w4(32'hbb313e2c),
	.w5(32'h3920d511),
	.w6(32'h3b602d02),
	.w7(32'h3b3b37e9),
	.w8(32'h3910c518),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a79d51),
	.w1(32'h3a1cebde),
	.w2(32'hba3bcc14),
	.w3(32'h3a1ae548),
	.w4(32'h3a5883f7),
	.w5(32'hb9e045bc),
	.w6(32'h3a200f48),
	.w7(32'h3a3cbdf9),
	.w8(32'h3a08517d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52ec57),
	.w1(32'h3a808025),
	.w2(32'h39c1f49b),
	.w3(32'h3a513b64),
	.w4(32'h3af073e7),
	.w5(32'hb984cf9f),
	.w6(32'h3ad2c60a),
	.w7(32'h3b2bafa0),
	.w8(32'h38dc77e5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3929d3b6),
	.w1(32'hb9b689e6),
	.w2(32'h3a847c9d),
	.w3(32'h37ffd7b7),
	.w4(32'hba89e0ef),
	.w5(32'hba8a220d),
	.w6(32'hb8dabd50),
	.w7(32'hba3f5662),
	.w8(32'h3a83a3ee),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb1708),
	.w1(32'hbb196a4d),
	.w2(32'h3b1e458a),
	.w3(32'hbb65a2ea),
	.w4(32'hbae1af39),
	.w5(32'h3b0cf14f),
	.w6(32'hba5ef6c8),
	.w7(32'h39b2c02b),
	.w8(32'h3abce345),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09990d),
	.w1(32'h3addfb22),
	.w2(32'h3a8e82a1),
	.w3(32'h3a94c7d0),
	.w4(32'h3a38d38a),
	.w5(32'hb96deb2c),
	.w6(32'h3a300aba),
	.w7(32'h3a2dacaf),
	.w8(32'hba4b9b4a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b4db69),
	.w1(32'hb9a66162),
	.w2(32'hb97e44ba),
	.w3(32'h39ea21f1),
	.w4(32'hbaa08bfa),
	.w5(32'hba0dfff3),
	.w6(32'hbac39936),
	.w7(32'hbb124902),
	.w8(32'h3b021023),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cc8cc),
	.w1(32'hb8032b2f),
	.w2(32'hb97b6b34),
	.w3(32'hbb42d68c),
	.w4(32'hbb0e9c57),
	.w5(32'h37c1a090),
	.w6(32'hbb12b4ce),
	.w7(32'hbaddb89f),
	.w8(32'h3aab0a46),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15bafd),
	.w1(32'h3acf27df),
	.w2(32'h3b27a171),
	.w3(32'h3a3e0e65),
	.w4(32'h3b2dab61),
	.w5(32'h3b1b7348),
	.w6(32'h3aaa993c),
	.w7(32'h3b42a1c9),
	.w8(32'h3b60c188),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47c9d),
	.w1(32'h3b04bab1),
	.w2(32'h3abee0f0),
	.w3(32'h3b259b96),
	.w4(32'h3b18d237),
	.w5(32'h3ae1170c),
	.w6(32'h3b9a9bda),
	.w7(32'h3b88d381),
	.w8(32'hba4811f4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd81a9),
	.w1(32'h3952a31d),
	.w2(32'h397fab9f),
	.w3(32'h3b1ac1d8),
	.w4(32'h3a97bd92),
	.w5(32'hba1b7d19),
	.w6(32'hba1f7d40),
	.w7(32'h38cadaf0),
	.w8(32'hba2c7bfd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ac45e),
	.w1(32'hba7e0235),
	.w2(32'hb9b02493),
	.w3(32'hbac652c8),
	.w4(32'hbae74f65),
	.w5(32'hb9b9fcc9),
	.w6(32'hbaeb3d70),
	.w7(32'hbadf8eeb),
	.w8(32'hba4a0650),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3817becf),
	.w1(32'h3b1476c8),
	.w2(32'h3a2da95a),
	.w3(32'h3ae9125e),
	.w4(32'h3ae262d8),
	.w5(32'h3a1e8986),
	.w6(32'h3a83611b),
	.w7(32'h3aa5fd0c),
	.w8(32'hb858dc9e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cefbf),
	.w1(32'h394fe210),
	.w2(32'h3aa5e07e),
	.w3(32'hbaf4a9bb),
	.w4(32'hbb0d434c),
	.w5(32'h3a3f0b79),
	.w6(32'hbb2672be),
	.w7(32'hbb1505aa),
	.w8(32'hb92d5659),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab68b4),
	.w1(32'h3a0d6365),
	.w2(32'h3a0a3e5e),
	.w3(32'h3b06eb70),
	.w4(32'h392be3f7),
	.w5(32'hba45f000),
	.w6(32'h3a96eea1),
	.w7(32'hb94fbf5f),
	.w8(32'h3a836c76),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a861d4),
	.w1(32'hb797ae9e),
	.w2(32'hb9a0d4d2),
	.w3(32'hba18eb95),
	.w4(32'hba8f8bd9),
	.w5(32'hba46fb14),
	.w6(32'h3a691477),
	.w7(32'h3a873d90),
	.w8(32'hba8cb3b6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab53209),
	.w1(32'hbad07f74),
	.w2(32'hba468b8e),
	.w3(32'hbb045148),
	.w4(32'hbb13f27f),
	.w5(32'hbabf0f9b),
	.w6(32'hbb116429),
	.w7(32'hbb19f519),
	.w8(32'h3a2c6f63),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e25210),
	.w1(32'hba4ade68),
	.w2(32'hbb4af7a2),
	.w3(32'h3a34a77b),
	.w4(32'hba124a4f),
	.w5(32'hbb349c74),
	.w6(32'h3a0b2318),
	.w7(32'hb87f3a0c),
	.w8(32'hba94682f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba811f66),
	.w1(32'hbaa4f192),
	.w2(32'h3b159cca),
	.w3(32'hb9769871),
	.w4(32'h39254cd9),
	.w5(32'h3adb6a32),
	.w6(32'h3854618a),
	.w7(32'hb986c45b),
	.w8(32'hb9e39c4f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a295cf9),
	.w1(32'h37f8e153),
	.w2(32'hba2a13f0),
	.w3(32'hbaac4cb8),
	.w4(32'h3aa17ddc),
	.w5(32'hb8b497d0),
	.w6(32'hba86d0b7),
	.w7(32'hb989ff37),
	.w8(32'hb9c1167c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3135b3),
	.w1(32'h396f6c9c),
	.w2(32'hb9d0da51),
	.w3(32'hb94b17ee),
	.w4(32'h3a9a436f),
	.w5(32'h3985d6f0),
	.w6(32'h3ac3df24),
	.w7(32'h39f8cceb),
	.w8(32'hb8daa005),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4c4b7),
	.w1(32'hb98e1506),
	.w2(32'hb809354d),
	.w3(32'hb9821d09),
	.w4(32'h3a7c8311),
	.w5(32'hbb0211d0),
	.w6(32'h3a1bd5c9),
	.w7(32'h3ad6e01a),
	.w8(32'hbade8bdc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6f180),
	.w1(32'h399b9681),
	.w2(32'hb9e0292d),
	.w3(32'hbb3a044f),
	.w4(32'hbb438eff),
	.w5(32'hbb1ff4d1),
	.w6(32'hbab95bdd),
	.w7(32'hbabca13c),
	.w8(32'hba580a6e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa5b46),
	.w1(32'hb9ce3f88),
	.w2(32'hbaa3d215),
	.w3(32'hbb24280b),
	.w4(32'hbb3dd228),
	.w5(32'h3aff9be8),
	.w6(32'hba95373b),
	.w7(32'h39e6c938),
	.w8(32'hb98fbd92),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba478d41),
	.w1(32'hbb2c923c),
	.w2(32'h3a3be418),
	.w3(32'h39f778d2),
	.w4(32'hbaf4fac4),
	.w5(32'h3953931b),
	.w6(32'h3a069a27),
	.w7(32'hbad0bb18),
	.w8(32'h3a1670a0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d5414),
	.w1(32'hbaf68fce),
	.w2(32'h39ac8171),
	.w3(32'hba64162d),
	.w4(32'hbb145eb4),
	.w5(32'hb9e99d79),
	.w6(32'hba0146b5),
	.w7(32'hbae856a8),
	.w8(32'hbafd59ee),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5b177),
	.w1(32'h3abb4c4d),
	.w2(32'h39b6017e),
	.w3(32'hbaba05aa),
	.w4(32'h3a5d906d),
	.w5(32'h3a19d530),
	.w6(32'hbb21954f),
	.w7(32'hb9333094),
	.w8(32'h3aeacd99),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dec4a),
	.w1(32'h3939fdb4),
	.w2(32'h3b24116a),
	.w3(32'hb884b7e4),
	.w4(32'h3a0c2966),
	.w5(32'hba345825),
	.w6(32'h3a5c7a8e),
	.w7(32'h3a3dc12c),
	.w8(32'h3af06d77),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a961df6),
	.w1(32'h3ac449fa),
	.w2(32'hbae30505),
	.w3(32'hbb1db6ce),
	.w4(32'hbadd8377),
	.w5(32'hbade3785),
	.w6(32'hba545527),
	.w7(32'hba505af7),
	.w8(32'hba3aae18),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc7b47),
	.w1(32'hba94b3b0),
	.w2(32'h3b388eb6),
	.w3(32'hbb09499d),
	.w4(32'hbab8f479),
	.w5(32'h3aad96af),
	.w6(32'hbb0b3d81),
	.w7(32'hba897c46),
	.w8(32'h3a287534),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3404c0),
	.w1(32'h399f2d61),
	.w2(32'hba292b54),
	.w3(32'h3b2ff07e),
	.w4(32'h3a0af22e),
	.w5(32'hba8de99c),
	.w6(32'h3afd96f7),
	.w7(32'h36e1c9c2),
	.w8(32'h3a012d4d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc6f81),
	.w1(32'hba899968),
	.w2(32'hba9b1415),
	.w3(32'hbb3dd356),
	.w4(32'hbaf32820),
	.w5(32'h3ad770ab),
	.w6(32'hb9268d16),
	.w7(32'h39813fe7),
	.w8(32'h3a555f2d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82a322),
	.w1(32'h3940ca92),
	.w2(32'hba88b4cf),
	.w3(32'h3a6586dc),
	.w4(32'h3aff4005),
	.w5(32'hba85f201),
	.w6(32'hb85d5b36),
	.w7(32'h3abdce7e),
	.w8(32'hb964588f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11e91),
	.w1(32'hbacac4f3),
	.w2(32'h3a889cec),
	.w3(32'hba9f36ad),
	.w4(32'hbb042165),
	.w5(32'hb915ff2c),
	.w6(32'hb9f3515f),
	.w7(32'hba982866),
	.w8(32'hb73281e5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2e18a),
	.w1(32'h39d6d920),
	.w2(32'hb899e858),
	.w3(32'hba929062),
	.w4(32'hba1741ab),
	.w5(32'hba2ba84a),
	.w6(32'hba89d409),
	.w7(32'hb963b43d),
	.w8(32'h38634da3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fa9ea),
	.w1(32'h3a62d4ac),
	.w2(32'hba9b093d),
	.w3(32'hba4e8f9c),
	.w4(32'h3a2cc90e),
	.w5(32'hba195993),
	.w6(32'hb9c3c6e0),
	.w7(32'h39add5d8),
	.w8(32'hba16ccea),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beb49d),
	.w1(32'hb5427094),
	.w2(32'hb9cda7c3),
	.w3(32'hb9c9dc4d),
	.w4(32'h3971ccec),
	.w5(32'hba7a3998),
	.w6(32'hba6257f9),
	.w7(32'hb9a9c4f6),
	.w8(32'hb9e5ddb4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d5e18),
	.w1(32'h399de053),
	.w2(32'h3a31188a),
	.w3(32'hba99a1b3),
	.w4(32'hb9853fa0),
	.w5(32'h39d68660),
	.w6(32'hba6d8f91),
	.w7(32'hb8dc15bc),
	.w8(32'h3ae27908),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37874775),
	.w1(32'h3b6c5dac),
	.w2(32'h38167d58),
	.w3(32'hba65dd05),
	.w4(32'h3b85d2b8),
	.w5(32'h39917abe),
	.w6(32'h3a8d3230),
	.w7(32'h3ba82fb9),
	.w8(32'hb9acaa1b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28d0b3),
	.w1(32'h3aba1945),
	.w2(32'h3975768a),
	.w3(32'h3a74245d),
	.w4(32'hb90a46e4),
	.w5(32'h388ce0ca),
	.w6(32'h39789b9b),
	.w7(32'hba0d71ea),
	.w8(32'hba803466),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a5813),
	.w1(32'h3a23cf90),
	.w2(32'hba0eb27c),
	.w3(32'hba2abc33),
	.w4(32'h395e9b73),
	.w5(32'h3b0108f1),
	.w6(32'hbabbef52),
	.w7(32'h3a07205f),
	.w8(32'h3ac392a0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb314763),
	.w1(32'hbac3ff01),
	.w2(32'h3ae8a84b),
	.w3(32'hba681de2),
	.w4(32'hb75ad2e3),
	.w5(32'h3b037b58),
	.w6(32'hbaccbd7c),
	.w7(32'hb997507e),
	.w8(32'h3af2a12a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b183540),
	.w1(32'h3a91bc4c),
	.w2(32'hb8c35b0d),
	.w3(32'h3b1e693b),
	.w4(32'h3aa60f0d),
	.w5(32'h3b126456),
	.w6(32'h3b1db718),
	.w7(32'h3a9d1ffc),
	.w8(32'h3a2c428b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae87c21),
	.w1(32'h3a75e67a),
	.w2(32'hba60f147),
	.w3(32'h3b89a5e8),
	.w4(32'h3b657ac2),
	.w5(32'h3a61fc9c),
	.w6(32'h3b6097d0),
	.w7(32'h3b1d3d62),
	.w8(32'h395621dc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7860d12),
	.w1(32'h3953e28d),
	.w2(32'hba29aa34),
	.w3(32'h39865878),
	.w4(32'h3b024255),
	.w5(32'h3aa8754d),
	.w6(32'hb9f87c8e),
	.w7(32'h39dea45d),
	.w8(32'h39fc0526),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7214a),
	.w1(32'h3aae9a70),
	.w2(32'h3b0983c7),
	.w3(32'h3a22ae40),
	.w4(32'h3b2ae1ec),
	.w5(32'h3b10d61d),
	.w6(32'h3a87ad8e),
	.w7(32'h39ddbb03),
	.w8(32'h3ae361b3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b285ed9),
	.w1(32'h3afafd3f),
	.w2(32'hb9c24a28),
	.w3(32'h3b8c7ccc),
	.w4(32'h3b76d2bd),
	.w5(32'hb9ad869c),
	.w6(32'h3b13c722),
	.w7(32'h3b1e831c),
	.w8(32'hb9d14d08),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f5cc9),
	.w1(32'hb9213239),
	.w2(32'hb9b6c222),
	.w3(32'h395d4934),
	.w4(32'h3948959e),
	.w5(32'hba7c67a2),
	.w6(32'hb6b9aac1),
	.w7(32'hb90d4dbf),
	.w8(32'hb9394eac),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e4e71),
	.w1(32'h3a69f29e),
	.w2(32'h39c3c578),
	.w3(32'hbad25230),
	.w4(32'h3aae158f),
	.w5(32'h391cd7e5),
	.w6(32'h39cc4b11),
	.w7(32'h3b10b9b2),
	.w8(32'h38e1169b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa1ec6),
	.w1(32'hb8a146cc),
	.w2(32'h3b2377cf),
	.w3(32'h39230dbc),
	.w4(32'h383402e6),
	.w5(32'h3ae3ff4d),
	.w6(32'h398bee56),
	.w7(32'h3883da9e),
	.w8(32'h3ab04f44),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5776d),
	.w1(32'h3b1e2ebd),
	.w2(32'hbb80a46f),
	.w3(32'h3a90b24b),
	.w4(32'h3aecfc21),
	.w5(32'hbbacb82f),
	.w6(32'h39839aaf),
	.w7(32'h3b0fac03),
	.w8(32'hbb9dd15e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2e2e2),
	.w1(32'hb9b3a982),
	.w2(32'h3b118fb7),
	.w3(32'hbb86e280),
	.w4(32'hbb1d2eb9),
	.w5(32'h397a738a),
	.w6(32'hbb74dba5),
	.w7(32'hbb75b128),
	.w8(32'h3a0f0b46),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8787),
	.w1(32'h3a6bbfc0),
	.w2(32'hba80c285),
	.w3(32'h3aeaacbe),
	.w4(32'h3800d3dd),
	.w5(32'hb9da9180),
	.w6(32'h3b07563e),
	.w7(32'h3a82695f),
	.w8(32'h38e11d8f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb18e2),
	.w1(32'hba67865d),
	.w2(32'hb8e388f4),
	.w3(32'h3b383abd),
	.w4(32'hba419753),
	.w5(32'h37bcd0bd),
	.w6(32'h3b337189),
	.w7(32'hb9c9960f),
	.w8(32'h386fa1ab),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f43c),
	.w1(32'h387bc691),
	.w2(32'hb9f0ecbb),
	.w3(32'hbb208379),
	.w4(32'hba21c8c3),
	.w5(32'hb8fa7ca5),
	.w6(32'hbb2687aa),
	.w7(32'hb9ebd0f6),
	.w8(32'hb9da94d7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0beca9),
	.w1(32'hba57d6e2),
	.w2(32'hbaded1d4),
	.w3(32'hb9a5d875),
	.w4(32'hb9e7d148),
	.w5(32'h39c2d6b9),
	.w6(32'hb8e17cb5),
	.w7(32'hba05949d),
	.w8(32'hb8bbb395),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4b3a6),
	.w1(32'h39d4a2f5),
	.w2(32'hb9a8dfbe),
	.w3(32'h3b1709b1),
	.w4(32'h3a72c0df),
	.w5(32'h3a7729e2),
	.w6(32'h3a98bd86),
	.w7(32'h3a8cddee),
	.w8(32'hbab019e4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f6cca),
	.w1(32'h399308bf),
	.w2(32'hbb08555d),
	.w3(32'h3ae0bd33),
	.w4(32'h3aa3dd76),
	.w5(32'hbb0e1e06),
	.w6(32'hbaa9f467),
	.w7(32'hba89838d),
	.w8(32'hbab7d2b7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74e7aa),
	.w1(32'hbb443435),
	.w2(32'h3aad73f0),
	.w3(32'hbb4f3273),
	.w4(32'hbb5860a5),
	.w5(32'hbb5b10dc),
	.w6(32'hbb075559),
	.w7(32'hbad82154),
	.w8(32'hbb07da1e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad35d67),
	.w1(32'hbae3db00),
	.w2(32'hbb529e3a),
	.w3(32'hbbd6ed0f),
	.w4(32'hbbd4f04f),
	.w5(32'hbb7970d6),
	.w6(32'hbbc27d93),
	.w7(32'hbbb4a004),
	.w8(32'hbb5bd034),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83158b),
	.w1(32'hbb6d71ce),
	.w2(32'h39f5324e),
	.w3(32'hbb8fa56f),
	.w4(32'hbb814dbb),
	.w5(32'hb822f686),
	.w6(32'hbb7f20bf),
	.w7(32'hbb685e79),
	.w8(32'h39d4c631),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c27511),
	.w1(32'h38ec20bf),
	.w2(32'hba28d842),
	.w3(32'hba7a1f11),
	.w4(32'hb8c16a70),
	.w5(32'hba9bcba3),
	.w6(32'hb9ac7156),
	.w7(32'h39846c85),
	.w8(32'h3a3be357),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928c20f),
	.w1(32'hb7c3958d),
	.w2(32'hb9b56638),
	.w3(32'hba4b0c14),
	.w4(32'hba177b12),
	.w5(32'h3b0ad35b),
	.w6(32'h39120c02),
	.w7(32'hba109ea1),
	.w8(32'hb8f32c96),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104b0c),
	.w1(32'hba6a55e2),
	.w2(32'hba83254e),
	.w3(32'h3a5f15e4),
	.w4(32'h3b247978),
	.w5(32'h3ac3fdb0),
	.w6(32'hbaf7aa31),
	.w7(32'hbad2920a),
	.w8(32'hba9dc69d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba881cbf),
	.w1(32'hbac2c048),
	.w2(32'h3ae7e09b),
	.w3(32'h3aee7272),
	.w4(32'h39ce33f6),
	.w5(32'h3b13053f),
	.w6(32'hbab5a7c0),
	.w7(32'hbab989e9),
	.w8(32'hb980fe22),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c39514),
	.w1(32'hba84a10e),
	.w2(32'hba59cd2d),
	.w3(32'h3b91560d),
	.w4(32'hb902df5e),
	.w5(32'h39e41393),
	.w6(32'h39ce6921),
	.w7(32'hb9b1c8a8),
	.w8(32'hb9c449a0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39708f2f),
	.w1(32'h3892067d),
	.w2(32'h39e42ca2),
	.w3(32'h3b099478),
	.w4(32'h3ae9897d),
	.w5(32'hbac686a2),
	.w6(32'h39f44088),
	.w7(32'h3a8b425f),
	.w8(32'hba429cfe),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96bd6c7),
	.w1(32'h3ada1585),
	.w2(32'hba81ab57),
	.w3(32'hbb0bb63f),
	.w4(32'h3a7d9cf2),
	.w5(32'h3afa1427),
	.w6(32'hbb130d14),
	.w7(32'h39e3c879),
	.w8(32'hb9092985),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ae8ba),
	.w1(32'hba955198),
	.w2(32'hbab08b37),
	.w3(32'h3b164da9),
	.w4(32'h3b162544),
	.w5(32'h3b1361d1),
	.w6(32'hba304f1c),
	.w7(32'hba5bc419),
	.w8(32'h3a5f9e07),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0359c2),
	.w1(32'hbab4fe57),
	.w2(32'hb9a6f73f),
	.w3(32'h3abe9426),
	.w4(32'h3b1e770d),
	.w5(32'h39f802ca),
	.w6(32'h3a483048),
	.w7(32'h3afd42f0),
	.w8(32'h3a8541b8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba411412),
	.w1(32'hb9f59e65),
	.w2(32'hba6e7f68),
	.w3(32'hb9acaa18),
	.w4(32'h3a2f37c0),
	.w5(32'hba9e364c),
	.w6(32'h391d26f5),
	.w7(32'h39c32471),
	.w8(32'hbaab5357),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe23e3),
	.w1(32'hba1b65db),
	.w2(32'hba2fc7bf),
	.w3(32'hbae920c5),
	.w4(32'h3ac09022),
	.w5(32'hba8d3fb4),
	.w6(32'h38ed0bc4),
	.w7(32'h3b4861d1),
	.w8(32'h393facc8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40b081),
	.w1(32'hbaf70521),
	.w2(32'hb9756102),
	.w3(32'hba28cf4a),
	.w4(32'hbb0f3b18),
	.w5(32'hb97a6167),
	.w6(32'hb9840fa4),
	.w7(32'hb9eb4d48),
	.w8(32'h3954f1e8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38717b9d),
	.w1(32'hb97e399c),
	.w2(32'hbaba9141),
	.w3(32'h38495371),
	.w4(32'h3987060e),
	.w5(32'hba9a1e00),
	.w6(32'h3aab710d),
	.w7(32'h3a3785b5),
	.w8(32'hba13c840),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36bce9),
	.w1(32'hba9ef2b1),
	.w2(32'hbb0a77af),
	.w3(32'h3891edf6),
	.w4(32'hbac3ab21),
	.w5(32'hb967ed7b),
	.w6(32'h3a5a2d66),
	.w7(32'hb9f59153),
	.w8(32'hb9cdecca),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ed12),
	.w1(32'hb8c649c2),
	.w2(32'h38632d68),
	.w3(32'hba626e55),
	.w4(32'h3aaa2cc7),
	.w5(32'h39d434a3),
	.w6(32'hbaca2440),
	.w7(32'h3908f680),
	.w8(32'hb9460bf9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa966),
	.w1(32'hba479c8c),
	.w2(32'hbb05ddf4),
	.w3(32'hbad6fed3),
	.w4(32'hba5502ca),
	.w5(32'h3ac9a1dd),
	.w6(32'hbb106ed2),
	.w7(32'hbb24db7a),
	.w8(32'hba76b3e9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061909),
	.w1(32'hbac309bd),
	.w2(32'h39f12f80),
	.w3(32'h3a5d1316),
	.w4(32'h3aab5700),
	.w5(32'h3a1f3a08),
	.w6(32'hba2749cc),
	.w7(32'hb81f3e53),
	.w8(32'h39eaa893),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6e056),
	.w1(32'hba78d258),
	.w2(32'h3a38cfa0),
	.w3(32'h3a79c697),
	.w4(32'h39f5cfaf),
	.w5(32'h3b052109),
	.w6(32'h38ea8568),
	.w7(32'h3aae586b),
	.w8(32'h3a7b3a78),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10be57),
	.w1(32'h396f715b),
	.w2(32'hbb053ee2),
	.w3(32'hb9eeeaf5),
	.w4(32'h3aaed598),
	.w5(32'hbb1d1a70),
	.w6(32'h38872d4f),
	.w7(32'h39fb3f59),
	.w8(32'hbac8af3e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb356616),
	.w1(32'hbb6f7180),
	.w2(32'hba26b2c6),
	.w3(32'hbb38c6cd),
	.w4(32'hbb3c521a),
	.w5(32'h3aa32b57),
	.w6(32'hbb35c294),
	.w7(32'hbb04f9bb),
	.w8(32'hba283055),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0af279),
	.w1(32'h3aa289a9),
	.w2(32'hbabbb4c5),
	.w3(32'h3a521e48),
	.w4(32'h3a93d9ef),
	.w5(32'hbb1f6886),
	.w6(32'h3a6fe19c),
	.w7(32'hba28100b),
	.w8(32'h3a12d614),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c6b9f),
	.w1(32'hbb132c2f),
	.w2(32'h3832e79f),
	.w3(32'hbb418b27),
	.w4(32'hbb48f974),
	.w5(32'h3953eed8),
	.w6(32'h3a4c7ff9),
	.w7(32'h3aae5727),
	.w8(32'hbadaf0bc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb752f381),
	.w1(32'h3a1940ef),
	.w2(32'h3b7248c6),
	.w3(32'hb90554b2),
	.w4(32'h39ab7ad4),
	.w5(32'h3ae4b7c4),
	.w6(32'hbb2e10ae),
	.w7(32'hbb120bfd),
	.w8(32'h3b1d03fb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b2e75),
	.w1(32'h3b643722),
	.w2(32'hb9fad88a),
	.w3(32'h3a832d6b),
	.w4(32'h3aefc883),
	.w5(32'hbae31b0e),
	.w6(32'h3aeb48f4),
	.w7(32'h3b5af30b),
	.w8(32'hba0d9e97),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04acaf),
	.w1(32'hba149d08),
	.w2(32'h3a90f7f2),
	.w3(32'hbb181406),
	.w4(32'hbb01ccb4),
	.w5(32'h3b80c78f),
	.w6(32'hba8f91cd),
	.w7(32'hba4c07c6),
	.w8(32'h393ce0de),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b3ca0),
	.w1(32'h39f6dd68),
	.w2(32'hba67df98),
	.w3(32'h3b015d21),
	.w4(32'h3b63589a),
	.w5(32'h3a4c8c96),
	.w6(32'hbabcf6fc),
	.w7(32'h38b5c86f),
	.w8(32'hb9ed62ea),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a82f),
	.w1(32'hba81b690),
	.w2(32'h3b13027c),
	.w3(32'hb8482ace),
	.w4(32'h39d92618),
	.w5(32'h3a85d948),
	.w6(32'hbb13e8c2),
	.w7(32'hb97e6f52),
	.w8(32'h3a7b2719),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3237e4),
	.w1(32'h3aab17e4),
	.w2(32'h3a7b66c8),
	.w3(32'h3adaecbb),
	.w4(32'h3a572b21),
	.w5(32'h3a959d5f),
	.w6(32'h3a895867),
	.w7(32'h3a81d58b),
	.w8(32'h3aae83db),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a463164),
	.w1(32'h3a7c7356),
	.w2(32'h3a991dcc),
	.w3(32'h3a8b5790),
	.w4(32'h3a8278f5),
	.w5(32'h3b05f785),
	.w6(32'h3a90d7f9),
	.w7(32'h3aad4d03),
	.w8(32'h3b034271),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcdbc3),
	.w1(32'h3b0e8928),
	.w2(32'hba779fd1),
	.w3(32'h3b553f5e),
	.w4(32'h3b68af66),
	.w5(32'hbb06846c),
	.w6(32'h3b427c98),
	.w7(32'h3b50e4da),
	.w8(32'hba57748c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749e29),
	.w1(32'hba190d38),
	.w2(32'h398ceb5f),
	.w3(32'hbb956e07),
	.w4(32'h398b45a9),
	.w5(32'h3752e9b7),
	.w6(32'hbafb2a96),
	.w7(32'h3a1070a5),
	.w8(32'hba0aa5c7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ea103),
	.w1(32'hbae4c0b1),
	.w2(32'hbb2448e4),
	.w3(32'hb984c3a0),
	.w4(32'hbb1add53),
	.w5(32'hbb0a79df),
	.w6(32'hba9df584),
	.w7(32'hbb326d6a),
	.w8(32'hba9019ec),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba472e76),
	.w1(32'hba4042a5),
	.w2(32'hba6c4175),
	.w3(32'hb995896f),
	.w4(32'hba974853),
	.w5(32'hbaf45c9c),
	.w6(32'hbac1fc3d),
	.w7(32'hbad4f072),
	.w8(32'hbaf1db63),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1f2b1),
	.w1(32'h39768cbd),
	.w2(32'h3aa5cfba),
	.w3(32'h39bc1c2f),
	.w4(32'hb953ab49),
	.w5(32'h3a272d05),
	.w6(32'h3a6de2e0),
	.w7(32'h3a125e99),
	.w8(32'h3a703ccf),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae828f),
	.w1(32'h3b3025ff),
	.w2(32'h395b74ef),
	.w3(32'h3b076626),
	.w4(32'h3b0b72bd),
	.w5(32'h39fa6ad8),
	.w6(32'h3af70eb1),
	.w7(32'h3af3ce33),
	.w8(32'hba8e6e9a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule