module layer_8_featuremap_174(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacafd54),
	.w1(32'hbc713516),
	.w2(32'hbc45b3e2),
	.w3(32'h3b00c7cb),
	.w4(32'h3b9e7dc0),
	.w5(32'hbc032447),
	.w6(32'hbc4ef61a),
	.w7(32'hbae6199d),
	.w8(32'h3aad931e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b51a8),
	.w1(32'hbb4250a6),
	.w2(32'hbb7d935b),
	.w3(32'hbc7b4d5d),
	.w4(32'hbb6e9254),
	.w5(32'hbbc05062),
	.w6(32'hbb6882a0),
	.w7(32'hbb77a59c),
	.w8(32'hbba2dae3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae69d74),
	.w1(32'hbbc5e552),
	.w2(32'h3af7bfeb),
	.w3(32'hbb66c14e),
	.w4(32'hbba8b321),
	.w5(32'h39e7a036),
	.w6(32'hbc01d472),
	.w7(32'hbc33679b),
	.w8(32'hbc237319),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25232b),
	.w1(32'hbb9f9263),
	.w2(32'hbb252b49),
	.w3(32'hb9b72b0f),
	.w4(32'hbc2e26cd),
	.w5(32'hba04c842),
	.w6(32'hbbd160d4),
	.w7(32'hbc3322fa),
	.w8(32'hbc01ea6f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d411),
	.w1(32'hbbca4393),
	.w2(32'hbbbbb3d1),
	.w3(32'hbb5edc72),
	.w4(32'hbbed363c),
	.w5(32'hbc004851),
	.w6(32'h3afc46d9),
	.w7(32'hbb7883c4),
	.w8(32'hbb2ba61c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85c315),
	.w1(32'h3c46ab99),
	.w2(32'hbbc0915f),
	.w3(32'h3af35e70),
	.w4(32'h3b3b154f),
	.w5(32'hbbb8654c),
	.w6(32'h3b38e510),
	.w7(32'hbb8406a2),
	.w8(32'hbc6e1a32),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ac655),
	.w1(32'h3ab26cb7),
	.w2(32'h39f66226),
	.w3(32'h3aec0713),
	.w4(32'h36b075ef),
	.w5(32'h39f4327a),
	.w6(32'h3a9aca95),
	.w7(32'hbacbad73),
	.w8(32'h39c2ca25),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed030),
	.w1(32'hbc4bac37),
	.w2(32'hbb21411d),
	.w3(32'hbc7a206b),
	.w4(32'hbcc7f8f4),
	.w5(32'hbcab7d36),
	.w6(32'hbb4a5773),
	.w7(32'hbc2ef9e7),
	.w8(32'hbc10e30d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc369f72),
	.w1(32'hbc1cf1e7),
	.w2(32'hbb8d786f),
	.w3(32'hbcad27a4),
	.w4(32'hbc56665a),
	.w5(32'hbc232d78),
	.w6(32'h3a6af576),
	.w7(32'hbbdb0079),
	.w8(32'hbb736fcb),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ccbe8),
	.w1(32'h3be05d15),
	.w2(32'hbc346590),
	.w3(32'h3acb0f9c),
	.w4(32'h3c1b4aaf),
	.w5(32'h3c534421),
	.w6(32'h3ac95c30),
	.w7(32'hbbb11ba4),
	.w8(32'hbb99aa3f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4aaea),
	.w1(32'hbb4dc55d),
	.w2(32'hbc664d58),
	.w3(32'h3c3e163f),
	.w4(32'hbc3c8056),
	.w5(32'hbc5eb59d),
	.w6(32'h3ac30d77),
	.w7(32'hbbb49608),
	.w8(32'hbbd0e1bd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03132f),
	.w1(32'hbc031811),
	.w2(32'hbc45b824),
	.w3(32'hbc417263),
	.w4(32'hbc1b5e35),
	.w5(32'hbc191ca6),
	.w6(32'h3a94db1b),
	.w7(32'h3a94138b),
	.w8(32'hbb905515),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf39b13),
	.w1(32'hbbc7bca8),
	.w2(32'hbc28fac3),
	.w3(32'hbbc2e79a),
	.w4(32'hbc1364ac),
	.w5(32'hbc06bfca),
	.w6(32'hbc1ae5f0),
	.w7(32'hbc07be7a),
	.w8(32'hbbd2e9a9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02309c),
	.w1(32'h3b3f24dc),
	.w2(32'h3bde8186),
	.w3(32'hbbd02d1d),
	.w4(32'h3c9d63b8),
	.w5(32'h3c709ac1),
	.w6(32'hbc1a256d),
	.w7(32'hba2ed6d1),
	.w8(32'hbad22d9c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a674fcf),
	.w1(32'h3b5763e6),
	.w2(32'h3a5a2854),
	.w3(32'hbaec8679),
	.w4(32'h3b8cef97),
	.w5(32'h3ae96b07),
	.w6(32'h3b95bd52),
	.w7(32'hba21ed1f),
	.w8(32'h3a7b850e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ea24d),
	.w1(32'hbb98b847),
	.w2(32'hbad59b95),
	.w3(32'hb982b4f1),
	.w4(32'hbb8d87dd),
	.w5(32'hbc80dfe4),
	.w6(32'hbb81497a),
	.w7(32'h3bd38456),
	.w8(32'h3b394e06),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafbfa3),
	.w1(32'hbad05b6e),
	.w2(32'hbc0d141e),
	.w3(32'hbc9402ef),
	.w4(32'hbc101681),
	.w5(32'h3b3052e2),
	.w6(32'h3c1107e2),
	.w7(32'hbb66910a),
	.w8(32'hbc1ea81a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35d58b),
	.w1(32'hbadd1830),
	.w2(32'h3af28dca),
	.w3(32'h3c21d89d),
	.w4(32'h3ab3b558),
	.w5(32'h3b30d3bd),
	.w6(32'h3a674c51),
	.w7(32'h3a914ff9),
	.w8(32'hbbb8b1c0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc1a25),
	.w1(32'hbc3ffaf3),
	.w2(32'hbca5cf2b),
	.w3(32'hbc0879db),
	.w4(32'hbca68820),
	.w5(32'hbcb8648c),
	.w6(32'h3c8fa92e),
	.w7(32'hbb9f1f2b),
	.w8(32'h3bcc9af9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4de3f8),
	.w1(32'hba8c9ce4),
	.w2(32'hbbe85a44),
	.w3(32'hbbe76edb),
	.w4(32'hbb0846bd),
	.w5(32'hbb8b9a52),
	.w6(32'h3c60fb65),
	.w7(32'h3c186baa),
	.w8(32'h3ac7ae16),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce9bc),
	.w1(32'h3b3473e4),
	.w2(32'h3b01c22c),
	.w3(32'h3bdf8f20),
	.w4(32'hb92e3aa6),
	.w5(32'h3ae10aa6),
	.w6(32'h3b95f475),
	.w7(32'h3c39d1f4),
	.w8(32'hbb3eda0f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44ad79),
	.w1(32'hbc08d435),
	.w2(32'h3b7aefb5),
	.w3(32'hba112ac7),
	.w4(32'hbc14c087),
	.w5(32'hbbbda25d),
	.w6(32'hbc299716),
	.w7(32'hbb16cc38),
	.w8(32'h3a91c2d1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8f157),
	.w1(32'hbb8ec03f),
	.w2(32'hbac8a922),
	.w3(32'h3ca2d4a9),
	.w4(32'hbcdd327c),
	.w5(32'hbccea610),
	.w6(32'h3cf820b9),
	.w7(32'h3b69ab62),
	.w8(32'hbb05127f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd67d0),
	.w1(32'hbbc5e09e),
	.w2(32'hbb80bed5),
	.w3(32'h3bb4532e),
	.w4(32'hbc14f48f),
	.w5(32'hbbbb0ab9),
	.w6(32'hbb98fb15),
	.w7(32'hbb9e1f6b),
	.w8(32'hbbbbec67),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b6bea),
	.w1(32'hbb17422d),
	.w2(32'hbb7a07c6),
	.w3(32'hba944136),
	.w4(32'h3be8afc7),
	.w5(32'h3bd53d26),
	.w6(32'hba9f53f6),
	.w7(32'hbb03d8df),
	.w8(32'hbb6b3456),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb4552),
	.w1(32'hbc8c4ffb),
	.w2(32'hbc50cd65),
	.w3(32'h3c90a57a),
	.w4(32'h3a43f01d),
	.w5(32'hbc492131),
	.w6(32'h3ad4d19d),
	.w7(32'h3c5f70bd),
	.w8(32'hbaf8333d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e43e2),
	.w1(32'hbb935538),
	.w2(32'hbb7237a6),
	.w3(32'h39df4769),
	.w4(32'hbb17ef76),
	.w5(32'h3b58711d),
	.w6(32'h3a36fe04),
	.w7(32'hbb598b5d),
	.w8(32'hbb335493),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01c376),
	.w1(32'hbc9efcea),
	.w2(32'hbd68c6c2),
	.w3(32'h3bbf6fd4),
	.w4(32'hbd6213eb),
	.w5(32'hbd8c0fdb),
	.w6(32'h3b314f02),
	.w7(32'hbcba9a62),
	.w8(32'hbd40a627),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ffd70),
	.w1(32'hba15b1fc),
	.w2(32'hbb115972),
	.w3(32'hbbad896f),
	.w4(32'hbbe44e85),
	.w5(32'hbc391120),
	.w6(32'h3bdd5e0d),
	.w7(32'h3b9e8bf8),
	.w8(32'h3a84d8c9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb386a6b),
	.w1(32'hbb00ede6),
	.w2(32'hbb9b142a),
	.w3(32'hbbe2d96a),
	.w4(32'h3cc118b8),
	.w5(32'h3c93ff97),
	.w6(32'hbb304c5c),
	.w7(32'hbb97bbf0),
	.w8(32'hbc844974),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56b380),
	.w1(32'h3c33320f),
	.w2(32'h3b7db80e),
	.w3(32'h3c6ad174),
	.w4(32'h3c4956f9),
	.w5(32'h3c09dd13),
	.w6(32'h3a8dad66),
	.w7(32'h3a8474fd),
	.w8(32'hbb301221),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d09a),
	.w1(32'h3a80423f),
	.w2(32'hbb9003b9),
	.w3(32'h3bba7933),
	.w4(32'h3b4567f6),
	.w5(32'hbb3c5077),
	.w6(32'h3ba52e68),
	.w7(32'h3b035d39),
	.w8(32'hbbd5f7e0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c6f42),
	.w1(32'h3c06ab1e),
	.w2(32'h3b926ff9),
	.w3(32'h3af53890),
	.w4(32'h3c154e59),
	.w5(32'h39e00f03),
	.w6(32'h3b77de04),
	.w7(32'hbb181f4a),
	.w8(32'hbb2ec58a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae84e73),
	.w1(32'h3c210bd1),
	.w2(32'h3b0dc339),
	.w3(32'h38af093a),
	.w4(32'h3c63e95a),
	.w5(32'h3c460dc7),
	.w6(32'h3b00653b),
	.w7(32'h3992768f),
	.w8(32'h3b8e7a89),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7da0b0),
	.w1(32'h3b20dd44),
	.w2(32'h3ab5ea1e),
	.w3(32'h3b3c3800),
	.w4(32'h3bc16bd0),
	.w5(32'h3bb901d1),
	.w6(32'h3b7a453f),
	.w7(32'h3b9b3606),
	.w8(32'h390db68e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cc03f),
	.w1(32'hbc11898c),
	.w2(32'hbbe44129),
	.w3(32'h3aa76de1),
	.w4(32'hbc4e000c),
	.w5(32'hbc267df4),
	.w6(32'hbac8c98a),
	.w7(32'h3b1ad87a),
	.w8(32'h3b5a3bdf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69219f),
	.w1(32'h3b26b493),
	.w2(32'h3a80ce0f),
	.w3(32'h3b82a6ac),
	.w4(32'hb7eaf807),
	.w5(32'h3ae80eb4),
	.w6(32'h3b18c7a1),
	.w7(32'h3b1c4186),
	.w8(32'h3b8b3cb4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b942f),
	.w1(32'h3b29683b),
	.w2(32'hba157f0f),
	.w3(32'h3b2ddcf7),
	.w4(32'hbabb1294),
	.w5(32'hbb66a7b0),
	.w6(32'h3bc602a7),
	.w7(32'h3a4ccb3f),
	.w8(32'h3b38c482),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a343844),
	.w1(32'hbbc02b1c),
	.w2(32'hbbc82dd8),
	.w3(32'hbb305dfb),
	.w4(32'hbc2ae7b2),
	.w5(32'hbc030410),
	.w6(32'hbb9b1e9e),
	.w7(32'hbaa58955),
	.w8(32'hbbf94d9f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edde97),
	.w1(32'hbb92da2f),
	.w2(32'hbb02e420),
	.w3(32'h3ade17c8),
	.w4(32'hbb4b4a71),
	.w5(32'hbb9a2b1a),
	.w6(32'hba10b670),
	.w7(32'hbb3e2445),
	.w8(32'h3a46d3dc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d15cd1),
	.w1(32'hbc1a3930),
	.w2(32'hbc8db86c),
	.w3(32'hbc3cac7e),
	.w4(32'hbc852dc2),
	.w5(32'hbcaec085),
	.w6(32'hbbcaeabf),
	.w7(32'hbb944825),
	.w8(32'hbc4c6d9a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1e15d),
	.w1(32'h3b61cf9f),
	.w2(32'hbb8dae2d),
	.w3(32'hbc080c1d),
	.w4(32'hb9e35c46),
	.w5(32'hbb8d8a52),
	.w6(32'h3ba00892),
	.w7(32'hbad571c1),
	.w8(32'hbb44616f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e383),
	.w1(32'hbacd3103),
	.w2(32'hbaded3b2),
	.w3(32'h3b1eae02),
	.w4(32'h3c0d85bd),
	.w5(32'h3bde7977),
	.w6(32'hba0d9768),
	.w7(32'h39c893b7),
	.w8(32'h3b1e699a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde0796),
	.w1(32'h3b9a5975),
	.w2(32'hbba18840),
	.w3(32'h3c439512),
	.w4(32'hbb9352c3),
	.w5(32'hbc4ead88),
	.w6(32'h3c07d38b),
	.w7(32'h3b1f342b),
	.w8(32'hbbc86c93),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af174b8),
	.w1(32'hbc98af4b),
	.w2(32'hbb9a645b),
	.w3(32'hbbd745ec),
	.w4(32'hbc965965),
	.w5(32'hbbaaf9b9),
	.w6(32'h3b009182),
	.w7(32'h3bbd31af),
	.w8(32'h3c04a9d4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b850e5e),
	.w1(32'hbb8d06ce),
	.w2(32'hbb591d43),
	.w3(32'h3c24f555),
	.w4(32'hba443169),
	.w5(32'h3a911d9e),
	.w6(32'h3ac70f7d),
	.w7(32'h3acc4ff7),
	.w8(32'h3a3891f3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bc033),
	.w1(32'hbc2e0645),
	.w2(32'hbc4ce83a),
	.w3(32'h3a867a17),
	.w4(32'hbbbc9580),
	.w5(32'hbc56a309),
	.w6(32'hbb8a5ee8),
	.w7(32'hbc0c8bdf),
	.w8(32'hbaf75e17),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87013f),
	.w1(32'hbc4a209b),
	.w2(32'hbbf5d11a),
	.w3(32'hbb6b7117),
	.w4(32'hbc8f8083),
	.w5(32'hbc5cffae),
	.w6(32'h3ac01494),
	.w7(32'hbb2c5485),
	.w8(32'h3b9fd2e2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801a39),
	.w1(32'hbbe36d17),
	.w2(32'hbbca8e39),
	.w3(32'hbb3f51ed),
	.w4(32'hbc1b9218),
	.w5(32'hbbbbcaff),
	.w6(32'hbbfb48ef),
	.w7(32'h3b7d2e6c),
	.w8(32'hbbd1aac2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e50e6),
	.w1(32'hba32c853),
	.w2(32'hbc35d464),
	.w3(32'h3ad6764b),
	.w4(32'h3b8c0b19),
	.w5(32'hbc0f87f5),
	.w6(32'h3a6c758f),
	.w7(32'h384604c6),
	.w8(32'hbb333333),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b115233),
	.w1(32'h3ba138a6),
	.w2(32'hbb51d8ee),
	.w3(32'hba1f338d),
	.w4(32'h3bf9af96),
	.w5(32'h3ae10748),
	.w6(32'h3beca2d7),
	.w7(32'h3c2693f7),
	.w8(32'h3bda9247),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3595c9),
	.w1(32'h3c144530),
	.w2(32'hba84f05c),
	.w3(32'hbbe6433e),
	.w4(32'hbcb65a1f),
	.w5(32'hbc53ccc1),
	.w6(32'h3b9bee6b),
	.w7(32'hbc958468),
	.w8(32'hbc3a3ebe),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ff22d),
	.w1(32'hbb0be558),
	.w2(32'hbbc8c446),
	.w3(32'hbc2c7dea),
	.w4(32'hbc466eb8),
	.w5(32'hbc293fe9),
	.w6(32'hbb6befb9),
	.w7(32'hbc39674a),
	.w8(32'hbbce81ea),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88640b),
	.w1(32'h3b8182be),
	.w2(32'hbb8a98c6),
	.w3(32'h3a5032cc),
	.w4(32'h3a1fecf8),
	.w5(32'hbc1cbf22),
	.w6(32'h3c8e38ec),
	.w7(32'h3c0fecdd),
	.w8(32'h3c2ff119),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bba40),
	.w1(32'h3c226ca2),
	.w2(32'h395d9a0d),
	.w3(32'hbba53e7a),
	.w4(32'h3c21919c),
	.w5(32'h3ba5c434),
	.w6(32'h3b8ba73f),
	.w7(32'hbb188ad3),
	.w8(32'h3b0b7542),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b19c2),
	.w1(32'hbbcea7ce),
	.w2(32'hbc8f95af),
	.w3(32'h3bd2a765),
	.w4(32'hbc343c82),
	.w5(32'hbc8cd65c),
	.w6(32'h3c6bd90a),
	.w7(32'hbb15e496),
	.w8(32'hb9512d1d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7dd4a),
	.w1(32'h3c090ccb),
	.w2(32'h3c108503),
	.w3(32'h3b4460ae),
	.w4(32'h3c0f8e38),
	.w5(32'h3bae4f39),
	.w6(32'h3c2db924),
	.w7(32'h3bd3f166),
	.w8(32'h3bbf806f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08e6c),
	.w1(32'h3a2ad33f),
	.w2(32'h3b7fce69),
	.w3(32'hb98181e1),
	.w4(32'hbc1564fa),
	.w5(32'hbacb6fc5),
	.w6(32'hbb96b21a),
	.w7(32'hbc29dc63),
	.w8(32'hbc1cb525),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83318f),
	.w1(32'hbb8e7c59),
	.w2(32'hbc026f84),
	.w3(32'h3bb0ce8f),
	.w4(32'hbbd4854b),
	.w5(32'hbc1bde1e),
	.w6(32'hbafec7d7),
	.w7(32'hbbd938a8),
	.w8(32'hbbaa1600),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995e3f9),
	.w1(32'hbba19740),
	.w2(32'hbb587082),
	.w3(32'hbad9a6f6),
	.w4(32'hbbacf94b),
	.w5(32'hb9deb778),
	.w6(32'hbbb4732c),
	.w7(32'hbc289518),
	.w8(32'hbb6c713b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eba95),
	.w1(32'hb967422d),
	.w2(32'hbbd0f718),
	.w3(32'hbbaf5ba6),
	.w4(32'hbbdeceb1),
	.w5(32'hbc13f5cf),
	.w6(32'hb8ce144f),
	.w7(32'hbb5ff0ae),
	.w8(32'hbc356cef),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a7d97),
	.w1(32'h3bd0202a),
	.w2(32'h3bba5b45),
	.w3(32'hba83dd8f),
	.w4(32'hbb7bcc2c),
	.w5(32'hbbdec7e4),
	.w6(32'h3c1665a0),
	.w7(32'h3bb84741),
	.w8(32'h3bd5aa2e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09f54a),
	.w1(32'h39a6aac5),
	.w2(32'hbc0134a4),
	.w3(32'hbc7264a1),
	.w4(32'hbbeb8552),
	.w5(32'hbbfd09c0),
	.w6(32'h3c216bcd),
	.w7(32'h3ae35046),
	.w8(32'hbc5964e8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ef61f),
	.w1(32'hbb9fd3d1),
	.w2(32'hbb584cb1),
	.w3(32'hbb26825c),
	.w4(32'hbc528deb),
	.w5(32'hbc31b4d3),
	.w6(32'hbc09a54e),
	.w7(32'hbc1703a4),
	.w8(32'hbb7a5a05),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af70944),
	.w1(32'h3b1e6126),
	.w2(32'h38c3539e),
	.w3(32'hbb9e0f21),
	.w4(32'hba3feeff),
	.w5(32'hbb5235d1),
	.w6(32'h3a7c003f),
	.w7(32'hb96c1e45),
	.w8(32'hb9cc41cb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986134e),
	.w1(32'hbbe61a48),
	.w2(32'hbbefebb0),
	.w3(32'hbb52e669),
	.w4(32'hbc4b5168),
	.w5(32'hbc374aa2),
	.w6(32'hbb4cbc5c),
	.w7(32'hbbd2546a),
	.w8(32'hbc0a5c14),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b379a),
	.w1(32'hbbd84e6d),
	.w2(32'hbb8d3f44),
	.w3(32'hbad3d9b0),
	.w4(32'hbc292fde),
	.w5(32'hbb32fad4),
	.w6(32'hbb32276d),
	.w7(32'h3b02484c),
	.w8(32'hbb9e5c04),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6dee1),
	.w1(32'hbc10fd3b),
	.w2(32'hbc5a1d19),
	.w3(32'h3c0a901c),
	.w4(32'hbb06716c),
	.w5(32'hbbe7558f),
	.w6(32'h3b434987),
	.w7(32'h3b93bef9),
	.w8(32'h3b581f1d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc57a64),
	.w1(32'h3b64670c),
	.w2(32'h3b2a153e),
	.w3(32'hbb896ca3),
	.w4(32'h3c7d7197),
	.w5(32'hba9d5f8e),
	.w6(32'h38030f4a),
	.w7(32'h3a847610),
	.w8(32'hbbe6fd47),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9640ef),
	.w1(32'hbb8d6178),
	.w2(32'hbc58d450),
	.w3(32'h3c8235b2),
	.w4(32'hbce94526),
	.w5(32'hbccf6acc),
	.w6(32'hbb958e59),
	.w7(32'hbc5ca81b),
	.w8(32'hbca5936a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96930a),
	.w1(32'h3b002b02),
	.w2(32'h3a1c2317),
	.w3(32'h3b4c181e),
	.w4(32'h3b856473),
	.w5(32'h3b9f071a),
	.w6(32'hbac1e406),
	.w7(32'hbb4bfb45),
	.w8(32'hbb05d03c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae41cef),
	.w1(32'hbb1e0759),
	.w2(32'h3b35b5df),
	.w3(32'hbbe37e36),
	.w4(32'hbb69661a),
	.w5(32'h3b504579),
	.w6(32'h3b7d725a),
	.w7(32'hbb9a7828),
	.w8(32'hbbe1381b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3ae2),
	.w1(32'hbac01298),
	.w2(32'h3c09d415),
	.w3(32'h3bf99556),
	.w4(32'hbbb383b1),
	.w5(32'h3a941739),
	.w6(32'hbba97cc3),
	.w7(32'h3b3f7b06),
	.w8(32'h3b7a06b2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc3507),
	.w1(32'hbc0a1a72),
	.w2(32'hbbc20f46),
	.w3(32'h3bea6ed5),
	.w4(32'hbc443229),
	.w5(32'hbc1d1472),
	.w6(32'hbb92a29f),
	.w7(32'hbbfb9b99),
	.w8(32'hbc03ae91),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ea9ce),
	.w1(32'hbb884efe),
	.w2(32'h3b8d953c),
	.w3(32'h3b989585),
	.w4(32'hbbcb11f4),
	.w5(32'hbaa0005c),
	.w6(32'hba81ccf7),
	.w7(32'hbab44ca5),
	.w8(32'h3b5da91c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47c9b3),
	.w1(32'h3a9f2781),
	.w2(32'h3c01b7d5),
	.w3(32'h3c306c65),
	.w4(32'hbbc685d5),
	.w5(32'hbaee2b4c),
	.w6(32'h3c54911e),
	.w7(32'h3b886e18),
	.w8(32'hbb1b6a3b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32848c),
	.w1(32'hbb71f8d1),
	.w2(32'h3aab4f34),
	.w3(32'hbb66eca4),
	.w4(32'hb8fdaf05),
	.w5(32'h3b47b586),
	.w6(32'hbb05946c),
	.w7(32'hbac59cd2),
	.w8(32'hbb14d788),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd8494),
	.w1(32'hbb988eef),
	.w2(32'hbbf82785),
	.w3(32'h3b67b016),
	.w4(32'hbc6982ec),
	.w5(32'hbc538e11),
	.w6(32'h3b6c4a7d),
	.w7(32'hb85847e2),
	.w8(32'hbbc0cb1d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23d88c),
	.w1(32'hbb869746),
	.w2(32'hbc10a585),
	.w3(32'hbb026f8a),
	.w4(32'h3ad0bc90),
	.w5(32'hba47369d),
	.w6(32'hbb401805),
	.w7(32'hbb0797fb),
	.w8(32'hbad95727),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14773e),
	.w1(32'h3bc0631e),
	.w2(32'hbb0c09d8),
	.w3(32'hbb4aa1f3),
	.w4(32'h3bb2eebb),
	.w5(32'hb921b134),
	.w6(32'h388bb226),
	.w7(32'hbb54d858),
	.w8(32'hbc06f18e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefb5a1),
	.w1(32'hbb9e361c),
	.w2(32'h3bf6887b),
	.w3(32'hbc181ca2),
	.w4(32'h3b94d59d),
	.w5(32'h3c277f51),
	.w6(32'hbbb3ae8d),
	.w7(32'hba4fb37b),
	.w8(32'hbbbee474),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12bbe),
	.w1(32'h39527a36),
	.w2(32'h3c1df147),
	.w3(32'h3b4c70d6),
	.w4(32'h3c3cb0d0),
	.w5(32'h3bc05e44),
	.w6(32'hba000885),
	.w7(32'hbb50fa49),
	.w8(32'hbbdacbbd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6e71b),
	.w1(32'hbbfd926a),
	.w2(32'hbc195ac1),
	.w3(32'hbb783a62),
	.w4(32'hbc4d1177),
	.w5(32'hbc2704b6),
	.w6(32'hbbb15941),
	.w7(32'h3935dc0a),
	.w8(32'h3a725597),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d419d1),
	.w1(32'hbbc910e3),
	.w2(32'hbc642b27),
	.w3(32'hbc9125af),
	.w4(32'hbc2731a1),
	.w5(32'hbc5e89e7),
	.w6(32'hbc021089),
	.w7(32'h394c2cc9),
	.w8(32'hbbd6abf6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf59cdd),
	.w1(32'hbc835cec),
	.w2(32'hbc35e89e),
	.w3(32'hb9c0d420),
	.w4(32'hbcb09fc0),
	.w5(32'hbcae155e),
	.w6(32'h3aa1519e),
	.w7(32'hbbe5e6ef),
	.w8(32'hba1871ec),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d31a),
	.w1(32'hbbad55f5),
	.w2(32'hbc0a7ed6),
	.w3(32'h3b93566b),
	.w4(32'hbc8e4d56),
	.w5(32'hbc03a724),
	.w6(32'h38a4c55f),
	.w7(32'hbc4644ef),
	.w8(32'hbc55b076),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847110),
	.w1(32'h3b3428f0),
	.w2(32'hbb239155),
	.w3(32'h3bd13a6f),
	.w4(32'h3bb8b8c3),
	.w5(32'h3baefc85),
	.w6(32'h39e9c938),
	.w7(32'hbb136c01),
	.w8(32'hbb8769e5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c6a6),
	.w1(32'hbbb6dcc1),
	.w2(32'hbbef5241),
	.w3(32'hbad22639),
	.w4(32'hbb9c1830),
	.w5(32'hbb1bdb85),
	.w6(32'h3ac1939a),
	.w7(32'hbace6af2),
	.w8(32'hbacf7b1c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf32392),
	.w1(32'h39187632),
	.w2(32'hbaeb9bd7),
	.w3(32'hbabbc127),
	.w4(32'h3c0cf449),
	.w5(32'h3c40704c),
	.w6(32'hbafd5d9c),
	.w7(32'hbbcbb3c8),
	.w8(32'hbb96aed9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e292),
	.w1(32'hbbd66e9e),
	.w2(32'hbb8d5e08),
	.w3(32'h3c267e2d),
	.w4(32'hbc31dbce),
	.w5(32'hbb3e299c),
	.w6(32'hbb97adae),
	.w7(32'hbaf52600),
	.w8(32'hbb9dbb77),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce12d5),
	.w1(32'hbb43b5cd),
	.w2(32'h3c05f9e2),
	.w3(32'h3bd8e35c),
	.w4(32'hbaf60b24),
	.w5(32'h3b65cfab),
	.w6(32'h3b691134),
	.w7(32'hbb79db67),
	.w8(32'hbbadf371),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2360b3),
	.w1(32'h3b405985),
	.w2(32'h3984f354),
	.w3(32'h3c5624e5),
	.w4(32'h3c5fef22),
	.w5(32'h3b10c782),
	.w6(32'h3a8969cd),
	.w7(32'hbbee165d),
	.w8(32'hbba33ef0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a34f5),
	.w1(32'h3b01d830),
	.w2(32'h3b764dcb),
	.w3(32'h39fed6b4),
	.w4(32'h395efb66),
	.w5(32'h3b8d7e59),
	.w6(32'hbc0d1b2a),
	.w7(32'hbb65b5f6),
	.w8(32'hbb102fe0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59b2d2),
	.w1(32'hbb87aa63),
	.w2(32'hbbc15a42),
	.w3(32'hbb599714),
	.w4(32'hbc2b2b63),
	.w5(32'hbc5d3f09),
	.w6(32'hbb1a44d9),
	.w7(32'hbbc08920),
	.w8(32'hbbd2f344),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb672391),
	.w1(32'hbc47d30f),
	.w2(32'hbc28cc8b),
	.w3(32'hba8daef9),
	.w4(32'hbb2f141e),
	.w5(32'h3a14e952),
	.w6(32'hb8ea655a),
	.w7(32'h3bf55163),
	.w8(32'h3c4d3e42),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055a85),
	.w1(32'h3a9b94b1),
	.w2(32'hbb3a0144),
	.w3(32'h3c6ff29f),
	.w4(32'h3b65d578),
	.w5(32'hba6df8ac),
	.w6(32'h3c3ba87c),
	.w7(32'h3b4d74c6),
	.w8(32'hbab91c1a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beefe7b),
	.w1(32'hb9d9e7f6),
	.w2(32'h3bf18491),
	.w3(32'h3b8d36ce),
	.w4(32'hbc941d70),
	.w5(32'hbbe08570),
	.w6(32'h3ba236d5),
	.w7(32'h3bbfcd93),
	.w8(32'h3aebabce),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d3366),
	.w1(32'hbb1d9290),
	.w2(32'h3a891af4),
	.w3(32'h3b54b879),
	.w4(32'hbc1f30ac),
	.w5(32'hbbe2ea5f),
	.w6(32'h3bda2eae),
	.w7(32'hbaa8b25e),
	.w8(32'hbaeb7ba4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fa76c),
	.w1(32'hbb118b47),
	.w2(32'h3b041303),
	.w3(32'h3b0c1eb7),
	.w4(32'hbbcf57cf),
	.w5(32'hbb829354),
	.w6(32'h3b51e4d5),
	.w7(32'h3a4aefd1),
	.w8(32'h3b13809b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6f25),
	.w1(32'hbb2223a6),
	.w2(32'hbc7a7cd7),
	.w3(32'hbac71460),
	.w4(32'h3c1fe925),
	.w5(32'h3c22e8f5),
	.w6(32'hba581802),
	.w7(32'hbc17e379),
	.w8(32'hbb9b27f5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4365e7),
	.w1(32'h3cde152f),
	.w2(32'h3c91ea29),
	.w3(32'h3be51edf),
	.w4(32'h3cbe33be),
	.w5(32'h3cb2a424),
	.w6(32'h3c2fefda),
	.w7(32'h3b9aa011),
	.w8(32'hba844726),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a140),
	.w1(32'h3b82be16),
	.w2(32'hbb97b529),
	.w3(32'h3c0b0f5e),
	.w4(32'hbb4e56bc),
	.w5(32'h3aa079c7),
	.w6(32'h3b6c264c),
	.w7(32'h3b1783f4),
	.w8(32'h3beaa84b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3a0b3),
	.w1(32'h3b890aca),
	.w2(32'h3c255471),
	.w3(32'h3bb7188a),
	.w4(32'h3c4cec2e),
	.w5(32'hb76980e4),
	.w6(32'hbbcee299),
	.w7(32'hb9f1ebc0),
	.w8(32'hbb8829ab),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb979b8),
	.w1(32'h3aeb0112),
	.w2(32'h3a7841fc),
	.w3(32'hbb9359aa),
	.w4(32'h3b813afe),
	.w5(32'h3c0c3268),
	.w6(32'hba45f8b4),
	.w7(32'hbae3a36c),
	.w8(32'hbab4aa30),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee762),
	.w1(32'h3b1e0236),
	.w2(32'hbb002a33),
	.w3(32'h3b7b5dfb),
	.w4(32'hbabc6c71),
	.w5(32'hbb703bc5),
	.w6(32'h3b587c77),
	.w7(32'h3a8006c4),
	.w8(32'h3a7acf12),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdcea9),
	.w1(32'hbb31b699),
	.w2(32'hbbcf8f70),
	.w3(32'h3a3f11b4),
	.w4(32'hbc82ec55),
	.w5(32'hbc4cc355),
	.w6(32'hbb9b29c2),
	.w7(32'hbc766159),
	.w8(32'hbc22e1cb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb773151),
	.w1(32'hbb4d7002),
	.w2(32'hbb741730),
	.w3(32'hbb0bff13),
	.w4(32'h39fb2786),
	.w5(32'h3bbda42a),
	.w6(32'h37b741c2),
	.w7(32'hbbd78a59),
	.w8(32'h3a239c5b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2a3a0),
	.w1(32'h39d79c4d),
	.w2(32'hbad286e6),
	.w3(32'h3b1d2e21),
	.w4(32'h3af8d851),
	.w5(32'hbaa0e8a5),
	.w6(32'h3ac66816),
	.w7(32'h3ae05b32),
	.w8(32'hb9a9f9e6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156c56),
	.w1(32'h3bd5f91c),
	.w2(32'hba8c692a),
	.w3(32'hba114c5f),
	.w4(32'h3c4231d1),
	.w5(32'h3bb58ee2),
	.w6(32'h3b54220d),
	.w7(32'h3b1df72a),
	.w8(32'h3b4fa96f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306157),
	.w1(32'hbc23204a),
	.w2(32'hbbbb0d47),
	.w3(32'hbb35e8ac),
	.w4(32'hbc0c02a7),
	.w5(32'hbbdd215b),
	.w6(32'hba5eeecc),
	.w7(32'hbba10b48),
	.w8(32'hbb8e757a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e5b9),
	.w1(32'hbaa6bdd6),
	.w2(32'hba6fdeb2),
	.w3(32'hbbbc8f37),
	.w4(32'hba6f3d08),
	.w5(32'h3ba8f338),
	.w6(32'hbb45187b),
	.w7(32'h3b1da0d3),
	.w8(32'h3bd20976),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e4c2e),
	.w1(32'h3bac6c1d),
	.w2(32'h3ade1f9a),
	.w3(32'h39b21afc),
	.w4(32'h3b2b29fa),
	.w5(32'hb9aaba9d),
	.w6(32'h3b0f3037),
	.w7(32'h3c07d291),
	.w8(32'h3b8896c1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78b3670),
	.w1(32'h3c6a9764),
	.w2(32'h3c3a4b72),
	.w3(32'h3aeaa42e),
	.w4(32'h3c69b99f),
	.w5(32'h3c465e56),
	.w6(32'h3c130c82),
	.w7(32'h3aa4c93a),
	.w8(32'h3c2cb3d8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47c500),
	.w1(32'h3a3f3ae6),
	.w2(32'h39a54069),
	.w3(32'h3ba4b28d),
	.w4(32'h3c9d24fb),
	.w5(32'h3c4cf3e8),
	.w6(32'hbb80617a),
	.w7(32'h3bda0e6b),
	.w8(32'h3aded402),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2479c),
	.w1(32'h3be76408),
	.w2(32'h3a38e284),
	.w3(32'h3c1c8032),
	.w4(32'h3c2dfb69),
	.w5(32'h3bffb009),
	.w6(32'hb9dd4d94),
	.w7(32'hbb9c7bec),
	.w8(32'hbc0ae62f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b116c33),
	.w1(32'h389580b0),
	.w2(32'hbb53edb9),
	.w3(32'h3ba97226),
	.w4(32'h3a7a8538),
	.w5(32'hbb8da10a),
	.w6(32'h3ab62498),
	.w7(32'hb8419566),
	.w8(32'hbb5a9dae),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1115),
	.w1(32'h3ab8cd05),
	.w2(32'hb9a5a3b9),
	.w3(32'hbaf2b89c),
	.w4(32'h3b66c417),
	.w5(32'h393ab885),
	.w6(32'h396f49a5),
	.w7(32'h3aa201b2),
	.w8(32'hbc007610),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf488b),
	.w1(32'h3be07b56),
	.w2(32'hba15e953),
	.w3(32'hbbead196),
	.w4(32'h3b9095a6),
	.w5(32'hb9b6e2c0),
	.w6(32'h3b8d3903),
	.w7(32'h3a97144b),
	.w8(32'hbb0bdf4d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b661709),
	.w1(32'hba986748),
	.w2(32'hbb9fea34),
	.w3(32'h3b37bb57),
	.w4(32'h3c3af4ea),
	.w5(32'h3b8f36be),
	.w6(32'h3a93f564),
	.w7(32'h3a7f748b),
	.w8(32'h39b46ba5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170446),
	.w1(32'h3a03f7a7),
	.w2(32'h3b2253b5),
	.w3(32'hbba6148c),
	.w4(32'h3bb4098f),
	.w5(32'h3beca6c7),
	.w6(32'h3b8e731f),
	.w7(32'h3a802e6c),
	.w8(32'h3a1d4dc5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae887e8),
	.w1(32'h3b6eaf90),
	.w2(32'hbae7c436),
	.w3(32'h3c6761c2),
	.w4(32'h3c4db2b0),
	.w5(32'h3bbdf2b7),
	.w6(32'h3b3843c1),
	.w7(32'hbab55a67),
	.w8(32'hbabf24e0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b140),
	.w1(32'hbc284fac),
	.w2(32'hbc7509e6),
	.w3(32'hbba031cb),
	.w4(32'hbc2dd9ba),
	.w5(32'hbc2f429c),
	.w6(32'hbacd4948),
	.w7(32'hbb78f305),
	.w8(32'h3ab289eb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7dba0),
	.w1(32'hbb8d6936),
	.w2(32'hbbd25656),
	.w3(32'hbaae05c9),
	.w4(32'hbb27e897),
	.w5(32'hbb8b4bc2),
	.w6(32'hbaf7cbf9),
	.w7(32'hbb2dc3ea),
	.w8(32'hbb5ecf09),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf64fef),
	.w1(32'h3c327024),
	.w2(32'h3b42404d),
	.w3(32'hb9450a8a),
	.w4(32'h3c072aad),
	.w5(32'h3bd077cb),
	.w6(32'h3bafe8c2),
	.w7(32'h39e79096),
	.w8(32'hba1c0dac),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0f02),
	.w1(32'h3bd47f9e),
	.w2(32'hbbb05b6b),
	.w3(32'h3ab6dcd8),
	.w4(32'h3c5ba86a),
	.w5(32'h3cd95526),
	.w6(32'hbb7d806a),
	.w7(32'hba82dbe3),
	.w8(32'h376c644f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfd603),
	.w1(32'hbbcd3b96),
	.w2(32'h3b1fd6c6),
	.w3(32'h3baacbe0),
	.w4(32'hbc0aa1aa),
	.w5(32'hbb6967fc),
	.w6(32'hbc3a0858),
	.w7(32'h39b69239),
	.w8(32'h3c00207d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d9874),
	.w1(32'hbb032540),
	.w2(32'h3af656de),
	.w3(32'hba29904c),
	.w4(32'h3a7784f8),
	.w5(32'hb9608525),
	.w6(32'h3b642e56),
	.w7(32'h3b8be9c4),
	.w8(32'h3b383e1a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53e15a),
	.w1(32'h3be5288e),
	.w2(32'hbbd3b0fa),
	.w3(32'h3b57e8d5),
	.w4(32'hba11126e),
	.w5(32'hbc57f795),
	.w6(32'h3a6476aa),
	.w7(32'hbb8ce6eb),
	.w8(32'hbba2d26a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule