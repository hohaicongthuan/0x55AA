module layer_10_featuremap_134(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3820a672),
	.w1(32'h39c04a19),
	.w2(32'hbaefc04d),
	.w3(32'h3950e94b),
	.w4(32'h39be0d87),
	.w5(32'h39174e2b),
	.w6(32'h3a2e0465),
	.w7(32'h3a346e7e),
	.w8(32'h3a768206),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dc07e),
	.w1(32'hba20f2ac),
	.w2(32'hb9ed2902),
	.w3(32'hb938f1cf),
	.w4(32'hba525f2f),
	.w5(32'hba1bae35),
	.w6(32'hbab46566),
	.w7(32'hba8dc173),
	.w8(32'hba9ab6e3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d1e8e),
	.w1(32'hb986da90),
	.w2(32'hb9784810),
	.w3(32'hb91a5579),
	.w4(32'hb98a4b64),
	.w5(32'hb95656e1),
	.w6(32'hb9eace0f),
	.w7(32'hba06f3c6),
	.w8(32'hb9b6e6a9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3845a5d1),
	.w1(32'h3a1d67f2),
	.w2(32'h38fd2bfb),
	.w3(32'hb88fd0b0),
	.w4(32'h3aa9c499),
	.w5(32'h3a5c2ef7),
	.w6(32'h39682191),
	.w7(32'h3a6c9f12),
	.w8(32'h3a3e0f23),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9d0f9),
	.w1(32'h39e5fbda),
	.w2(32'hb9523a94),
	.w3(32'h39bb38ab),
	.w4(32'h3a3b8cf4),
	.w5(32'hb92ccbbe),
	.w6(32'h3a5642a4),
	.w7(32'h3a25eef5),
	.w8(32'h388e7a64),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38476689),
	.w1(32'hb92d72a2),
	.w2(32'hb962e98f),
	.w3(32'h39b5a647),
	.w4(32'h381ef56c),
	.w5(32'hb91e93ad),
	.w6(32'h38c53d03),
	.w7(32'hb806f9f2),
	.w8(32'h3822b9c8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b379371),
	.w1(32'hba936cab),
	.w2(32'hbb1aaa02),
	.w3(32'h3b667a7c),
	.w4(32'hb9e5e3a0),
	.w5(32'hbb33214e),
	.w6(32'h3afd774a),
	.w7(32'hba4310ba),
	.w8(32'hbb021b8c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9996baa),
	.w1(32'hbafd1241),
	.w2(32'hbb85636f),
	.w3(32'h3ab8716a),
	.w4(32'h3a63b6ff),
	.w5(32'hbadf55b3),
	.w6(32'hbb1558b6),
	.w7(32'hbac8f45f),
	.w8(32'hbaffe50c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9090a),
	.w1(32'h39e155ed),
	.w2(32'hb8946501),
	.w3(32'h39f74bf2),
	.w4(32'h39cff12f),
	.w5(32'h39ab009d),
	.w6(32'h39bd0c2f),
	.w7(32'h3a0b513b),
	.w8(32'h3a02679e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82a34b),
	.w1(32'hbb4d73bf),
	.w2(32'hbb534cb1),
	.w3(32'h3907b6b8),
	.w4(32'hbae6c1b4),
	.w5(32'hbb3d137c),
	.w6(32'hba400af3),
	.w7(32'hbafa27ce),
	.w8(32'hbb2ab68b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86a7ed),
	.w1(32'hba5941fb),
	.w2(32'hba4adeb1),
	.w3(32'hba51eefe),
	.w4(32'hb97d7913),
	.w5(32'hb9868022),
	.w6(32'h380ab5a4),
	.w7(32'hba264bf7),
	.w8(32'hb9336394),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398cb0),
	.w1(32'h3ab03f0c),
	.w2(32'hbb5f5606),
	.w3(32'h3b88b52a),
	.w4(32'h3b29bc49),
	.w5(32'hbb1d1203),
	.w6(32'h3b2f1e5c),
	.w7(32'h3afdf18d),
	.w8(32'hbaeb6cb8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba186fc5),
	.w1(32'hbb258c8f),
	.w2(32'hbb51b4a7),
	.w3(32'h3a5cf6e8),
	.w4(32'hbad586b6),
	.w5(32'hbb214337),
	.w6(32'h391eea05),
	.w7(32'hbb0bd38d),
	.w8(32'hbb1e1f7c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a88c4),
	.w1(32'hbae1b353),
	.w2(32'hbb0e0d40),
	.w3(32'h387f0668),
	.w4(32'hbaa1ecaa),
	.w5(32'hbb02c1db),
	.w6(32'h3a06ffdb),
	.w7(32'hbaa7c457),
	.w8(32'hba988c3b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ccb98),
	.w1(32'h3a4e4de0),
	.w2(32'hba11062f),
	.w3(32'hba4f05a3),
	.w4(32'h3a2e580d),
	.w5(32'h3a882045),
	.w6(32'hb986535e),
	.w7(32'hb8b21fd2),
	.w8(32'hb8e570d6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b00012),
	.w1(32'hbb1a3045),
	.w2(32'hbb5e7c6c),
	.w3(32'h39e9a909),
	.w4(32'hbaca2d6a),
	.w5(32'hbb3e0b58),
	.w6(32'hbaf889a1),
	.w7(32'hbb3184df),
	.w8(32'hbb4d6b44),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d5891),
	.w1(32'hb71f5071),
	.w2(32'hb8a99249),
	.w3(32'h38d7a5db),
	.w4(32'hb8e17435),
	.w5(32'hb98d871a),
	.w6(32'h39704465),
	.w7(32'h395a3840),
	.w8(32'hb95cfb0d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9607e9),
	.w1(32'hbb3507f1),
	.w2(32'hbb89e0f9),
	.w3(32'h3ae25e6c),
	.w4(32'hbb14173b),
	.w5(32'hbb9f2613),
	.w6(32'hb90b4472),
	.w7(32'hbaf1b7ce),
	.w8(32'hbb86a791),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0da4d0),
	.w1(32'hbad559ef),
	.w2(32'hbb0a3627),
	.w3(32'h3a6a7323),
	.w4(32'hbac8e1e9),
	.w5(32'hbb3467e9),
	.w6(32'hba466223),
	.w7(32'hbb08fc70),
	.w8(32'hbb387ea3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368d2744),
	.w1(32'h3994dc66),
	.w2(32'h397c91ba),
	.w3(32'h36fd0e2f),
	.w4(32'h39623415),
	.w5(32'h38c5d19d),
	.w6(32'h397085cc),
	.w7(32'h39333351),
	.w8(32'hb813d1b5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be6664),
	.w1(32'h38fb83cd),
	.w2(32'hb8c206d1),
	.w3(32'h395ef823),
	.w4(32'hb83ad5e4),
	.w5(32'hb9945aa0),
	.w6(32'h386dd359),
	.w7(32'hb8fe7fa5),
	.w8(32'hb7d33d4f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91258f2),
	.w1(32'h3a623d13),
	.w2(32'h398f538b),
	.w3(32'hb906010a),
	.w4(32'h3ac6046e),
	.w5(32'h3a7bc9be),
	.w6(32'hb9ac2df6),
	.w7(32'h395ca774),
	.w8(32'h395130ac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bcc251),
	.w1(32'hbb0cb366),
	.w2(32'hbba23b45),
	.w3(32'h3a93758d),
	.w4(32'h3a8c8335),
	.w5(32'hbb8da0c0),
	.w6(32'h3a5b1f47),
	.w7(32'hba0ae061),
	.w8(32'hbb9ef540),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacafb4f),
	.w1(32'hb930626c),
	.w2(32'hba3582b5),
	.w3(32'hba9cc6a6),
	.w4(32'h37cea17e),
	.w5(32'hb9f1ee56),
	.w6(32'hba8828b5),
	.w7(32'hba505c2d),
	.w8(32'hba634e8c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248e8e),
	.w1(32'h3affdbb3),
	.w2(32'h3b06b4bf),
	.w3(32'hbb740619),
	.w4(32'h39383b50),
	.w5(32'h3ab90f69),
	.w6(32'hbb67babc),
	.w7(32'hba3959c4),
	.w8(32'hba1c6dbb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949a7c9),
	.w1(32'h38e02b95),
	.w2(32'hb9a98347),
	.w3(32'h392dffbd),
	.w4(32'h37fe70e4),
	.w5(32'hb902be48),
	.w6(32'h3937ce0e),
	.w7(32'hb8fec29a),
	.w8(32'hb93389a6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be83aa),
	.w1(32'h3981ff6a),
	.w2(32'h392f84e7),
	.w3(32'hb9b75063),
	.w4(32'h391dbd02),
	.w5(32'h38810d01),
	.w6(32'h39c81f9a),
	.w7(32'h3962720a),
	.w8(32'h38cf400f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109b39),
	.w1(32'h3894372b),
	.w2(32'h3a57eea3),
	.w3(32'hb9db0a76),
	.w4(32'hb8d00e83),
	.w5(32'hb9a4dd3b),
	.w6(32'h3b321a3b),
	.w7(32'h3af41970),
	.w8(32'h3acefccd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a029de5),
	.w1(32'h39f40964),
	.w2(32'hb88fb4d6),
	.w3(32'h3a100a15),
	.w4(32'h3a880ef1),
	.w5(32'hb92ecba1),
	.w6(32'h39968983),
	.w7(32'h39f0529f),
	.w8(32'h3a0918f0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0723ab),
	.w1(32'h3b3df7fb),
	.w2(32'h3b8a6b00),
	.w3(32'hbb3d406b),
	.w4(32'hba383d67),
	.w5(32'h3a98d038),
	.w6(32'hba72cace),
	.w7(32'hb91f9d36),
	.w8(32'h3a917138),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b38d44),
	.w1(32'h3929d2a0),
	.w2(32'h36efc949),
	.w3(32'hba6394be),
	.w4(32'h38b08e86),
	.w5(32'hb78695ba),
	.w6(32'h3993f5bd),
	.w7(32'h385a712c),
	.w8(32'h38b0c7bb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3780ce23),
	.w1(32'h38b1c4d9),
	.w2(32'hb8816421),
	.w3(32'h390ac435),
	.w4(32'h38c13db1),
	.w5(32'h374acd76),
	.w6(32'h398185bb),
	.w7(32'h390f0156),
	.w8(32'h393ae47c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea45ba),
	.w1(32'hb9afc41a),
	.w2(32'hb9f8789b),
	.w3(32'h3a594ad2),
	.w4(32'h37cdbeef),
	.w5(32'hba816fc3),
	.w6(32'hb9e9fa5c),
	.w7(32'h35ca9e04),
	.w8(32'hba5bb196),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20f684),
	.w1(32'h39f0af57),
	.w2(32'hb8de40df),
	.w3(32'hbaa1ab1e),
	.w4(32'hb83f7d1f),
	.w5(32'hb8d283e2),
	.w6(32'hb920eca1),
	.w7(32'hb9e1cc73),
	.w8(32'hba338ea3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b58f8f),
	.w1(32'hba0e0762),
	.w2(32'hb9c979fd),
	.w3(32'h39193fdc),
	.w4(32'hb9527b93),
	.w5(32'hb9d10e1b),
	.w6(32'hb8b95758),
	.w7(32'hb869ec3a),
	.w8(32'hb9a518c3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb7000),
	.w1(32'h3a4087e9),
	.w2(32'hba9734a8),
	.w3(32'h3a95e1fa),
	.w4(32'h3a14bf8d),
	.w5(32'hba9be133),
	.w6(32'h39c3dfc4),
	.w7(32'h38460f10),
	.w8(32'hba811549),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68f654),
	.w1(32'h3b37b227),
	.w2(32'hbc066d6c),
	.w3(32'h3aa31e7a),
	.w4(32'h3b853ace),
	.w5(32'hbba0c6d6),
	.w6(32'hbb62c084),
	.w7(32'hb8137206),
	.w8(32'hbbf23733),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80b793),
	.w1(32'h3bb12375),
	.w2(32'h3b99988c),
	.w3(32'hbb37c77f),
	.w4(32'h3ba5b015),
	.w5(32'h3b9b12d5),
	.w6(32'hbb05b942),
	.w7(32'h3b99c85d),
	.w8(32'h3b4346aa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93eebb),
	.w1(32'h3af64818),
	.w2(32'h3b959d7d),
	.w3(32'hbb49644c),
	.w4(32'h3af94db0),
	.w5(32'h3b8eeeca),
	.w6(32'h3a41d4db),
	.w7(32'h3b91cfce),
	.w8(32'h3bb981b2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853d318),
	.w1(32'h3ac87f8f),
	.w2(32'h3a62b324),
	.w3(32'hb892104a),
	.w4(32'h3ab788f4),
	.w5(32'h3a6c5f0f),
	.w6(32'hb99e3425),
	.w7(32'h3a7a791a),
	.w8(32'h39a77268),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e085a9),
	.w1(32'hba00e451),
	.w2(32'hba127ad5),
	.w3(32'h3897be10),
	.w4(32'hba23502d),
	.w5(32'hba714eb7),
	.w6(32'hba09e083),
	.w7(32'hba116f45),
	.w8(32'hb948ce9f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15e1fa),
	.w1(32'hb8dad989),
	.w2(32'h381c2c0b),
	.w3(32'hba5ab2e1),
	.w4(32'hb8bcaff0),
	.w5(32'hb8989cde),
	.w6(32'hb99c6aa5),
	.w7(32'hb9ec89dc),
	.w8(32'hb95da5f5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9237b15),
	.w1(32'h3932926b),
	.w2(32'h3783eb03),
	.w3(32'hb8e3241d),
	.w4(32'h39c38274),
	.w5(32'h394dfdaf),
	.w6(32'h39c0b7ba),
	.w7(32'h3a158b8c),
	.w8(32'h3a001898),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ed554),
	.w1(32'hbaf835f4),
	.w2(32'hbb4c7af8),
	.w3(32'h3a949456),
	.w4(32'h38bc4c80),
	.w5(32'hbb67b6c0),
	.w6(32'h3a279179),
	.w7(32'hbaea060c),
	.w8(32'hbb7c2bea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b36c3),
	.w1(32'h39a288e8),
	.w2(32'hba049b25),
	.w3(32'hbae883b9),
	.w4(32'hb9380092),
	.w5(32'hb989733e),
	.w6(32'hbac92fdf),
	.w7(32'hb95dcdc6),
	.w8(32'hba656929),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc9fc7),
	.w1(32'hb8f40af8),
	.w2(32'hba2814fc),
	.w3(32'hbaed73db),
	.w4(32'hb9daeecd),
	.w5(32'hba6f8b84),
	.w6(32'hbb02c3f3),
	.w7(32'hbaf25ff0),
	.w8(32'hbb1093c5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144137),
	.w1(32'h39e8e993),
	.w2(32'hb9d79bcb),
	.w3(32'hbabb462a),
	.w4(32'h3a00a99a),
	.w5(32'h3a218f4a),
	.w6(32'hba44c696),
	.w7(32'hb6271267),
	.w8(32'hb98c7399),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b780a25),
	.w1(32'hbb074d12),
	.w2(32'hbbafc313),
	.w3(32'h3b7aeedc),
	.w4(32'hbac37a83),
	.w5(32'hbba9a920),
	.w6(32'hba6b2409),
	.w7(32'hbb70864b),
	.w8(32'hbbafecd8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386deb4d),
	.w1(32'hb79d6bfe),
	.w2(32'hb8c9c4dc),
	.w3(32'hb96ca552),
	.w4(32'h36c8c8d8),
	.w5(32'hb910b10c),
	.w6(32'h396f642d),
	.w7(32'h38bc1de1),
	.w8(32'hb902a62e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9165d23),
	.w1(32'h39de4f1f),
	.w2(32'h38e8894d),
	.w3(32'hb828a27e),
	.w4(32'h3a002141),
	.w5(32'h39cda450),
	.w6(32'h3992ecb9),
	.w7(32'h39043ba0),
	.w8(32'h39b356e3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e2acd),
	.w1(32'hb9b9304c),
	.w2(32'hb9a471ce),
	.w3(32'h39d96937),
	.w4(32'hb9c9d357),
	.w5(32'hb999739e),
	.w6(32'hb9342338),
	.w7(32'hb9caf059),
	.w8(32'hb9b89aa8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f893),
	.w1(32'hb9e850c7),
	.w2(32'h3a3a9d5b),
	.w3(32'hba445ec1),
	.w4(32'h3884e708),
	.w5(32'h38182f73),
	.w6(32'hb9e173ba),
	.w7(32'hba45bdc2),
	.w8(32'hba76aa11),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad79acc),
	.w1(32'hb9fafcc1),
	.w2(32'hba975c03),
	.w3(32'h3a19c644),
	.w4(32'hba2faaa1),
	.w5(32'hba8f9c89),
	.w6(32'hb8f3aef6),
	.w7(32'hba4f7a1f),
	.w8(32'hba1fe749),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2ce30),
	.w1(32'hbb0e82d4),
	.w2(32'hbb77fb11),
	.w3(32'h3b471e1a),
	.w4(32'hb94802bf),
	.w5(32'hbb8bc8e3),
	.w6(32'h3a82c538),
	.w7(32'hba9278e4),
	.w8(32'hbb6b71db),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1f621),
	.w1(32'hb902a214),
	.w2(32'hba57371b),
	.w3(32'hb8ac6f51),
	.w4(32'hb9e155a0),
	.w5(32'hba845b94),
	.w6(32'h381110e9),
	.w7(32'hb9e3154c),
	.w8(32'hba8a89e6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7ed09),
	.w1(32'hb87aa670),
	.w2(32'h382acbef),
	.w3(32'hb95c32d3),
	.w4(32'hb9a6b3c8),
	.w5(32'hba248bee),
	.w6(32'hba006225),
	.w7(32'hb948deb7),
	.w8(32'hb971d0a9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f48708),
	.w1(32'hba174529),
	.w2(32'hba331a0b),
	.w3(32'hba0ec349),
	.w4(32'hba582a25),
	.w5(32'hba6a2bd4),
	.w6(32'hba172d88),
	.w7(32'hba6fffd3),
	.w8(32'hba7613de),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b1f4d),
	.w1(32'h3a164f3f),
	.w2(32'h39cb5e55),
	.w3(32'hba90c02b),
	.w4(32'h3a41f431),
	.w5(32'h39d7a248),
	.w6(32'h3a23f48d),
	.w7(32'h39f85b4e),
	.w8(32'h39a80e73),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b6843),
	.w1(32'h398142f6),
	.w2(32'h3884e572),
	.w3(32'h3a1eedf3),
	.w4(32'h3a186d15),
	.w5(32'h39b5900d),
	.w6(32'h38d128ec),
	.w7(32'h39db920c),
	.w8(32'h39c1d39e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98386a7),
	.w1(32'hb7daa340),
	.w2(32'hb93597ba),
	.w3(32'h3911db5c),
	.w4(32'h393c6eeb),
	.w5(32'hb91ddea4),
	.w6(32'h376a8948),
	.w7(32'hb979d60d),
	.w8(32'hb779520a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06df7c),
	.w1(32'hbae2afe1),
	.w2(32'hbb15d94d),
	.w3(32'hb9b89803),
	.w4(32'hbaae344d),
	.w5(32'hbb0f5e3a),
	.w6(32'hbaa76ad4),
	.w7(32'hbab17ece),
	.w8(32'hbae5621c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba601b56),
	.w1(32'hb9f07111),
	.w2(32'hbb0c236d),
	.w3(32'h3929c5ad),
	.w4(32'h3a25567b),
	.w5(32'hbb156d9e),
	.w6(32'h3a8865c4),
	.w7(32'hb92f07ed),
	.w8(32'hbaa70bbe),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f75c7),
	.w1(32'h38124a61),
	.w2(32'hb9489531),
	.w3(32'h39abbccb),
	.w4(32'h389e5b5f),
	.w5(32'h3935a187),
	.w6(32'hb9624fc6),
	.w7(32'h3909cde7),
	.w8(32'hb7b956b0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c15d99),
	.w1(32'hb900f21c),
	.w2(32'hb8b6b849),
	.w3(32'h37e7bb59),
	.w4(32'h391b7936),
	.w5(32'h38121379),
	.w6(32'h3932cf5e),
	.w7(32'h38ad8fd0),
	.w8(32'hb7612c6c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f0a5f),
	.w1(32'hb7d56efd),
	.w2(32'hb90c8b88),
	.w3(32'hb78cfc2a),
	.w4(32'h38ca99c2),
	.w5(32'hb86bea3b),
	.w6(32'hb806c016),
	.w7(32'hb7ace5cf),
	.w8(32'h38dba755),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d831ed),
	.w1(32'hb924e316),
	.w2(32'h397dda8c),
	.w3(32'h38099d51),
	.w4(32'h399ceed7),
	.w5(32'hb9aa010e),
	.w6(32'hb907e938),
	.w7(32'hb9d64c1f),
	.w8(32'hb92dc51f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a774fbe),
	.w1(32'hbbbdb7c6),
	.w2(32'hbbd7ab63),
	.w3(32'h3b94d315),
	.w4(32'hbae46678),
	.w5(32'hbbde6299),
	.w6(32'h399f3178),
	.w7(32'hbb2f9fcb),
	.w8(32'hbb54b4bb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7976),
	.w1(32'h39db7da9),
	.w2(32'hbb773b62),
	.w3(32'hbb00fa51),
	.w4(32'hba7d10e6),
	.w5(32'hbb5f66f8),
	.w6(32'hbb4da81c),
	.w7(32'hbb85ce2a),
	.w8(32'hbba0d8d6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97d5153),
	.w1(32'hbaa95e86),
	.w2(32'hbb2a5fb1),
	.w3(32'hb9d03a76),
	.w4(32'hbaa2d54d),
	.w5(32'hbb33595a),
	.w6(32'h39a99924),
	.w7(32'hbaa9206a),
	.w8(32'hbb421d74),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93cd89),
	.w1(32'h3b1d9c07),
	.w2(32'h3b2fbfa8),
	.w3(32'hbbb1a896),
	.w4(32'h3a8f1580),
	.w5(32'h3b0138cc),
	.w6(32'hbba9b793),
	.w7(32'hba4e64f1),
	.w8(32'hb9d2cd85),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e961d),
	.w1(32'hb9711415),
	.w2(32'hb8a2f125),
	.w3(32'hb7f77d48),
	.w4(32'hb9a710db),
	.w5(32'hb8a8fb89),
	.w6(32'hb88d0f20),
	.w7(32'hb8c17b86),
	.w8(32'hb961554f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c7172),
	.w1(32'h3964e17c),
	.w2(32'hb76a0376),
	.w3(32'hb93779ff),
	.w4(32'h39700740),
	.w5(32'h38911e0a),
	.w6(32'h39945947),
	.w7(32'hb60f900e),
	.w8(32'h3919340b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379068e9),
	.w1(32'h394902aa),
	.w2(32'hb82c5a03),
	.w3(32'h38def7e4),
	.w4(32'h39933dea),
	.w5(32'h393e2e01),
	.w6(32'h39228882),
	.w7(32'h37dd6299),
	.w8(32'h39302a95),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2bbd4),
	.w1(32'hb9308fd2),
	.w2(32'hba9155d6),
	.w3(32'h3a09c8b0),
	.w4(32'h37250717),
	.w5(32'hba592bb4),
	.w6(32'h39bd9cb8),
	.w7(32'hb897233b),
	.w8(32'hba05a47c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0b2be),
	.w1(32'hb990ba8c),
	.w2(32'hb8dfdf2d),
	.w3(32'h399367a4),
	.w4(32'hb9238b36),
	.w5(32'hb9443d08),
	.w6(32'hb9036811),
	.w7(32'hb9302cb3),
	.w8(32'h3875349a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82a556),
	.w1(32'hb905f497),
	.w2(32'hba23ba24),
	.w3(32'h3aee1003),
	.w4(32'h3a00c570),
	.w5(32'hba515adb),
	.w6(32'hb8a7fe4e),
	.w7(32'h39c909c1),
	.w8(32'hbae3b12f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bb14a),
	.w1(32'h3a4dc9af),
	.w2(32'hbb82983b),
	.w3(32'h3ad6a759),
	.w4(32'h3ae64760),
	.w5(32'hbb3a520a),
	.w6(32'hba27991b),
	.w7(32'hb9c8a13d),
	.w8(32'hbb1fb906),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fc983),
	.w1(32'hba0077ab),
	.w2(32'h366d49a3),
	.w3(32'hbb15447f),
	.w4(32'hba8e9c82),
	.w5(32'hb9f51bd5),
	.w6(32'hbb2c7c83),
	.w7(32'hba841220),
	.w8(32'hbaa60530),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb7496),
	.w1(32'hbab8c067),
	.w2(32'hbb3f7f51),
	.w3(32'h389d3d4d),
	.w4(32'hba952e61),
	.w5(32'hbb1da026),
	.w6(32'h386ef2f7),
	.w7(32'hbab25718),
	.w8(32'hbb0ee78e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4864bc),
	.w1(32'hba0f77dc),
	.w2(32'hbafe3dce),
	.w3(32'h3b0026e2),
	.w4(32'h39dc537a),
	.w5(32'hbb0b503a),
	.w6(32'h3aa0714d),
	.w7(32'hba01c697),
	.w8(32'hba4f9385),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5566d6),
	.w1(32'hba0872f2),
	.w2(32'hbaa7ea12),
	.w3(32'hb9b950b2),
	.w4(32'hb9a3fcbd),
	.w5(32'hbaaa9463),
	.w6(32'hba3c3582),
	.w7(32'hba9e4f55),
	.w8(32'hba8f7188),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31aced),
	.w1(32'hba5153df),
	.w2(32'hbaec38d8),
	.w3(32'h39f0d43e),
	.w4(32'hb9aa36ce),
	.w5(32'hbacd8e24),
	.w6(32'hb9d149e0),
	.w7(32'hba720be8),
	.w8(32'hbabcd3ec),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90dae2a),
	.w1(32'hb9bc7c75),
	.w2(32'hb9a1b22d),
	.w3(32'hb909bdc0),
	.w4(32'hb9951273),
	.w5(32'hb9e3fe8b),
	.w6(32'hb9ac631e),
	.w7(32'hb9f20ead),
	.w8(32'hb98ec83e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bec20),
	.w1(32'hb901b554),
	.w2(32'hb8c3ef1a),
	.w3(32'hb9bedf06),
	.w4(32'hb84348fc),
	.w5(32'hb80b48d7),
	.w6(32'hb83ea789),
	.w7(32'h390deac5),
	.w8(32'h38f9ee51),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e14afe),
	.w1(32'h39cc098b),
	.w2(32'hb985546a),
	.w3(32'h3912055b),
	.w4(32'h38f3df02),
	.w5(32'h382085bc),
	.w6(32'h396c0cea),
	.w7(32'hb899ee26),
	.w8(32'hb98b6fff),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cb1f8),
	.w1(32'hb95f7f63),
	.w2(32'h39e6f5ba),
	.w3(32'hba1914bc),
	.w4(32'hb9d86c0f),
	.w5(32'hb8df53fc),
	.w6(32'hba89e54b),
	.w7(32'hb97ac536),
	.w8(32'hb8e8e277),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef5689),
	.w1(32'h3a23d38e),
	.w2(32'hb9603128),
	.w3(32'hbaccd75f),
	.w4(32'h3a30ef26),
	.w5(32'h38c8477a),
	.w6(32'hba86cd15),
	.w7(32'h3a017ed6),
	.w8(32'hbabe4107),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d8820),
	.w1(32'h3a083ff1),
	.w2(32'h3973a02b),
	.w3(32'hb8f1c194),
	.w4(32'h39c323c5),
	.w5(32'h38dbc6f3),
	.w6(32'h391948e9),
	.w7(32'h39d623db),
	.w8(32'h39aaf0f4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89da3db),
	.w1(32'h3a476498),
	.w2(32'hb8b532c0),
	.w3(32'hbaf6cf05),
	.w4(32'hba1f1ab8),
	.w5(32'hba069e48),
	.w6(32'hbb009150),
	.w7(32'hba9ee82b),
	.w8(32'hbadad951),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae923b9),
	.w1(32'hba692305),
	.w2(32'hbb694394),
	.w3(32'h3ace6e66),
	.w4(32'h37d7dd15),
	.w5(32'hbb304b36),
	.w6(32'h39422c9b),
	.w7(32'hba830a18),
	.w8(32'hbb1d73f0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ac378),
	.w1(32'h3ac327ec),
	.w2(32'h3b32677f),
	.w3(32'hbaa19a64),
	.w4(32'h3af92e9f),
	.w5(32'h3b26d569),
	.w6(32'h3a7af7ea),
	.w7(32'h3b778023),
	.w8(32'h3b648034),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01fe5e),
	.w1(32'hbad2aeba),
	.w2(32'hbbc6986d),
	.w3(32'h3b523ac2),
	.w4(32'h3a51e093),
	.w5(32'hbb961706),
	.w6(32'h3b0ec8c5),
	.w7(32'hb97db07a),
	.w8(32'hbb48d423),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa51c59),
	.w1(32'h3acfe09e),
	.w2(32'h3ae44bf6),
	.w3(32'hbaa5c43f),
	.w4(32'h3ad8481d),
	.w5(32'h3aa1c8b1),
	.w6(32'hba39b7f5),
	.w7(32'h3ad11776),
	.w8(32'h3a9a80d6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69a575),
	.w1(32'hbb400716),
	.w2(32'hbba717c4),
	.w3(32'h3951ae93),
	.w4(32'hbb45fe14),
	.w5(32'hbba96ec5),
	.w6(32'hba86c72f),
	.w7(32'hbb5ea511),
	.w8(32'hbb714348),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eecadc),
	.w1(32'hba2e3c89),
	.w2(32'hba924977),
	.w3(32'h39e4762b),
	.w4(32'hba26a664),
	.w5(32'hba6443cf),
	.w6(32'h39270ec1),
	.w7(32'hba68c251),
	.w8(32'hba8bd2dd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26a307),
	.w1(32'h3b0adeeb),
	.w2(32'h3b461e51),
	.w3(32'hbb0db53b),
	.w4(32'h3a808b04),
	.w5(32'h3abb4df9),
	.w6(32'hb9329d72),
	.w7(32'h3ade49c7),
	.w8(32'h3acdf4e8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a1071),
	.w1(32'h3a1498df),
	.w2(32'h395e57a7),
	.w3(32'h381e054c),
	.w4(32'h39e49fdc),
	.w5(32'h38ce7f15),
	.w6(32'h39a4dbf7),
	.w7(32'h37dc6b7e),
	.w8(32'hb8f71814),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39084591),
	.w1(32'hbab77e1a),
	.w2(32'hbb4ac969),
	.w3(32'h3a14cf8a),
	.w4(32'hbaa41c44),
	.w5(32'hbb3a64ad),
	.w6(32'hba28b21f),
	.w7(32'hbb1e6655),
	.w8(32'hbb301c7a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed4760),
	.w1(32'hbaf0472f),
	.w2(32'hbb8fc083),
	.w3(32'h3b5b02e7),
	.w4(32'h3a3e83c1),
	.w5(32'hbb426c55),
	.w6(32'h3b4eb89c),
	.w7(32'h3a6572a3),
	.w8(32'hbaf0cf44),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ae51),
	.w1(32'h3b78cd08),
	.w2(32'hbbb3e91a),
	.w3(32'hba441ef5),
	.w4(32'h3b544ccd),
	.w5(32'hbb90a425),
	.w6(32'hbbb55506),
	.w7(32'hba1e0f85),
	.w8(32'hbbe55dc9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec52a5),
	.w1(32'h3bc402c0),
	.w2(32'h3b86e3e2),
	.w3(32'hb9bec923),
	.w4(32'h3bdd95c8),
	.w5(32'h3ba04006),
	.w6(32'h3b3cd98d),
	.w7(32'h3bf06939),
	.w8(32'h3bbc72c1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97568b),
	.w1(32'h3abfa964),
	.w2(32'h3b2989ad),
	.w3(32'hbb129e5f),
	.w4(32'h39f0b26a),
	.w5(32'h3a2b1c15),
	.w6(32'hbb07f6a8),
	.w7(32'hba8f1acd),
	.w8(32'hba6b7efd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020a13),
	.w1(32'hb900b488),
	.w2(32'hbbce9643),
	.w3(32'h3b16e7ed),
	.w4(32'h3acbbbad),
	.w5(32'hbb98677a),
	.w6(32'h3aa54072),
	.w7(32'h3969ca18),
	.w8(32'hbb83b01d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a28b1),
	.w1(32'h390e7a9f),
	.w2(32'hb99a839a),
	.w3(32'h3a30eac1),
	.w4(32'h38466d29),
	.w5(32'hb985f22b),
	.w6(32'h393469e5),
	.w7(32'hb803a248),
	.w8(32'hb8406fa4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46f38),
	.w1(32'hba827946),
	.w2(32'hbbc2cd3f),
	.w3(32'hbb3d4797),
	.w4(32'h3afca94c),
	.w5(32'hbb23560c),
	.w6(32'hbb88a9bd),
	.w7(32'hb97f9233),
	.w8(32'hbba8785e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a621b80),
	.w1(32'h3a812cb1),
	.w2(32'hbb1b50a6),
	.w3(32'h3b1ce0b0),
	.w4(32'h3aea113b),
	.w5(32'hbaa19c07),
	.w6(32'h3b0d2751),
	.w7(32'h3af5627c),
	.w8(32'hbab0aacf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3606853f),
	.w1(32'hb9c9deb9),
	.w2(32'hb9f73c0d),
	.w3(32'hb857ebed),
	.w4(32'hb9c89d20),
	.w5(32'hb94d9882),
	.w6(32'hb9e4fbaf),
	.w7(32'hb991e551),
	.w8(32'hb968bb16),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ef61e),
	.w1(32'hb9b688f6),
	.w2(32'hba2b6fc9),
	.w3(32'hb9329be3),
	.w4(32'h37926c5e),
	.w5(32'hba2a41e9),
	.w6(32'hba3b3726),
	.w7(32'hba87a5ab),
	.w8(32'hbabe901a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5817d),
	.w1(32'hb9ebf47a),
	.w2(32'hbb061c7d),
	.w3(32'h39d2a851),
	.w4(32'hb9a02d81),
	.w5(32'hbafabba9),
	.w6(32'hb97d3318),
	.w7(32'hbacf8a8b),
	.w8(32'hbb10a6bb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba088f21),
	.w1(32'h3a869d70),
	.w2(32'h3a3b6ac0),
	.w3(32'hba897383),
	.w4(32'h3992cd02),
	.w5(32'h39ea23b7),
	.w6(32'hbadfbd2c),
	.w7(32'h38e1f0a2),
	.w8(32'hb8b5be65),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e762),
	.w1(32'h3a36bfdd),
	.w2(32'h3ada7669),
	.w3(32'hbaa62bc0),
	.w4(32'h3a9bdb92),
	.w5(32'h3b1d8608),
	.w6(32'h3a0f44ca),
	.w7(32'h3b11d795),
	.w8(32'h3b2a9d74),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf7e23),
	.w1(32'hba0bcdf9),
	.w2(32'hba7e7bd6),
	.w3(32'hba84d894),
	.w4(32'hb6f1a798),
	.w5(32'hb71a3ebb),
	.w6(32'hba9c4baf),
	.w7(32'hb7b9be64),
	.w8(32'h39a2a3e3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f8a7),
	.w1(32'h3b615fce),
	.w2(32'h3a84ece1),
	.w3(32'hba311e10),
	.w4(32'h3abe3409),
	.w5(32'h399f87e6),
	.w6(32'hbadcf7ca),
	.w7(32'hba34da16),
	.w8(32'hba9ce3c2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1f0e3),
	.w1(32'hbb783a73),
	.w2(32'hbb6a8a06),
	.w3(32'hba358583),
	.w4(32'hbb39ca8f),
	.w5(32'hbb400e44),
	.w6(32'hbadfb2a6),
	.w7(32'hbb52fb43),
	.w8(32'hbb50e3b7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c57813),
	.w1(32'h3a3aecb7),
	.w2(32'h39a31427),
	.w3(32'hb9d682b9),
	.w4(32'h38d822a2),
	.w5(32'hb93a347c),
	.w6(32'hb985f8a5),
	.w7(32'h3964d96b),
	.w8(32'hb9c23ee2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4e0bf),
	.w1(32'h39d484e4),
	.w2(32'h374ba256),
	.w3(32'h38d9f8ff),
	.w4(32'h3a3b3f28),
	.w5(32'h39894e6a),
	.w6(32'h3a2d966d),
	.w7(32'h399ad4f1),
	.w8(32'h3a04fe7b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d28baa),
	.w1(32'hb875a049),
	.w2(32'hba285fef),
	.w3(32'h3a56b3e3),
	.w4(32'hb7d7dcd6),
	.w5(32'hb9f37428),
	.w6(32'h38ca6a8e),
	.w7(32'hb9c71ef0),
	.w8(32'hb9afa0d5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39040186),
	.w1(32'h392bc582),
	.w2(32'hb8902bb0),
	.w3(32'h39a400c0),
	.w4(32'h399ddec6),
	.w5(32'h379661d6),
	.w6(32'h39b406b1),
	.w7(32'h38d5c0c0),
	.w8(32'h396e3e0d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8587c04),
	.w1(32'hb9503b14),
	.w2(32'hba1c2b99),
	.w3(32'h392f5f4c),
	.w4(32'h39cdeab7),
	.w5(32'h38502bd4),
	.w6(32'h39bda95e),
	.w7(32'h3903e4e2),
	.w8(32'h3a1b4cf4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6811f8),
	.w1(32'h39fdf031),
	.w2(32'h39686a4b),
	.w3(32'hba2561c5),
	.w4(32'hb898d693),
	.w5(32'hb8a11849),
	.w6(32'hba856660),
	.w7(32'hba476daf),
	.w8(32'hba3a7174),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a773d9),
	.w1(32'hb99805cf),
	.w2(32'hba09e6ef),
	.w3(32'hb9a59c00),
	.w4(32'hb9805111),
	.w5(32'hb9d77b5e),
	.w6(32'hb89c8f10),
	.w7(32'hb986a957),
	.w8(32'hb9be8db6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1dde6),
	.w1(32'hba561292),
	.w2(32'hbb1fcb36),
	.w3(32'h3a456c32),
	.w4(32'hba28af49),
	.w5(32'hbad5e6d7),
	.w6(32'h38c504d4),
	.w7(32'hba8eb599),
	.w8(32'hbac6bc1e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2192ca),
	.w1(32'h3aa82b0d),
	.w2(32'h3aab5c70),
	.w3(32'hbb25839b),
	.w4(32'h39c59e2e),
	.w5(32'h3a9b943c),
	.w6(32'hbab91a90),
	.w7(32'hb9acb119),
	.w8(32'hba14ca41),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39878f43),
	.w1(32'h3a1a3481),
	.w2(32'h3a2f6730),
	.w3(32'h39c4ffd2),
	.w4(32'h3a4ae313),
	.w5(32'h39a426ce),
	.w6(32'h3a1dfc2b),
	.w7(32'h3a63da88),
	.w8(32'h3a34bd13),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d249e),
	.w1(32'hb9b4cf4e),
	.w2(32'hb9e732fa),
	.w3(32'h39a8442e),
	.w4(32'hb9d6be66),
	.w5(32'hba3fd74c),
	.w6(32'hb5fe1ea9),
	.w7(32'hb918e188),
	.w8(32'hb9725401),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dac14d),
	.w1(32'h38d5105e),
	.w2(32'hb8925640),
	.w3(32'hba01296f),
	.w4(32'h39258712),
	.w5(32'hb8855223),
	.w6(32'h397f8f9b),
	.w7(32'hb8858842),
	.w8(32'hb809417a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38283007),
	.w1(32'hb8fee7cb),
	.w2(32'hb7d69339),
	.w3(32'h38e1a458),
	.w4(32'hb9512b54),
	.w5(32'hb6b6ccd5),
	.w6(32'hb8d55bc8),
	.w7(32'hb994606d),
	.w8(32'hb863926d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8a33a),
	.w1(32'h3b2bfb3a),
	.w2(32'hbab2892c),
	.w3(32'h3ab700a6),
	.w4(32'hbaa6c5dc),
	.w5(32'hbb46897a),
	.w6(32'hba65ed2a),
	.w7(32'hbb0dde18),
	.w8(32'hbb34c8d2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9694eb),
	.w1(32'hbae95358),
	.w2(32'hbb150700),
	.w3(32'h3af626a0),
	.w4(32'hba45ac37),
	.w5(32'hbb1c0d98),
	.w6(32'hb9e0a511),
	.w7(32'hbadaf807),
	.w8(32'hbafc26f6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15815a),
	.w1(32'hb79aae7b),
	.w2(32'hba11db01),
	.w3(32'h3a275896),
	.w4(32'h3973d13e),
	.w5(32'hb9b5d400),
	.w6(32'h39f9c548),
	.w7(32'h3958b411),
	.w8(32'hb96844d5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb62b5),
	.w1(32'hba24f60e),
	.w2(32'hbab1d045),
	.w3(32'h38c45be5),
	.w4(32'hb9c8f8c2),
	.w5(32'hba399da6),
	.w6(32'hb9d6404f),
	.w7(32'hba3e73b4),
	.w8(32'hbaa09e11),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0de77),
	.w1(32'h3981cb76),
	.w2(32'hb81e9d00),
	.w3(32'hb98b1975),
	.w4(32'h393a7b70),
	.w5(32'hb9208ea9),
	.w6(32'hb91c1c8e),
	.w7(32'h39349f0f),
	.w8(32'hb9885960),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70cfdd4),
	.w1(32'hb9e533df),
	.w2(32'hbaafbbdb),
	.w3(32'h3982540b),
	.w4(32'hb9a2b8ee),
	.w5(32'hba8977b2),
	.w6(32'hb96a4791),
	.w7(32'hba5e6da0),
	.w8(32'hba9c0901),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e0268),
	.w1(32'hba826532),
	.w2(32'hbabc463f),
	.w3(32'hb86dc24e),
	.w4(32'hba3e7aa0),
	.w5(32'hbac9bb6e),
	.w6(32'hba0a4ba0),
	.w7(32'hba85f61c),
	.w8(32'hbab3e138),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab53ff8),
	.w1(32'hbb0c9367),
	.w2(32'hbb6f4a6f),
	.w3(32'h3b5361e4),
	.w4(32'hb99e85c9),
	.w5(32'hbb5519ec),
	.w6(32'h3a5b393f),
	.w7(32'hbaddb268),
	.w8(32'hbb291359),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba702732),
	.w1(32'h3aa3e221),
	.w2(32'h3aad26bf),
	.w3(32'hbaa271e6),
	.w4(32'h3a1b75e4),
	.w5(32'h3a3f9dfd),
	.w6(32'hba6d1986),
	.w7(32'h39ae766f),
	.w8(32'hb8a4a29b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a50593),
	.w1(32'hba64a964),
	.w2(32'hbad4af3f),
	.w3(32'h3a974660),
	.w4(32'hb92ac9a8),
	.w5(32'hba8b78b1),
	.w6(32'h39a4f344),
	.w7(32'hba91b8f6),
	.w8(32'hbaaf7e23),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc5f52),
	.w1(32'hba790b04),
	.w2(32'hbb374e6c),
	.w3(32'h3b1ff539),
	.w4(32'hb6cd8f03),
	.w5(32'hbb1c2fee),
	.w6(32'h3acd29c2),
	.w7(32'hb9b572b7),
	.w8(32'hbb048339),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb5726),
	.w1(32'h3ab78d60),
	.w2(32'h3a03a7d4),
	.w3(32'hba779714),
	.w4(32'h3a1cf636),
	.w5(32'h38dc58c6),
	.w6(32'hbab45f5c),
	.w7(32'hba29a2bf),
	.w8(32'hba9be938),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41e9bc),
	.w1(32'hbaaeb92b),
	.w2(32'hbb180ed1),
	.w3(32'h3aaa5739),
	.w4(32'hba228780),
	.w5(32'hbb0bc1fc),
	.w6(32'hb815c0bc),
	.w7(32'hbab07f06),
	.w8(32'hbafb9d38),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a63952),
	.w1(32'hb89a7d51),
	.w2(32'hb90acfb9),
	.w3(32'hb9a0fe8e),
	.w4(32'hb8d892a5),
	.w5(32'hb954cdff),
	.w6(32'hb9b86a59),
	.w7(32'hb96c09a1),
	.w8(32'hb9bd43e9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec5a9),
	.w1(32'h3b714d3f),
	.w2(32'h3bba747a),
	.w3(32'hbb454cd8),
	.w4(32'h3ad1b4be),
	.w5(32'h3b5d4701),
	.w6(32'h3a08e89c),
	.w7(32'h3b480b3f),
	.w8(32'h3b3520d1),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a952b3),
	.w1(32'h3910ad13),
	.w2(32'hb997b1a8),
	.w3(32'h398b6a45),
	.w4(32'hb884faea),
	.w5(32'hb9fc2e13),
	.w6(32'hb85e6743),
	.w7(32'h395cc1de),
	.w8(32'hb9aed756),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831b337),
	.w1(32'hb6d12586),
	.w2(32'hb81cf80d),
	.w3(32'h384ae935),
	.w4(32'hb721f2e2),
	.w5(32'hb888fd9d),
	.w6(32'h3859f735),
	.w7(32'hb784d7a3),
	.w8(32'hb7c0f0ab),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce0a9c),
	.w1(32'h36e9816c),
	.w2(32'h386667b1),
	.w3(32'hb75c57ce),
	.w4(32'h3783b275),
	.w5(32'h38803d92),
	.w6(32'h38159cf8),
	.w7(32'h37f51d41),
	.w8(32'h386801f0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39325309),
	.w1(32'h392eba65),
	.w2(32'hb9db5723),
	.w3(32'h3a0d33b6),
	.w4(32'h39d89af7),
	.w5(32'hb7d872d0),
	.w6(32'h39a131f3),
	.w7(32'h3a4f1859),
	.w8(32'h39d3b053),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab496f6),
	.w1(32'h39b32491),
	.w2(32'hb8aa0789),
	.w3(32'hba7405d9),
	.w4(32'h39a0acc4),
	.w5(32'h3a182f83),
	.w6(32'hba70028d),
	.w7(32'h39daec72),
	.w8(32'hb984de21),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2adcc),
	.w1(32'hbaec0cca),
	.w2(32'hbb1bf3a3),
	.w3(32'hbab29b73),
	.w4(32'hbaa83044),
	.w5(32'hbadfc9cf),
	.w6(32'hba67a7a7),
	.w7(32'hba56113e),
	.w8(32'hbaa8ac9a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ca3ea6),
	.w1(32'hb6cbf0b7),
	.w2(32'hb68162af),
	.w3(32'hb6b26323),
	.w4(32'hb6f0572a),
	.w5(32'hb59f1444),
	.w6(32'hb53a4aaa),
	.w7(32'hb734eb13),
	.w8(32'hb5bf9ec4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99108c4),
	.w1(32'hbadfaa3a),
	.w2(32'hbb1fec50),
	.w3(32'h38f2bb90),
	.w4(32'hba95b2d6),
	.w5(32'hbafa9d8c),
	.w6(32'hba3989f7),
	.w7(32'hbad9b255),
	.w8(32'hbb07549c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9954ccc),
	.w1(32'hb79b05e2),
	.w2(32'hb776ab89),
	.w3(32'hba027441),
	.w4(32'hba00e08f),
	.w5(32'hb96e6732),
	.w6(32'hba8e186e),
	.w7(32'hba8af8a7),
	.w8(32'hba5b96a7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b7fb),
	.w1(32'hb9590bfa),
	.w2(32'hbb751c43),
	.w3(32'h3aef3172),
	.w4(32'hb903e09b),
	.w5(32'hbb4e2cb8),
	.w6(32'h3a588fde),
	.w7(32'hbaa2f653),
	.w8(32'hbb2ba6b5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb584a49),
	.w1(32'h3a30d6e2),
	.w2(32'h3a177ce7),
	.w3(32'hbaed087a),
	.w4(32'hb8b74767),
	.w5(32'h3a24a8f5),
	.w6(32'hb9f5becd),
	.w7(32'h394645bd),
	.w8(32'h39305080),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169295),
	.w1(32'h39bd1f43),
	.w2(32'hb9f47e09),
	.w3(32'h3999383e),
	.w4(32'h381a714e),
	.w5(32'hba55437b),
	.w6(32'h393e3481),
	.w7(32'hb93de771),
	.w8(32'hba839375),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0d279),
	.w1(32'h384dfb58),
	.w2(32'hb8fbd737),
	.w3(32'hb9998270),
	.w4(32'hb8e2e4a6),
	.w5(32'hb8e52298),
	.w6(32'hb903b406),
	.w7(32'hb8635e2d),
	.w8(32'hb82b2cee),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60f096),
	.w1(32'h3a8e78cd),
	.w2(32'h3a8885a6),
	.w3(32'hba8d5e59),
	.w4(32'h3a1fa520),
	.w5(32'h3a50617e),
	.w6(32'hba7713f5),
	.w7(32'h3859fd84),
	.w8(32'h389d1dcb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979bf70),
	.w1(32'h3aad316f),
	.w2(32'h386b3ff5),
	.w3(32'h3a4b4962),
	.w4(32'h3adbf877),
	.w5(32'h39438e44),
	.w6(32'h3acbee97),
	.w7(32'h3b06533c),
	.w8(32'hb7adc23b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc0543),
	.w1(32'h3ae78ab5),
	.w2(32'h3aa77526),
	.w3(32'hb9ee2a70),
	.w4(32'h3abeb51b),
	.w5(32'h3a96e3ec),
	.w6(32'hb9a80daa),
	.w7(32'h3aa7b61c),
	.w8(32'h3a27a308),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39138f),
	.w1(32'hb91f591a),
	.w2(32'hba7df6d4),
	.w3(32'h39ea4a65),
	.w4(32'h366e5882),
	.w5(32'hb9f42740),
	.w6(32'h394efc49),
	.w7(32'hb8bf429e),
	.w8(32'hba1f9f8e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38167c82),
	.w1(32'hb93e6fc0),
	.w2(32'hb95db990),
	.w3(32'hb8d4f54c),
	.w4(32'hb92b004c),
	.w5(32'hb93930ef),
	.w6(32'hb9131abc),
	.w7(32'hb98114ea),
	.w8(32'hb95e2bb8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf31c),
	.w1(32'hba9029da),
	.w2(32'hbb10504c),
	.w3(32'h3acd4b79),
	.w4(32'hb9831bb7),
	.w5(32'hbb0dba90),
	.w6(32'hb797bbb8),
	.w7(32'hba4faad4),
	.w8(32'hbac9ba1a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c100a1),
	.w1(32'h3984fbcc),
	.w2(32'hb9ee9db1),
	.w3(32'h3a116c5a),
	.w4(32'h39dd98db),
	.w5(32'hb8f6561c),
	.w6(32'h39b53472),
	.w7(32'h3a1153ff),
	.w8(32'h3943c874),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba038150),
	.w1(32'h399b7ace),
	.w2(32'h3a7a0fe7),
	.w3(32'hba935504),
	.w4(32'hb9db53d5),
	.w5(32'h399ac843),
	.w6(32'hba5b4eb2),
	.w7(32'hba421aff),
	.w8(32'hb9a571ef),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e26c9),
	.w1(32'h3710b0d8),
	.w2(32'hb84efc82),
	.w3(32'h37a74696),
	.w4(32'h386068a4),
	.w5(32'hb81280b2),
	.w6(32'h36df22d1),
	.w7(32'h381f5013),
	.w8(32'hb7decd60),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa019f7),
	.w1(32'h3a07f912),
	.w2(32'hb98a5692),
	.w3(32'h3a2207dc),
	.w4(32'h3a0ba3cd),
	.w5(32'hb8d45db8),
	.w6(32'hb9bf3e97),
	.w7(32'h398ec2a3),
	.w8(32'h392b7fc0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81d5560),
	.w1(32'hb822ddd8),
	.w2(32'hb799f31b),
	.w3(32'hb8449e61),
	.w4(32'hb81ff752),
	.w5(32'hb7d749a2),
	.w6(32'hb821ff78),
	.w7(32'hb82f7a6b),
	.w8(32'hb83567d6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e272b),
	.w1(32'hb889d396),
	.w2(32'hb88828ec),
	.w3(32'hb841ced4),
	.w4(32'hb84d3bdb),
	.w5(32'hb8975c1c),
	.w6(32'hb873ad56),
	.w7(32'hb80a87e7),
	.w8(32'hb86fc8de),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaca7e9),
	.w1(32'hb9839b81),
	.w2(32'h39a05a44),
	.w3(32'hbaa7b86e),
	.w4(32'hba739540),
	.w5(32'hb908e9ca),
	.w6(32'hba8872aa),
	.w7(32'hba61e5f6),
	.w8(32'hba11c445),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d3a4),
	.w1(32'h3b1755c9),
	.w2(32'hba96a712),
	.w3(32'h39f0af18),
	.w4(32'h3a8ecb93),
	.w5(32'hbad0e1ed),
	.w6(32'hbae0f25c),
	.w7(32'hba6b637d),
	.w8(32'hbb1b7f3e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac3520),
	.w1(32'h3a16f459),
	.w2(32'h39713d4d),
	.w3(32'h39cc2e5e),
	.w4(32'h3a74cdee),
	.w5(32'h39e6367e),
	.w6(32'h39a61a26),
	.w7(32'h3a391359),
	.w8(32'h39ccbb93),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bb8fd),
	.w1(32'h3a196a89),
	.w2(32'h392f23c3),
	.w3(32'hba871b33),
	.w4(32'hba3afb0c),
	.w5(32'hba18c4e0),
	.w6(32'hba69f73b),
	.w7(32'hba81694b),
	.w8(32'hba96f7d1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9131690),
	.w1(32'hb7f65ad8),
	.w2(32'hb9927df5),
	.w3(32'hb869fc62),
	.w4(32'hb9aba3bd),
	.w5(32'hba39ffb1),
	.w6(32'h3a229625),
	.w7(32'h368722f5),
	.w8(32'hb74a0627),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf80d75),
	.w1(32'hbb77ce3d),
	.w2(32'hbb713743),
	.w3(32'h396b86cf),
	.w4(32'hbad04f47),
	.w5(32'hbb8287ec),
	.w6(32'h3a057325),
	.w7(32'hbaea7f13),
	.w8(32'hbb6f13e8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b67130),
	.w1(32'hb9a64025),
	.w2(32'hbb026161),
	.w3(32'h3a11bf68),
	.w4(32'hb806b3a9),
	.w5(32'hba9f87d2),
	.w6(32'h39729c28),
	.w7(32'hba0a51dc),
	.w8(32'hba6a99e8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a164b42),
	.w1(32'hbaaf1913),
	.w2(32'hbad39efc),
	.w3(32'h3a846bab),
	.w4(32'hba8032bb),
	.w5(32'hbaf14d26),
	.w6(32'hba017e1e),
	.w7(32'hbaea57ae),
	.w8(32'hbaffef2b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ad1146),
	.w1(32'hb770c32e),
	.w2(32'h38637354),
	.w3(32'hb7b7dd5e),
	.w4(32'h37d557b9),
	.w5(32'h38f66309),
	.w6(32'h370372c2),
	.w7(32'h38ad0784),
	.w8(32'h391c844f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b5b55),
	.w1(32'hba2b3013),
	.w2(32'hba9de22b),
	.w3(32'h38c3ae96),
	.w4(32'hba8d46cf),
	.w5(32'hbad26881),
	.w6(32'hb91f8e4b),
	.w7(32'hbac3dc3b),
	.w8(32'hbad0f15c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4eff6),
	.w1(32'h36d3dccf),
	.w2(32'h36b532ad),
	.w3(32'h37bdd77b),
	.w4(32'h361d384f),
	.w5(32'h34ae2251),
	.w6(32'h37d98fe5),
	.w7(32'h371c74ea),
	.w8(32'h371d581d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91390a6),
	.w1(32'h37a2febe),
	.w2(32'h384d7bba),
	.w3(32'h3890d0b4),
	.w4(32'h39a220de),
	.w5(32'h396f3a27),
	.w6(32'h36e48196),
	.w7(32'h39b2df59),
	.w8(32'h393cd416),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8460d07),
	.w1(32'h399313e1),
	.w2(32'h39698c47),
	.w3(32'h370c4aa3),
	.w4(32'h396737f4),
	.w5(32'h397d6a29),
	.w6(32'hb8b32408),
	.w7(32'h38bf51f3),
	.w8(32'hb8a5b8ca),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1f1fd),
	.w1(32'hbaa4b3ce),
	.w2(32'hbafd6339),
	.w3(32'h39577a1e),
	.w4(32'hba8352c7),
	.w5(32'hbb1409a9),
	.w6(32'hb960d810),
	.w7(32'hbac3e0b0),
	.w8(32'hbb11333a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371b8934),
	.w1(32'h3704f930),
	.w2(32'h36cb1b9c),
	.w3(32'h347309a4),
	.w4(32'h363049d6),
	.w5(32'h366853ea),
	.w6(32'h35d29394),
	.w7(32'h352cbad7),
	.w8(32'hb528e1f6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380997f4),
	.w1(32'h377b2857),
	.w2(32'h36934677),
	.w3(32'h3803c50a),
	.w4(32'h36ff6caf),
	.w5(32'h3676774c),
	.w6(32'h3841669d),
	.w7(32'h379279bf),
	.w8(32'hb4d39a71),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c3faf),
	.w1(32'h393139d8),
	.w2(32'h399607dd),
	.w3(32'hb8fbb2c2),
	.w4(32'h3952e364),
	.w5(32'h399bc488),
	.w6(32'hba295ad1),
	.w7(32'hb952f719),
	.w8(32'hb95df94d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82bbc3b),
	.w1(32'hba643a7f),
	.w2(32'hbb142d6a),
	.w3(32'h3b010b58),
	.w4(32'hb92388f0),
	.w5(32'hbb1aef93),
	.w6(32'h3b2aa19c),
	.w7(32'hb966bfc6),
	.w8(32'hbb2e9773),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0b922),
	.w1(32'h3ad90594),
	.w2(32'hbb079c94),
	.w3(32'hb898b54a),
	.w4(32'h3b250ed1),
	.w5(32'hba6f7a5b),
	.w6(32'hbac604b9),
	.w7(32'h3a83017a),
	.w8(32'hbafaa4b5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d6aa2),
	.w1(32'hb8925e33),
	.w2(32'hb852bb81),
	.w3(32'hb823e0b0),
	.w4(32'hb3adca21),
	.w5(32'hb76fdb73),
	.w6(32'h3783a346),
	.w7(32'h38251c5d),
	.w8(32'hb7327f00),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02db24),
	.w1(32'hbb95fb45),
	.w2(32'hbba38193),
	.w3(32'hbabc4612),
	.w4(32'hbb62be43),
	.w5(32'hbb97a712),
	.w6(32'hbb1878de),
	.w7(32'hbb5998ca),
	.w8(32'hbb93f5a8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09cf94),
	.w1(32'h3a5cd948),
	.w2(32'hbab1e57a),
	.w3(32'hb9cc5862),
	.w4(32'h3a7a65d9),
	.w5(32'hbaf41732),
	.w6(32'h39b98847),
	.w7(32'h3a80175f),
	.w8(32'hba93f5d4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33db46),
	.w1(32'h37b4a18c),
	.w2(32'hbab5bd67),
	.w3(32'h3aabbc54),
	.w4(32'h3a039d59),
	.w5(32'hba80d7ce),
	.w6(32'hb883ba29),
	.w7(32'h39671fbb),
	.w8(32'hba4a4e84),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a4b618),
	.w1(32'hb80e99c5),
	.w2(32'hb7cb2384),
	.w3(32'hb7ec719e),
	.w4(32'hb804d090),
	.w5(32'hb7c31af6),
	.w6(32'hb72f6b55),
	.w7(32'hb77fffe6),
	.w8(32'hb7b56c0e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c48523),
	.w1(32'h370fab99),
	.w2(32'h36b4dca3),
	.w3(32'h38354846),
	.w4(32'h37ee1ac2),
	.w5(32'h37585f23),
	.w6(32'h3885b203),
	.w7(32'h3869f8c7),
	.w8(32'h369b3a81),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376ed626),
	.w1(32'hb4067326),
	.w2(32'hb5a5bfef),
	.w3(32'h373b01ea),
	.w4(32'hb62aa735),
	.w5(32'hb5f7328d),
	.w6(32'h3738da50),
	.w7(32'hb628b05b),
	.w8(32'hb5f20f63),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad59b95),
	.w1(32'h3a032004),
	.w2(32'hbab72a42),
	.w3(32'h3ae53c2b),
	.w4(32'h3a2010e0),
	.w5(32'hbaa47f59),
	.w6(32'h39f5e1ab),
	.w7(32'hb9806edd),
	.w8(32'hba8c9fed),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc629),
	.w1(32'h3988d173),
	.w2(32'hba5cadc0),
	.w3(32'h3a8cb51b),
	.w4(32'h39968887),
	.w5(32'hba8acf14),
	.w6(32'h3a4e1501),
	.w7(32'hb917bd1b),
	.w8(32'hba8b2cea),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0608a2),
	.w1(32'hb802d887),
	.w2(32'hba39a569),
	.w3(32'hbb260a3c),
	.w4(32'hba20abf2),
	.w5(32'hba3bff40),
	.w6(32'hbb26747d),
	.w7(32'hba72bc59),
	.w8(32'hbac408b8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949e3cd),
	.w1(32'h3956ef92),
	.w2(32'h395fdb36),
	.w3(32'hba096154),
	.w4(32'h387c2225),
	.w5(32'h396ee32c),
	.w6(32'hb9ef54c6),
	.w7(32'hb917cd3c),
	.w8(32'hb87f106e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdb880),
	.w1(32'hbb1ab9f2),
	.w2(32'hbb284a7d),
	.w3(32'h39521d2b),
	.w4(32'hba84348e),
	.w5(32'hbb1e47b3),
	.w6(32'hba8805c8),
	.w7(32'hbaf24aa6),
	.w8(32'hbb0fa11f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8291b9d),
	.w1(32'hb987a46b),
	.w2(32'hbabb9cf8),
	.w3(32'hb869d8e0),
	.w4(32'hb9a9f7cd),
	.w5(32'hba6b15db),
	.w6(32'hb99f492d),
	.w7(32'hba079fbb),
	.w8(32'hba99bee0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379d129e),
	.w1(32'h374e13e2),
	.w2(32'h37bd914e),
	.w3(32'h378da081),
	.w4(32'h370c127e),
	.w5(32'h37903b81),
	.w6(32'h378f7f2a),
	.w7(32'h37273f3d),
	.w8(32'h378a856a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd4d6b),
	.w1(32'hbaf24c8d),
	.w2(32'hbadfc493),
	.w3(32'hba36c525),
	.w4(32'hba4e0881),
	.w5(32'hba98ec90),
	.w6(32'hba23fd90),
	.w7(32'hba9a2e4d),
	.w8(32'hba952bc5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3808b0d5),
	.w1(32'h37a7e51e),
	.w2(32'h381625c6),
	.w3(32'h37b60f51),
	.w4(32'h344df776),
	.w5(32'h37a3cdd0),
	.w6(32'h37e21351),
	.w7(32'h37407161),
	.w8(32'h37a3c7b6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de0970),
	.w1(32'hba5e184d),
	.w2(32'hbabb2296),
	.w3(32'hb96a9699),
	.w4(32'hba116126),
	.w5(32'hba9af480),
	.w6(32'hba2e0228),
	.w7(32'hba554c6a),
	.w8(32'hba9a2bf7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fabf8),
	.w1(32'h3b0b8080),
	.w2(32'h3a5c9133),
	.w3(32'hb98eb7da),
	.w4(32'h3aeaeb4c),
	.w5(32'h3a1a628e),
	.w6(32'hba287bdf),
	.w7(32'h3a8fd5c3),
	.w8(32'hba0bbf12),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55e361),
	.w1(32'h396fd28b),
	.w2(32'hb99db353),
	.w3(32'hba787de2),
	.w4(32'hb90d2bf0),
	.w5(32'hb9ce01de),
	.w6(32'hba8d025a),
	.w7(32'hba239455),
	.w8(32'hba90ef5a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d6868),
	.w1(32'h38323188),
	.w2(32'hb802559e),
	.w3(32'h38c8f510),
	.w4(32'h3950874e),
	.w5(32'h38b0c064),
	.w6(32'h38b51fac),
	.w7(32'h3939eb4d),
	.w8(32'h38327fed),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d77ba),
	.w1(32'hba347275),
	.w2(32'hb9b84def),
	.w3(32'hbb3062ed),
	.w4(32'hba9d20ad),
	.w5(32'hba3a077c),
	.w6(32'hbb04db77),
	.w7(32'hbaa7cd68),
	.w8(32'hbab24879),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a221f),
	.w1(32'hba8e2685),
	.w2(32'hbab8b5f3),
	.w3(32'h3a032373),
	.w4(32'hba1f7b88),
	.w5(32'hbac34b98),
	.w6(32'hb9ca825b),
	.w7(32'hba8cde3e),
	.w8(32'hba9fbfe2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab81b96),
	.w1(32'hb9e33c33),
	.w2(32'hbad2b312),
	.w3(32'hba3f44c8),
	.w4(32'h38aa599d),
	.w5(32'hba7ff948),
	.w6(32'hba143cbf),
	.w7(32'hb8ad0842),
	.w8(32'hba82bcb3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc3d80),
	.w1(32'hb63e682d),
	.w2(32'h378ffd12),
	.w3(32'h37a97de2),
	.w4(32'hb60e5f03),
	.w5(32'h3733d663),
	.w6(32'h37e07430),
	.w7(32'h37cbb998),
	.w8(32'h380c6786),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363512db),
	.w1(32'hb45bd2ed),
	.w2(32'hb7b2526d),
	.w3(32'hb85edb48),
	.w4(32'hb87f045d),
	.w5(32'hb8c7d992),
	.w6(32'hb85a8102),
	.w7(32'hb80f8638),
	.w8(32'hb82819e6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae064e2),
	.w1(32'h3aa11ad9),
	.w2(32'hbb1c9e57),
	.w3(32'h373a862f),
	.w4(32'h3a6f04c7),
	.w5(32'hbadbedad),
	.w6(32'hbab63eba),
	.w7(32'hbaa649ef),
	.w8(32'hbb4485c4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b4374),
	.w1(32'h39dfe4cc),
	.w2(32'hba7bbd91),
	.w3(32'hb843f6d1),
	.w4(32'hb7b05aa6),
	.w5(32'hba9ad404),
	.w6(32'hb9d3edad),
	.w7(32'hba2b6562),
	.w8(32'hbae94a8d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace7c97),
	.w1(32'h380a333a),
	.w2(32'hba0383ec),
	.w3(32'hbae55435),
	.w4(32'hba17c0c4),
	.w5(32'hba095b93),
	.w6(32'hbaffc48f),
	.w7(32'hbaa0e12d),
	.w8(32'hbab8acde),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c5b1e),
	.w1(32'hbae1336d),
	.w2(32'hbb58f558),
	.w3(32'h3b704fe9),
	.w4(32'h39a4eba7),
	.w5(32'hbb38489e),
	.w6(32'h3b176c96),
	.w7(32'hb9ad143e),
	.w8(32'hbae681bc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399594db),
	.w1(32'hb90e9c11),
	.w2(32'h37439853),
	.w3(32'h3983594c),
	.w4(32'hb7364c14),
	.w5(32'h38561fe1),
	.w6(32'h37600f31),
	.w7(32'hb812ef1b),
	.w8(32'h381003b6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02ca1c),
	.w1(32'hb8f9fcbe),
	.w2(32'hba1322eb),
	.w3(32'h38630127),
	.w4(32'hb9570bf1),
	.w5(32'hb9b097bb),
	.w6(32'h38e12229),
	.w7(32'hb9e32fbb),
	.w8(32'hb9cd6e4c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf736),
	.w1(32'h3baf3b2a),
	.w2(32'hbb252f52),
	.w3(32'h3b266365),
	.w4(32'h3b8d873f),
	.w5(32'hbb28877f),
	.w6(32'hbb04d85b),
	.w7(32'h3abaa1e9),
	.w8(32'hbb1b6594),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3dcf9),
	.w1(32'hbb188561),
	.w2(32'hbb757349),
	.w3(32'h3a0c9e6a),
	.w4(32'hbab453a2),
	.w5(32'hbb46053a),
	.w6(32'hba0d578d),
	.w7(32'hba561674),
	.w8(32'hbb06d3f2),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0984ce),
	.w1(32'h38c02e03),
	.w2(32'hbb574a47),
	.w3(32'h3a8cc02b),
	.w4(32'h3a1c0416),
	.w5(32'hbb3b4121),
	.w6(32'hba3b6c06),
	.w7(32'hb98c33fc),
	.w8(32'hbb665ad6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f88bb),
	.w1(32'h3b0d9e1e),
	.w2(32'h3b0080ff),
	.w3(32'hba8d83b8),
	.w4(32'h3ac78fc1),
	.w5(32'h3ad96f24),
	.w6(32'hba252cf5),
	.w7(32'h3ac50aed),
	.w8(32'h3a9aaeee),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb385d41),
	.w1(32'h39b38991),
	.w2(32'h3a4af48c),
	.w3(32'hbb3f1861),
	.w4(32'hb9d71655),
	.w5(32'h3a34280c),
	.w6(32'hbb0581e0),
	.w7(32'hb9e6b40d),
	.w8(32'hba014f62),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c96a07),
	.w1(32'h36e18224),
	.w2(32'h36f48bab),
	.w3(32'h360b2887),
	.w4(32'h3687fc64),
	.w5(32'h36b16f38),
	.w6(32'h368d4fd4),
	.w7(32'h369fb52f),
	.w8(32'h36960739),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b8c6a),
	.w1(32'h36a3e1e0),
	.w2(32'h3718151c),
	.w3(32'h371226c3),
	.w4(32'h36a29342),
	.w5(32'h37101037),
	.w6(32'h373ef076),
	.w7(32'h36d1be99),
	.w8(32'h3728d871),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd271e),
	.w1(32'h392b014e),
	.w2(32'hb95b5966),
	.w3(32'h38f55ed6),
	.w4(32'hb9d7ee1c),
	.w5(32'hba26cad8),
	.w6(32'hb9cd60d3),
	.w7(32'hb9db30dc),
	.w8(32'hb9d4af25),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3749c198),
	.w1(32'hb64cb85d),
	.w2(32'h36f35979),
	.w3(32'h36b9a406),
	.w4(32'hb6cea229),
	.w5(32'h3632f5f5),
	.w6(32'h3706e0b5),
	.w7(32'hb6887637),
	.w8(32'h3668d857),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aeaa0),
	.w1(32'h370d68d8),
	.w2(32'hba5c5618),
	.w3(32'h3a9cd1b0),
	.w4(32'h38b00716),
	.w5(32'hba4fb3fe),
	.w6(32'h3a0bd710),
	.w7(32'hb9fc7658),
	.w8(32'hba177b7c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeca036),
	.w1(32'hb9de3aa1),
	.w2(32'hbac1579e),
	.w3(32'hb974bf99),
	.w4(32'hba815738),
	.w5(32'hbac46544),
	.w6(32'hb96ca795),
	.w7(32'hbaaa3dfa),
	.w8(32'hbb15e911),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bde41),
	.w1(32'h39361747),
	.w2(32'hb91b3ba1),
	.w3(32'hb9f6cd26),
	.w4(32'hb9f7579b),
	.w5(32'hb9bce80a),
	.w6(32'hba3b5ee4),
	.w7(32'hba6d31cd),
	.w8(32'hba6757eb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b1bf5),
	.w1(32'h378d5908),
	.w2(32'h37c8280d),
	.w3(32'h372082b8),
	.w4(32'h376d534f),
	.w5(32'h37be72d1),
	.w6(32'h36f8d331),
	.w7(32'h37a6cd90),
	.w8(32'h37c30a85),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a8d3a),
	.w1(32'h3a39e5d4),
	.w2(32'hbbb6c691),
	.w3(32'h3b20d4ab),
	.w4(32'h3ab7601f),
	.w5(32'hbb9a00d5),
	.w6(32'hba88bccb),
	.w7(32'hb9ac2d76),
	.w8(32'hbb9f2953),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a69eb),
	.w1(32'hb9e95048),
	.w2(32'hba9920b6),
	.w3(32'h3a79bbd0),
	.w4(32'hb86de3fd),
	.w5(32'hba9af3e0),
	.w6(32'hb7e3651c),
	.w7(32'hba0f8492),
	.w8(32'hba995ad3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817df6d),
	.w1(32'h38e8be96),
	.w2(32'h3939c0fd),
	.w3(32'hb8b897bd),
	.w4(32'h38529de8),
	.w5(32'h3953c5c1),
	.w6(32'hb7d72688),
	.w7(32'h38b5e929),
	.w8(32'h398a70a0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac95b84),
	.w1(32'hb86d9991),
	.w2(32'hbad9a37a),
	.w3(32'h3ac60187),
	.w4(32'h399ca10f),
	.w5(32'hbaae1e8f),
	.w6(32'h3a01f137),
	.w7(32'hb84adb21),
	.w8(32'hba70f80b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37675383),
	.w1(32'h37e337ac),
	.w2(32'h377fb33c),
	.w3(32'h37565ca8),
	.w4(32'h37cf6a84),
	.w5(32'h37625ae5),
	.w6(32'hb76ef684),
	.w7(32'h3770c12e),
	.w8(32'h376cf70c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949815b),
	.w1(32'h391d0d63),
	.w2(32'h38207e19),
	.w3(32'h39559500),
	.w4(32'h391fb147),
	.w5(32'h38a136a5),
	.w6(32'hb743e887),
	.w7(32'hb6e8de10),
	.w8(32'hb76b705b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379933ae),
	.w1(32'h36bd0254),
	.w2(32'h363dced7),
	.w3(32'h3683814a),
	.w4(32'hb5f63359),
	.w5(32'h35319694),
	.w6(32'hb6a408d0),
	.w7(32'h36715706),
	.w8(32'hb7527ea9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383e0a8c),
	.w1(32'hb7b36a2b),
	.w2(32'hb79369a4),
	.w3(32'h37752a95),
	.w4(32'hb7efb039),
	.w5(32'hb7f81f91),
	.w6(32'hb7bc9128),
	.w7(32'hb852315b),
	.w8(32'hb83e6604),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95fd6a8),
	.w1(32'h3a571d64),
	.w2(32'h3a265f57),
	.w3(32'hb9defc3e),
	.w4(32'h3a0422d7),
	.w5(32'h3a160734),
	.w6(32'hb814b9e1),
	.w7(32'h3a1f1856),
	.w8(32'h399a2a43),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888c815),
	.w1(32'hbb45cabe),
	.w2(32'hbb6db776),
	.w3(32'h3aea77ef),
	.w4(32'hbac5dbb5),
	.w5(32'hbb5b15bd),
	.w6(32'h3a86d4fd),
	.w7(32'hbb2300de),
	.w8(32'hbb238323),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacea38),
	.w1(32'hba4b3b02),
	.w2(32'hbaf996b5),
	.w3(32'h3a9f1731),
	.w4(32'hba217719),
	.w5(32'hbadce274),
	.w6(32'h398a02f9),
	.w7(32'hba58007b),
	.w8(32'hbab3386e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba312a9c),
	.w1(32'hbb268d8d),
	.w2(32'hbb28d658),
	.w3(32'h39e4edb7),
	.w4(32'hba7a4fb4),
	.w5(32'hbb205cda),
	.w6(32'h38c61bca),
	.w7(32'hbaa48568),
	.w8(32'hbab7708c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803904c),
	.w1(32'h3849834d),
	.w2(32'h38703863),
	.w3(32'h3738b766),
	.w4(32'h381d6463),
	.w5(32'h37efe3af),
	.w6(32'hb7ba58d2),
	.w7(32'hb67dd9cc),
	.w8(32'hb7af5d9f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc59c3),
	.w1(32'hb887e63f),
	.w2(32'hb974b6d2),
	.w3(32'h39315677),
	.w4(32'hb91a420b),
	.w5(32'hb969269d),
	.w6(32'hb873969b),
	.w7(32'hb940ed80),
	.w8(32'hb969848f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e70a7a),
	.w1(32'hb7003e7c),
	.w2(32'hb5ccc3b3),
	.w3(32'hb6c18c4a),
	.w4(32'hb7830931),
	.w5(32'hb6215e49),
	.w6(32'hb62b3e06),
	.w7(32'hb766d6a8),
	.w8(32'hb7694bfc),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a0cca9),
	.w1(32'h374cf571),
	.w2(32'h37130102),
	.w3(32'h37959ccf),
	.w4(32'h37656448),
	.w5(32'h36052ae6),
	.w6(32'h37c4de7a),
	.w7(32'h3761827a),
	.w8(32'hb56a0f4d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91615d0),
	.w1(32'hbb001831),
	.w2(32'hbb520bcd),
	.w3(32'h39aeee16),
	.w4(32'hbac5b531),
	.w5(32'hbb4d498d),
	.w6(32'hba1f19d9),
	.w7(32'hbb20a09b),
	.w8(32'hbb5584ba),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7db789e),
	.w1(32'hb8412926),
	.w2(32'hb77ce530),
	.w3(32'h36cacf22),
	.w4(32'hb81ecfde),
	.w5(32'hb7697cdb),
	.w6(32'h37a906d9),
	.w7(32'hb5797a69),
	.w8(32'hb5907cf1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68072ba),
	.w1(32'h39641c01),
	.w2(32'hb9278d22),
	.w3(32'h3913c8d1),
	.w4(32'h39ca9d10),
	.w5(32'hb864f65e),
	.w6(32'h391f8b18),
	.w7(32'h396c9c95),
	.w8(32'hb938fe6d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79c1e3b),
	.w1(32'hb8619692),
	.w2(32'hb9fada43),
	.w3(32'h35fa2a30),
	.w4(32'hb4daaaf4),
	.w5(32'hb9ab464a),
	.w6(32'h37a08088),
	.w7(32'hb88128e8),
	.w8(32'hb9317e57),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb706428f),
	.w1(32'hb7c5f6ef),
	.w2(32'hb778b51e),
	.w3(32'h36479f9a),
	.w4(32'hb7d3edb3),
	.w5(32'hb7e403eb),
	.w6(32'h37d0a668),
	.w7(32'hb4735434),
	.w8(32'hb7a6d1d4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930c068),
	.w1(32'hba3d123e),
	.w2(32'hba72e530),
	.w3(32'h386c956a),
	.w4(32'hba04025f),
	.w5(32'hba4080c3),
	.w6(32'hb994532d),
	.w7(32'hba12c4cf),
	.w8(32'hba5082ef),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835e839),
	.w1(32'hb9707962),
	.w2(32'hb96a9178),
	.w3(32'h37a90cca),
	.w4(32'hb935d453),
	.w5(32'hb9270628),
	.w6(32'hb9398985),
	.w7(32'hb958fbee),
	.w8(32'hb94fc48b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b2caf),
	.w1(32'hbb500dc1),
	.w2(32'hbbb31648),
	.w3(32'h3aa722e4),
	.w4(32'hba100f9d),
	.w5(32'hbba02b9f),
	.w6(32'hba85a819),
	.w7(32'hbb300c5c),
	.w8(32'hbb67a1e8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d8825),
	.w1(32'hbaa8b08c),
	.w2(32'hbaeb2511),
	.w3(32'h378f930f),
	.w4(32'hba9d3c38),
	.w5(32'hbab8b025),
	.w6(32'hba8d9bb6),
	.w7(32'hbaddc6a6),
	.w8(32'hba392d46),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ba9d),
	.w1(32'hba074f5f),
	.w2(32'hbb07e01c),
	.w3(32'hb9c86925),
	.w4(32'hba703600),
	.w5(32'hbaf81985),
	.w6(32'hbb587ca4),
	.w7(32'hbb4b1a91),
	.w8(32'hbb36c77c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule