module layer_10_featuremap_101(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e165c),
	.w1(32'hbb1ed495),
	.w2(32'hbb95017f),
	.w3(32'hb9393e8b),
	.w4(32'h3b6079f2),
	.w5(32'hba50ad49),
	.w6(32'hbbb1ea1a),
	.w7(32'hbac15465),
	.w8(32'hba02a9b4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5538e1),
	.w1(32'h3af0c2cf),
	.w2(32'h3b2c3126),
	.w3(32'hba4fd8b5),
	.w4(32'hba83e38e),
	.w5(32'h3ab62649),
	.w6(32'h391c7149),
	.w7(32'h3a810f3d),
	.w8(32'h3af59a82),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c4f91),
	.w1(32'hba1aca11),
	.w2(32'h3bb534d6),
	.w3(32'h39246234),
	.w4(32'hbac3888c),
	.w5(32'hb974aba9),
	.w6(32'hb90125dc),
	.w7(32'h38db78fc),
	.w8(32'hb7fbd1aa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a695f37),
	.w1(32'h3aa62cfe),
	.w2(32'hbb79acb7),
	.w3(32'hbb2a3239),
	.w4(32'hbb102bc2),
	.w5(32'h39856266),
	.w6(32'h3a2ddf60),
	.w7(32'hbb71f475),
	.w8(32'hbba16f97),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19bdcd),
	.w1(32'hba6c1cb7),
	.w2(32'h3a5a5629),
	.w3(32'hbb58506a),
	.w4(32'h398ee9d8),
	.w5(32'hbaa229d7),
	.w6(32'h3910bab8),
	.w7(32'h3a349d44),
	.w8(32'hba67ef57),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94a771),
	.w1(32'h396e0470),
	.w2(32'hbae5c9dc),
	.w3(32'h3b1a6fe5),
	.w4(32'hba62fc16),
	.w5(32'hba7a9894),
	.w6(32'hb99ab642),
	.w7(32'hb907284d),
	.w8(32'h39e1fbd5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba817762),
	.w1(32'h3b1b7ffe),
	.w2(32'h3b2bab09),
	.w3(32'hba303502),
	.w4(32'h3a20a60a),
	.w5(32'h391d24e7),
	.w6(32'hba055b12),
	.w7(32'h396d5767),
	.w8(32'hba9f63ae),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0f540),
	.w1(32'h39b4c4bd),
	.w2(32'hba99a261),
	.w3(32'hbac32815),
	.w4(32'hb9f84f7d),
	.w5(32'hbab8e3b2),
	.w6(32'hbaa9dfde),
	.w7(32'hbb825563),
	.w8(32'hbb2d02b9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a536a9d),
	.w1(32'h3846b740),
	.w2(32'h36dbef38),
	.w3(32'h3ad05054),
	.w4(32'h38f2672f),
	.w5(32'h3a5b6157),
	.w6(32'h3980a7e9),
	.w7(32'h39a3b051),
	.w8(32'hb99d845e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd25a5),
	.w1(32'hbbab268f),
	.w2(32'hbb34e22a),
	.w3(32'hbbb07ea7),
	.w4(32'hbb6d4534),
	.w5(32'h384197d2),
	.w6(32'hbb820c20),
	.w7(32'hbbc73448),
	.w8(32'hbbb26b31),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89eb54),
	.w1(32'h3c1ea87b),
	.w2(32'h3ca10896),
	.w3(32'h3a989ab1),
	.w4(32'hbb22d8c0),
	.w5(32'h3b027821),
	.w6(32'h3c2f2b2d),
	.w7(32'h3bc8631c),
	.w8(32'h3c1c0b78),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c754987),
	.w1(32'h3b56629c),
	.w2(32'h3bdcb65b),
	.w3(32'h3ac0198f),
	.w4(32'h37b84d37),
	.w5(32'h3bc10409),
	.w6(32'h3b41615b),
	.w7(32'h3ab851b1),
	.w8(32'h3a813fc4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9ec6),
	.w1(32'hbb851dfe),
	.w2(32'h3aa6b7fc),
	.w3(32'hbba38cfe),
	.w4(32'hbba15601),
	.w5(32'hba54fc0e),
	.w6(32'hbbe6415d),
	.w7(32'hbbe07c1b),
	.w8(32'hbb4dda08),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eac56),
	.w1(32'h3a0dab76),
	.w2(32'h3b2e8773),
	.w3(32'hbb302aab),
	.w4(32'hba052d1f),
	.w5(32'h3b56fba5),
	.w6(32'hbace1204),
	.w7(32'hbb6cc7ec),
	.w8(32'hba8980c6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad025e7),
	.w1(32'hbb6d5775),
	.w2(32'hba5e508a),
	.w3(32'h3a5b416e),
	.w4(32'hbb793334),
	.w5(32'hbb064978),
	.w6(32'h3b452b5c),
	.w7(32'hb9b3a204),
	.w8(32'hbac79efb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e57cd),
	.w1(32'hbb0e6f8d),
	.w2(32'hba3b4f31),
	.w3(32'hbb85a376),
	.w4(32'hbb25ed05),
	.w5(32'hba0ba5a9),
	.w6(32'hbb50f8a4),
	.w7(32'hbb82bcdc),
	.w8(32'hbb6a928a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9542693),
	.w1(32'hbaa27468),
	.w2(32'h3bf817d0),
	.w3(32'h398fcd9f),
	.w4(32'hbb1d764a),
	.w5(32'h3bb32136),
	.w6(32'hb9e2b725),
	.w7(32'h3ba50829),
	.w8(32'hbab82974),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e4a5b),
	.w1(32'hb961e022),
	.w2(32'h3ad0fe96),
	.w3(32'hbb440278),
	.w4(32'hbb8fdf43),
	.w5(32'hbb4c5d62),
	.w6(32'hbb77d86a),
	.w7(32'hbbccd025),
	.w8(32'hbc105842),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11460c),
	.w1(32'hb9da9b85),
	.w2(32'h3b0a1aeb),
	.w3(32'hbb02f097),
	.w4(32'hbb42ee41),
	.w5(32'hba3a1cbd),
	.w6(32'hbb6c7b8f),
	.w7(32'hbb3063fd),
	.w8(32'hbb92012b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3abe57),
	.w1(32'h3a545325),
	.w2(32'h3a00f281),
	.w3(32'hba9fdd14),
	.w4(32'h39ef8562),
	.w5(32'h39f2d927),
	.w6(32'h3a01dc9e),
	.w7(32'h3aaded99),
	.w8(32'hba1070a0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b83554),
	.w1(32'hbb19bd94),
	.w2(32'hbb352e65),
	.w3(32'hb8d71045),
	.w4(32'hbb106c88),
	.w5(32'h3a2b6ff2),
	.w6(32'hbaeae912),
	.w7(32'hb9da92cb),
	.w8(32'hbaf08edd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf840e7),
	.w1(32'hb9f2c90d),
	.w2(32'h3c5f8a37),
	.w3(32'hbaee3aa4),
	.w4(32'hb9e12344),
	.w5(32'hb9f45460),
	.w6(32'h38e2715f),
	.w7(32'hb9985f4b),
	.w8(32'h3c0793f3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceeb89),
	.w1(32'h3bac7f1d),
	.w2(32'h3c85ccb4),
	.w3(32'hbb593b9c),
	.w4(32'hbbad4f97),
	.w5(32'h3c4a03a8),
	.w6(32'h3b8e24d4),
	.w7(32'h3c2a1f2d),
	.w8(32'h3bcaf2d6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a4ebd),
	.w1(32'hbb2a1b60),
	.w2(32'hba06c10e),
	.w3(32'hbbc9186d),
	.w4(32'hbb6fb77a),
	.w5(32'hb94b6ec3),
	.w6(32'hbb07e406),
	.w7(32'hbb5cedb4),
	.w8(32'hb984b067),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6ba8),
	.w1(32'h3b19d6cc),
	.w2(32'h3b781e98),
	.w3(32'hb9ddb8f1),
	.w4(32'hbac0728f),
	.w5(32'h3b172c73),
	.w6(32'hba3e55c1),
	.w7(32'h39d738c7),
	.w8(32'h3b7f52e2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98598a0),
	.w1(32'hbb6f412a),
	.w2(32'h3b534c05),
	.w3(32'hbaed3014),
	.w4(32'hbb9d0ff5),
	.w5(32'h3a574005),
	.w6(32'hba92989f),
	.w7(32'hb81a0179),
	.w8(32'hbad6d464),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852d66f),
	.w1(32'h3ab14d16),
	.w2(32'h3a43ba0f),
	.w3(32'hbb82448b),
	.w4(32'h3a831e90),
	.w5(32'h3a9d78f9),
	.w6(32'h3a8f8bb9),
	.w7(32'h3ad61393),
	.w8(32'hb7608f30),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a478d76),
	.w1(32'h39fa2303),
	.w2(32'hbb0a6f86),
	.w3(32'h3a8cfb1c),
	.w4(32'hb93f8f93),
	.w5(32'hbab955c7),
	.w6(32'h3b2872ef),
	.w7(32'hbaabbfdb),
	.w8(32'hbaca2930),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef4289),
	.w1(32'h3a05e960),
	.w2(32'h3bb824dc),
	.w3(32'hbb204861),
	.w4(32'hbbbb4509),
	.w5(32'h3b15dfc2),
	.w6(32'hb9b582d7),
	.w7(32'h3b033f33),
	.w8(32'h3b84d41b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30b452),
	.w1(32'hbc559479),
	.w2(32'hbb77200f),
	.w3(32'hbb966570),
	.w4(32'hbc2850e6),
	.w5(32'h3a558c1d),
	.w6(32'hbbbe126d),
	.w7(32'h3948ba49),
	.w8(32'h3b275971),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b482297),
	.w1(32'hba9519be),
	.w2(32'hb9d28d3b),
	.w3(32'h3b58fd9c),
	.w4(32'hba3f10a0),
	.w5(32'h39a0fd16),
	.w6(32'hb8d4fc53),
	.w7(32'h3a010245),
	.w8(32'hb8846b5b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f7003),
	.w1(32'h3a83c383),
	.w2(32'h3ab97e7a),
	.w3(32'hba34ae29),
	.w4(32'hb9d70c78),
	.w5(32'h39517830),
	.w6(32'h3a3829b0),
	.w7(32'h3a3f64eb),
	.w8(32'h38d657f5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b162c),
	.w1(32'h3a40d10a),
	.w2(32'h3bab8ba5),
	.w3(32'hbb08145b),
	.w4(32'hba8e812c),
	.w5(32'h3ab3d1a4),
	.w6(32'h3b0081af),
	.w7(32'h3b94dd44),
	.w8(32'hb7c5630d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89e8a6),
	.w1(32'h388f016e),
	.w2(32'hbb6530d3),
	.w3(32'h3b926e6e),
	.w4(32'h3af376c9),
	.w5(32'hbb872de4),
	.w6(32'hbafdc84e),
	.w7(32'hba443db9),
	.w8(32'hb8a024c1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1dec8),
	.w1(32'h3a25e003),
	.w2(32'hb9de8b30),
	.w3(32'hbb9f7e2b),
	.w4(32'h39cb0284),
	.w5(32'hba0c1bb0),
	.w6(32'hba5bf5f3),
	.w7(32'hbaca8e4c),
	.w8(32'hbb0fcd15),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9727cb5),
	.w1(32'h3b10b3ee),
	.w2(32'h3b4a98c2),
	.w3(32'hba4aa29a),
	.w4(32'h39a77953),
	.w5(32'h3a5cd869),
	.w6(32'h3a757c48),
	.w7(32'h3a99a644),
	.w8(32'hba4a09aa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984933d),
	.w1(32'hbac9eafa),
	.w2(32'h3aaa2a6f),
	.w3(32'hba64f3fd),
	.w4(32'hbb483365),
	.w5(32'h3b50f71b),
	.w6(32'hbb0f40fc),
	.w7(32'hbb685694),
	.w8(32'hbad20365),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebe9c0),
	.w1(32'h3bf71456),
	.w2(32'h3c2ecccb),
	.w3(32'h398a39ca),
	.w4(32'hba6943e0),
	.w5(32'h3b7ccb8c),
	.w6(32'h3bbf1cdf),
	.w7(32'h3bb794aa),
	.w8(32'h3c1513ea),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b99d0),
	.w1(32'h3bc8ba73),
	.w2(32'h3c38a6f0),
	.w3(32'hbb80855e),
	.w4(32'h3a8cb98f),
	.w5(32'h3be5918b),
	.w6(32'h3b46b8f2),
	.w7(32'h3bd4976f),
	.w8(32'h3c332bd6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00f880),
	.w1(32'h3b054f60),
	.w2(32'h3aaf6adc),
	.w3(32'h399c524e),
	.w4(32'h3a6c2cf8),
	.w5(32'h3a38c653),
	.w6(32'h3b055313),
	.w7(32'h3a900bc8),
	.w8(32'h39041f51),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957a510),
	.w1(32'hbc35b064),
	.w2(32'hbb6e3744),
	.w3(32'h39bca98c),
	.w4(32'hbbd54079),
	.w5(32'h3a680218),
	.w6(32'hbad2aa3d),
	.w7(32'h3bdd166c),
	.w8(32'h3c1b6bdc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3d952),
	.w1(32'h398a4982),
	.w2(32'h3b0ef7fa),
	.w3(32'h3b14a161),
	.w4(32'hbb7224ba),
	.w5(32'hb6f8da5d),
	.w6(32'h3b6d5349),
	.w7(32'h3a2ec622),
	.w8(32'hba39814f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895eb0e),
	.w1(32'hbb406e99),
	.w2(32'h3aa0894b),
	.w3(32'hbb2b5283),
	.w4(32'hbb15ac0e),
	.w5(32'h3b9061d2),
	.w6(32'hba0a440c),
	.w7(32'h3a1bc7a1),
	.w8(32'h3ad2a30b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82d93b),
	.w1(32'hbb126993),
	.w2(32'hbb6268f7),
	.w3(32'hbbfaa177),
	.w4(32'h39963d08),
	.w5(32'hba0b0316),
	.w6(32'hbbcfa845),
	.w7(32'hbc2ed2c6),
	.w8(32'hbc1a5b96),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace19de),
	.w1(32'hbb0a408e),
	.w2(32'h3b4e2710),
	.w3(32'hba34c0b9),
	.w4(32'hbb378eb4),
	.w5(32'hb94266e6),
	.w6(32'hba4e1866),
	.w7(32'hba32d8bc),
	.w8(32'hba2ecea9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994dd3),
	.w1(32'hbac437f9),
	.w2(32'h3b9c58fb),
	.w3(32'hbbaf3e8f),
	.w4(32'hbb8da4e5),
	.w5(32'hbae3424a),
	.w6(32'hbba19e5f),
	.w7(32'hbba224ad),
	.w8(32'hbadba6ac),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a541654),
	.w1(32'hba1000f8),
	.w2(32'hba3ccb57),
	.w3(32'hba8a4744),
	.w4(32'hba4ced09),
	.w5(32'h3be60312),
	.w6(32'h3b9c1ffb),
	.w7(32'h3b4f9da6),
	.w8(32'h3b51104a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba027e6),
	.w1(32'h39d6a45b),
	.w2(32'h3b9a8cd6),
	.w3(32'hbb9ca1e0),
	.w4(32'hbbec8348),
	.w5(32'hb99be16c),
	.w6(32'hbbad5ed9),
	.w7(32'hbb77395c),
	.w8(32'hbbe2728f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b498c67),
	.w1(32'h3ab1031d),
	.w2(32'h3b1d4c30),
	.w3(32'hbb47a1c7),
	.w4(32'h396c9b6a),
	.w5(32'h3b0b0f94),
	.w6(32'h393fdb4a),
	.w7(32'h3b41b16a),
	.w8(32'h3a38eed4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8625ee),
	.w1(32'h3b073a7c),
	.w2(32'h3a2ec699),
	.w3(32'hb7a2a87e),
	.w4(32'h3b340dac),
	.w5(32'h3b34c8e2),
	.w6(32'h3ad008a7),
	.w7(32'h3a8979e3),
	.w8(32'h3b32802b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397741ba),
	.w1(32'h3ae03388),
	.w2(32'h3b1746c4),
	.w3(32'h39415b7a),
	.w4(32'h3aa106fb),
	.w5(32'h3abac869),
	.w6(32'hba87a687),
	.w7(32'hbae7ecfa),
	.w8(32'hbb015c07),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cbca6),
	.w1(32'h3a78545d),
	.w2(32'hbb89b76b),
	.w3(32'hbb09865f),
	.w4(32'hba566804),
	.w5(32'hbb205dc1),
	.w6(32'h379c0fa5),
	.w7(32'hbb5e690e),
	.w8(32'hbbd97f4b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36d084),
	.w1(32'hba094876),
	.w2(32'hba807cc2),
	.w3(32'h3b3237bc),
	.w4(32'hbb1f8641),
	.w5(32'h39b7812d),
	.w6(32'h3a96ae6f),
	.w7(32'h3abef048),
	.w8(32'h3b0e67c5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364522),
	.w1(32'hbb02ce4f),
	.w2(32'h39f28459),
	.w3(32'hbb55357f),
	.w4(32'hbad98031),
	.w5(32'hbb826b33),
	.w6(32'hbb9b6471),
	.w7(32'hbbceb506),
	.w8(32'hbbdfa6bf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926ac55),
	.w1(32'hbaad1983),
	.w2(32'h3a763060),
	.w3(32'h3b1ca4fd),
	.w4(32'hbb17a513),
	.w5(32'h3a1be41d),
	.w6(32'h3a765f1c),
	.w7(32'h3b91572d),
	.w8(32'h3b6accb0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44226a),
	.w1(32'hbc196b7b),
	.w2(32'hb9cfc149),
	.w3(32'hbac44034),
	.w4(32'hbbb57a60),
	.w5(32'h3a93087e),
	.w6(32'h3af4c71f),
	.w7(32'h3bcda3be),
	.w8(32'h3c3675fb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d018b),
	.w1(32'hb99740b1),
	.w2(32'h3b5ae91c),
	.w3(32'h3ba7b1b3),
	.w4(32'hbb6f6159),
	.w5(32'hbaad0884),
	.w6(32'h3ab7304a),
	.w7(32'h3b542094),
	.w8(32'h3b982482),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6eaaa),
	.w1(32'h3a377508),
	.w2(32'h3b127151),
	.w3(32'hbaba7acc),
	.w4(32'h39ec04ba),
	.w5(32'hbb017d4a),
	.w6(32'hba4c05ca),
	.w7(32'hbaa509fe),
	.w8(32'h392e171e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb9658),
	.w1(32'h39cb2654),
	.w2(32'hb96cfaa2),
	.w3(32'hb9965775),
	.w4(32'hba54b281),
	.w5(32'hba0f79e6),
	.w6(32'hb934d4ce),
	.w7(32'hbae6513a),
	.w8(32'hbabb03c3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba759c3d),
	.w1(32'hb97db321),
	.w2(32'hbad50c8c),
	.w3(32'hba5e07a8),
	.w4(32'hba1bce05),
	.w5(32'hba8471a9),
	.w6(32'h3a0933b9),
	.w7(32'hba1a708f),
	.w8(32'hbab205d5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadde299),
	.w1(32'hb9f51af9),
	.w2(32'h3a950277),
	.w3(32'hbaa88ef0),
	.w4(32'hbad73a80),
	.w5(32'hba4e538d),
	.w6(32'hbb4eabbd),
	.w7(32'hbb2d59c5),
	.w8(32'hbb358ad2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b19288),
	.w1(32'hbb2cb6fe),
	.w2(32'hbb1c8495),
	.w3(32'hba8273e4),
	.w4(32'hbb121c09),
	.w5(32'hbb3e1a32),
	.w6(32'h37a17f1b),
	.w7(32'hbb30d1e5),
	.w8(32'hbb35c4e8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21fbc),
	.w1(32'hb924f07e),
	.w2(32'h39480627),
	.w3(32'hba4735d6),
	.w4(32'hb991bf86),
	.w5(32'hbb79d914),
	.w6(32'h3bd7c19a),
	.w7(32'h3b127a00),
	.w8(32'hbac42213),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bdec0a),
	.w1(32'h3b2b798c),
	.w2(32'h398772f4),
	.w3(32'h3a1ad1c2),
	.w4(32'h3b83a598),
	.w5(32'h3af8f6c8),
	.w6(32'h3a65c502),
	.w7(32'hba874544),
	.w8(32'hba8b5594),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e9e45),
	.w1(32'hb98f79b0),
	.w2(32'h3a53eb6b),
	.w3(32'h3b1a09ad),
	.w4(32'hbacc9c5a),
	.w5(32'h3982516d),
	.w6(32'hba5ba960),
	.w7(32'h3a0abc4b),
	.w8(32'h380d95e4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5619a),
	.w1(32'h39762c64),
	.w2(32'h3a2adbab),
	.w3(32'hba2a1c69),
	.w4(32'h3a4f3ead),
	.w5(32'hbb92935e),
	.w6(32'hbb6bf973),
	.w7(32'hbb8cb60a),
	.w8(32'hb98eb88e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadedd7e),
	.w1(32'hbb89fe27),
	.w2(32'h3adf5046),
	.w3(32'h39be4afd),
	.w4(32'hbba40966),
	.w5(32'hbab56015),
	.w6(32'hba34b26f),
	.w7(32'h3aea3243),
	.w8(32'h3bb29e49),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e0aa8),
	.w1(32'hbb643fc9),
	.w2(32'hba07a0c2),
	.w3(32'h39da58d5),
	.w4(32'hbba5b95b),
	.w5(32'h3b9b6d61),
	.w6(32'h3bbcf81f),
	.w7(32'h3c3ea92b),
	.w8(32'h3c274890),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3ced8),
	.w1(32'h3b4d53cb),
	.w2(32'h3ba4ff61),
	.w3(32'hbab207f8),
	.w4(32'hbb2c6ac7),
	.w5(32'h3ad5cbc6),
	.w6(32'h3a1ca039),
	.w7(32'hb99d4c50),
	.w8(32'h3aed5e45),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa97138),
	.w1(32'h3b91d9a6),
	.w2(32'h3c0ec6c2),
	.w3(32'hbac72a87),
	.w4(32'h3b23699a),
	.w5(32'h3be57431),
	.w6(32'h3aa3dd2f),
	.w7(32'hbb12fd97),
	.w8(32'h3bb47505),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d8e5a),
	.w1(32'h3a8b5ecf),
	.w2(32'h3a3e335c),
	.w3(32'h3a870560),
	.w4(32'hba8050e1),
	.w5(32'hba3517f3),
	.w6(32'h39a0137d),
	.w7(32'h39861976),
	.w8(32'hba8675ac),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829c4a6),
	.w1(32'h38b33373),
	.w2(32'hba07176b),
	.w3(32'hbab911f2),
	.w4(32'hba12a570),
	.w5(32'h38cb40ca),
	.w6(32'h3a596309),
	.w7(32'hb7470c68),
	.w8(32'h395af335),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba546241),
	.w1(32'h398f6b75),
	.w2(32'hba3aa62b),
	.w3(32'h371a0bb6),
	.w4(32'h3913e5a7),
	.w5(32'h38996bcc),
	.w6(32'h3a14c5d0),
	.w7(32'hb91cd600),
	.w8(32'hba551e71),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9176e1a),
	.w1(32'h3b1e4e97),
	.w2(32'h3b545a7c),
	.w3(32'hb8a41d47),
	.w4(32'hb9e1f00e),
	.w5(32'h3a945e01),
	.w6(32'h3ac8c398),
	.w7(32'h3ad1bf48),
	.w8(32'hba26e87d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9327d5),
	.w1(32'hb9855e1d),
	.w2(32'hba9ba895),
	.w3(32'hbaa8ec28),
	.w4(32'hba1efdf4),
	.w5(32'hbab18c92),
	.w6(32'hba777e45),
	.w7(32'hba204ccf),
	.w8(32'hba21f1d4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d7cc3),
	.w1(32'h3afd8064),
	.w2(32'h3a51f4e9),
	.w3(32'hba24b41a),
	.w4(32'hbbfde36e),
	.w5(32'h3b61ecd8),
	.w6(32'h3bbf4310),
	.w7(32'h3a535d93),
	.w8(32'hbbe82e9a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee0831),
	.w1(32'h3ac6c70d),
	.w2(32'h3a697aab),
	.w3(32'h399e2885),
	.w4(32'hbad589de),
	.w5(32'hba504206),
	.w6(32'hbb3c7b01),
	.w7(32'hbbc8f35b),
	.w8(32'hbb9fa793),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64016e),
	.w1(32'hbb96ae23),
	.w2(32'hba9b2a3e),
	.w3(32'hbb2bfc12),
	.w4(32'hbbc96bd1),
	.w5(32'hbb1ac707),
	.w6(32'hbb8d683f),
	.w7(32'hbb81113d),
	.w8(32'hbb845411),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf901c),
	.w1(32'hbab80de6),
	.w2(32'h3bee0dc5),
	.w3(32'hbb4ac7c9),
	.w4(32'hbb47b4a5),
	.w5(32'h3bad4d61),
	.w6(32'hba33b4b8),
	.w7(32'h3bfbdb4e),
	.w8(32'hbad044e9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0717ee),
	.w1(32'hbb4a587b),
	.w2(32'hbb3a7b8c),
	.w3(32'hbb15b72f),
	.w4(32'hbb4e642f),
	.w5(32'hb9c8596d),
	.w6(32'hbb188054),
	.w7(32'hba9c76cb),
	.w8(32'hba928bfe),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698336),
	.w1(32'hbc06d66d),
	.w2(32'hbb9598ee),
	.w3(32'hbb63e89c),
	.w4(32'hbbe0db66),
	.w5(32'hb981d542),
	.w6(32'h3bbe3b50),
	.w7(32'h3c060a87),
	.w8(32'h3c3830ad),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f58903),
	.w1(32'hbae2e496),
	.w2(32'hbab1cf72),
	.w3(32'hb9d38bfa),
	.w4(32'hbb95fb2b),
	.w5(32'hbb6388be),
	.w6(32'hbb9130cf),
	.w7(32'hbbcb08ca),
	.w8(32'hbbb70971),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6347d0),
	.w1(32'hb9e2594f),
	.w2(32'h3b13ee92),
	.w3(32'hbacb25dd),
	.w4(32'hbb34ef3d),
	.w5(32'hb957c270),
	.w6(32'h3a839aa9),
	.w7(32'h3b02ef83),
	.w8(32'h3ae4646e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36aa01),
	.w1(32'hba182b86),
	.w2(32'hb98c9208),
	.w3(32'hb968ae13),
	.w4(32'hba10dec5),
	.w5(32'hbada1ba9),
	.w6(32'hba42658c),
	.w7(32'h39d97649),
	.w8(32'h39f991ca),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24cda7),
	.w1(32'h3c1ae4fb),
	.w2(32'h3c5af666),
	.w3(32'hba395fdf),
	.w4(32'hbb809a81),
	.w5(32'hb86db0a8),
	.w6(32'h3c14ca5e),
	.w7(32'h3c11efeb),
	.w8(32'h3c0a5336),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77afdb),
	.w1(32'hbb091a5d),
	.w2(32'h3a073601),
	.w3(32'hbafa76e5),
	.w4(32'hbb49668c),
	.w5(32'hba2eb1d7),
	.w6(32'hb91985be),
	.w7(32'h3ab122fe),
	.w8(32'h3b4739d8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab36c29),
	.w1(32'h399d356b),
	.w2(32'hbaec6926),
	.w3(32'h3a993dbd),
	.w4(32'hb97ed597),
	.w5(32'h3a7e1298),
	.w6(32'h3aa38b2d),
	.w7(32'hba652483),
	.w8(32'hbb3bcaf5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a515edf),
	.w1(32'hba95697c),
	.w2(32'hb9565069),
	.w3(32'hbab29221),
	.w4(32'hbaef31ea),
	.w5(32'h3982c61f),
	.w6(32'h3a380066),
	.w7(32'h3a476d39),
	.w8(32'h38b666a6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75362a),
	.w1(32'hbb91ee60),
	.w2(32'hbb2c9ecc),
	.w3(32'hbb6aa7ef),
	.w4(32'hbba3f199),
	.w5(32'hbaae7fa8),
	.w6(32'hba9ab6ee),
	.w7(32'h3ab8f9ea),
	.w8(32'h3b312c4e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a440460),
	.w1(32'hbb3cb408),
	.w2(32'hbab171b8),
	.w3(32'hbb2c6533),
	.w4(32'hbb8eda0d),
	.w5(32'hbabb7002),
	.w6(32'hbbbc43c1),
	.w7(32'hbb8f3eb8),
	.w8(32'hbb932923),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5223dc),
	.w1(32'h3b1151bc),
	.w2(32'h3b902278),
	.w3(32'hbadb94d6),
	.w4(32'hba92d8d7),
	.w5(32'h3aee1f90),
	.w6(32'h3b0c1ee8),
	.w7(32'h3b06710b),
	.w8(32'h3b6f5f13),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c4fcf),
	.w1(32'h3b0728e8),
	.w2(32'h3b84bf3f),
	.w3(32'hbaa0342c),
	.w4(32'hbb627b54),
	.w5(32'h3990dd24),
	.w6(32'hbb00e052),
	.w7(32'hb9b530ea),
	.w8(32'h391a9a81),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbc394),
	.w1(32'hbaae1ee6),
	.w2(32'hba06f7af),
	.w3(32'hbabccdb4),
	.w4(32'hbb6badf4),
	.w5(32'hbac868d2),
	.w6(32'h39b51816),
	.w7(32'hb99a7f78),
	.w8(32'h3b17dd16),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38829492),
	.w1(32'hbbd0eabf),
	.w2(32'hbb1c9bc9),
	.w3(32'hbb53fd59),
	.w4(32'hbbbd1e90),
	.w5(32'h3a80a7c9),
	.w6(32'h3b76c038),
	.w7(32'h3c08a12b),
	.w8(32'h3c624962),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa39d13),
	.w1(32'hb9ada7b7),
	.w2(32'h3b81b0ef),
	.w3(32'h3b01aa46),
	.w4(32'hbb09d9d8),
	.w5(32'hbaab6c56),
	.w6(32'h392e249b),
	.w7(32'h3ac9b218),
	.w8(32'h3afca8ae),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78e851),
	.w1(32'hba175a27),
	.w2(32'h3a181422),
	.w3(32'hbb3e7b0f),
	.w4(32'h388be206),
	.w5(32'hb9192e44),
	.w6(32'hba057f94),
	.w7(32'hbac87d95),
	.w8(32'h3aa7c677),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bdb44),
	.w1(32'hbb4adaf1),
	.w2(32'h3b5b6764),
	.w3(32'h3a3e6510),
	.w4(32'hbae48d67),
	.w5(32'h3bfd8553),
	.w6(32'h39e72a25),
	.w7(32'h3baa41ef),
	.w8(32'h395bc2b5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5003c2),
	.w1(32'h3a361110),
	.w2(32'hb9ee3f77),
	.w3(32'hbb79ae98),
	.w4(32'hb7d37f2e),
	.w5(32'hb9d3ce32),
	.w6(32'hbb2a6e06),
	.w7(32'hbb3d0d5f),
	.w8(32'hbbbded62),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34fa52),
	.w1(32'h3b69c316),
	.w2(32'h3b98cded),
	.w3(32'hb9eff7c7),
	.w4(32'hba88b07b),
	.w5(32'h3ae9ba8a),
	.w6(32'h3b41c6c5),
	.w7(32'h3b34d9e5),
	.w8(32'h3b8a40a1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f3f77),
	.w1(32'hb97254e2),
	.w2(32'h3ae6bd01),
	.w3(32'hbae05ca6),
	.w4(32'hbb6663a8),
	.w5(32'hb9816530),
	.w6(32'hbbbc55db),
	.w7(32'hbb5670cb),
	.w8(32'hb998de8f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6405ac),
	.w1(32'h3c356f9c),
	.w2(32'h3c95e1cc),
	.w3(32'h3ab8adca),
	.w4(32'h3ad532a6),
	.w5(32'h3b6137a7),
	.w6(32'h3c2e1b17),
	.w7(32'h3c3650e8),
	.w8(32'h3c6b2884),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad421c),
	.w1(32'hbbe6b0f9),
	.w2(32'hba48fe05),
	.w3(32'hbbaa49b8),
	.w4(32'hbb3cfcd4),
	.w5(32'hba029c54),
	.w6(32'hbba82455),
	.w7(32'hbbd248e6),
	.w8(32'hbac80dd4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2a14),
	.w1(32'h3a4356b9),
	.w2(32'hb91d1812),
	.w3(32'hba763f2c),
	.w4(32'h3aac1c89),
	.w5(32'h3b28a915),
	.w6(32'hbaf12685),
	.w7(32'hbb71eba2),
	.w8(32'h394e6dbd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00803e),
	.w1(32'hba39fc07),
	.w2(32'hb9cd8328),
	.w3(32'hb9b3d3b8),
	.w4(32'hbb49dfaa),
	.w5(32'hbac60e56),
	.w6(32'hba162bed),
	.w7(32'h38061daa),
	.w8(32'hba815895),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74eda8),
	.w1(32'h392b390e),
	.w2(32'hbb012586),
	.w3(32'hba1402b0),
	.w4(32'hb9a65a4b),
	.w5(32'h39d9520d),
	.w6(32'hbb5abbee),
	.w7(32'hbb7ecc90),
	.w8(32'hba6a1e99),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b63bcc),
	.w1(32'h3ab2971c),
	.w2(32'h3a75d5dd),
	.w3(32'h3a99fadb),
	.w4(32'h37dba4ea),
	.w5(32'h3a3c6fa3),
	.w6(32'h3a8e2ef2),
	.w7(32'h3ae98b0e),
	.w8(32'hba1bb5fd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba172a3d),
	.w1(32'hb951d464),
	.w2(32'h3b66deda),
	.w3(32'hb9f9cb3f),
	.w4(32'hbb300e86),
	.w5(32'hbb27a834),
	.w6(32'hb910e0ff),
	.w7(32'h39d1421d),
	.w8(32'h3a199b67),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c62c7),
	.w1(32'h3a68948f),
	.w2(32'h3ab764fa),
	.w3(32'hbb2ac405),
	.w4(32'hba876ed2),
	.w5(32'h3ab5d779),
	.w6(32'h397f7e7e),
	.w7(32'h3afebc45),
	.w8(32'hb8dca0c0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaecec),
	.w1(32'hbb5aa62e),
	.w2(32'hbb0161f7),
	.w3(32'hbbe99486),
	.w4(32'hbb0dd56a),
	.w5(32'h38df1c8a),
	.w6(32'hbba27bab),
	.w7(32'hbbd184c0),
	.w8(32'hbb77d306),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dba28),
	.w1(32'hbb526f79),
	.w2(32'hb9b6697c),
	.w3(32'hbb454c2a),
	.w4(32'hbb563ecb),
	.w5(32'hb8d99665),
	.w6(32'hbb890b8c),
	.w7(32'hbb2a7426),
	.w8(32'hbb05451e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b175f7c),
	.w1(32'h3b04806b),
	.w2(32'h3a83b254),
	.w3(32'h393b8427),
	.w4(32'hb9824d71),
	.w5(32'h37afa721),
	.w6(32'h3b4bb566),
	.w7(32'h3b39b777),
	.w8(32'h3acdd05d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc07f2),
	.w1(32'hbb347b0b),
	.w2(32'hbb71bf13),
	.w3(32'hbb15c41e),
	.w4(32'hbae46a95),
	.w5(32'hbab5cc4d),
	.w6(32'h3a39acd0),
	.w7(32'h3b09bce3),
	.w8(32'hba693ed8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91caddd),
	.w1(32'h3abadb30),
	.w2(32'h3b32ea51),
	.w3(32'hb933e06f),
	.w4(32'hbb22144b),
	.w5(32'hba066409),
	.w6(32'hbac78427),
	.w7(32'hbabd3414),
	.w8(32'hb9bd4b45),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6cb7),
	.w1(32'hbbc5689b),
	.w2(32'hbb27dfcd),
	.w3(32'hbb053b42),
	.w4(32'hbba7e2b0),
	.w5(32'hbb601cbe),
	.w6(32'hbb83cc88),
	.w7(32'hbbb508f9),
	.w8(32'hbba96567),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cca71),
	.w1(32'hbac5def4),
	.w2(32'hbaaa924f),
	.w3(32'hbbc01737),
	.w4(32'hbb1c5b1a),
	.w5(32'hbb00a948),
	.w6(32'hb896e34a),
	.w7(32'hb8be20cc),
	.w8(32'hba0c2041),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0275a),
	.w1(32'h3ab81bde),
	.w2(32'hba7ddbc1),
	.w3(32'hba95264c),
	.w4(32'h3b3881a2),
	.w5(32'h3a8dc56f),
	.w6(32'h3af1e3a2),
	.w7(32'hba12f885),
	.w8(32'h3a0d4186),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d9ae5),
	.w1(32'h39eb3946),
	.w2(32'hb9e1b496),
	.w3(32'h3a846e43),
	.w4(32'h39fe4a89),
	.w5(32'h3a232363),
	.w6(32'h3a5198b1),
	.w7(32'hb97b9c36),
	.w8(32'h397a98d1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0bfb9),
	.w1(32'h39d6d956),
	.w2(32'hba663525),
	.w3(32'h39199ba7),
	.w4(32'h3a5a792a),
	.w5(32'h39f6d9af),
	.w6(32'h39e45795),
	.w7(32'hba45f566),
	.w8(32'hb980db66),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b09ba),
	.w1(32'hbb12ec90),
	.w2(32'h3b7888d4),
	.w3(32'h38df40c0),
	.w4(32'h3a78067e),
	.w5(32'hba0f6f0d),
	.w6(32'hbb3ff182),
	.w7(32'hbb8a202c),
	.w8(32'hba8f10b1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b265e),
	.w1(32'h38e4ae7b),
	.w2(32'h3b3eb3c8),
	.w3(32'hbba8f96c),
	.w4(32'hbb3cff0f),
	.w5(32'hbb1c554f),
	.w6(32'hbaae6a7a),
	.w7(32'hb9d57e20),
	.w8(32'hbb907757),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f1cd1),
	.w1(32'h3b02debe),
	.w2(32'h3adc24f0),
	.w3(32'hbaff8f27),
	.w4(32'hb949d5d2),
	.w5(32'h39d31ec5),
	.w6(32'h3ada5b31),
	.w7(32'h3b241bfe),
	.w8(32'h3ac3d8d8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6cd2c),
	.w1(32'h39b5ed58),
	.w2(32'h3832ca89),
	.w3(32'h3aaf1014),
	.w4(32'h39d9072f),
	.w5(32'h3a24ef11),
	.w6(32'hba9c62ce),
	.w7(32'hba86c7e3),
	.w8(32'hba5cbb90),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013c73),
	.w1(32'h39e456ca),
	.w2(32'h398fb45d),
	.w3(32'hba68069b),
	.w4(32'hb9dce457),
	.w5(32'h39b7b64d),
	.w6(32'h3ab4ace6),
	.w7(32'hb7aa8b91),
	.w8(32'h3a8cbb6c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba407321),
	.w1(32'hbb542d21),
	.w2(32'hbb4848e9),
	.w3(32'hb813184d),
	.w4(32'h39f66b34),
	.w5(32'hbb3e3e38),
	.w6(32'hbb9082cc),
	.w7(32'hbb616100),
	.w8(32'hb91dd5cc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc101d29),
	.w1(32'hba2a5fe3),
	.w2(32'hbb5ca328),
	.w3(32'hbb522307),
	.w4(32'hbb53c655),
	.w5(32'hbac2cc37),
	.w6(32'h398bf7c2),
	.w7(32'h39ada4d7),
	.w8(32'h3b485150),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae140cb),
	.w1(32'hba3c7d0d),
	.w2(32'hbab245aa),
	.w3(32'hbaaef536),
	.w4(32'hbabc5011),
	.w5(32'h3a3be798),
	.w6(32'h394dfe3d),
	.w7(32'h395353cb),
	.w8(32'hba17e2c5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9230dca),
	.w1(32'hb9cb8cac),
	.w2(32'hb98a54d0),
	.w3(32'hba4f8e22),
	.w4(32'hba22703f),
	.w5(32'hb9d9ed17),
	.w6(32'hba05097e),
	.w7(32'hba3715fa),
	.w8(32'hb892f883),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5d0e4),
	.w1(32'hba7daaae),
	.w2(32'h38267ad9),
	.w3(32'hbb3d4cde),
	.w4(32'hbb2321ce),
	.w5(32'hbad692e5),
	.w6(32'hbbad49a1),
	.w7(32'hbb9bc585),
	.w8(32'hbb80ede8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac403c0),
	.w1(32'hbb0741dc),
	.w2(32'hbabb8cb1),
	.w3(32'hba4aa1ce),
	.w4(32'hba998dd2),
	.w5(32'hba8bfa8b),
	.w6(32'hbb1c4ce5),
	.w7(32'hbb70687a),
	.w8(32'hbb6a2e2e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921dfb5),
	.w1(32'h3984dbc6),
	.w2(32'h399a75d6),
	.w3(32'h3a4d7248),
	.w4(32'h3917d996),
	.w5(32'h38f9abec),
	.w6(32'hb9a33a26),
	.w7(32'hb966bd19),
	.w8(32'hb9107196),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39d293),
	.w1(32'h39b5f97e),
	.w2(32'h3a5a9320),
	.w3(32'hba2579c6),
	.w4(32'hba6300cc),
	.w5(32'hb8c43dd6),
	.w6(32'hb95828ba),
	.w7(32'hb9e45ed1),
	.w8(32'h395ab3e0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c3886),
	.w1(32'hba35c85e),
	.w2(32'hba04f4e6),
	.w3(32'hb99df20d),
	.w4(32'hb9fb7364),
	.w5(32'hb9f4f52b),
	.w6(32'h383169fa),
	.w7(32'hb8806b3b),
	.w8(32'h399ab1e4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86cd73),
	.w1(32'hbacf485e),
	.w2(32'hba78933e),
	.w3(32'hbae96932),
	.w4(32'hbb06a335),
	.w5(32'hba838be6),
	.w6(32'hbb0f7ce7),
	.w7(32'hbb35c5e1),
	.w8(32'hbaeb4005),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca94bc),
	.w1(32'hb9f3c0f0),
	.w2(32'hb984cc27),
	.w3(32'h3922e332),
	.w4(32'hba5f7aad),
	.w5(32'hba2aae10),
	.w6(32'h39649d63),
	.w7(32'hba18de3e),
	.w8(32'h3a08d6d5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffb7c2),
	.w1(32'hb9c7f8cc),
	.w2(32'h396d7e10),
	.w3(32'hba4cdfe3),
	.w4(32'hbab85471),
	.w5(32'hba3b7ab6),
	.w6(32'hbb627cba),
	.w7(32'hbb6494e2),
	.w8(32'hbb20b45d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05333b),
	.w1(32'hbb0f1d65),
	.w2(32'hba71519d),
	.w3(32'hbb05cac5),
	.w4(32'hbace8274),
	.w5(32'h395a1737),
	.w6(32'hbaad1c40),
	.w7(32'hbab7b687),
	.w8(32'hb9b0f0bd),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba8b3c),
	.w1(32'hba843716),
	.w2(32'hba5f9c97),
	.w3(32'hba85ffdd),
	.w4(32'hbacc9263),
	.w5(32'hba8a4651),
	.w6(32'hba8a5876),
	.w7(32'hba00c9f9),
	.w8(32'hb9a2418d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29bbb6),
	.w1(32'hbb081339),
	.w2(32'hbabe2f10),
	.w3(32'hbb4da2d6),
	.w4(32'hbb768227),
	.w5(32'hb9ce081c),
	.w6(32'hbba79e78),
	.w7(32'hbbbe9fef),
	.w8(32'hbb5dee87),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cbfad),
	.w1(32'hb9fa425b),
	.w2(32'h397f362c),
	.w3(32'hbaa73970),
	.w4(32'hba8657d5),
	.w5(32'h37ea0af6),
	.w6(32'hba8b9df3),
	.w7(32'hb9b0a9a7),
	.w8(32'h3a06eb4e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13dcfa),
	.w1(32'hbae467b9),
	.w2(32'hb984b32e),
	.w3(32'hbaf04da5),
	.w4(32'hbaa6cf6d),
	.w5(32'h398802f3),
	.w6(32'hb9b3616b),
	.w7(32'hba52bbe1),
	.w8(32'hb9501988),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1063cd),
	.w1(32'hbac3ad6c),
	.w2(32'hba556675),
	.w3(32'hbab4b63a),
	.w4(32'hbac41bc7),
	.w5(32'hba6455ce),
	.w6(32'hbac403d3),
	.w7(32'hbade652f),
	.w8(32'hbaa372c9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba552a0c),
	.w1(32'hbafc2ee1),
	.w2(32'hba82a659),
	.w3(32'hba1deb57),
	.w4(32'hba6e2317),
	.w5(32'h3a18c76c),
	.w6(32'h3b11f658),
	.w7(32'h3a15b56e),
	.w8(32'h3ab2083c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802c0bd),
	.w1(32'h39a6074e),
	.w2(32'hb9b95452),
	.w3(32'h391ea1db),
	.w4(32'hb998ec6f),
	.w5(32'hbab7e68e),
	.w6(32'h3aa0df46),
	.w7(32'h3aa75131),
	.w8(32'h3a110768),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d1a06),
	.w1(32'h375101b9),
	.w2(32'h378c45e2),
	.w3(32'h38845a63),
	.w4(32'h3904774d),
	.w5(32'h38bcb175),
	.w6(32'hb8a740db),
	.w7(32'hb8a6b761),
	.w8(32'h38074caf),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39159971),
	.w1(32'hb89c3e4f),
	.w2(32'hb9b0331a),
	.w3(32'h390ce733),
	.w4(32'hb8c283cf),
	.w5(32'hb9e63b23),
	.w6(32'hb9c4f1b0),
	.w7(32'hb991523e),
	.w8(32'hb9d38144),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b81ea9),
	.w1(32'h38e702c4),
	.w2(32'hb996e068),
	.w3(32'hb914e9e7),
	.w4(32'h39238eb9),
	.w5(32'hb6969d72),
	.w6(32'hb8d68d51),
	.w7(32'h3a0a6314),
	.w8(32'h396bb89d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0a6dc),
	.w1(32'h39d540a7),
	.w2(32'h3a5ff992),
	.w3(32'h3ac06baf),
	.w4(32'h3a4ee910),
	.w5(32'h3aa06531),
	.w6(32'h3b268b6c),
	.w7(32'h3b468be9),
	.w8(32'h3b355ac6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70003b),
	.w1(32'hbb78e312),
	.w2(32'hba6f6bce),
	.w3(32'hbbc8f483),
	.w4(32'hbb94e44f),
	.w5(32'hbb234862),
	.w6(32'hbc051d47),
	.w7(32'hbbe8733e),
	.w8(32'hbbaa4b2c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9839a07),
	.w1(32'hba1ac6be),
	.w2(32'hba1f4198),
	.w3(32'hb9623285),
	.w4(32'hb992c4d9),
	.w5(32'hb9c53d68),
	.w6(32'hb9a4ccec),
	.w7(32'hb99cf6f2),
	.w8(32'hb8630142),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c9583),
	.w1(32'hbb3b650a),
	.w2(32'hbaea78d0),
	.w3(32'hbb1f6ef7),
	.w4(32'hbb0a9c2e),
	.w5(32'hba2543f5),
	.w6(32'hbb3ce647),
	.w7(32'hbb63a24b),
	.w8(32'hbb3067e3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41aed5),
	.w1(32'hbb17abc0),
	.w2(32'hbaab6b03),
	.w3(32'hbac67974),
	.w4(32'hba5faa29),
	.w5(32'h39d681e3),
	.w6(32'hbaae7cb1),
	.w7(32'hba22e377),
	.w8(32'h3a04adab),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf3cc3),
	.w1(32'hba6f5617),
	.w2(32'hba6410ad),
	.w3(32'hbaec9e94),
	.w4(32'hbb0fcf81),
	.w5(32'hba109eae),
	.w6(32'hbb62b1a1),
	.w7(32'hbb7daa26),
	.w8(32'hbb279b8a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac73480),
	.w1(32'h3a60d661),
	.w2(32'h3a79808c),
	.w3(32'h3a7fc122),
	.w4(32'h391a9cb1),
	.w5(32'h3a1cef96),
	.w6(32'h3b2a4dfb),
	.w7(32'h3a9c8fdd),
	.w8(32'h3b331cd7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab124ff),
	.w1(32'h3aa47baf),
	.w2(32'h3a909b77),
	.w3(32'h3a4b5f96),
	.w4(32'h3a6f9a01),
	.w5(32'h3a5c547f),
	.w6(32'h3a3247d7),
	.w7(32'h3acb14e5),
	.w8(32'h3ad00be6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c63995),
	.w1(32'hbabbfc86),
	.w2(32'hba511845),
	.w3(32'hba165ec9),
	.w4(32'hbae9579e),
	.w5(32'hbaef019b),
	.w6(32'hbae0c7c2),
	.w7(32'hbb2677c2),
	.w8(32'hbab2af0d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39db72),
	.w1(32'hbae28608),
	.w2(32'hba35963b),
	.w3(32'hbb015bc7),
	.w4(32'hba68de14),
	.w5(32'h3a4fc099),
	.w6(32'hb95341f2),
	.w7(32'h398e0b28),
	.w8(32'h3acb1536),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8a86f),
	.w1(32'h3a552b42),
	.w2(32'h3b082753),
	.w3(32'h39a2fc11),
	.w4(32'h398bcdec),
	.w5(32'h3aa69388),
	.w6(32'h3ab8dc40),
	.w7(32'h3b0e15a1),
	.w8(32'h3b8d4ca7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82b087),
	.w1(32'h379e4e97),
	.w2(32'h3aacf2fd),
	.w3(32'hba52cad1),
	.w4(32'hb9e029ba),
	.w5(32'h3a6521f6),
	.w6(32'h3a8a6c9d),
	.w7(32'h3a42ac08),
	.w8(32'h3ae70487),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c5f6bf),
	.w1(32'hb9d8a115),
	.w2(32'hb9a6c586),
	.w3(32'hb9607d27),
	.w4(32'hba1d9fb3),
	.w5(32'hba21511e),
	.w6(32'hba8c0308),
	.w7(32'hbaa04340),
	.w8(32'hba62581c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0df1a),
	.w1(32'hb9c4c50a),
	.w2(32'hba00e0fe),
	.w3(32'hb99e3591),
	.w4(32'hb9c9e26d),
	.w5(32'hb9e5376a),
	.w6(32'hba0a6bbd),
	.w7(32'hba01b036),
	.w8(32'hb9c0e863),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d1f3d),
	.w1(32'h3ada0173),
	.w2(32'h3ae58581),
	.w3(32'h38c6e77a),
	.w4(32'hb83c1e7f),
	.w5(32'h3a536981),
	.w6(32'hb9de7156),
	.w7(32'hba829bf8),
	.w8(32'hb9f3b2ad),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e7834),
	.w1(32'hba112445),
	.w2(32'hb8553c4f),
	.w3(32'hba15e3e6),
	.w4(32'hba17a8f6),
	.w5(32'hba378344),
	.w6(32'hb95b4868),
	.w7(32'hb90c7c85),
	.w8(32'hb81dc284),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2cf1),
	.w1(32'hbb0fb56d),
	.w2(32'hbad0b11d),
	.w3(32'hbb191b86),
	.w4(32'hbb1116ae),
	.w5(32'hb9e492ee),
	.w6(32'hb9bf3d11),
	.w7(32'hbac72b15),
	.w8(32'hba667da3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34a3e0),
	.w1(32'hb9e20bf3),
	.w2(32'hb98f2e6f),
	.w3(32'h3a38eb38),
	.w4(32'hba3f3784),
	.w5(32'hba09fe19),
	.w6(32'hba46d805),
	.w7(32'hba770b1a),
	.w8(32'hb9d12450),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d27a3),
	.w1(32'h3a798105),
	.w2(32'h3b5e0214),
	.w3(32'hba9e193e),
	.w4(32'hba5ae956),
	.w5(32'h3ac6d480),
	.w6(32'hba7ac2b0),
	.w7(32'hb981f8a1),
	.w8(32'h3abdf4a5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04e5a3),
	.w1(32'hb9631584),
	.w2(32'hb89bb9a1),
	.w3(32'h39eb13aa),
	.w4(32'hb9a95025),
	.w5(32'hb8ddc377),
	.w6(32'hb7527624),
	.w7(32'hb99352fd),
	.w8(32'hb85e26c8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b079e),
	.w1(32'hb937ee64),
	.w2(32'h38db9cf2),
	.w3(32'hb9247c9d),
	.w4(32'hb99ec8c7),
	.w5(32'h37c4dc3d),
	.w6(32'hb98bfa3c),
	.w7(32'hb98f21c8),
	.w8(32'h3961cd83),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce20d),
	.w1(32'hbae98cf3),
	.w2(32'hb9bd8cb5),
	.w3(32'hba5d8bb3),
	.w4(32'hbadea68b),
	.w5(32'h398d5c30),
	.w6(32'hb9912dec),
	.w7(32'hba39d87e),
	.w8(32'h3a816b10),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5bed),
	.w1(32'hbb5e53a7),
	.w2(32'hbae4428b),
	.w3(32'hbb066f23),
	.w4(32'hbb2ee1d4),
	.w5(32'hbae03e7e),
	.w6(32'hbb483d73),
	.w7(32'hbae33e27),
	.w8(32'hbacd9367),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43c945),
	.w1(32'h3a2e1929),
	.w2(32'h3b30a555),
	.w3(32'hbad13e12),
	.w4(32'hba42346b),
	.w5(32'h3a573b1c),
	.w6(32'hba009707),
	.w7(32'hba43c819),
	.w8(32'h3a5058ba),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e5cac),
	.w1(32'hbbacd118),
	.w2(32'hbb7794f1),
	.w3(32'hbb7739ae),
	.w4(32'hbb8a7219),
	.w5(32'hbaaf1ecb),
	.w6(32'hbb3a04f7),
	.w7(32'hbb7bf9f9),
	.w8(32'hbb34386b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a01f9),
	.w1(32'h3a0015ea),
	.w2(32'hb8f5a477),
	.w3(32'hba0e320f),
	.w4(32'h3a3005ec),
	.w5(32'hb861eb5f),
	.w6(32'h3ad0c06c),
	.w7(32'h3a89bda6),
	.w8(32'h3a481289),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943b742),
	.w1(32'hb9de4d6c),
	.w2(32'h3b05b999),
	.w3(32'hbac1f295),
	.w4(32'hbb04be72),
	.w5(32'h3808b65d),
	.w6(32'hba4e532c),
	.w7(32'hbb1a03bd),
	.w8(32'hba8cfe35),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068181),
	.w1(32'h3b09ca19),
	.w2(32'h3b85f6d2),
	.w3(32'h38576c98),
	.w4(32'hb9f18c34),
	.w5(32'h3a9e7eae),
	.w6(32'h397da801),
	.w7(32'hba68c567),
	.w8(32'h3ab381f6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a7c85),
	.w1(32'hbb3ce17c),
	.w2(32'hba739a58),
	.w3(32'hbb52e16b),
	.w4(32'hbb0d142b),
	.w5(32'hbaa04abe),
	.w6(32'hbb636579),
	.w7(32'hbb494800),
	.w8(32'hbb410601),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa38ff),
	.w1(32'hba65d0ef),
	.w2(32'hbad5b43d),
	.w3(32'h39106522),
	.w4(32'hba5b4153),
	.w5(32'hbaac2d60),
	.w6(32'hbac9c21e),
	.w7(32'hbab72c6b),
	.w8(32'hbab905fe),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf142a8),
	.w1(32'hbad8601b),
	.w2(32'hbaed3cfd),
	.w3(32'hba33322d),
	.w4(32'hba83d69e),
	.w5(32'hba852c58),
	.w6(32'hba0f1b8a),
	.w7(32'hba32a371),
	.w8(32'hba406529),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11b249),
	.w1(32'hb8c6ab8e),
	.w2(32'hb9a3bab6),
	.w3(32'hb9eb33b5),
	.w4(32'hb60ca962),
	.w5(32'hb9b01a59),
	.w6(32'hb7b91705),
	.w7(32'hb937053b),
	.w8(32'hb9244c83),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9807676),
	.w1(32'hb9a9bea8),
	.w2(32'h3987ef03),
	.w3(32'hba71ed8f),
	.w4(32'hba804f1f),
	.w5(32'hb98d2e6d),
	.w6(32'hb9cf7c76),
	.w7(32'hba5e4cce),
	.w8(32'h3935f16d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bfc24),
	.w1(32'h39ef64e0),
	.w2(32'h3abaab82),
	.w3(32'hba184806),
	.w4(32'h3a3a62aa),
	.w5(32'h3a8120e5),
	.w6(32'h39c7a582),
	.w7(32'h3924565c),
	.w8(32'h375f8dc5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad46447),
	.w1(32'h3987d1d9),
	.w2(32'h3a6df878),
	.w3(32'h39b565a3),
	.w4(32'hb707200a),
	.w5(32'h3a9671d5),
	.w6(32'hba223dcd),
	.w7(32'hba2e4352),
	.w8(32'h39e2f9c0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d7e59),
	.w1(32'h37417405),
	.w2(32'h3964ff63),
	.w3(32'h39e2ad0b),
	.w4(32'hb8b1258c),
	.w5(32'h39307b7e),
	.w6(32'h38882094),
	.w7(32'h39918ebc),
	.w8(32'h3894eb01),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e730d),
	.w1(32'h3a111063),
	.w2(32'h39e74ce2),
	.w3(32'h39d6ca5b),
	.w4(32'h399a45e9),
	.w5(32'h39ebb4f0),
	.w6(32'h3920e744),
	.w7(32'h3994af48),
	.w8(32'h3937c9fd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951d2d3),
	.w1(32'hba9fef54),
	.w2(32'hbab60d08),
	.w3(32'hba046f6d),
	.w4(32'hbacfb9af),
	.w5(32'hbacb09c1),
	.w6(32'hbabc1d4f),
	.w7(32'hbb03641f),
	.w8(32'hbac0b5ad),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cda28),
	.w1(32'h3ab7c67a),
	.w2(32'h3b1e1247),
	.w3(32'hba80ce54),
	.w4(32'h3a02dec3),
	.w5(32'h3b282f39),
	.w6(32'hb6b53b2e),
	.w7(32'h395c3395),
	.w8(32'h3b08f32b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b029e),
	.w1(32'hb965ffbc),
	.w2(32'hba034ee9),
	.w3(32'h3a185682),
	.w4(32'h39e3fde6),
	.w5(32'h389e5c6d),
	.w6(32'hbad51311),
	.w7(32'hba1c9ddc),
	.w8(32'h38604c4f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5224e),
	.w1(32'h39ad24f2),
	.w2(32'h3a830269),
	.w3(32'hb9d566f7),
	.w4(32'hb90d892e),
	.w5(32'h3a008ffc),
	.w6(32'hb968dfa4),
	.w7(32'hb7b44010),
	.w8(32'h3806827b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85fcc1),
	.w1(32'hbb760b5e),
	.w2(32'hba230ec1),
	.w3(32'hbbe34cad),
	.w4(32'hbb84a79a),
	.w5(32'hba8e761f),
	.w6(32'hbc23f561),
	.w7(32'hbbfc42f1),
	.w8(32'hbbba3772),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae61015),
	.w1(32'h3b0874fe),
	.w2(32'h3a8127b3),
	.w3(32'h3ab8f867),
	.w4(32'h3a9e39d3),
	.w5(32'h3ab089cf),
	.w6(32'h3b76c792),
	.w7(32'h3b671bb4),
	.w8(32'h3b447f4a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390489e8),
	.w1(32'hb98ebd1f),
	.w2(32'hb963b6cb),
	.w3(32'hb94fdef8),
	.w4(32'hb9c58ea6),
	.w5(32'hb94113ce),
	.w6(32'hba1fc027),
	.w7(32'hba6a0694),
	.w8(32'hba1d829f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa8bda),
	.w1(32'h3a800055),
	.w2(32'h39e6d2f4),
	.w3(32'hb9332136),
	.w4(32'h3ab97be3),
	.w5(32'h3a43d381),
	.w6(32'h3a12e66c),
	.w7(32'h38d0c5e4),
	.w8(32'hba814f21),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fee195),
	.w1(32'h3a9bfa36),
	.w2(32'h3a95610e),
	.w3(32'hba0597a8),
	.w4(32'h3a8319f9),
	.w5(32'h3a905446),
	.w6(32'h3a4e6cc1),
	.w7(32'h3a68bd4c),
	.w8(32'h3a9c742c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398641db),
	.w1(32'h3825537b),
	.w2(32'hb845ff3f),
	.w3(32'h3a01d863),
	.w4(32'h38395494),
	.w5(32'hb8068931),
	.w6(32'h391b3c3d),
	.w7(32'hb873ab86),
	.w8(32'h392eb326),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d785d5),
	.w1(32'h37b31b2d),
	.w2(32'h39f0afab),
	.w3(32'hb8401cce),
	.w4(32'hb96ea851),
	.w5(32'h362858f0),
	.w6(32'hba9095aa),
	.w7(32'hba34e765),
	.w8(32'hb9badd4e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a528de3),
	.w1(32'hbb18f145),
	.w2(32'hbae0d71a),
	.w3(32'hbaf0db4f),
	.w4(32'hbb8ae089),
	.w5(32'hbb157ee7),
	.w6(32'hb9397479),
	.w7(32'hba8d08af),
	.w8(32'hbaa56f3b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1396d5),
	.w1(32'hbb09e537),
	.w2(32'hbab01cb8),
	.w3(32'hbb5a5208),
	.w4(32'hbb0219e2),
	.w5(32'hbaad0f26),
	.w6(32'hbb24c689),
	.w7(32'hbb00eda9),
	.w8(32'hba9e8778),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba707623),
	.w1(32'hba539da0),
	.w2(32'h394eda65),
	.w3(32'hbab40415),
	.w4(32'hbab90da0),
	.w5(32'hb88ddd17),
	.w6(32'hb8d6d53a),
	.w7(32'hb9e629d7),
	.w8(32'h3a053eae),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7470ed),
	.w1(32'h37059da3),
	.w2(32'h3b21f3a9),
	.w3(32'hbb375bab),
	.w4(32'hbac71beb),
	.w5(32'h3b1ad72d),
	.w6(32'hbb6c60b4),
	.w7(32'hbb3724c3),
	.w8(32'h39931cc2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965215b),
	.w1(32'hb9ae610a),
	.w2(32'h38bc6909),
	.w3(32'hba442e63),
	.w4(32'hb9e44404),
	.w5(32'h39052505),
	.w6(32'hba5233e2),
	.w7(32'hba39e4a3),
	.w8(32'hb75653af),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39667949),
	.w1(32'hb928aac3),
	.w2(32'hb9150d11),
	.w3(32'h398cc98e),
	.w4(32'h378e7930),
	.w5(32'hb8a84655),
	.w6(32'hb8c72a06),
	.w7(32'hb89c56e1),
	.w8(32'h38b4f558),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38788005),
	.w1(32'hba8a6f32),
	.w2(32'hba5547f9),
	.w3(32'h38d8e703),
	.w4(32'hb8b78964),
	.w5(32'hb8a33c57),
	.w6(32'hba453e32),
	.w7(32'hba1468aa),
	.w8(32'hba031bc4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddb112),
	.w1(32'hba2e789d),
	.w2(32'hba58002f),
	.w3(32'h3980ea56),
	.w4(32'hb9d2ad77),
	.w5(32'hba282393),
	.w6(32'hba1ce69e),
	.w7(32'hba185a40),
	.w8(32'hba0114d0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b75bd),
	.w1(32'h3a82e5bd),
	.w2(32'h3abf8705),
	.w3(32'hba84f0f3),
	.w4(32'hb99b5636),
	.w5(32'h391eb3d7),
	.w6(32'hba74737a),
	.w7(32'hba96411c),
	.w8(32'hba0e5094),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab54867),
	.w1(32'h3baa36d8),
	.w2(32'h3c0ed083),
	.w3(32'hb910e651),
	.w4(32'h3aee10b0),
	.w5(32'h3b846ed4),
	.w6(32'h3b3bfe97),
	.w7(32'h3b8b73cd),
	.w8(32'h3bcfe301),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886e275),
	.w1(32'hb9a23015),
	.w2(32'h3aac376c),
	.w3(32'hbad203b8),
	.w4(32'hb9e15e39),
	.w5(32'h3abd7f05),
	.w6(32'hb884b519),
	.w7(32'h388a11f9),
	.w8(32'h3b24af7e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5d84b),
	.w1(32'h3a2f2e46),
	.w2(32'h3ab519bd),
	.w3(32'hb963c22d),
	.w4(32'h39c87993),
	.w5(32'h3a86c8c8),
	.w6(32'h3a004fad),
	.w7(32'h3a095643),
	.w8(32'h3a39a595),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbf8ba),
	.w1(32'hba5362cd),
	.w2(32'hb7e41177),
	.w3(32'hbad04158),
	.w4(32'hba1e2e2d),
	.w5(32'h394fb502),
	.w6(32'h3956a460),
	.w7(32'h38d937ff),
	.w8(32'h3a4f24c9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e85f5),
	.w1(32'hbb4a044f),
	.w2(32'hbb03da65),
	.w3(32'hbb0c6e6e),
	.w4(32'hbb367b60),
	.w5(32'hbaacfbf7),
	.w6(32'hbb5d932b),
	.w7(32'hbb6137f6),
	.w8(32'hbb13c039),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb765fd0),
	.w1(32'hbb8991c8),
	.w2(32'hbb2d065c),
	.w3(32'hbb748f20),
	.w4(32'hbb74a2a9),
	.w5(32'hbb2ec59c),
	.w6(32'hbb9d5473),
	.w7(32'hbb6a610f),
	.w8(32'hbb6278b8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f7ad4),
	.w1(32'h39c0fd9e),
	.w2(32'h3a1d0f4d),
	.w3(32'hba043bc0),
	.w4(32'h399db73d),
	.w5(32'h3a05b129),
	.w6(32'h39431058),
	.w7(32'h39baec29),
	.w8(32'h39b8f678),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10e3e4),
	.w1(32'h391f3dee),
	.w2(32'h38834f02),
	.w3(32'h39f75751),
	.w4(32'h392ff636),
	.w5(32'hb712eae2),
	.w6(32'h38d25181),
	.w7(32'h38341f43),
	.w8(32'h36982f96),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32a563),
	.w1(32'h3b508499),
	.w2(32'h3b9152ff),
	.w3(32'hba4d7a10),
	.w4(32'hb87391b4),
	.w5(32'h3b0071b3),
	.w6(32'h39c25809),
	.w7(32'h3a2ed813),
	.w8(32'h3b03d3ec),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29d611),
	.w1(32'hbb213ce3),
	.w2(32'hba40ed44),
	.w3(32'hbab52a5f),
	.w4(32'hbb4abc28),
	.w5(32'hba2ce467),
	.w6(32'hbb05a35c),
	.w7(32'hbb22ca2b),
	.w8(32'hba82c91f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab65bcf),
	.w1(32'hba6f8c0d),
	.w2(32'h3ab694ff),
	.w3(32'hbb2ab25e),
	.w4(32'hbad5bbce),
	.w5(32'h39aefebe),
	.w6(32'hba958ae6),
	.w7(32'hba8433f7),
	.w8(32'h3a24a566),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a4bb1),
	.w1(32'h3907ed30),
	.w2(32'h3a7f1128),
	.w3(32'hb8d07861),
	.w4(32'h38166b56),
	.w5(32'h3a29755d),
	.w6(32'hb98465c3),
	.w7(32'h3a46fa8a),
	.w8(32'h39516d96),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39695854),
	.w1(32'hb9dc856f),
	.w2(32'hba1bbf67),
	.w3(32'hb8b46599),
	.w4(32'hb98711cc),
	.w5(32'hb9f72dc4),
	.w6(32'hb9cc99ec),
	.w7(32'hb9bb1b63),
	.w8(32'hb9b961bb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f9a4b),
	.w1(32'h39deae0d),
	.w2(32'h38c7030e),
	.w3(32'h38d5e0f9),
	.w4(32'h398a254b),
	.w5(32'h3995edf6),
	.w6(32'h392f6960),
	.w7(32'h38fe14b5),
	.w8(32'hb8d08c43),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60d11e),
	.w1(32'h382b6bd9),
	.w2(32'h3b00c118),
	.w3(32'hba5c6b23),
	.w4(32'hb9e0a6a0),
	.w5(32'h393a0652),
	.w6(32'hbb0ffd3d),
	.w7(32'hba93b3c5),
	.w8(32'h38a952c9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a790970),
	.w1(32'hbad2d4b7),
	.w2(32'hb99327a3),
	.w3(32'hbae3f88c),
	.w4(32'hbb728601),
	.w5(32'hba7be3c5),
	.w6(32'hbb8f1a57),
	.w7(32'hbb8005e0),
	.w8(32'hbb8f51c5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b84b4),
	.w1(32'h3a2fb1d6),
	.w2(32'h3a752f00),
	.w3(32'hb9412f38),
	.w4(32'hb990942a),
	.w5(32'h38a88064),
	.w6(32'hbb575098),
	.w7(32'hbb29e284),
	.w8(32'hbb025e1f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80d0ef),
	.w1(32'h3afa0bd2),
	.w2(32'h3b51c25b),
	.w3(32'hba306d13),
	.w4(32'h3887e866),
	.w5(32'h3ac19958),
	.w6(32'h3aa8391c),
	.w7(32'h3a89a546),
	.w8(32'h3b1ecf65),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5cb89),
	.w1(32'hbacc092e),
	.w2(32'hbac1ae18),
	.w3(32'hba59e561),
	.w4(32'hbada87a3),
	.w5(32'hba52daac),
	.w6(32'h38fce361),
	.w7(32'h38143199),
	.w8(32'h3ad69122),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba240410),
	.w1(32'h38107012),
	.w2(32'hb8c2eefb),
	.w3(32'hb9fe2d1d),
	.w4(32'hb89e9fc4),
	.w5(32'hb87715e9),
	.w6(32'h38f69409),
	.w7(32'h38b58bbf),
	.w8(32'h3869e63f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367e450f),
	.w1(32'hba1acad9),
	.w2(32'hb981377c),
	.w3(32'h37c1fe5c),
	.w4(32'hb942c3c1),
	.w5(32'hb7c44737),
	.w6(32'hb9ee97d4),
	.w7(32'hb9dabe8e),
	.w8(32'hba1f3627),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aeda41),
	.w1(32'hb8103298),
	.w2(32'hb991c87e),
	.w3(32'h38733452),
	.w4(32'hb976bd98),
	.w5(32'hb975079a),
	.w6(32'hb99f2a7d),
	.w7(32'hb9f37272),
	.w8(32'hba2ddde0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae1b42),
	.w1(32'h38e8d337),
	.w2(32'hb98a2682),
	.w3(32'hba0d3766),
	.w4(32'h39cf62a5),
	.w5(32'hb8effd23),
	.w6(32'h391675c1),
	.w7(32'hb9812c64),
	.w8(32'hb9719c60),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38798fbc),
	.w1(32'h3a049b56),
	.w2(32'h3a750696),
	.w3(32'hb9f2e957),
	.w4(32'h38c042bf),
	.w5(32'h3a235370),
	.w6(32'h391a828f),
	.w7(32'h39106ae5),
	.w8(32'h398fec05),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19515e),
	.w1(32'hba11282d),
	.w2(32'h3abdf303),
	.w3(32'hb993867c),
	.w4(32'hbab06745),
	.w5(32'h3ad56ac8),
	.w6(32'hbab74c2b),
	.w7(32'hbb0b81ed),
	.w8(32'h3963a736),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26d9fd),
	.w1(32'hbb1bcd16),
	.w2(32'hbaa74fc9),
	.w3(32'hb9df11ee),
	.w4(32'hbb2a2081),
	.w5(32'hba6647ec),
	.w6(32'hba96a84b),
	.w7(32'hbad5d204),
	.w8(32'hb982a2a3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fdc6e1),
	.w1(32'hb9b8f867),
	.w2(32'h3a3a1292),
	.w3(32'hb8011596),
	.w4(32'hb99bd8d7),
	.w5(32'hb965daf2),
	.w6(32'hb9dad7f6),
	.w7(32'hb9f4fa76),
	.w8(32'hba5e0db9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e94f2),
	.w1(32'h3a2bf077),
	.w2(32'h3b1f8882),
	.w3(32'hbab9af7f),
	.w4(32'hb9e046f4),
	.w5(32'h3aa8731e),
	.w6(32'hbb940c9c),
	.w7(32'hbb7c195d),
	.w8(32'hbab5e40e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b43aa9),
	.w1(32'hba77d58a),
	.w2(32'hba6dc2f0),
	.w3(32'hba7a0cae),
	.w4(32'hba930332),
	.w5(32'hbaa8e054),
	.w6(32'hbb05bf6a),
	.w7(32'hbb0bd50e),
	.w8(32'hbb0eadb2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d6395),
	.w1(32'h395213fe),
	.w2(32'hb904b4c1),
	.w3(32'h39fb8256),
	.w4(32'h399f2d6b),
	.w5(32'h388f5f71),
	.w6(32'h399706f6),
	.w7(32'hb8965ffb),
	.w8(32'h3951a397),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0fcfa),
	.w1(32'hbad28742),
	.w2(32'hba408815),
	.w3(32'hbaeb3d48),
	.w4(32'hbb121da8),
	.w5(32'hba561e1c),
	.w6(32'hbb490e1d),
	.w7(32'hbb4a33fe),
	.w8(32'hbb26d03e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dd602),
	.w1(32'hb92a85d5),
	.w2(32'hb96b5e60),
	.w3(32'hb9f97530),
	.w4(32'hb8da101b),
	.w5(32'hb88e22f4),
	.w6(32'h391c1982),
	.w7(32'hb825c071),
	.w8(32'h3740962e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7882671),
	.w1(32'hba0714b6),
	.w2(32'hb99f2c89),
	.w3(32'h38ae90af),
	.w4(32'hb9c38183),
	.w5(32'hb98f90f8),
	.w6(32'hb97edfe1),
	.w7(32'hb8f9ac22),
	.w8(32'h38746cdf),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c850f3),
	.w1(32'hb8b50058),
	.w2(32'hb9c69b29),
	.w3(32'hb95d64aa),
	.w4(32'h38d01e33),
	.w5(32'hb94a589d),
	.w6(32'h39397c13),
	.w7(32'hb861dab3),
	.w8(32'h38bc61bf),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e8429),
	.w1(32'h3a01fc03),
	.w2(32'h38f60051),
	.w3(32'hb7465579),
	.w4(32'h39e86cf5),
	.w5(32'h3910072b),
	.w6(32'h39ffbf8c),
	.w7(32'h394f1e9d),
	.w8(32'h3757c278),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c21b9),
	.w1(32'h3aae4243),
	.w2(32'h3b33957b),
	.w3(32'h3914c65c),
	.w4(32'h3a8d6b76),
	.w5(32'h3b2c697c),
	.w6(32'h3b095e72),
	.w7(32'h3aa7c25c),
	.w8(32'h3b2e4d70),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7714de),
	.w1(32'hbb75c0ad),
	.w2(32'hbb246aaa),
	.w3(32'hbb1f79be),
	.w4(32'hbae764a6),
	.w5(32'hba45bd28),
	.w6(32'hbb0a7719),
	.w7(32'hbb55f1d4),
	.w8(32'hbb7ba258),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45743f),
	.w1(32'hbb4c8504),
	.w2(32'hbb0deabf),
	.w3(32'hbb3db2d1),
	.w4(32'hbb2d2913),
	.w5(32'hbacf42cf),
	.w6(32'hbb802c2d),
	.w7(32'hbb8622d1),
	.w8(32'hbb6afb6e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb018ee0),
	.w1(32'hbb14c645),
	.w2(32'hba7d788a),
	.w3(32'hba959109),
	.w4(32'hbb0b851d),
	.w5(32'hbabb4374),
	.w6(32'hbb2aa485),
	.w7(32'hbb38c978),
	.w8(32'hbb1ccb68),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0e08d),
	.w1(32'h39804d21),
	.w2(32'h39e49f1f),
	.w3(32'hb9a637e1),
	.w4(32'h38e3f208),
	.w5(32'h394ddc1a),
	.w6(32'h3994dbc5),
	.w7(32'h39206dc0),
	.w8(32'h38ab9ad5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38034c6b),
	.w1(32'h38853ad9),
	.w2(32'hb9c0f09f),
	.w3(32'h3881e715),
	.w4(32'h39bbec15),
	.w5(32'hb8db99f0),
	.w6(32'h39b8dfca),
	.w7(32'h37367b7f),
	.w8(32'h3922ff43),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb756a4fd),
	.w1(32'h37557de4),
	.w2(32'hb79f9b12),
	.w3(32'h39447734),
	.w4(32'h3960798a),
	.w5(32'h38a0b6e9),
	.w6(32'h390fde6d),
	.w7(32'h38a87233),
	.w8(32'h3947126a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ef202),
	.w1(32'h364fca7a),
	.w2(32'h34b0cff6),
	.w3(32'h3979cf70),
	.w4(32'h39542f9c),
	.w5(32'h3935b02d),
	.w6(32'h38a4be5c),
	.w7(32'h38ad4f0f),
	.w8(32'h39b5c791),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0130),
	.w1(32'h3b009c2c),
	.w2(32'h3ab387fa),
	.w3(32'h3b448e8a),
	.w4(32'h3a86386e),
	.w5(32'h3a37eb3b),
	.w6(32'h3b152586),
	.w7(32'h39b3cb8a),
	.w8(32'hbaacf2dc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ffabd),
	.w1(32'h3991d500),
	.w2(32'hb6f58387),
	.w3(32'h3a587231),
	.w4(32'h394e3f09),
	.w5(32'h390ebe5e),
	.w6(32'h37eaef9b),
	.w7(32'h39c1bd39),
	.w8(32'h3a29ddfe),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b6d3e),
	.w1(32'hba801779),
	.w2(32'h391f24b1),
	.w3(32'hba3a447b),
	.w4(32'hbac41364),
	.w5(32'hb93961d4),
	.w6(32'hba0214d8),
	.w7(32'hbaab3840),
	.w8(32'h390ca601),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3935e28e),
	.w1(32'h37ce0088),
	.w2(32'h39bcfa04),
	.w3(32'h3971e46e),
	.w4(32'h39366679),
	.w5(32'h3a249228),
	.w6(32'hb9131c3a),
	.w7(32'hb97d6a8f),
	.w8(32'h39c30a12),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899eed7),
	.w1(32'h39a29c38),
	.w2(32'h3929fd1a),
	.w3(32'h390f7878),
	.w4(32'h39cbe789),
	.w5(32'h391f361b),
	.w6(32'hb8929255),
	.w7(32'h38a1a1fe),
	.w8(32'h3969408e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af0be4),
	.w1(32'h392e489c),
	.w2(32'h3937a3f0),
	.w3(32'h3796336d),
	.w4(32'h390ea392),
	.w5(32'h37efc714),
	.w6(32'hba83be81),
	.w7(32'hba8fcb03),
	.w8(32'hbad23873),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eaf9fe),
	.w1(32'hba205c53),
	.w2(32'hb98e2138),
	.w3(32'h3984c4f9),
	.w4(32'hb8a889b4),
	.w5(32'h3980b8bb),
	.w6(32'hba01ba73),
	.w7(32'hb9e0a4a2),
	.w8(32'hb96f62ca),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a009d5e),
	.w1(32'hba8002c1),
	.w2(32'hbb04c62c),
	.w3(32'h3a8bbd3c),
	.w4(32'hbb4fabba),
	.w5(32'hbb58246c),
	.w6(32'hbac1b782),
	.w7(32'hbb6d39e7),
	.w8(32'hbb83d54f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad5c5f),
	.w1(32'hbcea0b21),
	.w2(32'hbc0fed66),
	.w3(32'hb9610d44),
	.w4(32'hbc55710c),
	.w5(32'hbb62ae22),
	.w6(32'hbc9fb96c),
	.w7(32'hbbb5bc65),
	.w8(32'h3b6fc83f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12fdb8),
	.w1(32'hbce9af25),
	.w2(32'h3b4a7835),
	.w3(32'h3a2cbee0),
	.w4(32'hbc939cad),
	.w5(32'hbbb3e7a0),
	.w6(32'hbc7e780f),
	.w7(32'h3b5b40f3),
	.w8(32'h3c338340),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule