module layer_10_featuremap_70(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5ea5),
	.w1(32'hbbc6a972),
	.w2(32'hba754d2c),
	.w3(32'h3c0c4cf3),
	.w4(32'h3c85ee5c),
	.w5(32'hba772d15),
	.w6(32'h3c2d452c),
	.w7(32'h3cf7a3de),
	.w8(32'hbc19b738),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6017c),
	.w1(32'h3c0c0d22),
	.w2(32'h3bcaa69f),
	.w3(32'h3c64438a),
	.w4(32'h3c9b5268),
	.w5(32'h3b8e988a),
	.w6(32'hbbbb60ce),
	.w7(32'h3ca009d1),
	.w8(32'h37d3a98d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371d1aa2),
	.w1(32'hbb09657e),
	.w2(32'h3b697ea8),
	.w3(32'h3b456f3f),
	.w4(32'h3b2c8609),
	.w5(32'h3bc47a3f),
	.w6(32'hb773138a),
	.w7(32'h3c084bf2),
	.w8(32'h3b96c91d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4422f2),
	.w1(32'h3ba87d83),
	.w2(32'hbc950fee),
	.w3(32'h39e0d017),
	.w4(32'h3be363de),
	.w5(32'hbcb04ac4),
	.w6(32'h3b43f64f),
	.w7(32'h3b2b7d68),
	.w8(32'hbcbb90c9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d196e),
	.w1(32'h3d0b6f72),
	.w2(32'hbaeb388e),
	.w3(32'hbc6b4264),
	.w4(32'h3c190680),
	.w5(32'hbc39b0eb),
	.w6(32'hbc86cff9),
	.w7(32'hbb614f11),
	.w8(32'hbc15f2aa),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1cf1),
	.w1(32'h3aca7c2d),
	.w2(32'h3bdda866),
	.w3(32'h3b1c403c),
	.w4(32'hbc144604),
	.w5(32'h3b933ed4),
	.w6(32'h3b078d9e),
	.w7(32'hbc16b915),
	.w8(32'h3b896e52),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62ce91),
	.w1(32'h3b38de47),
	.w2(32'hbc2685b3),
	.w3(32'hbb0eac38),
	.w4(32'hbb6152d3),
	.w5(32'hbbd252a9),
	.w6(32'hba1f25d8),
	.w7(32'hba35c037),
	.w8(32'hbbee9a2e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d914),
	.w1(32'h3c3bb4df),
	.w2(32'hbb5538c4),
	.w3(32'hbbfedb3d),
	.w4(32'h3c17d596),
	.w5(32'hbb8912f6),
	.w6(32'hbc223182),
	.w7(32'hba6391bb),
	.w8(32'hba053a05),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4ea69),
	.w1(32'hbc088de2),
	.w2(32'h3c1abb86),
	.w3(32'h3ba791ef),
	.w4(32'h3c0bd2d7),
	.w5(32'h3be5e667),
	.w6(32'h3c18d252),
	.w7(32'h3c70eecf),
	.w8(32'h3c2124fc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae5658),
	.w1(32'hbb9c4854),
	.w2(32'hbb25bbec),
	.w3(32'h3b3d3d4e),
	.w4(32'hbc0f2521),
	.w5(32'hbb5166dd),
	.w6(32'h3bd3fe81),
	.w7(32'hbb8c8366),
	.w8(32'hbbade21e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9503c2),
	.w1(32'hbb3708ad),
	.w2(32'h3a16f2a7),
	.w3(32'hba37807b),
	.w4(32'hbaf2f0b3),
	.w5(32'h3ad3ab7a),
	.w6(32'hbb172b7b),
	.w7(32'hbb1e070c),
	.w8(32'h3a96428a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ba8c),
	.w1(32'h3b4fde41),
	.w2(32'hbac21171),
	.w3(32'h3b0eeaf6),
	.w4(32'h3b7e758f),
	.w5(32'hbb7e966f),
	.w6(32'hbb1f3d32),
	.w7(32'h3c1c25ce),
	.w8(32'hbacf3140),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f9a8e),
	.w1(32'h3bae8003),
	.w2(32'h3aef42a5),
	.w3(32'hbb9300d4),
	.w4(32'h3b96916e),
	.w5(32'h3a3fe25e),
	.w6(32'hbb014a15),
	.w7(32'h3b9928f8),
	.w8(32'h3bd971a4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6a63),
	.w1(32'h3c01e2a9),
	.w2(32'h3c0b2398),
	.w3(32'h3c8480c6),
	.w4(32'h3b31d3d2),
	.w5(32'h3b48e166),
	.w6(32'h3c39736c),
	.w7(32'h3a20cbd7),
	.w8(32'hba105dc9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac50ff7),
	.w1(32'h3c602204),
	.w2(32'hbb145ed2),
	.w3(32'hbab345c1),
	.w4(32'h3cb0f7fb),
	.w5(32'hba22bf44),
	.w6(32'hbae8cdba),
	.w7(32'h3c8b9a7e),
	.w8(32'h3bbe5a64),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4f5c8),
	.w1(32'hbaeb350d),
	.w2(32'h3a03d17f),
	.w3(32'hbb85c16c),
	.w4(32'hbbd22958),
	.w5(32'h39517186),
	.w6(32'h3bb77a12),
	.w7(32'h3aa30546),
	.w8(32'hba5699d0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a109d25),
	.w1(32'hbac55c65),
	.w2(32'h3a874f13),
	.w3(32'h3a863eb9),
	.w4(32'h392ba6a5),
	.w5(32'h3b9643cc),
	.w6(32'hba067efb),
	.w7(32'hba45a93a),
	.w8(32'h3c1210be),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb703291),
	.w1(32'hbbe5a722),
	.w2(32'h3b59e94b),
	.w3(32'hba6e1bff),
	.w4(32'hbc135945),
	.w5(32'hb985c164),
	.w6(32'h3bebe26a),
	.w7(32'hbb8a4efb),
	.w8(32'h3a5790a0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf94da),
	.w1(32'h3b5014c2),
	.w2(32'hbc070204),
	.w3(32'h3c1fd081),
	.w4(32'h3b8ba1c0),
	.w5(32'hbc27d39a),
	.w6(32'h3b8480a2),
	.w7(32'h3b28e5f8),
	.w8(32'hbc684f80),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b219),
	.w1(32'h39e52a8f),
	.w2(32'h3b52f301),
	.w3(32'hbad36476),
	.w4(32'h3cb5a088),
	.w5(32'hbb0f26a6),
	.w6(32'hbc0b782f),
	.w7(32'h3ccaace4),
	.w8(32'hbaa86f73),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395cb5bf),
	.w1(32'h3b7dcfb7),
	.w2(32'h3a28914d),
	.w3(32'hbbbf0494),
	.w4(32'hbbb011ec),
	.w5(32'hbb14f3a3),
	.w6(32'hbbca0368),
	.w7(32'hbb4079b6),
	.w8(32'h39c4cee9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67fb1e),
	.w1(32'h3b6e0e33),
	.w2(32'hba5c7d43),
	.w3(32'hbbae6a19),
	.w4(32'h3be7d671),
	.w5(32'hbb7b4893),
	.w6(32'hbb8b10bc),
	.w7(32'h3c016622),
	.w8(32'hbb8d68d2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ad531),
	.w1(32'hbc14b227),
	.w2(32'h393b8a30),
	.w3(32'hbc1ebada),
	.w4(32'hbc47a01c),
	.w5(32'hbb120351),
	.w6(32'hbbfb6ad0),
	.w7(32'hbc04e7c5),
	.w8(32'hbae7deac),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c5c9d),
	.w1(32'h3a6ee108),
	.w2(32'h3ba3a463),
	.w3(32'hb951524b),
	.w4(32'h3a1d8558),
	.w5(32'h3adc9326),
	.w6(32'hbb454370),
	.w7(32'hb7017171),
	.w8(32'h3bbefb9d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff0e9),
	.w1(32'h3be34869),
	.w2(32'hbc25dcda),
	.w3(32'h3c23f590),
	.w4(32'h3bc784e2),
	.w5(32'hbc6ba188),
	.w6(32'h3bbc4351),
	.w7(32'h3a34e6af),
	.w8(32'hbc243cbc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa4c81),
	.w1(32'h3c1194c2),
	.w2(32'hbac3e103),
	.w3(32'hbc137fa2),
	.w4(32'h3ca5c8e0),
	.w5(32'h3aaf6aed),
	.w6(32'hbc3ddb02),
	.w7(32'h3c678fdb),
	.w8(32'hbb9be4d1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ee5b1),
	.w1(32'h3a675024),
	.w2(32'h3a8e73d2),
	.w3(32'hbbfd4b2b),
	.w4(32'h3b6c066f),
	.w5(32'h3ade475b),
	.w6(32'hbb38d997),
	.w7(32'h3b27576a),
	.w8(32'h3aae3adf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a353c8a),
	.w1(32'hbacd2e94),
	.w2(32'h3c1e43b4),
	.w3(32'h3b7f79c8),
	.w4(32'hbb212ec6),
	.w5(32'h3c0ac941),
	.w6(32'h3b3995c0),
	.w7(32'hba642d7f),
	.w8(32'h3c6537cb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a2dab),
	.w1(32'h3bb13fde),
	.w2(32'hba539259),
	.w3(32'hb69736e7),
	.w4(32'h3c4e5eee),
	.w5(32'hbbd26b6e),
	.w6(32'hbb1b4d62),
	.w7(32'h3c20a876),
	.w8(32'hbc1fce40),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b888042),
	.w1(32'h3b9d021e),
	.w2(32'hba877172),
	.w3(32'hba0172d1),
	.w4(32'h3b9f518e),
	.w5(32'hbc4bfcc0),
	.w6(32'h3a976603),
	.w7(32'h3b79a43c),
	.w8(32'hbbbd4015),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb04da4),
	.w1(32'h3a5450b9),
	.w2(32'hbb2485cc),
	.w3(32'hbabce4f8),
	.w4(32'hbae5a95d),
	.w5(32'h39f6cc4d),
	.w6(32'h3aa20d70),
	.w7(32'h38878126),
	.w8(32'hbbb5cde5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d1b58),
	.w1(32'h3a9ec39f),
	.w2(32'h3a836852),
	.w3(32'h3b5d5d6b),
	.w4(32'h3b34e158),
	.w5(32'hbb9e43ce),
	.w6(32'hba05f8bb),
	.w7(32'h3babb8e3),
	.w8(32'hbba9a096),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e0cb),
	.w1(32'hbb6ebba1),
	.w2(32'h3b7776d8),
	.w3(32'h3bbe40e4),
	.w4(32'hbb48e10a),
	.w5(32'hbba1836f),
	.w6(32'h3a83dffc),
	.w7(32'h3b061e87),
	.w8(32'h3a36ac9d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945bbd),
	.w1(32'hbaac4b5a),
	.w2(32'hbbc2eb96),
	.w3(32'h3b75317b),
	.w4(32'hbb9d93f7),
	.w5(32'h3c825ae3),
	.w6(32'h3b19eda4),
	.w7(32'hbb47fe51),
	.w8(32'h3c6ce6e6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e5b2c),
	.w1(32'h3b3b7306),
	.w2(32'h3b7d3046),
	.w3(32'h3c16fe47),
	.w4(32'h3bc917f2),
	.w5(32'h3c02cee7),
	.w6(32'h3c2754db),
	.w7(32'h3c1b22a2),
	.w8(32'h3bce49a9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ace23),
	.w1(32'hbb7bb36b),
	.w2(32'h3a7444c5),
	.w3(32'h3a14b8fe),
	.w4(32'hbbe2c0db),
	.w5(32'hbc790ff4),
	.w6(32'hbb27684d),
	.w7(32'hbbde2d61),
	.w8(32'hbca173ea),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd42e6),
	.w1(32'hbb7dfac3),
	.w2(32'hbb5f3452),
	.w3(32'h3b212c9c),
	.w4(32'hb84b79e9),
	.w5(32'hbc8f5e90),
	.w6(32'hba6e5de1),
	.w7(32'h3b1867bd),
	.w8(32'hbc1eb5cc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf20fe0),
	.w1(32'hb92ce7b1),
	.w2(32'hbbe190be),
	.w3(32'h3aa47c6f),
	.w4(32'hbb276979),
	.w5(32'h3acd3067),
	.w6(32'h3b63b342),
	.w7(32'hb9c32f34),
	.w8(32'h3bda3d3a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb0d08),
	.w1(32'h3c094193),
	.w2(32'hbc17a09e),
	.w3(32'h3b99930f),
	.w4(32'h3bb8091d),
	.w5(32'hbc5bc005),
	.w6(32'h3b8d8426),
	.w7(32'h3b1c40b5),
	.w8(32'hbca2e210),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bab88),
	.w1(32'hbc900ed3),
	.w2(32'h3b10a147),
	.w3(32'hbc4b3e8b),
	.w4(32'hbcbbcfa6),
	.w5(32'h3b157e35),
	.w6(32'hbc924df7),
	.w7(32'hbcb10083),
	.w8(32'hbb154910),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f2045),
	.w1(32'h3b80afd9),
	.w2(32'h3ba522d1),
	.w3(32'h3ba2effc),
	.w4(32'h3bf45fb2),
	.w5(32'h3c524dc0),
	.w6(32'hba92f01d),
	.w7(32'h3c245172),
	.w8(32'h3b24f771),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be52e3c),
	.w1(32'h3a7fe341),
	.w2(32'hbbe15071),
	.w3(32'h3c6f2888),
	.w4(32'hbb987479),
	.w5(32'h3b7664fe),
	.w6(32'h3bd25d42),
	.w7(32'h3ab1d117),
	.w8(32'h3b02d0d0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f740e),
	.w1(32'h3af23b7a),
	.w2(32'h3b4acf6a),
	.w3(32'h39034918),
	.w4(32'h3b3ff1f2),
	.w5(32'h3c228e38),
	.w6(32'h3bba2cd8),
	.w7(32'h3bb90aae),
	.w8(32'h3b977e09),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85eb70c),
	.w1(32'hbba16e5d),
	.w2(32'h39a28aea),
	.w3(32'h3b147751),
	.w4(32'hbbabd364),
	.w5(32'hb72c4d32),
	.w6(32'h3b6cc35a),
	.w7(32'hbb985bf1),
	.w8(32'hba7883ac),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c1e5d),
	.w1(32'h3c84bfce),
	.w2(32'h3a6003e4),
	.w3(32'h3c112467),
	.w4(32'h3c6388ae),
	.w5(32'hbc2e6a64),
	.w6(32'h3bfc12d6),
	.w7(32'h3c8510f7),
	.w8(32'hbb924fc7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8779fd),
	.w1(32'hbae684ab),
	.w2(32'hbc012f32),
	.w3(32'hbbbf475d),
	.w4(32'hbc35cefe),
	.w5(32'hbb0472c6),
	.w6(32'hbb78225e),
	.w7(32'h3b75d098),
	.w8(32'hbb5bb977),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9980c20),
	.w1(32'h3b27a90f),
	.w2(32'h3b949ed7),
	.w3(32'h3b204257),
	.w4(32'h3a613af1),
	.w5(32'h3b073650),
	.w6(32'h3c21c632),
	.w7(32'h3a2b93cd),
	.w8(32'h3b0d546a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4974e),
	.w1(32'h3ba6b8c6),
	.w2(32'h3bfd285b),
	.w3(32'h3c1fd409),
	.w4(32'h3bb39109),
	.w5(32'h3c8d5852),
	.w6(32'h3bb340ed),
	.w7(32'h3bd9addd),
	.w8(32'h3c4b0988),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41291b),
	.w1(32'hbb9f1561),
	.w2(32'hb9b67412),
	.w3(32'h3b8da533),
	.w4(32'hbbc5f6ef),
	.w5(32'h3bc27381),
	.w6(32'h3bbdde47),
	.w7(32'hbbe6da33),
	.w8(32'h3c5e7771),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51da03),
	.w1(32'h39ef7187),
	.w2(32'hbb0e06d7),
	.w3(32'hbb09bc45),
	.w4(32'hbc647b1a),
	.w5(32'hbc0a6331),
	.w6(32'hba5438c5),
	.w7(32'hbbef98a8),
	.w8(32'hbb88c6c8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab020e1),
	.w1(32'h3b571791),
	.w2(32'hbc661f26),
	.w3(32'hbaf48d41),
	.w4(32'h3b858669),
	.w5(32'hbc9a9faa),
	.w6(32'hbb5d3c9e),
	.w7(32'h3a878a41),
	.w8(32'hbc2c6e85),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83fa11),
	.w1(32'hbc66516c),
	.w2(32'hbb404d98),
	.w3(32'hbc739ea6),
	.w4(32'hbcccb28a),
	.w5(32'hbbda8285),
	.w6(32'hbbdde625),
	.w7(32'hbc12e0fa),
	.w8(32'hbc0e0ede),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14edbe),
	.w1(32'hbb90f54b),
	.w2(32'h3bb72707),
	.w3(32'hbac38eca),
	.w4(32'h3ae91b57),
	.w5(32'h3c33321c),
	.w6(32'hbbe28997),
	.w7(32'h3b593312),
	.w8(32'h3b0625e8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37adb4),
	.w1(32'hbc38d177),
	.w2(32'h3bd17cdf),
	.w3(32'hbb66c7ba),
	.w4(32'hbc926630),
	.w5(32'hb992ad3a),
	.w6(32'hba80009c),
	.w7(32'hbbae370d),
	.w8(32'hbb9a3f1c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cb348c),
	.w1(32'hbbd9f781),
	.w2(32'hbbe8a905),
	.w3(32'hbc09de4d),
	.w4(32'hbb290bac),
	.w5(32'h3af0fe3e),
	.w6(32'hbc23d75e),
	.w7(32'hbb62dda7),
	.w8(32'h3b535080),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99617a),
	.w1(32'h390062d1),
	.w2(32'hbb35e1a5),
	.w3(32'h3b6e83cb),
	.w4(32'h3b8c4f9d),
	.w5(32'hb8f6a8f9),
	.w6(32'h39a7a760),
	.w7(32'hba85a6ac),
	.w8(32'h3b462147),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c226f8e),
	.w1(32'h3c092601),
	.w2(32'h3cc85661),
	.w3(32'h3c154994),
	.w4(32'h3c4aa608),
	.w5(32'h3d33da33),
	.w6(32'h3c707338),
	.w7(32'h3c10158e),
	.w8(32'h3d2fcfe4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0f501),
	.w1(32'h3d1a3328),
	.w2(32'h3a446f6c),
	.w3(32'h3d2c7270),
	.w4(32'h3d4927e2),
	.w5(32'h3af93aac),
	.w6(32'h3d0c2d0c),
	.w7(32'h3d3c3b28),
	.w8(32'hbb9991b5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfb5b),
	.w1(32'h3c6514bf),
	.w2(32'hbbf52528),
	.w3(32'h3c056ddb),
	.w4(32'h3c46f0fd),
	.w5(32'h3ad7cb03),
	.w6(32'h3bccb6e5),
	.w7(32'h3c5a1669),
	.w8(32'h3bb507c6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a850c70),
	.w1(32'hbb096166),
	.w2(32'h3bf04fb3),
	.w3(32'h3a78fd3e),
	.w4(32'hbc2f22ec),
	.w5(32'h3bebfe23),
	.w6(32'h3b1e8796),
	.w7(32'hbbdb360c),
	.w8(32'h3c17eb79),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c359105),
	.w1(32'h3bffbca8),
	.w2(32'hbbc3b2bd),
	.w3(32'h3b98bd0c),
	.w4(32'h3b711904),
	.w5(32'hbc54561a),
	.w6(32'h3b81fe06),
	.w7(32'hbb0c4810),
	.w8(32'hbbba9706),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc233d92),
	.w1(32'hbc020fc2),
	.w2(32'hbc300745),
	.w3(32'hbc203894),
	.w4(32'hbbbf22ce),
	.w5(32'hbc2125fd),
	.w6(32'hbc3d0fd9),
	.w7(32'hbb4bf2e6),
	.w8(32'hbb951d86),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc117d2),
	.w1(32'h3a1cf46a),
	.w2(32'hb9c3d5ab),
	.w3(32'hbadce901),
	.w4(32'h3ab2000d),
	.w5(32'h3bd332f4),
	.w6(32'hbae4ed62),
	.w7(32'hb90ab22e),
	.w8(32'hbb9c2a5a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d5e4),
	.w1(32'h3be44e9f),
	.w2(32'hbbba4dda),
	.w3(32'h3c340fac),
	.w4(32'h3bd086ff),
	.w5(32'h395127e6),
	.w6(32'h3bab80f1),
	.w7(32'h3c0d8502),
	.w8(32'hb9b53448),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e268e5),
	.w1(32'hbae3f563),
	.w2(32'h3c871f95),
	.w3(32'h3b676f81),
	.w4(32'h3a87242d),
	.w5(32'h3cafaf59),
	.w6(32'h39c4f2ce),
	.w7(32'h3b83b3f5),
	.w8(32'h3c8f3e35),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49a074),
	.w1(32'h3c706629),
	.w2(32'hbb778780),
	.w3(32'h3c60be05),
	.w4(32'h3ca60b08),
	.w5(32'hbb29df7f),
	.w6(32'h3c7201ab),
	.w7(32'h3cbaadb8),
	.w8(32'hbb036b61),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf465d9),
	.w1(32'h3bc49f92),
	.w2(32'h3af9e066),
	.w3(32'h3c4f1b53),
	.w4(32'h3c3d3a3b),
	.w5(32'hbb2fe555),
	.w6(32'h3c4743bc),
	.w7(32'h3c1f3666),
	.w8(32'hb9ac68f7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97878d),
	.w1(32'hbb2bb94a),
	.w2(32'h39187096),
	.w3(32'h3c2ca57b),
	.w4(32'hbb52823b),
	.w5(32'hbb8649b1),
	.w6(32'h3b7d203a),
	.w7(32'h3b6beba3),
	.w8(32'hbb128028),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a590),
	.w1(32'h3afa3972),
	.w2(32'h3bf67bbd),
	.w3(32'hbb42adcc),
	.w4(32'h3aa091b4),
	.w5(32'h3c0bc895),
	.w6(32'hbb8001c8),
	.w7(32'hb9f23e68),
	.w8(32'h3c06a41a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d2b3f),
	.w1(32'h3abf8154),
	.w2(32'hbd3ddbb7),
	.w3(32'h3b8b2c01),
	.w4(32'h3abc5048),
	.w5(32'hbd83e067),
	.w6(32'h3b30f4cf),
	.w7(32'h3afad195),
	.w8(32'hbd464bfa),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd410b19),
	.w1(32'hbcca62dd),
	.w2(32'h3bbfb16d),
	.w3(32'hbd5ec5b0),
	.w4(32'hbd19b541),
	.w5(32'h3c3b2213),
	.w6(32'hbd2dd380),
	.w7(32'hbd1ce4da),
	.w8(32'h3c1aab11),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c9236),
	.w1(32'hb92b2a64),
	.w2(32'h3b152d9b),
	.w3(32'h3c11d778),
	.w4(32'h3b575cde),
	.w5(32'hb8cbd39f),
	.w6(32'h3ac43a7f),
	.w7(32'h3b9cb3b4),
	.w8(32'hbb6132f9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8069af),
	.w1(32'h3962d489),
	.w2(32'hbbb21b99),
	.w3(32'h3c22d838),
	.w4(32'hbb815b68),
	.w5(32'hbc1eea88),
	.w6(32'h3b4f8cf0),
	.w7(32'hbb81e125),
	.w8(32'hbc4ddd65),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85a061),
	.w1(32'h3b282f9c),
	.w2(32'h3bf28d8e),
	.w3(32'h3b3bbc57),
	.w4(32'h39b5a30f),
	.w5(32'h3b90b869),
	.w6(32'h3ae44374),
	.w7(32'h3bf352a1),
	.w8(32'h3b974809),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a063129),
	.w1(32'hbb82ac5d),
	.w2(32'h3c3652fb),
	.w3(32'hbbd9135d),
	.w4(32'hbc746a64),
	.w5(32'h3c473c3c),
	.w6(32'hbb434c0c),
	.w7(32'hbc32b575),
	.w8(32'h3c1d9efa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985b735),
	.w1(32'hbc85f513),
	.w2(32'hbbce0298),
	.w3(32'hba8c93a6),
	.w4(32'hbcbf6c86),
	.w5(32'hbb789326),
	.w6(32'h3a55f040),
	.w7(32'hbcac0261),
	.w8(32'hbb3ca961),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931f423),
	.w1(32'h3b8c7107),
	.w2(32'hbb9ca7e4),
	.w3(32'hbb86ca15),
	.w4(32'h3bdb2caa),
	.w5(32'hbb6b84d5),
	.w6(32'hbb642646),
	.w7(32'hbb6c0970),
	.w8(32'hbbea08ab),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e8f01),
	.w1(32'h3b027a3c),
	.w2(32'h3c2c3862),
	.w3(32'h3c027425),
	.w4(32'h3bade906),
	.w5(32'h3c664352),
	.w6(32'h3be31185),
	.w7(32'hba87450f),
	.w8(32'h3c19d126),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd2671),
	.w1(32'hba1aa1bc),
	.w2(32'h3b6d5e8a),
	.w3(32'h3c073263),
	.w4(32'h3c7329b0),
	.w5(32'h3b53bbe3),
	.w6(32'h3b941b00),
	.w7(32'h3c3ad703),
	.w8(32'h3b8362cb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc475e87),
	.w1(32'hbab877dd),
	.w2(32'hbc07010d),
	.w3(32'hbc676add),
	.w4(32'hbb461ba9),
	.w5(32'hbc904e78),
	.w6(32'hbc6db22b),
	.w7(32'hba56f297),
	.w8(32'hbc828d31),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47d071),
	.w1(32'hbc0ba0ee),
	.w2(32'h3bc54d7d),
	.w3(32'hbc6f2330),
	.w4(32'hbc6c024e),
	.w5(32'hb89e77f0),
	.w6(32'hbc36ab84),
	.w7(32'hbc8ca0ad),
	.w8(32'h3aedb1ec),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27cdc8),
	.w1(32'hbb01f9a5),
	.w2(32'hbb6730da),
	.w3(32'h3c11d164),
	.w4(32'hbb61f32e),
	.w5(32'hbbb5f07c),
	.w6(32'h3c25ce05),
	.w7(32'hbb26ba2a),
	.w8(32'hbb22ed13),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb13d1e),
	.w1(32'h3b65907b),
	.w2(32'hbcbbe527),
	.w3(32'hbb953be2),
	.w4(32'h3b1d3e98),
	.w5(32'hbcd2a484),
	.w6(32'hbb52f06f),
	.w7(32'hbb0643e6),
	.w8(32'hbca1de25),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a937e),
	.w1(32'h398744b2),
	.w2(32'hbb16c2b7),
	.w3(32'hbc6fa8ab),
	.w4(32'hbbbdb33a),
	.w5(32'hbb4e026e),
	.w6(32'hbbfba7c0),
	.w7(32'hb6c3b32d),
	.w8(32'hbb9f6566),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c2fc9),
	.w1(32'h3ad92ec0),
	.w2(32'hba0ea460),
	.w3(32'hbb16b8e5),
	.w4(32'hba802390),
	.w5(32'h3a9c80e0),
	.w6(32'h3b0c3e33),
	.w7(32'hbaeb071d),
	.w8(32'h3ab1c077),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77087d),
	.w1(32'h3bbf223a),
	.w2(32'h3cbb971d),
	.w3(32'h3c0889e4),
	.w4(32'h3c091e29),
	.w5(32'h3cfe2931),
	.w6(32'h3c4d9143),
	.w7(32'h3c2d5cde),
	.w8(32'h3ceacd05),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1101f),
	.w1(32'h3ca0f473),
	.w2(32'h3a9d9eaa),
	.w3(32'h3d17bb7e),
	.w4(32'h3d0c29b6),
	.w5(32'h3b8ad51d),
	.w6(32'h3d0dd9ca),
	.w7(32'h3d0b77d8),
	.w8(32'h3a1a6bbe),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0cfd0),
	.w1(32'hbb40d8af),
	.w2(32'h3b73b24f),
	.w3(32'hba4d3c66),
	.w4(32'hbb88b414),
	.w5(32'hbbe1e834),
	.w6(32'hbb4b73cf),
	.w7(32'hbba8621b),
	.w8(32'hbb2bd6fe),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf84ad),
	.w1(32'hb7b88391),
	.w2(32'hbc22398f),
	.w3(32'hbb7c125c),
	.w4(32'hba96e685),
	.w5(32'hbaa47660),
	.w6(32'hb973b7c1),
	.w7(32'hbbd20b93),
	.w8(32'h3bbe78f8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba784e9),
	.w1(32'h3c1cf3a0),
	.w2(32'hbb666c64),
	.w3(32'h38ddcc77),
	.w4(32'hba9c0d7c),
	.w5(32'hbbd0e809),
	.w6(32'h3bef3d41),
	.w7(32'hbc013e91),
	.w8(32'hbb7e055d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3fdb5),
	.w1(32'h3bd9851c),
	.w2(32'hbc984a6b),
	.w3(32'h3b93f331),
	.w4(32'h3b5aa243),
	.w5(32'hbcb9ce0b),
	.w6(32'h3b96675c),
	.w7(32'hba9976bd),
	.w8(32'hbc8b53e0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ce78d),
	.w1(32'h3cd5d7df),
	.w2(32'h3bb042ae),
	.w3(32'h3bc8003f),
	.w4(32'h3cea8544),
	.w5(32'h3bf8c911),
	.w6(32'h3bed36af),
	.w7(32'h3cc6d8e9),
	.w8(32'h3b991d4a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0f707),
	.w1(32'hbc3dd1f5),
	.w2(32'hbbb0d19c),
	.w3(32'hbc1fe444),
	.w4(32'hbc5e0041),
	.w5(32'hbb174ad7),
	.w6(32'hbc16c1a7),
	.w7(32'hbc55bc72),
	.w8(32'hbb6281f1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba211acf),
	.w1(32'hbb069010),
	.w2(32'hbb43ee09),
	.w3(32'h3b1a7a03),
	.w4(32'h3ace4a4f),
	.w5(32'hbbae7e09),
	.w6(32'h3b27ee0b),
	.w7(32'h3a3c9b49),
	.w8(32'hbb8edb12),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9458ec),
	.w1(32'hbb59beac),
	.w2(32'hbc020c05),
	.w3(32'hba1c240e),
	.w4(32'hbba558a4),
	.w5(32'hbb39ddf8),
	.w6(32'hb98d34b2),
	.w7(32'h3b47797d),
	.w8(32'hbbd23b3e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0f838),
	.w1(32'h3c2cb88b),
	.w2(32'h3ad96c40),
	.w3(32'hbb1cdefd),
	.w4(32'h3c6a22c1),
	.w5(32'hb7a72c36),
	.w6(32'h3ba04e0d),
	.w7(32'h3c3ab855),
	.w8(32'hba879af3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16313),
	.w1(32'hbc89418c),
	.w2(32'h393393e9),
	.w3(32'hbacf77ea),
	.w4(32'hbc933a90),
	.w5(32'hbaed2962),
	.w6(32'hbb9c1c49),
	.w7(32'hbc1022df),
	.w8(32'h3ba5dc50),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1182ed),
	.w1(32'hbac9b90a),
	.w2(32'h3b2df934),
	.w3(32'h3b020ebd),
	.w4(32'h3ba1971d),
	.w5(32'h3c4dff85),
	.w6(32'h3b5374a8),
	.w7(32'h3af7ba63),
	.w8(32'h3c5591e9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2744c),
	.w1(32'h3b35c774),
	.w2(32'hbcb555b1),
	.w3(32'h3c45031a),
	.w4(32'h3b777dbb),
	.w5(32'hbd2e47c6),
	.w6(32'h3c1f827c),
	.w7(32'h3a460d5b),
	.w8(32'hbd287f08),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d23bd),
	.w1(32'hbb4857a4),
	.w2(32'hba8fe324),
	.w3(32'hbbd2a3a2),
	.w4(32'hbc145fb1),
	.w5(32'hbbb5bdcc),
	.w6(32'hbc24290b),
	.w7(32'hbc4c890b),
	.w8(32'hbc221091),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002b83),
	.w1(32'hba552fa8),
	.w2(32'hbc2b2fe8),
	.w3(32'h3b05d76e),
	.w4(32'hbb0985f7),
	.w5(32'hbc089e47),
	.w6(32'hbbcb1c25),
	.w7(32'h3a76a3fa),
	.w8(32'hbc1e427e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074d27),
	.w1(32'hba1f3d1b),
	.w2(32'hbb11e9e0),
	.w3(32'h3af48f8c),
	.w4(32'h38ec3b1c),
	.w5(32'h3b86cc80),
	.w6(32'h3b1660a8),
	.w7(32'h3bb85333),
	.w8(32'h3b6cdf5a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad981cd),
	.w1(32'hbbed8c08),
	.w2(32'hbc99bc7b),
	.w3(32'h3c6eb581),
	.w4(32'hbc254be7),
	.w5(32'hbc8501c3),
	.w6(32'h3c1fb7e7),
	.w7(32'hbc2e7d90),
	.w8(32'hbc9d54c8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb6dac),
	.w1(32'hbb87d62a),
	.w2(32'hba91c68e),
	.w3(32'hbc7f2b36),
	.w4(32'hbc47fb2a),
	.w5(32'h3a5b9521),
	.w6(32'hbbf0d861),
	.w7(32'hbc493414),
	.w8(32'h3b3292b5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02b7db),
	.w1(32'h3b06804d),
	.w2(32'hb963b425),
	.w3(32'h3bb11d18),
	.w4(32'hba444eb7),
	.w5(32'h3b198c20),
	.w6(32'h3b11bd7b),
	.w7(32'hbabf42fa),
	.w8(32'h3b96b6c2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391efd77),
	.w1(32'h3af5aa8d),
	.w2(32'h3c69da28),
	.w3(32'h3b8de77e),
	.w4(32'h3bc265cb),
	.w5(32'h3cb5dc8f),
	.w6(32'h3b12ba1f),
	.w7(32'h39802fe1),
	.w8(32'h3cac0838),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4ae9d),
	.w1(32'hbb140cbf),
	.w2(32'hbb667795),
	.w3(32'h3c2f9eb8),
	.w4(32'h3bed0dac),
	.w5(32'hbc712839),
	.w6(32'h3c0f77ee),
	.w7(32'h3bb8aa7f),
	.w8(32'hbbfce10f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae64ae3),
	.w1(32'hb78e4d47),
	.w2(32'hbb8d7a89),
	.w3(32'hbb87b906),
	.w4(32'hbb739a89),
	.w5(32'hbb054027),
	.w6(32'hbaf0e483),
	.w7(32'h3a53e893),
	.w8(32'hbbe26752),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ff2a),
	.w1(32'hbc084052),
	.w2(32'h3a9f84ad),
	.w3(32'hbb48cd83),
	.w4(32'hb8a97317),
	.w5(32'hb7dab76e),
	.w6(32'hba88a9d7),
	.w7(32'h3aa2cee7),
	.w8(32'h3ab1f5cf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa508),
	.w1(32'hbb07ccb4),
	.w2(32'hbba8e8e8),
	.w3(32'hbac896a5),
	.w4(32'hbc315d46),
	.w5(32'hbc446d6d),
	.w6(32'hbb8535d8),
	.w7(32'hba34395e),
	.w8(32'hb9334b5f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3f9cb),
	.w1(32'hbbb197ab),
	.w2(32'hbaf1def7),
	.w3(32'hbbf5cf48),
	.w4(32'hba3f148e),
	.w5(32'hbb504188),
	.w6(32'h3b926409),
	.w7(32'h3985ef4f),
	.w8(32'hba9514fc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec1a1),
	.w1(32'hbc1b1e99),
	.w2(32'hbc4fb113),
	.w3(32'h3a59a29d),
	.w4(32'hbbc5eb4c),
	.w5(32'hbc9f8fee),
	.w6(32'h3bb47d22),
	.w7(32'hbc592d73),
	.w8(32'hbcb59547),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc891365),
	.w1(32'hbbf091c1),
	.w2(32'hb98d62d1),
	.w3(32'hbc7b8a38),
	.w4(32'hbc5d9ca9),
	.w5(32'hbb5a981d),
	.w6(32'hbca17b86),
	.w7(32'hbc0035b5),
	.w8(32'hbac8d618),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6b87),
	.w1(32'h3a49617d),
	.w2(32'hbc48654d),
	.w3(32'h3b4b08e1),
	.w4(32'hbb54e90a),
	.w5(32'hbb26d5ed),
	.w6(32'hbacd1312),
	.w7(32'hbb0faccd),
	.w8(32'h39fd2616),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7d10c),
	.w1(32'h3a8da929),
	.w2(32'hbba64c60),
	.w3(32'hbb1e6a56),
	.w4(32'h3b2c31d0),
	.w5(32'hbc3d9c98),
	.w6(32'h3ba344db),
	.w7(32'h3c43f231),
	.w8(32'hbb9e9f65),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80556c),
	.w1(32'hbb1d4002),
	.w2(32'h3b723ef5),
	.w3(32'hbba9ed36),
	.w4(32'hbbce737f),
	.w5(32'hbc27f5bb),
	.w6(32'hb927709f),
	.w7(32'h394e9e56),
	.w8(32'hbcb7c269),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e3b13),
	.w1(32'hba19503c),
	.w2(32'h3b33f752),
	.w3(32'h3b7b0568),
	.w4(32'hbb9d546f),
	.w5(32'h3c006407),
	.w6(32'h3b2c6530),
	.w7(32'h3be9d79d),
	.w8(32'h3b424f48),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7375),
	.w1(32'h3ad016ed),
	.w2(32'hbc1804a8),
	.w3(32'h3a451413),
	.w4(32'hbb2e9c0c),
	.w5(32'h3ace34c6),
	.w6(32'h3b7816c6),
	.w7(32'h3ba544ba),
	.w8(32'hbc01643f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57be95),
	.w1(32'hb9b9d171),
	.w2(32'hbbda0282),
	.w3(32'h3beb7302),
	.w4(32'h3a7922cb),
	.w5(32'hbbb06176),
	.w6(32'hbb355086),
	.w7(32'h3c1f2161),
	.w8(32'hbbf85bea),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48b020),
	.w1(32'h3b19631d),
	.w2(32'hbbe6df3c),
	.w3(32'hba6ea2a2),
	.w4(32'hbb902b98),
	.w5(32'hbb850a22),
	.w6(32'hb9b54f03),
	.w7(32'h3a3bd10e),
	.w8(32'hbac0c8a4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d932f),
	.w1(32'hb8bcbd93),
	.w2(32'hba91e470),
	.w3(32'hbb8b44f1),
	.w4(32'h399bb74f),
	.w5(32'hbbae1996),
	.w6(32'hbb806757),
	.w7(32'hbbb60fa8),
	.w8(32'hbb898953),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22ca86),
	.w1(32'hbb0a7d7c),
	.w2(32'hbab6fbcb),
	.w3(32'hbb8f4f66),
	.w4(32'hbbc5c354),
	.w5(32'hbbf23000),
	.w6(32'hbb848f33),
	.w7(32'hbb6f88f7),
	.w8(32'hbbabde99),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89caf0),
	.w1(32'h3ada0348),
	.w2(32'h3b7b4135),
	.w3(32'h3a82ce5a),
	.w4(32'hb9df6f41),
	.w5(32'h3c811ecd),
	.w6(32'hba52a349),
	.w7(32'hb9dab419),
	.w8(32'h3c8a67ee),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fddb17),
	.w1(32'hbbfe48c5),
	.w2(32'h3c9544fb),
	.w3(32'h3b982057),
	.w4(32'h3b3eee26),
	.w5(32'h3cf20bba),
	.w6(32'h3b140cd7),
	.w7(32'hb99d2105),
	.w8(32'h3cd16bbb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c585e25),
	.w1(32'h3caf5ab9),
	.w2(32'hbbab515d),
	.w3(32'h3c8fa13e),
	.w4(32'h3cc17634),
	.w5(32'hbb329fa6),
	.w6(32'h3c8beaeb),
	.w7(32'h3cb530a0),
	.w8(32'hbc06e724),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6f882),
	.w1(32'hbc31020c),
	.w2(32'hbc03b7e7),
	.w3(32'h394df1d1),
	.w4(32'h3a0a8273),
	.w5(32'hbbb16e07),
	.w6(32'hbb73fec3),
	.w7(32'h3b151686),
	.w8(32'hbc1066f7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9988b9),
	.w1(32'h38d5c051),
	.w2(32'hbbaeb972),
	.w3(32'h3b2eda43),
	.w4(32'hbb8eae8c),
	.w5(32'hbbc86fff),
	.w6(32'h3ae2ac6c),
	.w7(32'hbbb2fd2f),
	.w8(32'hbb997b69),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef7689),
	.w1(32'hbbea8413),
	.w2(32'hba745b27),
	.w3(32'h3b83896b),
	.w4(32'hbbd80ad5),
	.w5(32'hbb93369f),
	.w6(32'h3aacbafc),
	.w7(32'hba27417a),
	.w8(32'h3b260cbd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c87d5),
	.w1(32'h3a6c134b),
	.w2(32'hba2d1b0b),
	.w3(32'h3c4b0692),
	.w4(32'hbabbd0be),
	.w5(32'hbc5b96ca),
	.w6(32'h3be2fb49),
	.w7(32'h3a2ff1f4),
	.w8(32'hbc0d3087),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb9de),
	.w1(32'hbc06658a),
	.w2(32'hbc0e24cb),
	.w3(32'hbad19c2a),
	.w4(32'hbbe9ad2e),
	.w5(32'h3b554f6d),
	.w6(32'hbb78e4ac),
	.w7(32'hbbfe71a3),
	.w8(32'hbba2511b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b709cc1),
	.w1(32'h3b384bbc),
	.w2(32'hbaa0647e),
	.w3(32'h3bf96c0a),
	.w4(32'hbb1b2736),
	.w5(32'hbaf09af2),
	.w6(32'h3bb3bcf3),
	.w7(32'h3bae5430),
	.w8(32'hbb9f9851),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93569),
	.w1(32'h3ba475cc),
	.w2(32'hbc54f775),
	.w3(32'h3a08ab8d),
	.w4(32'h3b90123d),
	.w5(32'hbbdf5fc0),
	.w6(32'h3c0a6b0c),
	.w7(32'hbba321cd),
	.w8(32'hbb8e4325),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93b4d6),
	.w1(32'h3ad73f97),
	.w2(32'hbb99c53d),
	.w3(32'h3a05907f),
	.w4(32'h3aef667b),
	.w5(32'hbb94fec8),
	.w6(32'h3b30ee6b),
	.w7(32'hbb2f4f60),
	.w8(32'hbb2ec88c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394673e6),
	.w1(32'hbbad6035),
	.w2(32'hb9e3301e),
	.w3(32'h3bd66954),
	.w4(32'hbb6c2e9c),
	.w5(32'hbb9a54b9),
	.w6(32'hb99508d4),
	.w7(32'hbae03e52),
	.w8(32'hbb562d2c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d455e),
	.w1(32'h3a442320),
	.w2(32'h3bdc2c1b),
	.w3(32'hba86a805),
	.w4(32'hbbe0eaa9),
	.w5(32'h3c243a29),
	.w6(32'h3acdf72d),
	.w7(32'hbac895a6),
	.w8(32'h3ba7d5f1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32dbce),
	.w1(32'hbc0c4797),
	.w2(32'h3c1ebe9f),
	.w3(32'hbb0bd999),
	.w4(32'hbc3db69a),
	.w5(32'h3c915e52),
	.w6(32'hbb1a2d61),
	.w7(32'hbc2a2f4b),
	.w8(32'h3c85b9b6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f1796),
	.w1(32'hbc2fa844),
	.w2(32'h3b139a0e),
	.w3(32'h3b04e5f6),
	.w4(32'hbba2f934),
	.w5(32'hbb7d10a6),
	.w6(32'h3997d97b),
	.w7(32'hbb51b740),
	.w8(32'hba93bbdd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dfba4),
	.w1(32'h3c313582),
	.w2(32'hbc5eeea6),
	.w3(32'h3c43e541),
	.w4(32'h3c44fae3),
	.w5(32'hbca8b89f),
	.w6(32'h3c2f8d21),
	.w7(32'h3c6421e4),
	.w8(32'hbc7e13ea),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae49e28),
	.w1(32'h3b0fedc3),
	.w2(32'hba8035a1),
	.w3(32'hbaf05b44),
	.w4(32'h3b4b51f6),
	.w5(32'hb8cb71ba),
	.w6(32'hbb60153d),
	.w7(32'h3aecf3c0),
	.w8(32'hbad54e97),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393915c9),
	.w1(32'h3b8206a5),
	.w2(32'hbb2b42c8),
	.w3(32'h3a4f241b),
	.w4(32'h3b9f1555),
	.w5(32'hbb79a6a8),
	.w6(32'h3b95b594),
	.w7(32'h3a4bb9b1),
	.w8(32'hbb5ab66f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007775),
	.w1(32'hbb65fb97),
	.w2(32'hb84ccd7f),
	.w3(32'hbb8da3ff),
	.w4(32'hbbe90447),
	.w5(32'hbab4d187),
	.w6(32'hbb175fb7),
	.w7(32'hbbb28dea),
	.w8(32'h3b1a2065),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4ef55),
	.w1(32'h3b1b4596),
	.w2(32'hba99421a),
	.w3(32'h3bbcf30c),
	.w4(32'h3b4bcd44),
	.w5(32'hbbed0079),
	.w6(32'hb952cb3c),
	.w7(32'h3b25add5),
	.w8(32'hbbb29147),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c781),
	.w1(32'hbb9262bb),
	.w2(32'hbc57bf8e),
	.w3(32'h3b8badfe),
	.w4(32'hbb0e91ca),
	.w5(32'hbcbab3ca),
	.w6(32'h3b5000da),
	.w7(32'hbb3d14d0),
	.w8(32'hbc9b8ee5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13d0ae),
	.w1(32'hbc1519a3),
	.w2(32'hbb7f3c10),
	.w3(32'hbcae6357),
	.w4(32'hbc83bf25),
	.w5(32'hbbdf4324),
	.w6(32'hbc80ef6b),
	.w7(32'hbc16d491),
	.w8(32'hbbaff70e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b496eae),
	.w1(32'h3a9ea54f),
	.w2(32'hbbc8bf9d),
	.w3(32'h3b59409f),
	.w4(32'h3b4a3ef8),
	.w5(32'hbbcda556),
	.w6(32'h3b14ad93),
	.w7(32'h3a6e02de),
	.w8(32'hba8d80d6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f8f9a),
	.w1(32'h399dd4c4),
	.w2(32'hb9f61633),
	.w3(32'h3b65b7d2),
	.w4(32'hbb970a66),
	.w5(32'h3a807e80),
	.w6(32'h3b49ba82),
	.w7(32'hbc152cfe),
	.w8(32'h3a6d4904),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53ff2b),
	.w1(32'h3b74c087),
	.w2(32'h3b964fa7),
	.w3(32'hb97f0da1),
	.w4(32'h3bc26846),
	.w5(32'h3b55ef5f),
	.w6(32'hba8eeacf),
	.w7(32'h3b1ac39a),
	.w8(32'hbaa182e2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16349b),
	.w1(32'h3bf820d3),
	.w2(32'hbbeaa6cd),
	.w3(32'h3ba600b0),
	.w4(32'h3b5d7043),
	.w5(32'hbc0ba874),
	.w6(32'h3a48234f),
	.w7(32'h3b05a856),
	.w8(32'hbc01255b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7360),
	.w1(32'hb9b5bf9a),
	.w2(32'hbb9f1029),
	.w3(32'hbc3e1467),
	.w4(32'hbbd61a71),
	.w5(32'hbc519e15),
	.w6(32'hbbd26512),
	.w7(32'hbace9f87),
	.w8(32'hbb8d517d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7225c),
	.w1(32'h3a0267d4),
	.w2(32'hbba2ee65),
	.w3(32'hbb33b7ec),
	.w4(32'hbb3fdfb8),
	.w5(32'h3814bd9e),
	.w6(32'hbade2750),
	.w7(32'h3a4f9a63),
	.w8(32'hbb8ef26c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b230395),
	.w1(32'hbbfb0fc9),
	.w2(32'h3be8a0ef),
	.w3(32'hbb38dba5),
	.w4(32'hbc94cf50),
	.w5(32'hb96d906f),
	.w6(32'hba2baa66),
	.w7(32'hbc46602a),
	.w8(32'h3b9a268f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7343e),
	.w1(32'h3a98460c),
	.w2(32'hbacbd15e),
	.w3(32'h39fe4aec),
	.w4(32'hbb645dd0),
	.w5(32'h39370588),
	.w6(32'h3b0b40f0),
	.w7(32'hba5a5dad),
	.w8(32'hba894f86),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c69471),
	.w1(32'h3bb1fc3f),
	.w2(32'hbbc40815),
	.w3(32'h3b7085db),
	.w4(32'hb83ea786),
	.w5(32'hbad315e7),
	.w6(32'h3ae1013c),
	.w7(32'h3b9353cc),
	.w8(32'hba9219d4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bacb0),
	.w1(32'h3b7fd392),
	.w2(32'hbbf4f711),
	.w3(32'h3b5bfb6c),
	.w4(32'h3c3c1258),
	.w5(32'hbc276efd),
	.w6(32'h3b27422d),
	.w7(32'hbaa8e87e),
	.w8(32'hba1a99aa),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226dbe),
	.w1(32'hbb025ebc),
	.w2(32'h3b35a411),
	.w3(32'hbab9a3c3),
	.w4(32'h3bd86595),
	.w5(32'hbb25e290),
	.w6(32'hbba4ccbd),
	.w7(32'hbb1e1e3e),
	.w8(32'h3b069aa6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133de3),
	.w1(32'h3b4067ec),
	.w2(32'hba978eb5),
	.w3(32'hbc5520f5),
	.w4(32'hbb24eb55),
	.w5(32'h3c45e743),
	.w6(32'hbc22b388),
	.w7(32'h3b0e366a),
	.w8(32'hbacb1dc0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe004c),
	.w1(32'hbcc662d1),
	.w2(32'h39caa19b),
	.w3(32'hbc11ed1f),
	.w4(32'hbcfbb518),
	.w5(32'hba1bd8ad),
	.w6(32'hbca47f7b),
	.w7(32'hbcd48ea1),
	.w8(32'h3b71ba75),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6596fb),
	.w1(32'hbb5a55bd),
	.w2(32'hbbf5e82e),
	.w3(32'h3c0b837a),
	.w4(32'hbbd4a8e9),
	.w5(32'hbc3c768b),
	.w6(32'h3bf9b6fb),
	.w7(32'hbc0aadfe),
	.w8(32'hbc03b07e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cdd2c),
	.w1(32'hbc001743),
	.w2(32'hba36acf7),
	.w3(32'hbc6187d4),
	.w4(32'hbc0e6215),
	.w5(32'h3b9d5276),
	.w6(32'hbc274076),
	.w7(32'hbc0d3742),
	.w8(32'h3c2cedb0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79806),
	.w1(32'hbb9d18d1),
	.w2(32'hbb200e45),
	.w3(32'h3c0d049f),
	.w4(32'hbba1fcd2),
	.w5(32'hb9d214fe),
	.w6(32'h3c5dec6e),
	.w7(32'h39c26cfb),
	.w8(32'h3c88483e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe575),
	.w1(32'h3c03dfa2),
	.w2(32'hbb772a4a),
	.w3(32'h3c3266e7),
	.w4(32'h3c6608ea),
	.w5(32'hbb9ae9ad),
	.w6(32'h3ca1e976),
	.w7(32'h3bd325fa),
	.w8(32'hbb4d50eb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe2219),
	.w1(32'h3bcd6012),
	.w2(32'hbb477766),
	.w3(32'hbb1658c0),
	.w4(32'h3bf5a14f),
	.w5(32'hbb391ff7),
	.w6(32'h3b91543f),
	.w7(32'h3c29eded),
	.w8(32'hbb5ef0b3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9fbb0),
	.w1(32'h3a22822a),
	.w2(32'hbba846b4),
	.w3(32'h3a5127fb),
	.w4(32'hba66e797),
	.w5(32'hbabeb29f),
	.w6(32'h3b769b4b),
	.w7(32'hbaf4f6aa),
	.w8(32'hbb8d6bca),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58e6f5),
	.w1(32'hbb8a1e61),
	.w2(32'h3bbf1c7d),
	.w3(32'hbb2ea5fe),
	.w4(32'hba91157c),
	.w5(32'hba2b73d7),
	.w6(32'hba822fe6),
	.w7(32'h3adb34b8),
	.w8(32'hbc51081a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a367af5),
	.w1(32'hbb0b57e5),
	.w2(32'hbcafa82c),
	.w3(32'hba815d83),
	.w4(32'hbb8602a2),
	.w5(32'hbcc2c6b4),
	.w6(32'hbbcbd4b0),
	.w7(32'hbc06bcbe),
	.w8(32'hbc8867d9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc23b38),
	.w1(32'hbc61d1ec),
	.w2(32'hbc1e54e6),
	.w3(32'hbcee023d),
	.w4(32'hbc0cabc9),
	.w5(32'hbb925aaf),
	.w6(32'hbc6537ac),
	.w7(32'hbb5865b8),
	.w8(32'hbb58b21a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1258c7),
	.w1(32'hbc0d79b2),
	.w2(32'hbc2d842e),
	.w3(32'h3b3e484f),
	.w4(32'hbc2573af),
	.w5(32'hbb796e31),
	.w6(32'h3aa4f02e),
	.w7(32'h3ad4c8a7),
	.w8(32'hbc43fd24),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dad31),
	.w1(32'hbc2436e1),
	.w2(32'hbbcee96f),
	.w3(32'h3c3397b3),
	.w4(32'hbc4f9bf9),
	.w5(32'h3a9f2a55),
	.w6(32'h3ba9062f),
	.w7(32'hbb7461e1),
	.w8(32'hbb262d6e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c434c18),
	.w1(32'hbba6bd1f),
	.w2(32'hba9c922c),
	.w3(32'h3cc6cc1c),
	.w4(32'h391e5d3c),
	.w5(32'h3a1a28d2),
	.w6(32'h3c8fd3fa),
	.w7(32'h3992e682),
	.w8(32'h3adb1fa6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10ecc1),
	.w1(32'h3c43a8ef),
	.w2(32'hb9e0b183),
	.w3(32'h3bdb210a),
	.w4(32'h3bb72829),
	.w5(32'hbb9e8ec2),
	.w6(32'h3bab3162),
	.w7(32'h3c3b4fd3),
	.w8(32'h3bd412ff),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9163bf),
	.w1(32'h3ada08b6),
	.w2(32'hbc1d412a),
	.w3(32'h3c508af1),
	.w4(32'hbb33fbc2),
	.w5(32'hbc84f881),
	.w6(32'h3be0126d),
	.w7(32'hb9f50cdb),
	.w8(32'hbc3b28ed),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2acadf),
	.w1(32'hbb7285db),
	.w2(32'hbb864dad),
	.w3(32'hbc8d7e14),
	.w4(32'hbb969289),
	.w5(32'h3a265a7d),
	.w6(32'hbbe58e5c),
	.w7(32'h3a591e5c),
	.w8(32'h3c14f720),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e2165),
	.w1(32'hbb745eb6),
	.w2(32'h3c57f160),
	.w3(32'h3c61bc56),
	.w4(32'h3b849e68),
	.w5(32'h3b5679d3),
	.w6(32'h3c2d7dc4),
	.w7(32'hba8b1aee),
	.w8(32'h3ac752cc),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20a325),
	.w1(32'h3bae426b),
	.w2(32'h3b83489b),
	.w3(32'h3bc8e5ac),
	.w4(32'h3c872b5c),
	.w5(32'hba396e3b),
	.w6(32'h3b951b31),
	.w7(32'h3c0e37a1),
	.w8(32'hb94a9905),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0a909),
	.w1(32'h3a5490d4),
	.w2(32'h3ac84970),
	.w3(32'h3c319d9e),
	.w4(32'h3b761f00),
	.w5(32'h3bc7df5d),
	.w6(32'h3c061bc3),
	.w7(32'h3b1f6787),
	.w8(32'hbb20c54f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e52fd),
	.w1(32'h3bafbede),
	.w2(32'hbb573ccf),
	.w3(32'h3cc27201),
	.w4(32'h3c4e0c9a),
	.w5(32'hbae71637),
	.w6(32'h3c848502),
	.w7(32'h3bbdb49c),
	.w8(32'hb9224d62),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242b50),
	.w1(32'hbb4ea28f),
	.w2(32'h3b7bf599),
	.w3(32'hb9609798),
	.w4(32'hbab06a8c),
	.w5(32'h3c319d20),
	.w6(32'h3b12673e),
	.w7(32'hb9fa46e4),
	.w8(32'h3bcbb8fc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1a48d),
	.w1(32'h3bdc488f),
	.w2(32'hb872377e),
	.w3(32'h3c4d27ed),
	.w4(32'h3c19c7d1),
	.w5(32'hbbb78fd5),
	.w6(32'h3c096134),
	.w7(32'h3bfb68d1),
	.w8(32'hbbbdde18),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47427),
	.w1(32'hbb93e3d4),
	.w2(32'hbc34e8b9),
	.w3(32'hbc05005c),
	.w4(32'hbb8d84b4),
	.w5(32'hbc658b7c),
	.w6(32'hbbc56a44),
	.w7(32'hbb12d1e5),
	.w8(32'hbbe1b6bb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29eae1),
	.w1(32'hbc54337c),
	.w2(32'h3ae3277f),
	.w3(32'h3c68c308),
	.w4(32'hbbcff59b),
	.w5(32'hbb4d3b5e),
	.w6(32'h3c7aa62c),
	.w7(32'hbbbec036),
	.w8(32'h3b4993f4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc549c54),
	.w1(32'hbbebdf7e),
	.w2(32'hbc47efcf),
	.w3(32'hb8f9d1e8),
	.w4(32'h3b09b200),
	.w5(32'hbbb12d86),
	.w6(32'hba7be653),
	.w7(32'h3bb64e02),
	.w8(32'h38f64ce0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccd243),
	.w1(32'hbabdc760),
	.w2(32'h3b68be50),
	.w3(32'h3be3517e),
	.w4(32'h3c226257),
	.w5(32'h3c0c9e70),
	.w6(32'h3c0f7603),
	.w7(32'h3abdd8a9),
	.w8(32'h3ab9e78a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be33302),
	.w1(32'h3b2fe0d5),
	.w2(32'hb9f06854),
	.w3(32'h3b80b0c9),
	.w4(32'hba4eb456),
	.w5(32'hbc065330),
	.w6(32'h3adeb3e2),
	.w7(32'h3bdce2a8),
	.w8(32'h3bcb0c1d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175ab7),
	.w1(32'h3c28beda),
	.w2(32'h3b83fc2e),
	.w3(32'hbbc44fe3),
	.w4(32'h3b3bd206),
	.w5(32'h3c153c07),
	.w6(32'h3ba77f98),
	.w7(32'h3bc02927),
	.w8(32'h3c1e4584),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c85526),
	.w1(32'h3bc87b77),
	.w2(32'h3c3388de),
	.w3(32'hbb9c1296),
	.w4(32'h3bcd7f81),
	.w5(32'h3c1d3649),
	.w6(32'h3b9c677b),
	.w7(32'h3b26d609),
	.w8(32'hb9cfb5ec),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45e589),
	.w1(32'h3b876a54),
	.w2(32'h39f65e38),
	.w3(32'h3bb99fbb),
	.w4(32'h3b43bbc5),
	.w5(32'hba1b8dcc),
	.w6(32'hbb531780),
	.w7(32'h3c42dd90),
	.w8(32'h3b86b4b1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb684988),
	.w1(32'hba31a0f7),
	.w2(32'h3a57e2ae),
	.w3(32'hbb9f36ef),
	.w4(32'h3b8cf78b),
	.w5(32'h3c029cf4),
	.w6(32'h3c0e5210),
	.w7(32'h3ca4b96f),
	.w8(32'hbb247090),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a3645),
	.w1(32'h3b824a4e),
	.w2(32'h3b0d16be),
	.w3(32'h3c9c5759),
	.w4(32'h3bfc04d6),
	.w5(32'hbbb9ff61),
	.w6(32'h3ac81df5),
	.w7(32'hb9cc000a),
	.w8(32'hbb4359bc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd64aa),
	.w1(32'h3a8137e3),
	.w2(32'hbac1f062),
	.w3(32'h3c1ab15e),
	.w4(32'h3bfe26b8),
	.w5(32'hbad4cbf4),
	.w6(32'h3c230e84),
	.w7(32'h3baa4c42),
	.w8(32'h3b895e42),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd24bb),
	.w1(32'h3c512246),
	.w2(32'h3b3bf99c),
	.w3(32'hbb4e7512),
	.w4(32'h3b7870d9),
	.w5(32'h3c016a44),
	.w6(32'h3b6f1ea1),
	.w7(32'h37700a67),
	.w8(32'h3aa02051),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f4411),
	.w1(32'h3c1def83),
	.w2(32'h3ac8b365),
	.w3(32'h3cd06638),
	.w4(32'h3c7dd405),
	.w5(32'hbc2ea390),
	.w6(32'h3c9ed3b5),
	.w7(32'h3c0015ba),
	.w8(32'hba9eaa60),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc468315),
	.w1(32'hbb2acfde),
	.w2(32'hbb81b41b),
	.w3(32'hbcbfdc50),
	.w4(32'hbc2983b5),
	.w5(32'hba524adf),
	.w6(32'hbc4806e6),
	.w7(32'hbb404c1d),
	.w8(32'hbc083a7f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ea24d3),
	.w1(32'hbab80fd3),
	.w2(32'hba54778b),
	.w3(32'hbad5017c),
	.w4(32'h3b127080),
	.w5(32'h3badd0f8),
	.w6(32'hbbaafb57),
	.w7(32'hbc2dff92),
	.w8(32'h3c3d55cb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe60502),
	.w1(32'hbc811e65),
	.w2(32'hbc4c4beb),
	.w3(32'hbb07721a),
	.w4(32'hbc5c28ed),
	.w5(32'hbcb9ccee),
	.w6(32'h3befd217),
	.w7(32'hbbd03dba),
	.w8(32'hbc1e70d8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5021fc),
	.w1(32'h39b8dcf7),
	.w2(32'hba834f00),
	.w3(32'hbcc5dbf6),
	.w4(32'hb810158e),
	.w5(32'hbad9d0c6),
	.w6(32'hbbbf84d0),
	.w7(32'h3bfe0edc),
	.w8(32'hb93ddfbf),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd9f55),
	.w1(32'hbb068594),
	.w2(32'h3c193905),
	.w3(32'h3c4744ac),
	.w4(32'h39e544cf),
	.w5(32'h3bf0e341),
	.w6(32'h3c32c284),
	.w7(32'h39769f1d),
	.w8(32'h3bb46feb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9efdfb),
	.w1(32'h3c3e8c95),
	.w2(32'h3b1e402f),
	.w3(32'h3cadd27b),
	.w4(32'h3c006ee7),
	.w5(32'h3a82d8df),
	.w6(32'h3c28ba8b),
	.w7(32'h3c0e7a60),
	.w8(32'h39c065b6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66bcdf),
	.w1(32'hbb41999f),
	.w2(32'hbb2b8fdb),
	.w3(32'hbc84288e),
	.w4(32'hbb94a4d7),
	.w5(32'hb98300c8),
	.w6(32'hbc8930a6),
	.w7(32'hbb89f623),
	.w8(32'h3c155e9d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c869b2c),
	.w1(32'h3be414ec),
	.w2(32'h3b26c9de),
	.w3(32'h3cf9f26a),
	.w4(32'h3c6b49b1),
	.w5(32'h3bc42e8a),
	.w6(32'h3cf61183),
	.w7(32'h3be710e4),
	.w8(32'h3af8d59c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffecce),
	.w1(32'hbbdc9161),
	.w2(32'hbbb77611),
	.w3(32'h3c6bd8b4),
	.w4(32'hbbce3998),
	.w5(32'hbb69ea6a),
	.w6(32'h3c3a87f6),
	.w7(32'hbb8b2cb6),
	.w8(32'hbb495c77),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc04396),
	.w1(32'h38f57870),
	.w2(32'hbca68333),
	.w3(32'h3c245686),
	.w4(32'h3b0a3360),
	.w5(32'hbce3af6c),
	.w6(32'h3c50d5b3),
	.w7(32'h3b70ae14),
	.w8(32'hbc90098e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85000d),
	.w1(32'hbbd5f54e),
	.w2(32'hbafc6c8a),
	.w3(32'hbcfba8d8),
	.w4(32'hbc95c68b),
	.w5(32'hbbe800b9),
	.w6(32'hbcb244f5),
	.w7(32'hbc238704),
	.w8(32'h3a94e177),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9838b),
	.w1(32'hbbd94b86),
	.w2(32'hba8fb361),
	.w3(32'hbcf03ebb),
	.w4(32'hbc2d89f3),
	.w5(32'h3a44a84a),
	.w6(32'hbcad845d),
	.w7(32'hbb8259fb),
	.w8(32'hbbe03482),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c017776),
	.w1(32'hba042869),
	.w2(32'h3aa33b6e),
	.w3(32'h3ca375d5),
	.w4(32'h3bf18270),
	.w5(32'hba8cb85a),
	.w6(32'h3c5260fe),
	.w7(32'h3a101b68),
	.w8(32'h3a344ad3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a5629),
	.w1(32'h3a654639),
	.w2(32'hb8ecd49a),
	.w3(32'h3a09c4ed),
	.w4(32'hbb0995fa),
	.w5(32'hbb932b7b),
	.w6(32'h3ae82e03),
	.w7(32'hba61da30),
	.w8(32'h37c55795),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9602),
	.w1(32'hbb95c140),
	.w2(32'h3bd4ebd0),
	.w3(32'hbb5bfc35),
	.w4(32'hbb6d1aec),
	.w5(32'h3b6552eb),
	.w6(32'hbb82ac72),
	.w7(32'h3b032f16),
	.w8(32'h3aad416b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0e255),
	.w1(32'h3c681f48),
	.w2(32'h3b11b887),
	.w3(32'h3c54d768),
	.w4(32'h3c03f5bd),
	.w5(32'h3bec27ef),
	.w6(32'h3c936483),
	.w7(32'h3bbedc43),
	.w8(32'h3a9609f4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f2b6),
	.w1(32'h3b60d0dc),
	.w2(32'h3b3ca68a),
	.w3(32'h39c3e2a3),
	.w4(32'h3bb5c72e),
	.w5(32'hbbf48a6e),
	.w6(32'hbc148856),
	.w7(32'h3acc0da7),
	.w8(32'hb9e3fc1e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff8325),
	.w1(32'h3906b7f0),
	.w2(32'hbbc89cb8),
	.w3(32'h3c17475a),
	.w4(32'h3b4db363),
	.w5(32'hbca3aa37),
	.w6(32'h3c2f768f),
	.w7(32'h3bbe7438),
	.w8(32'hbc21f8c4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadd37e),
	.w1(32'h39954920),
	.w2(32'h3bf631cf),
	.w3(32'hbd13b360),
	.w4(32'hbbe3b418),
	.w5(32'h3bf385b7),
	.w6(32'hbcb7463d),
	.w7(32'hb82baebc),
	.w8(32'h3ac4785a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87ff83),
	.w1(32'h39da9594),
	.w2(32'h3b8c85a0),
	.w3(32'h3c3ff0e4),
	.w4(32'h3a5cf367),
	.w5(32'hb9e9f3e2),
	.w6(32'h3c526bf3),
	.w7(32'h38e79733),
	.w8(32'hbbeda014),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a779c7a),
	.w1(32'hbaadab90),
	.w2(32'hba1ab11e),
	.w3(32'h3c297b22),
	.w4(32'h3bbd2762),
	.w5(32'hbb49b6ba),
	.w6(32'h3c2bb3ae),
	.w7(32'h3c1cce4c),
	.w8(32'h3b9b8d54),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7b9ca),
	.w1(32'h3be99e52),
	.w2(32'h3b05d818),
	.w3(32'h3bb5e438),
	.w4(32'h3aa2116b),
	.w5(32'h3c275322),
	.w6(32'h392f7a64),
	.w7(32'hbbf3167a),
	.w8(32'h39de3757),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9025ee),
	.w1(32'h3aa0bdb9),
	.w2(32'h3ae203ee),
	.w3(32'h3bc2ad65),
	.w4(32'h391eb669),
	.w5(32'h3b9dfb3a),
	.w6(32'h3b1f405c),
	.w7(32'h3c546aa6),
	.w8(32'h3bbe1852),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28e22c),
	.w1(32'hbc9e3d71),
	.w2(32'hbc61faf1),
	.w3(32'hbc39ef76),
	.w4(32'hbcb867e0),
	.w5(32'hbc771add),
	.w6(32'hbb9255fe),
	.w7(32'hbc4b70f1),
	.w8(32'hbc8a0dfa),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc422c09),
	.w1(32'hbc1b0968),
	.w2(32'h3b44a727),
	.w3(32'hbc4429f0),
	.w4(32'hbc01f729),
	.w5(32'h3ab71cfd),
	.w6(32'hbc758ad3),
	.w7(32'hbc4a75cd),
	.w8(32'h3ba7a122),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb212b27),
	.w1(32'hbb9a876c),
	.w2(32'hbb8661a3),
	.w3(32'h3b793898),
	.w4(32'hba0b8bbb),
	.w5(32'hbb8147cc),
	.w6(32'h3b5aa3ee),
	.w7(32'h3b8688f4),
	.w8(32'h3b4bf66c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399558ad),
	.w1(32'hbb5cc720),
	.w2(32'hbcbdd5f6),
	.w3(32'h3c0cedff),
	.w4(32'hbb979ab0),
	.w5(32'hbc96b5b7),
	.w6(32'h3caaafb6),
	.w7(32'h3a9a306c),
	.w8(32'h3c208bbc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd206a83),
	.w1(32'hbca59037),
	.w2(32'hbc4cb222),
	.w3(32'hbc78fd3a),
	.w4(32'hbb6c8a9c),
	.w5(32'hbc57a119),
	.w6(32'h3cea0c79),
	.w7(32'h3ca8cad5),
	.w8(32'hbc23f226),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc705b7b),
	.w1(32'hbc76e0c4),
	.w2(32'hbb0c0476),
	.w3(32'hbc8c098c),
	.w4(32'hbc474a68),
	.w5(32'hbb45fc5c),
	.w6(32'hbc600035),
	.w7(32'hbc18969f),
	.w8(32'hbb60693a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcc1c2),
	.w1(32'hba8fb78b),
	.w2(32'h3aba91a2),
	.w3(32'hbc14c5d0),
	.w4(32'hbb649caf),
	.w5(32'h3a65f66f),
	.w6(32'hbbe92905),
	.w7(32'hbab7386f),
	.w8(32'hb95686db),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdce188),
	.w1(32'h3ba88c9a),
	.w2(32'h3ba75e69),
	.w3(32'h3c355746),
	.w4(32'h3c0d598e),
	.w5(32'h3bb334cc),
	.w6(32'h3bff11e6),
	.w7(32'h3bffe240),
	.w8(32'h3c23793c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237130),
	.w1(32'h3bd55460),
	.w2(32'hb99e9d4c),
	.w3(32'h3c84aade),
	.w4(32'h3c438019),
	.w5(32'hbbb9d81b),
	.w6(32'h3c1bf6bf),
	.w7(32'h3c1c94ca),
	.w8(32'hbb844aa0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f381),
	.w1(32'hbc33ff7e),
	.w2(32'h3c0ea8bc),
	.w3(32'h3bb02286),
	.w4(32'hbc41674e),
	.w5(32'h3c0961e6),
	.w6(32'hbb56c552),
	.w7(32'hbccea2de),
	.w8(32'h3b2ec1e6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41c91f),
	.w1(32'h3bf9ee81),
	.w2(32'hbc1e3fd7),
	.w3(32'h3c811cb6),
	.w4(32'h3bca8ca2),
	.w5(32'hbbb06cb1),
	.w6(32'h3c35fe21),
	.w7(32'h3bd28d14),
	.w8(32'hbbc2a575),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a03d),
	.w1(32'h3b190e11),
	.w2(32'h3b8228be),
	.w3(32'h3bc87cc9),
	.w4(32'h3a9a8d48),
	.w5(32'h3baf2ba6),
	.w6(32'h3a0ee287),
	.w7(32'hbaf73cca),
	.w8(32'h3b87256f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba100e8c),
	.w1(32'h3be82138),
	.w2(32'hbcb28c5e),
	.w3(32'h3b50a01a),
	.w4(32'h3c22a518),
	.w5(32'hbd08c813),
	.w6(32'h3ca5e906),
	.w7(32'h3c808847),
	.w8(32'hbcd8be6d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bed42),
	.w1(32'h3cb734a9),
	.w2(32'hbb53873f),
	.w3(32'hbbd6532e),
	.w4(32'h3d2989ab),
	.w5(32'h3b87c796),
	.w6(32'hbbb4cae0),
	.w7(32'h3cdc8003),
	.w8(32'hba9c1f01),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d12e6),
	.w1(32'hbb6df212),
	.w2(32'hbbed0e73),
	.w3(32'h3b6ddd4d),
	.w4(32'h3a015eda),
	.w5(32'hbb3fedaa),
	.w6(32'h3bb1b476),
	.w7(32'hbb9188cd),
	.w8(32'hbb5e5936),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9e842),
	.w1(32'hbb33786d),
	.w2(32'h3aa606fa),
	.w3(32'hbc28bfd0),
	.w4(32'hbb65ccf5),
	.w5(32'h3afd35f4),
	.w6(32'hbb994336),
	.w7(32'hbb2eef7e),
	.w8(32'h3b84f560),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242a04),
	.w1(32'hb9ed40bd),
	.w2(32'hbc20d65c),
	.w3(32'hbbbd3349),
	.w4(32'hbb055e42),
	.w5(32'hbc4ee9d3),
	.w6(32'hbb907303),
	.w7(32'hbbf402ad),
	.w8(32'hbbbf0df2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9f83a),
	.w1(32'hbab01834),
	.w2(32'h3ba8885e),
	.w3(32'h3b0e0063),
	.w4(32'h3c2a3bdd),
	.w5(32'h3ba06b01),
	.w6(32'h3c249c23),
	.w7(32'h3c903a79),
	.w8(32'h3c08e8af),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabbff1),
	.w1(32'h3c2fbf9c),
	.w2(32'h3b533077),
	.w3(32'h3af8922e),
	.w4(32'h3c8ea01c),
	.w5(32'h3b03aed7),
	.w6(32'h3c043875),
	.w7(32'h3c82f970),
	.w8(32'h3ae9be0c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14e729),
	.w1(32'hbb096801),
	.w2(32'h3c1b9daa),
	.w3(32'h3b5c0400),
	.w4(32'hbb90705a),
	.w5(32'h3c653303),
	.w6(32'h3c19e858),
	.w7(32'h3b89786e),
	.w8(32'h3c313966),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16e079),
	.w1(32'hbb24bfa6),
	.w2(32'hbc148561),
	.w3(32'h3c55cd87),
	.w4(32'hbb85acc1),
	.w5(32'h3b1cf705),
	.w6(32'h3c678e40),
	.w7(32'h3ab6e57f),
	.w8(32'hbc2d61ee),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c1373),
	.w1(32'h3c06c707),
	.w2(32'hbb14902a),
	.w3(32'h3c9dafe9),
	.w4(32'h3cb7c9dd),
	.w5(32'hbc66ee55),
	.w6(32'h3b35d9af),
	.w7(32'h3be8a9dd),
	.w8(32'hbbbdbce0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26c363),
	.w1(32'h3be6c8c9),
	.w2(32'h3bb6929f),
	.w3(32'h3b28f6a0),
	.w4(32'h3bcfd957),
	.w5(32'hbb842e45),
	.w6(32'hbb8f324f),
	.w7(32'hbba03c4b),
	.w8(32'hbadf51b3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0437cc),
	.w1(32'h3c00e5e9),
	.w2(32'hbb9ba87a),
	.w3(32'h3bdbcb06),
	.w4(32'h39f9c2e8),
	.w5(32'h396a9ad5),
	.w6(32'h3c04afdb),
	.w7(32'h3bb57f87),
	.w8(32'hbb6761ca),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60aac1),
	.w1(32'h3bb88998),
	.w2(32'hbb6ef195),
	.w3(32'hbacb98b2),
	.w4(32'hbb99b05f),
	.w5(32'hba20d98d),
	.w6(32'h3bbfa29e),
	.w7(32'hbbde7c57),
	.w8(32'h39e6aca0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52bf4e),
	.w1(32'h3b9230c7),
	.w2(32'h3a2af96f),
	.w3(32'h3bc7bbe9),
	.w4(32'h3b22747d),
	.w5(32'h3ae05ca8),
	.w6(32'h3c0098c8),
	.w7(32'h3ac9fe0d),
	.w8(32'h3ad5c243),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac86d4),
	.w1(32'h3b4f9e92),
	.w2(32'h3b07a94e),
	.w3(32'h3c83cd79),
	.w4(32'h3b833ac8),
	.w5(32'h3ac462bd),
	.w6(32'h3cb62154),
	.w7(32'h3bff464b),
	.w8(32'h3b8731f4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c292d6f),
	.w1(32'h3bffc216),
	.w2(32'h3bf17d59),
	.w3(32'h3c372908),
	.w4(32'h3c3dffc8),
	.w5(32'h3bceedf2),
	.w6(32'h3c37865b),
	.w7(32'h3bd4e1c0),
	.w8(32'h3bb6ac6f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b1e47),
	.w1(32'h3c07d622),
	.w2(32'h3bafcbfc),
	.w3(32'h3aa17cf4),
	.w4(32'h3bbd5047),
	.w5(32'h3b9ba785),
	.w6(32'hba9c7ad4),
	.w7(32'h3b5713bf),
	.w8(32'hbc5f25ce),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c487aff),
	.w1(32'h3c18f472),
	.w2(32'hbc4fccda),
	.w3(32'h3c177b7c),
	.w4(32'h3c2a7db7),
	.w5(32'h3be8f46b),
	.w6(32'hbc6daf8f),
	.w7(32'hbc351139),
	.w8(32'h3c13464a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcf849),
	.w1(32'hbb175126),
	.w2(32'h3b65c707),
	.w3(32'h3cccd321),
	.w4(32'h3c7e710d),
	.w5(32'hbb83e44d),
	.w6(32'h3cd933ff),
	.w7(32'h3c715efb),
	.w8(32'hbc6eb76d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c372c07),
	.w1(32'h3b71bf8a),
	.w2(32'h3aae37a4),
	.w3(32'h3b8d39ec),
	.w4(32'h3916db25),
	.w5(32'h3c07de5f),
	.w6(32'hbc33c641),
	.w7(32'hbc2b6e80),
	.w8(32'h3bcb24ce),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e4a11),
	.w1(32'hbad27699),
	.w2(32'hbb094e87),
	.w3(32'h3c3208ff),
	.w4(32'hba1a64c5),
	.w5(32'h3894c1c4),
	.w6(32'h3c4fdf7f),
	.w7(32'h3b05d01b),
	.w8(32'hbb309162),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807b24),
	.w1(32'h3b0adf9b),
	.w2(32'hbb20f115),
	.w3(32'h3b21cdf0),
	.w4(32'h3bcb1917),
	.w5(32'h3b85d675),
	.w6(32'hbb9dbcbc),
	.w7(32'hbb9b9614),
	.w8(32'h3b8b4911),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dc6ac),
	.w1(32'h3ba09143),
	.w2(32'hbc0534b2),
	.w3(32'h3c6087ef),
	.w4(32'h3c58ecc0),
	.w5(32'hbc2093a8),
	.w6(32'h3c5c6ed7),
	.w7(32'h3bb0b0d7),
	.w8(32'hbc1735f9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc447d7e),
	.w1(32'hbc2afc7c),
	.w2(32'h3b86495e),
	.w3(32'hbc5cd0dc),
	.w4(32'hbc5ecf95),
	.w5(32'h3bde8595),
	.w6(32'hbc54a952),
	.w7(32'hbc57000c),
	.w8(32'h3bb067a2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3cd1),
	.w1(32'h3b5f2be9),
	.w2(32'h3c06fe26),
	.w3(32'h3c63a258),
	.w4(32'h3bb757af),
	.w5(32'h3c5942b4),
	.w6(32'h3c196029),
	.w7(32'h3ae350e9),
	.w8(32'h3bb2b814),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62d0d3),
	.w1(32'h3c5ce3f8),
	.w2(32'h3c04ad98),
	.w3(32'h3b9dffc9),
	.w4(32'h3c002de3),
	.w5(32'h3c1f1f6f),
	.w6(32'h3bc005f1),
	.w7(32'h3c60a31f),
	.w8(32'hbaaeb0a7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33dfa6),
	.w1(32'hbc402793),
	.w2(32'hbb280429),
	.w3(32'h3b858eae),
	.w4(32'hbc57eabb),
	.w5(32'h3c266c58),
	.w6(32'hbbd34c0f),
	.w7(32'hbc870456),
	.w8(32'h3bb4a430),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09d706),
	.w1(32'h39866adf),
	.w2(32'hb9c5e034),
	.w3(32'h3c5d9683),
	.w4(32'h3c043cb2),
	.w5(32'h3ad6c5fd),
	.w6(32'h3c997339),
	.w7(32'h3b1ddef5),
	.w8(32'hbb308d69),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd385b),
	.w1(32'hbb2b6a06),
	.w2(32'hbbb3217e),
	.w3(32'hbb821372),
	.w4(32'h3ac37011),
	.w5(32'hbb13fcfb),
	.w6(32'hbb358709),
	.w7(32'h3ab0cb67),
	.w8(32'h3b2f0286),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba5cac),
	.w1(32'hbbaf9122),
	.w2(32'hbb409392),
	.w3(32'h3c81f2e2),
	.w4(32'h3b17367e),
	.w5(32'h3b64a0e3),
	.w6(32'h3bc795a2),
	.w7(32'h3a6c7489),
	.w8(32'hbba6bab6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule