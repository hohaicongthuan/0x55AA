module layer_10_featuremap_2(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a74c),
	.w1(32'h3acb79ca),
	.w2(32'h3b514fb2),
	.w3(32'h3c4cf427),
	.w4(32'h3be11214),
	.w5(32'h3c508a0f),
	.w6(32'h3cad2a88),
	.w7(32'h3c3539f8),
	.w8(32'h3c04342b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb384b1f),
	.w1(32'h3bc0a25b),
	.w2(32'hbaaf57ae),
	.w3(32'h3bbeaf51),
	.w4(32'h3bc391c4),
	.w5(32'hbba5f513),
	.w6(32'h3c949027),
	.w7(32'h3c4bd497),
	.w8(32'h3b9a3e69),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99a1df),
	.w1(32'hbc9d2c60),
	.w2(32'hbbf7a216),
	.w3(32'hbcce0763),
	.w4(32'hbd097273),
	.w5(32'hbbbeca6d),
	.w6(32'hbc83d59c),
	.w7(32'hbcaff97b),
	.w8(32'h3bdb54d1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0c34d),
	.w1(32'hba848bb6),
	.w2(32'h3ab4bf7e),
	.w3(32'h3c384eed),
	.w4(32'h3c938e99),
	.w5(32'hbb3e616a),
	.w6(32'h3ba20c98),
	.w7(32'h3c100997),
	.w8(32'hbba3291a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcace42),
	.w1(32'h3c26e65a),
	.w2(32'h3b32f5cc),
	.w3(32'hb971cf6a),
	.w4(32'h3c2ea54a),
	.w5(32'h3b45aacf),
	.w6(32'h3c65eb53),
	.w7(32'h3cb6314b),
	.w8(32'hbae02ec6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb69443),
	.w1(32'hbb4fea4e),
	.w2(32'hbc1578c3),
	.w3(32'h3bced2f8),
	.w4(32'h3a98b53b),
	.w5(32'hbc40ec01),
	.w6(32'h3b8998d6),
	.w7(32'h3b3c6801),
	.w8(32'hbb950605),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4246c2),
	.w1(32'h3be64671),
	.w2(32'h3c1fcac3),
	.w3(32'h3bd403a1),
	.w4(32'h3bf87c9f),
	.w5(32'h3a1b8f92),
	.w6(32'h3c437ae4),
	.w7(32'h3c4b4f7d),
	.w8(32'h3c2f8d45),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a138),
	.w1(32'hbc024c85),
	.w2(32'h3bd8954e),
	.w3(32'hbbc35941),
	.w4(32'hbc1d95ed),
	.w5(32'h3b63e899),
	.w6(32'h3b8fc677),
	.w7(32'h3c0c8b95),
	.w8(32'h3ba7968e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10305f),
	.w1(32'h3bad18b9),
	.w2(32'hbc246461),
	.w3(32'hba454e59),
	.w4(32'hbb3e5044),
	.w5(32'hbb29ff8f),
	.w6(32'hbbb02225),
	.w7(32'hbc17b44d),
	.w8(32'hbaa4e346),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51ff14),
	.w1(32'h3cd0c025),
	.w2(32'h3ada0191),
	.w3(32'h3d25c00c),
	.w4(32'h3d5d8a9c),
	.w5(32'h3b8eac78),
	.w6(32'h3d24be48),
	.w7(32'h3d43a642),
	.w8(32'h3b94a53f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8719b9),
	.w1(32'h3b1af672),
	.w2(32'hbbd1ac2b),
	.w3(32'h3c0ec465),
	.w4(32'h3b98410f),
	.w5(32'hbbe3483f),
	.w6(32'h3bfd4de7),
	.w7(32'h3b5914b3),
	.w8(32'hb9d00f8c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31c731),
	.w1(32'h3b390fad),
	.w2(32'hbb073c6d),
	.w3(32'h3b8a5ca3),
	.w4(32'h3c4e9285),
	.w5(32'hbba1eb95),
	.w6(32'h3c6bad29),
	.w7(32'h3c8569b5),
	.w8(32'hba252aa0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cc123),
	.w1(32'h3c00c6df),
	.w2(32'h3bc028a8),
	.w3(32'h3a1da404),
	.w4(32'h3bd570b9),
	.w5(32'h3b723911),
	.w6(32'h3b80b38d),
	.w7(32'h3c322c6f),
	.w8(32'h3bbfd715),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ab029),
	.w1(32'h3c978090),
	.w2(32'h3b406534),
	.w3(32'h3c6f72d9),
	.w4(32'h3c2760ec),
	.w5(32'h3b7d1308),
	.w6(32'h3c727d1c),
	.w7(32'h3c87dbbb),
	.w8(32'h3bccd0c1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1eb1e),
	.w1(32'h3bf223d3),
	.w2(32'hbb637f19),
	.w3(32'h3b5e0dc4),
	.w4(32'h3c83a0d4),
	.w5(32'hbb0729a1),
	.w6(32'h3b628e6a),
	.w7(32'h3bf4c949),
	.w8(32'h3ac78bd2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd080e),
	.w1(32'hb9846478),
	.w2(32'h3b976269),
	.w3(32'h3af42b0d),
	.w4(32'h3b935659),
	.w5(32'h3b8668fb),
	.w6(32'hbac69e3f),
	.w7(32'hb89a1f86),
	.w8(32'h3b624693),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cd687),
	.w1(32'hbab7dc24),
	.w2(32'h3bc57514),
	.w3(32'h3a599d54),
	.w4(32'hbbb4c0a5),
	.w5(32'h3b87e78d),
	.w6(32'hba17efc1),
	.w7(32'hbbec9aba),
	.w8(32'h3c32b0c4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63af2b),
	.w1(32'hbbd27f28),
	.w2(32'h3b458082),
	.w3(32'hbc16416e),
	.w4(32'hbc7529c7),
	.w5(32'hb91a1c6b),
	.w6(32'hb8d8e3c9),
	.w7(32'hbc5648bf),
	.w8(32'h3bb136bf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c073e81),
	.w1(32'h3c1c646d),
	.w2(32'hbb9c7116),
	.w3(32'h3c2c146c),
	.w4(32'h3c29cab4),
	.w5(32'hba68186a),
	.w6(32'h3b7bcd4f),
	.w7(32'h3bee1448),
	.w8(32'h3abda40d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56b325),
	.w1(32'h3b501b14),
	.w2(32'h3b2c5c39),
	.w3(32'hbb8d3533),
	.w4(32'hbc7563c5),
	.w5(32'hbb74323e),
	.w6(32'h372a4a07),
	.w7(32'hbc3c6ac0),
	.w8(32'hba82a70f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aa4c4),
	.w1(32'hbad0f7fb),
	.w2(32'hbb70f3b2),
	.w3(32'hbac3f074),
	.w4(32'h38b492d9),
	.w5(32'hbbf2dd21),
	.w6(32'h3a409364),
	.w7(32'h3b2d67ec),
	.w8(32'hbae7c7fa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676514),
	.w1(32'h3c0a0da7),
	.w2(32'hbb264f0f),
	.w3(32'h3bfe63da),
	.w4(32'h3c4d022d),
	.w5(32'hbb4942dd),
	.w6(32'h3c2c7f9d),
	.w7(32'h3bda8f51),
	.w8(32'hbb87b36a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac014c9),
	.w1(32'hbb6687aa),
	.w2(32'hbbc215b6),
	.w3(32'h3a9835c3),
	.w4(32'hbc1db8e6),
	.w5(32'hbb7e1351),
	.w6(32'hbac3f98f),
	.w7(32'hbbb3874e),
	.w8(32'hbba5781d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b974df3),
	.w1(32'h3c141bf4),
	.w2(32'h3b4e2891),
	.w3(32'h3c274fcd),
	.w4(32'h3c52f0a7),
	.w5(32'h3b87864c),
	.w6(32'h3c096cf8),
	.w7(32'h3c441ec0),
	.w8(32'h3bf3135d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa0b6a),
	.w1(32'h3ac666c5),
	.w2(32'hbb05f105),
	.w3(32'h3bf29bce),
	.w4(32'h3bb5bf17),
	.w5(32'h3b3e27a5),
	.w6(32'h3ba0dc38),
	.w7(32'h3be62650),
	.w8(32'h3b4d7f25),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba0f29),
	.w1(32'h3c146534),
	.w2(32'hbb8f7c3f),
	.w3(32'h3c30afa5),
	.w4(32'h3b5dc01a),
	.w5(32'hbb8d61fb),
	.w6(32'h3ba0d869),
	.w7(32'h3bca99fc),
	.w8(32'hbbbdc2eb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf70270),
	.w1(32'h3b3a00b7),
	.w2(32'hb82fd0bd),
	.w3(32'hbb872b6c),
	.w4(32'h3c30a84a),
	.w5(32'hbb03e0c6),
	.w6(32'h3b59ffaa),
	.w7(32'h3bd01025),
	.w8(32'hb85555fc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab63527),
	.w1(32'h375bca5d),
	.w2(32'hbc31e70a),
	.w3(32'h3ac7b8dd),
	.w4(32'hbade09ec),
	.w5(32'hbc5fee9c),
	.w6(32'h3ac20b7d),
	.w7(32'hb8cd02d6),
	.w8(32'h3bee875e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca594fe),
	.w1(32'h3ad67ab9),
	.w2(32'hbc40df13),
	.w3(32'h3a6e71e9),
	.w4(32'h3c9e15f0),
	.w5(32'h3bb331e5),
	.w6(32'h3c692e4d),
	.w7(32'h3c46855e),
	.w8(32'h3b95dbed),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc412acd),
	.w1(32'hbb595c1a),
	.w2(32'h3ab0ab99),
	.w3(32'h3bb09846),
	.w4(32'h3b6f30d3),
	.w5(32'hbb8d404b),
	.w6(32'h3cbc0b12),
	.w7(32'h3bf0b360),
	.w8(32'h3b5335ef),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62c3a9),
	.w1(32'h3ad41db6),
	.w2(32'h3bad96cd),
	.w3(32'hbbcd8d79),
	.w4(32'h3a2a9b2d),
	.w5(32'h3c94e961),
	.w6(32'h3b33e416),
	.w7(32'h3c27a600),
	.w8(32'hbb192a42),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51db2e),
	.w1(32'hbbc554ad),
	.w2(32'hbac7510c),
	.w3(32'h3c55692e),
	.w4(32'hbbba5946),
	.w5(32'h3cedfb9f),
	.w6(32'hbab21ae0),
	.w7(32'hbc0acbd5),
	.w8(32'h3bb045f3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1760eb),
	.w1(32'h3b5a4eb8),
	.w2(32'hbbb28170),
	.w3(32'h3ca4aec5),
	.w4(32'h3c5737aa),
	.w5(32'hbbc0bba0),
	.w6(32'h3b3dc9e6),
	.w7(32'hbb690157),
	.w8(32'h3b03d9cb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe112a1),
	.w1(32'hb8f64e75),
	.w2(32'h3c27871e),
	.w3(32'hbb449cbf),
	.w4(32'h3aed5409),
	.w5(32'hbb81d2ac),
	.w6(32'h3bac3c5f),
	.w7(32'h3b81a30e),
	.w8(32'hb9d41262),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b7e17),
	.w1(32'hbb45fc6f),
	.w2(32'hbb1ec744),
	.w3(32'hbac7bd61),
	.w4(32'hbc22d73c),
	.w5(32'hbb4a1c20),
	.w6(32'hbc1e4268),
	.w7(32'hbb7fc4f7),
	.w8(32'hbb7196d9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc050d),
	.w1(32'hbaccddfd),
	.w2(32'hbce84f2f),
	.w3(32'h3965f658),
	.w4(32'hbaa2192f),
	.w5(32'hbb194b09),
	.w6(32'hbb69233e),
	.w7(32'hbc0714d2),
	.w8(32'h3c17adc4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf173c6),
	.w1(32'hbc105e7a),
	.w2(32'hbc4d7393),
	.w3(32'h3c6e98be),
	.w4(32'h3cca9e67),
	.w5(32'hbc032400),
	.w6(32'h3bdc878b),
	.w7(32'h3c42b257),
	.w8(32'hbafb6237),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccede6),
	.w1(32'h3b970d59),
	.w2(32'hbaba6743),
	.w3(32'h3a54096c),
	.w4(32'h3aff10b6),
	.w5(32'h3b29d181),
	.w6(32'h39233152),
	.w7(32'hbb63ddc7),
	.w8(32'h3c596d16),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb490f85),
	.w1(32'hbb572c29),
	.w2(32'h3bbad871),
	.w3(32'h3c4a64dc),
	.w4(32'h3be39911),
	.w5(32'h3a497547),
	.w6(32'h3c9a5ade),
	.w7(32'h3c1551ed),
	.w8(32'h3c0b0a19),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d737),
	.w1(32'h3aef608c),
	.w2(32'hba179290),
	.w3(32'h3ab19206),
	.w4(32'hbc0b34d5),
	.w5(32'hbb46fcb7),
	.w6(32'h3c51398b),
	.w7(32'hb99086e7),
	.w8(32'h3b4c55a6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596b83),
	.w1(32'hbbec674b),
	.w2(32'hbc1886e9),
	.w3(32'hbbeb3e16),
	.w4(32'hbc0b143a),
	.w5(32'hbb33810f),
	.w6(32'h3aeae67c),
	.w7(32'hba8a6917),
	.w8(32'h3b7f7457),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8aeef9),
	.w1(32'hbc0c54fd),
	.w2(32'h3c0bffb5),
	.w3(32'h3a330dd4),
	.w4(32'h3bcd5357),
	.w5(32'hbb5c1d4a),
	.w6(32'h3c380e11),
	.w7(32'h3ba01700),
	.w8(32'h3b8bce3d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acde01c),
	.w1(32'hbbc5f08f),
	.w2(32'hbba8f6a0),
	.w3(32'hbb9a122c),
	.w4(32'hbb72419b),
	.w5(32'hbb25bba5),
	.w6(32'hbb7d4373),
	.w7(32'hbb05c1e4),
	.w8(32'hbc0817a8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8372e),
	.w1(32'hba13e1a5),
	.w2(32'h3c54d440),
	.w3(32'h3ba1f3d7),
	.w4(32'hbb4cf822),
	.w5(32'h3ba5cae0),
	.w6(32'hbbee916e),
	.w7(32'hbc748fe8),
	.w8(32'hbb21bd6f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c736b1e),
	.w1(32'h3bd24ba9),
	.w2(32'h3ba432d4),
	.w3(32'h3be99aef),
	.w4(32'hbb719eb5),
	.w5(32'hbbe79f71),
	.w6(32'h3ba1a3e0),
	.w7(32'h3b134859),
	.w8(32'hbbdaf555),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081094),
	.w1(32'hba6a2ccc),
	.w2(32'h3be8e17a),
	.w3(32'hbc6be4c0),
	.w4(32'h3a97d1ef),
	.w5(32'hbb08c8d6),
	.w6(32'h3bcab4c0),
	.w7(32'h3bc2965a),
	.w8(32'hbb310ca1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1a38b),
	.w1(32'hbab70791),
	.w2(32'h3be0c89c),
	.w3(32'h3a8c4b84),
	.w4(32'h3844c75c),
	.w5(32'hbc3c03f2),
	.w6(32'hbaa8f92c),
	.w7(32'h3c545dfd),
	.w8(32'hbc2e8fbb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fe3ac),
	.w1(32'h3b49ae77),
	.w2(32'h3a830b88),
	.w3(32'hbc500444),
	.w4(32'hbba45b44),
	.w5(32'h3b39d458),
	.w6(32'hbc25a534),
	.w7(32'hb926d7fc),
	.w8(32'hbbb0c78d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86ee71),
	.w1(32'h3b0b1957),
	.w2(32'h3bb9a9f9),
	.w3(32'h3bdbd83a),
	.w4(32'h3b37e8df),
	.w5(32'hbb54e1ac),
	.w6(32'hbb9de5af),
	.w7(32'hbbe26b4b),
	.w8(32'hbae7bcc5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3be414),
	.w1(32'h3ae74850),
	.w2(32'hbb85be6d),
	.w3(32'hbbc18fe9),
	.w4(32'hbba6be0a),
	.w5(32'h3b121bbc),
	.w6(32'hbb41a1c9),
	.w7(32'h3b035128),
	.w8(32'hba9cf277),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc794d),
	.w1(32'hbc17843d),
	.w2(32'h3c314ecc),
	.w3(32'h3aa87013),
	.w4(32'hbc0b1c3d),
	.w5(32'h3c0f4307),
	.w6(32'hbbf783d5),
	.w7(32'hb8f77135),
	.w8(32'hbc56498d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ea656),
	.w1(32'hbb813d1c),
	.w2(32'h3b0d0386),
	.w3(32'hbc5ec964),
	.w4(32'hbc90f80b),
	.w5(32'h3ba52fe1),
	.w6(32'hbb879873),
	.w7(32'hba388f65),
	.w8(32'hbb05d5d3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e7b0f),
	.w1(32'h3b1fe91d),
	.w2(32'h3c282a03),
	.w3(32'h393fbbc1),
	.w4(32'hbaffc540),
	.w5(32'h3cb76e99),
	.w6(32'hbb83790d),
	.w7(32'hbb358e28),
	.w8(32'hbbc186f7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad5509),
	.w1(32'h3be5ac48),
	.w2(32'hb9536571),
	.w3(32'h3c49a7cc),
	.w4(32'hbbb456fd),
	.w5(32'hbb39012f),
	.w6(32'hbc83d534),
	.w7(32'hbc2d8d7f),
	.w8(32'h3b7eb5a4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be34fc2),
	.w1(32'hbbbc5702),
	.w2(32'h3b8b4e69),
	.w3(32'h3b8d2b05),
	.w4(32'h3bb6daed),
	.w5(32'h3c40debb),
	.w6(32'h3bd5c88a),
	.w7(32'h3bc7a124),
	.w8(32'h3bf08858),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c800a5a),
	.w1(32'h3c36d9bd),
	.w2(32'h3b77ff73),
	.w3(32'h3c68f027),
	.w4(32'hbb9dab3b),
	.w5(32'hbc8451bc),
	.w6(32'hbaaf4903),
	.w7(32'hbc7f8eab),
	.w8(32'hbc35e881),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7b3d8),
	.w1(32'h3b255d76),
	.w2(32'h3b9f5c6e),
	.w3(32'hbc0d1cf3),
	.w4(32'h3bf2cdec),
	.w5(32'h3a11dd59),
	.w6(32'h3bdbecaf),
	.w7(32'h3c2234e9),
	.w8(32'h3b162230),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08454),
	.w1(32'h3b55e87c),
	.w2(32'hbba06a53),
	.w3(32'hbb7f1aa8),
	.w4(32'h3be7c951),
	.w5(32'hbba63cba),
	.w6(32'h3ba38a9e),
	.w7(32'h3c1013cc),
	.w8(32'h3b986560),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab055d),
	.w1(32'hbab0d212),
	.w2(32'hbbadba39),
	.w3(32'hbab3618c),
	.w4(32'hbb41dae6),
	.w5(32'hbb1da2b4),
	.w6(32'h3bb030d1),
	.w7(32'h3b21e3c1),
	.w8(32'h3c0b9281),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b4e8e),
	.w1(32'hba82cc40),
	.w2(32'h3ba17d5f),
	.w3(32'h38c3fe51),
	.w4(32'h3c0ef990),
	.w5(32'hbc242637),
	.w6(32'h3c92725e),
	.w7(32'h3c2e5b73),
	.w8(32'hb83d2967),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d443b),
	.w1(32'h3a4b1d85),
	.w2(32'h3a9c2012),
	.w3(32'hbc6697fc),
	.w4(32'hbb4631f1),
	.w5(32'hbbd5abe7),
	.w6(32'h3bf4c876),
	.w7(32'h3c6d56c7),
	.w8(32'hbb0aee24),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f32c),
	.w1(32'hbc16bfec),
	.w2(32'hb900604f),
	.w3(32'hbc0ff3d4),
	.w4(32'hbb94fe64),
	.w5(32'hb9fa6538),
	.w6(32'hbb12ec65),
	.w7(32'h3be609dc),
	.w8(32'h3c2096b9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a303ed1),
	.w1(32'h3b6f12d4),
	.w2(32'hbc1fafd6),
	.w3(32'h3bc99808),
	.w4(32'h3bb76fa9),
	.w5(32'h39e30f1c),
	.w6(32'h3c9ba0ed),
	.w7(32'h3c942817),
	.w8(32'h3bc85fa5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a3552),
	.w1(32'hbb20a604),
	.w2(32'hbb0cfa07),
	.w3(32'h3c2b4b99),
	.w4(32'h3c5d4f19),
	.w5(32'h3bb5b41e),
	.w6(32'h3c479b4c),
	.w7(32'h3c376e45),
	.w8(32'hbb286b52),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e89db),
	.w1(32'hbc08b5ea),
	.w2(32'h3c0fd9bf),
	.w3(32'h3c1f6999),
	.w4(32'h3b0b9de0),
	.w5(32'h3c3dbee3),
	.w6(32'hbb7b91fc),
	.w7(32'hbbe70100),
	.w8(32'h3ad94877),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b683b),
	.w1(32'h3acd3853),
	.w2(32'h39126b5d),
	.w3(32'h3b9ddb24),
	.w4(32'hb7b8c989),
	.w5(32'h3b59b945),
	.w6(32'hbb1751cb),
	.w7(32'hbadf9f14),
	.w8(32'h3b4abb30),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a2a52),
	.w1(32'h3ba21807),
	.w2(32'h3b41b8ed),
	.w3(32'h3c1ca740),
	.w4(32'h3b5d6f94),
	.w5(32'h3bad4739),
	.w6(32'h3b963fa0),
	.w7(32'hbb6bdca3),
	.w8(32'h3b47408e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16b78e),
	.w1(32'h391a5cbc),
	.w2(32'h3c01c90e),
	.w3(32'hbb4dd8c3),
	.w4(32'h3afd2182),
	.w5(32'h3b9c6b57),
	.w6(32'hbba64a4a),
	.w7(32'hbb22bb64),
	.w8(32'h3bdced68),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6136ee),
	.w1(32'h3c48a271),
	.w2(32'hba07968f),
	.w3(32'h3c2c6344),
	.w4(32'h3beef070),
	.w5(32'hbb243fb6),
	.w6(32'h3c0c9a4b),
	.w7(32'h3beafa6f),
	.w8(32'h3b4af325),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56691e),
	.w1(32'hbae6e4c3),
	.w2(32'h3bcdef46),
	.w3(32'hbb8689bf),
	.w4(32'hbb73f848),
	.w5(32'hbb12cd25),
	.w6(32'h3adb87f9),
	.w7(32'hba2bb99a),
	.w8(32'hbc297ff1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56cd13),
	.w1(32'h3a491480),
	.w2(32'h3c2d017d),
	.w3(32'hbb063575),
	.w4(32'hbbf797c0),
	.w5(32'h3ade839e),
	.w6(32'hbc24104a),
	.w7(32'h3b0feaa5),
	.w8(32'h3938f3ee),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be96bdc),
	.w1(32'hbb78a64e),
	.w2(32'hbbbe8e42),
	.w3(32'h3b5fffe1),
	.w4(32'hbb869de6),
	.w5(32'hbb5042a1),
	.w6(32'h3ad7f343),
	.w7(32'h3ab94d9d),
	.w8(32'hbb48f34a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af00ffa),
	.w1(32'hbba1a8af),
	.w2(32'h3b022327),
	.w3(32'hbb847019),
	.w4(32'h3955b43a),
	.w5(32'h3bb1954b),
	.w6(32'h3ada52cd),
	.w7(32'h3c00ff9f),
	.w8(32'h3b7aa96a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ff2ab),
	.w1(32'h3c146142),
	.w2(32'h3ba03250),
	.w3(32'h3bbfd83f),
	.w4(32'h3c04a763),
	.w5(32'h3ac612e9),
	.w6(32'hbac8e464),
	.w7(32'h3ac17837),
	.w8(32'h35deb035),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24b74f),
	.w1(32'h3bcb3890),
	.w2(32'hbaed2899),
	.w3(32'hb9baf099),
	.w4(32'h3ba13b30),
	.w5(32'hbc197156),
	.w6(32'hbba5b503),
	.w7(32'h3a07dd3d),
	.w8(32'hbc35b65d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba502a1),
	.w1(32'hbc3f65a2),
	.w2(32'hbc0269c2),
	.w3(32'hbc627f18),
	.w4(32'hbc322df3),
	.w5(32'hbb72db46),
	.w6(32'hbc230737),
	.w7(32'hbb3b6015),
	.w8(32'hbc0cd4a0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985d5c4),
	.w1(32'hbacf2425),
	.w2(32'hbc9e7161),
	.w3(32'hbb7d24fd),
	.w4(32'hbc45da77),
	.w5(32'h3a093281),
	.w6(32'hbbf0d672),
	.w7(32'hbc3b59a4),
	.w8(32'hbcb0dd0e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4261),
	.w1(32'hbbb1df6e),
	.w2(32'h38105f34),
	.w3(32'hbb6d755c),
	.w4(32'hbc9afebf),
	.w5(32'hbc8c8578),
	.w6(32'hbcc49907),
	.w7(32'hbca7abd5),
	.w8(32'hbb55300e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e0393),
	.w1(32'hbaaf13d9),
	.w2(32'h3b15c945),
	.w3(32'hbc17836a),
	.w4(32'h3b2d3df4),
	.w5(32'hbb7b909f),
	.w6(32'h3b838a38),
	.w7(32'h3c1f7405),
	.w8(32'h3b46ec3b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb668823),
	.w1(32'h3adc203a),
	.w2(32'h3c1519a5),
	.w3(32'hbc322659),
	.w4(32'hbbdf72b0),
	.w5(32'h3b2e40c9),
	.w6(32'hbb1fe178),
	.w7(32'h3ac1f04f),
	.w8(32'hbab982ad),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2af4b5),
	.w1(32'h3c0ae4b0),
	.w2(32'hbba8f5e9),
	.w3(32'h3b8f460c),
	.w4(32'hb98fe2c7),
	.w5(32'hbc26cab2),
	.w6(32'hbb944a42),
	.w7(32'hbb9cf701),
	.w8(32'hb903e5ff),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6b8d3),
	.w1(32'hbb25b20e),
	.w2(32'h3ad946f5),
	.w3(32'hbc098225),
	.w4(32'hbb49538c),
	.w5(32'h3a9953c9),
	.w6(32'h3b1c0ff5),
	.w7(32'h3b6f35d0),
	.w8(32'hba32f30d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51203e),
	.w1(32'h3b4948f9),
	.w2(32'hbb0d45c2),
	.w3(32'hbba155e0),
	.w4(32'h3c1e854f),
	.w5(32'h3a9825f4),
	.w6(32'hbc00159f),
	.w7(32'h3b9fe37e),
	.w8(32'h3c3eeeee),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa44aa8),
	.w1(32'hbac893b7),
	.w2(32'hbbdb22d7),
	.w3(32'hba3f2553),
	.w4(32'hbba16062),
	.w5(32'hbba5329d),
	.w6(32'h3b9e32b7),
	.w7(32'h3c043735),
	.w8(32'h3ba61c98),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeca10b),
	.w1(32'h3a9857ef),
	.w2(32'hbba394bb),
	.w3(32'hba809628),
	.w4(32'h3bcd5f1c),
	.w5(32'hbc188475),
	.w6(32'h3c2fbeb7),
	.w7(32'h3c814075),
	.w8(32'hbb30b748),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a39ff),
	.w1(32'hbc6e5f72),
	.w2(32'hbb3be4b6),
	.w3(32'hbc37d244),
	.w4(32'h3b9033fb),
	.w5(32'h38f7aaad),
	.w6(32'h3c28c19a),
	.w7(32'h3bb2f406),
	.w8(32'hba1cc73f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc135c09),
	.w1(32'hbc353454),
	.w2(32'h39c518a6),
	.w3(32'h38888e93),
	.w4(32'hbbf004a3),
	.w5(32'hbb52dbbe),
	.w6(32'h3b339eb9),
	.w7(32'hba83cc88),
	.w8(32'hbb772fbc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b64042),
	.w1(32'hba29b3ae),
	.w2(32'h3b048aea),
	.w3(32'hbb8c9d20),
	.w4(32'hb9f57617),
	.w5(32'h3b07cdde),
	.w6(32'hbac6752b),
	.w7(32'h39bfc845),
	.w8(32'h39a997f8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1de3b5),
	.w1(32'h3b716db3),
	.w2(32'h3bfe0d1f),
	.w3(32'h3b8e6015),
	.w4(32'hbbaab2d0),
	.w5(32'h3c8094e2),
	.w6(32'hbb957f2f),
	.w7(32'hbb120174),
	.w8(32'hbc615ab5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ddae6),
	.w1(32'hb987d217),
	.w2(32'h3c5bdb6d),
	.w3(32'h3be11f72),
	.w4(32'hbb845d13),
	.w5(32'h3c6e959b),
	.w6(32'hbcb091d6),
	.w7(32'hbca351ca),
	.w8(32'hbbd410c2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d9ca7),
	.w1(32'h3bca0c06),
	.w2(32'h3c510424),
	.w3(32'h3c7bbf5c),
	.w4(32'hbb85b8eb),
	.w5(32'h3c1754b9),
	.w6(32'hbcaaaf33),
	.w7(32'hbc5274f5),
	.w8(32'h3c7d40ec),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd53513),
	.w1(32'h3c2e3737),
	.w2(32'hbb8e865d),
	.w3(32'h3c0497fd),
	.w4(32'h3c705a8a),
	.w5(32'hbb959302),
	.w6(32'h3c9c7670),
	.w7(32'h3c8b5814),
	.w8(32'hbb1d3248),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963005),
	.w1(32'hbb48ca31),
	.w2(32'h3b0987e9),
	.w3(32'hbba4004e),
	.w4(32'hbb9875f4),
	.w5(32'hbbe1a146),
	.w6(32'hbb8b335f),
	.w7(32'hbb19c2d7),
	.w8(32'hbb303e62),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181fc0),
	.w1(32'h3b00eef8),
	.w2(32'h3bc985da),
	.w3(32'hbb8e3791),
	.w4(32'hba0bccc9),
	.w5(32'h3be301b4),
	.w6(32'h3b002807),
	.w7(32'h3b7cf57d),
	.w8(32'h3b0b533e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab76734),
	.w1(32'h3b43255f),
	.w2(32'h3bc62086),
	.w3(32'h3b95a391),
	.w4(32'h3b2cc2a6),
	.w5(32'h3c06f54b),
	.w6(32'h3b7bb153),
	.w7(32'h3b8f11b8),
	.w8(32'hbbd5b9d3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c745630),
	.w1(32'h3c28cba2),
	.w2(32'hbb4f9fc0),
	.w3(32'hbc009b92),
	.w4(32'hbc4fcc19),
	.w5(32'hbbe5611b),
	.w6(32'hbcbc1706),
	.w7(32'hbc5af4b6),
	.w8(32'hbc1b0532),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd69849),
	.w1(32'hbbc63483),
	.w2(32'h39943425),
	.w3(32'hbadcb903),
	.w4(32'h3bb2d5bd),
	.w5(32'h3b84534b),
	.w6(32'hbb3f453d),
	.w7(32'hbaef4a42),
	.w8(32'h3b63b6cf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe8519),
	.w1(32'hbc042dc7),
	.w2(32'hbac7f008),
	.w3(32'h3c44f855),
	.w4(32'h3ba5ac58),
	.w5(32'h3bc51eb2),
	.w6(32'h3c5bebb2),
	.w7(32'h3c91fef8),
	.w8(32'hbb8ada8b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67c490),
	.w1(32'h3b6de159),
	.w2(32'hbb091fe2),
	.w3(32'h3b8feed1),
	.w4(32'h3955ec5e),
	.w5(32'h3ae225e5),
	.w6(32'hbbe71068),
	.w7(32'hbc7f57c5),
	.w8(32'h3ba9c675),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c397095),
	.w1(32'h3c043eca),
	.w2(32'h3badd379),
	.w3(32'h3be6576b),
	.w4(32'hbb9e78c5),
	.w5(32'h3ac3dfa6),
	.w6(32'h3b0dc449),
	.w7(32'hbbefc780),
	.w8(32'h3af465cf),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac68c7),
	.w1(32'h3b384e0e),
	.w2(32'hbb01f137),
	.w3(32'h3afb42d2),
	.w4(32'h3a4cee1e),
	.w5(32'h3ba8da5f),
	.w6(32'hba091d1d),
	.w7(32'hbc01067f),
	.w8(32'hbc17840c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1bc4b),
	.w1(32'hba4136da),
	.w2(32'hbc96d09f),
	.w3(32'h3b954baa),
	.w4(32'hbb46c69f),
	.w5(32'hbaf44c67),
	.w6(32'hbbcf019f),
	.w7(32'hbc4c111f),
	.w8(32'h3bb08977),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03958d),
	.w1(32'h39ca45de),
	.w2(32'h3c4a592e),
	.w3(32'h3c9a62eb),
	.w4(32'h3c73c06d),
	.w5(32'h3c5a18c8),
	.w6(32'h3ca4ae01),
	.w7(32'h3b50349d),
	.w8(32'hbbea8517),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84358e),
	.w1(32'h3b1464da),
	.w2(32'h3b9df277),
	.w3(32'h3a0d5e6d),
	.w4(32'hbc5512e8),
	.w5(32'hba63ba36),
	.w6(32'hbca6b866),
	.w7(32'hbcbf7111),
	.w8(32'h3a40c392),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8850be1),
	.w1(32'hbb11fff1),
	.w2(32'h3b4d6908),
	.w3(32'hba42b3e4),
	.w4(32'h3b9ddcbc),
	.w5(32'h3b1f3214),
	.w6(32'hbc240ba6),
	.w7(32'hb91a0e19),
	.w8(32'h3b4a23e8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad03aa),
	.w1(32'h3b0a092e),
	.w2(32'h3b91905a),
	.w3(32'h3c3c4ff5),
	.w4(32'h3c062072),
	.w5(32'h3bdd7e3c),
	.w6(32'h3bf7d277),
	.w7(32'h3b978784),
	.w8(32'h3b9f7567),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98f8b3),
	.w1(32'hb929cb23),
	.w2(32'hbb99c62a),
	.w3(32'hb972c057),
	.w4(32'h3b1bfb0e),
	.w5(32'h3a3ca924),
	.w6(32'hb60ce6ba),
	.w7(32'h3a943ed6),
	.w8(32'h3b095432),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ea2f2),
	.w1(32'hbb4aa165),
	.w2(32'hbb7c7ebe),
	.w3(32'h3b64c2b8),
	.w4(32'h3b024e84),
	.w5(32'h3c053d0f),
	.w6(32'h3bca5c1c),
	.w7(32'h3bcb25c1),
	.w8(32'h3b81a6f3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fa785),
	.w1(32'h3bd4b469),
	.w2(32'h3c04e41b),
	.w3(32'h3a9bf458),
	.w4(32'hbb541cb2),
	.w5(32'h3bf38aa7),
	.w6(32'h3c218228),
	.w7(32'h3c282780),
	.w8(32'hbc6209d1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0295b),
	.w1(32'hbbcb7026),
	.w2(32'hbac65c6e),
	.w3(32'h3c31d1f4),
	.w4(32'h3b1d40a1),
	.w5(32'h3b2aa514),
	.w6(32'hbc3b379f),
	.w7(32'hbc137d04),
	.w8(32'h3bfde457),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934f48),
	.w1(32'hbbbb2212),
	.w2(32'h3ac89f22),
	.w3(32'h3ad96660),
	.w4(32'h3b89cb67),
	.w5(32'hbbc04b8e),
	.w6(32'h3c00246d),
	.w7(32'h3c1c5a15),
	.w8(32'hbbc97f84),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88c1b2),
	.w1(32'hb9b62c1b),
	.w2(32'hbbbb9d5c),
	.w3(32'hbc2b43bb),
	.w4(32'hbc06dd59),
	.w5(32'h3c103ddd),
	.w6(32'hbbc1d0c4),
	.w7(32'hbb8d08d8),
	.w8(32'h3c07ea51),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b9c5a),
	.w1(32'h3c1954d1),
	.w2(32'h3be2e992),
	.w3(32'h3c8453fd),
	.w4(32'h3afda304),
	.w5(32'hb9c58e2e),
	.w6(32'hbb944952),
	.w7(32'hbb513ed2),
	.w8(32'hbc027c96),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb527068),
	.w1(32'hbc1ec2e0),
	.w2(32'hbc7c9a42),
	.w3(32'h3a9a2b84),
	.w4(32'hbbcc2057),
	.w5(32'hbc54f5d9),
	.w6(32'hbb5fc1f3),
	.w7(32'hbbde7d57),
	.w8(32'h3ba28ca0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca1f1e),
	.w1(32'hbc527d65),
	.w2(32'hbc43b596),
	.w3(32'hbc7f932a),
	.w4(32'hbc009e1f),
	.w5(32'hbc0325c1),
	.w6(32'h3bd81efe),
	.w7(32'h3c037fdb),
	.w8(32'h3b5f7c3b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc709b9d),
	.w1(32'hbb67e789),
	.w2(32'h3c677d75),
	.w3(32'hbb898a4a),
	.w4(32'h3b377dc3),
	.w5(32'h3c0562a0),
	.w6(32'h3c0a3347),
	.w7(32'h3c1aaf00),
	.w8(32'hbb32c8c1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35643d),
	.w1(32'hbb3e5015),
	.w2(32'hbc8d7a52),
	.w3(32'hbab51c04),
	.w4(32'hbbe353a8),
	.w5(32'hbbac1cc3),
	.w6(32'hbba699b7),
	.w7(32'h3ba0be87),
	.w8(32'h3b75d57c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c2e92),
	.w1(32'hbc0bf0c7),
	.w2(32'h3b9888f4),
	.w3(32'hbb0c4342),
	.w4(32'h3b9e7f25),
	.w5(32'h3bd44244),
	.w6(32'h3c3425ca),
	.w7(32'h3c25b877),
	.w8(32'h3b020226),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90bf8d),
	.w1(32'h3c00a947),
	.w2(32'hb9c2fbfc),
	.w3(32'h3c5a86fa),
	.w4(32'h3bed72d8),
	.w5(32'h3c7f4cbd),
	.w6(32'h3ad4c76f),
	.w7(32'hbbdfb296),
	.w8(32'hba3070d8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395c5b),
	.w1(32'hba57a743),
	.w2(32'hbb1be590),
	.w3(32'h3c1ea749),
	.w4(32'h3bc0fe7a),
	.w5(32'h3af78d05),
	.w6(32'hbb081741),
	.w7(32'hbc10fa32),
	.w8(32'h3be97002),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab868fe),
	.w1(32'h3b8a78f8),
	.w2(32'h3aa058c3),
	.w3(32'h3bc5bbae),
	.w4(32'h3b2d4fab),
	.w5(32'hba492d2e),
	.w6(32'h3c6bcb7a),
	.w7(32'h3c7cfd91),
	.w8(32'hbaa17e29),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d6dd),
	.w1(32'h3a4701c5),
	.w2(32'h3ac459b0),
	.w3(32'hbb345389),
	.w4(32'h3ac2194c),
	.w5(32'hbb9ef750),
	.w6(32'hb913c107),
	.w7(32'h3b8316d9),
	.w8(32'hbb9bbbdf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801aaa),
	.w1(32'hbb4e8331),
	.w2(32'hbc59adfe),
	.w3(32'hbc1630cf),
	.w4(32'hbbc582af),
	.w5(32'h3b7a7397),
	.w6(32'hbbc54410),
	.w7(32'h3ad6191e),
	.w8(32'h3c4f66c7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd47724),
	.w1(32'hbbca276b),
	.w2(32'hbc351891),
	.w3(32'h3ca43210),
	.w4(32'h3c2ef527),
	.w5(32'hbb558032),
	.w6(32'h3c33bec2),
	.w7(32'h3c03695b),
	.w8(32'h3bc13fa2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dea00),
	.w1(32'hbb52565b),
	.w2(32'h3bf8bbe9),
	.w3(32'hbac68b6b),
	.w4(32'h3c019e2e),
	.w5(32'h3b5f5e01),
	.w6(32'h3c31ce19),
	.w7(32'h3c403bb2),
	.w8(32'hbba4c109),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8715df),
	.w1(32'h3bd21c15),
	.w2(32'h3b2c060d),
	.w3(32'hbba67244),
	.w4(32'h3ae443ff),
	.w5(32'hbaa3bfa2),
	.w6(32'hbb86b158),
	.w7(32'hbc049970),
	.w8(32'hbb453a22),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891e47),
	.w1(32'hba118a76),
	.w2(32'h3c216bd0),
	.w3(32'h39fb49c5),
	.w4(32'h3ad64028),
	.w5(32'hbaee87e2),
	.w6(32'hbb3b1342),
	.w7(32'hbba0b89c),
	.w8(32'hbc00b211),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfe6ad),
	.w1(32'hbb898b7f),
	.w2(32'h3bcb657c),
	.w3(32'hbc1e1738),
	.w4(32'hbb492d04),
	.w5(32'hbc00f343),
	.w6(32'hbbbbc27c),
	.w7(32'h3b609c07),
	.w8(32'hbafd3d6f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72e416),
	.w1(32'hbb3791a1),
	.w2(32'hbc18e3b5),
	.w3(32'hbc7617e5),
	.w4(32'hbc29c89f),
	.w5(32'h3b96cd2d),
	.w6(32'h3b85108a),
	.w7(32'h3b9ad950),
	.w8(32'h3b4cf4fb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0107b3),
	.w1(32'hba855325),
	.w2(32'hbbe7401a),
	.w3(32'h3bedb152),
	.w4(32'h3aeb5832),
	.w5(32'h3a4330c1),
	.w6(32'h393d252d),
	.w7(32'h3b792922),
	.w8(32'h3c4381e0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f3c1d),
	.w1(32'hbad88ff9),
	.w2(32'h3b9c83fd),
	.w3(32'hb9ca4aee),
	.w4(32'h3b8e44a9),
	.w5(32'h3b188323),
	.w6(32'h3a7679e6),
	.w7(32'hbb9610be),
	.w8(32'h3c1f2556),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb51974),
	.w1(32'hba3c7dba),
	.w2(32'hbc486520),
	.w3(32'h3bbe05e6),
	.w4(32'h3b429edd),
	.w5(32'hbbcddc9a),
	.w6(32'h3c319d42),
	.w7(32'h3c0885d1),
	.w8(32'h3c0c5abc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3edffa),
	.w1(32'hbb0829f4),
	.w2(32'h3bafdc17),
	.w3(32'hbbd3910a),
	.w4(32'hbc2be1de),
	.w5(32'hbb49994f),
	.w6(32'hbb0e8d47),
	.w7(32'hbbfb03d8),
	.w8(32'hbbcd99bd),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b7c12),
	.w1(32'hbac3387f),
	.w2(32'hbb2fc32c),
	.w3(32'hbb9e572c),
	.w4(32'hbc037319),
	.w5(32'hbc010275),
	.w6(32'hbb8343bd),
	.w7(32'hbbf25d7c),
	.w8(32'hbc1b8d73),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19d079),
	.w1(32'h3b43814c),
	.w2(32'hbc8f2af7),
	.w3(32'hbbf12755),
	.w4(32'hb9da1fe6),
	.w5(32'h3aca4cc0),
	.w6(32'hbbf7551e),
	.w7(32'hbb57a5cc),
	.w8(32'h3af36d23),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc928989),
	.w1(32'hbaf14162),
	.w2(32'h3c5d7f01),
	.w3(32'hbadc70a1),
	.w4(32'h3b948998),
	.w5(32'h3c9ac276),
	.w6(32'h3be272b5),
	.w7(32'h3b9362a5),
	.w8(32'hbbb1f51a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf05b85),
	.w1(32'hbbc2cfeb),
	.w2(32'hbc235088),
	.w3(32'h3c7bc468),
	.w4(32'h3846289a),
	.w5(32'hbc5f7eee),
	.w6(32'hbb951d25),
	.w7(32'hbac052a4),
	.w8(32'h396ca1bc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc308b4b),
	.w1(32'hbb84c54d),
	.w2(32'h3b7e75fe),
	.w3(32'hbc1400a6),
	.w4(32'hbb86550c),
	.w5(32'hb994ffaf),
	.w6(32'hb9f17e38),
	.w7(32'hbbc3fed2),
	.w8(32'h3b9180cc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a675b2e),
	.w1(32'h3aee95b8),
	.w2(32'h3c008000),
	.w3(32'hbb8d67c1),
	.w4(32'hb85ed704),
	.w5(32'h3c231dff),
	.w6(32'h3b88d3eb),
	.w7(32'h3be886ea),
	.w8(32'h3bbb8bfd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5fde2),
	.w1(32'h3b7de806),
	.w2(32'hbb238033),
	.w3(32'h3bd8efb9),
	.w4(32'h3ac38077),
	.w5(32'hbbef15c7),
	.w6(32'h3b4e5ecd),
	.w7(32'h3ba83443),
	.w8(32'hbbbe3660),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba31fee),
	.w1(32'hbb96faac),
	.w2(32'hbb34c0ca),
	.w3(32'hbc24681c),
	.w4(32'hbbd6ce84),
	.w5(32'hbc14df2b),
	.w6(32'hbbe12d65),
	.w7(32'hbb923b6a),
	.w8(32'hba56ddb7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1fcee),
	.w1(32'hbb7092e4),
	.w2(32'h3cbe417f),
	.w3(32'hbafddf68),
	.w4(32'hbac73348),
	.w5(32'hbbd39067),
	.w6(32'h3b9a7822),
	.w7(32'h3b34ea1e),
	.w8(32'hbb9caca0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca61ace),
	.w1(32'h39ecfe8b),
	.w2(32'hbc2bf4f0),
	.w3(32'hbccf60b4),
	.w4(32'hbc9a9797),
	.w5(32'hbbb7cc23),
	.w6(32'hbbc9a18b),
	.w7(32'hbc0850b2),
	.w8(32'h3c0758e9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d88f1),
	.w1(32'hbbc0c0b5),
	.w2(32'h3ab0e80e),
	.w3(32'hbae9f2ce),
	.w4(32'h3ad3b63c),
	.w5(32'hbb600ef4),
	.w6(32'h3c61f3ab),
	.w7(32'h3c36f4df),
	.w8(32'h3ad51b26),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd3f1),
	.w1(32'hbae8dc9d),
	.w2(32'h3ca0d712),
	.w3(32'hbbc69bd7),
	.w4(32'hbac24962),
	.w5(32'h3c66c636),
	.w6(32'h3b62fd2c),
	.w7(32'h3beb6c61),
	.w8(32'hbb163c02),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1074e),
	.w1(32'h3cc1ea79),
	.w2(32'hbbebb7cf),
	.w3(32'h3c1f834d),
	.w4(32'h3c2d2d68),
	.w5(32'hbbd30aba),
	.w6(32'hbc5a11af),
	.w7(32'hbc83e8cc),
	.w8(32'hbb996c10),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b81d8),
	.w1(32'h3a0370f8),
	.w2(32'h3bc709f2),
	.w3(32'h39b78800),
	.w4(32'h3b1ddd8a),
	.w5(32'h39bce530),
	.w6(32'h3be5560d),
	.w7(32'h3a0c1b9a),
	.w8(32'hbaf6f491),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9c8b6),
	.w1(32'hbbad99b1),
	.w2(32'h3c57a54d),
	.w3(32'h3bc94c57),
	.w4(32'h3a4577b2),
	.w5(32'h3c39965d),
	.w6(32'hbc1a1400),
	.w7(32'hbb829512),
	.w8(32'h3ac3a46e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e2a2e),
	.w1(32'h3ac570a6),
	.w2(32'hbb02b617),
	.w3(32'h3a0e2208),
	.w4(32'hbc2925f7),
	.w5(32'hbb7cc341),
	.w6(32'hbc24e163),
	.w7(32'hbc457be9),
	.w8(32'h3bac09dd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1833c),
	.w1(32'hbb10dc18),
	.w2(32'hbc3ca2df),
	.w3(32'hb900710d),
	.w4(32'hba737f9d),
	.w5(32'hba7f1808),
	.w6(32'h3c10d566),
	.w7(32'h3c99529f),
	.w8(32'h3b1d00e6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68571),
	.w1(32'hbbcef7b0),
	.w2(32'hbaf61da7),
	.w3(32'hbb72dc62),
	.w4(32'hbc1366db),
	.w5(32'hbbd85405),
	.w6(32'hbbc8fba2),
	.w7(32'hbbc6b0a6),
	.w8(32'hbb2ed333),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2c325),
	.w1(32'hbb150384),
	.w2(32'hbbb8e5f5),
	.w3(32'hbc48a017),
	.w4(32'hbb6a7fc4),
	.w5(32'hbba9388c),
	.w6(32'hbb5d12d2),
	.w7(32'h3b36ae71),
	.w8(32'hbb7571c7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb845fee),
	.w1(32'h3964fd9c),
	.w2(32'h3c7ac876),
	.w3(32'hb9beab8a),
	.w4(32'hbb51f044),
	.w5(32'h3be6b21c),
	.w6(32'h3bc382fe),
	.w7(32'hbbd2288e),
	.w8(32'h3bcf6cf1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5df0bd),
	.w1(32'h3adeed0f),
	.w2(32'hba71af27),
	.w3(32'h3c04b5e0),
	.w4(32'h3bb8f6f0),
	.w5(32'h3b858378),
	.w6(32'hbb29968c),
	.w7(32'hbbc03f22),
	.w8(32'hbb52d3fc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baac3d3),
	.w1(32'h3b576724),
	.w2(32'h3b2afd04),
	.w3(32'hbab65b07),
	.w4(32'hbca05de7),
	.w5(32'h3b84ba2b),
	.w6(32'hbc4d0133),
	.w7(32'hbc1fc99e),
	.w8(32'h3ad1b753),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dd1a2),
	.w1(32'h3a93a4e1),
	.w2(32'hbc8e243e),
	.w3(32'h3bd4e60d),
	.w4(32'h3b1b71e9),
	.w5(32'hbc244a97),
	.w6(32'h39aebcef),
	.w7(32'h394a0be8),
	.w8(32'hbc4ab158),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc897957),
	.w1(32'hbb412be5),
	.w2(32'h3bfe508e),
	.w3(32'h38380039),
	.w4(32'h3c35d153),
	.w5(32'h3c677458),
	.w6(32'hbc1438b3),
	.w7(32'h3b864476),
	.w8(32'h3b7bb46c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157030),
	.w1(32'h389f772d),
	.w2(32'hbb8bfe3a),
	.w3(32'hba832299),
	.w4(32'hbb4e66e9),
	.w5(32'hbbb1c393),
	.w6(32'h3aed3aca),
	.w7(32'hbba68676),
	.w8(32'h38b432df),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea6fcd),
	.w1(32'hbbc1f193),
	.w2(32'hbcb2b1e8),
	.w3(32'hbaa2d3e8),
	.w4(32'hbb93c23d),
	.w5(32'hbd1a13e0),
	.w6(32'h3b5c815a),
	.w7(32'h39f91b71),
	.w8(32'hbcb1efc2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd204a41),
	.w1(32'hbcde2394),
	.w2(32'hbc280048),
	.w3(32'hbd6da7d3),
	.w4(32'hbd3f8e4a),
	.w5(32'hbc95c13c),
	.w6(32'hbd271407),
	.w7(32'hbd0862b0),
	.w8(32'hbbf8f782),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0dcd),
	.w1(32'hbb975ca8),
	.w2(32'hbb54d040),
	.w3(32'hbca6de10),
	.w4(32'hbc85fcbe),
	.w5(32'hbbeaea7f),
	.w6(32'hbca7aa43),
	.w7(32'hbbd90f40),
	.w8(32'h396a5833),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44bb6d),
	.w1(32'hbbef608a),
	.w2(32'hba71be4d),
	.w3(32'hbc0866c2),
	.w4(32'hbc4da779),
	.w5(32'hbb14a222),
	.w6(32'h3a9ff33a),
	.w7(32'hbbcc0d61),
	.w8(32'h3b65efa5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8630ee),
	.w1(32'hbb90cf11),
	.w2(32'hbbd6d6e9),
	.w3(32'hbb0e8104),
	.w4(32'hbb1643a0),
	.w5(32'hbb9ea680),
	.w6(32'hba2a9d61),
	.w7(32'h3bb68f35),
	.w8(32'hbb96bb76),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf228c),
	.w1(32'hb81702fa),
	.w2(32'hbce88543),
	.w3(32'h3afd2535),
	.w4(32'h3b0e0b88),
	.w5(32'hbcdd55d4),
	.w6(32'h3908eefb),
	.w7(32'h36e14202),
	.w8(32'hbc782e53),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d816),
	.w1(32'hba35cfb3),
	.w2(32'hbc198b31),
	.w3(32'hbc4d7bb2),
	.w4(32'h3c0ac8d4),
	.w5(32'hbc06d951),
	.w6(32'hbb7ba77c),
	.w7(32'h3bd5b05c),
	.w8(32'hbb496185),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af27ac8),
	.w1(32'hbb36454b),
	.w2(32'h37698253),
	.w3(32'h3c5b4fe4),
	.w4(32'h3bbbd5a4),
	.w5(32'h3c044a21),
	.w6(32'h3ca291ce),
	.w7(32'h3c3ee209),
	.w8(32'h3bf58a34),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9c50),
	.w1(32'hbb01c360),
	.w2(32'hbb24d32d),
	.w3(32'h389b09e5),
	.w4(32'hbb847694),
	.w5(32'hbbc47fb0),
	.w6(32'h3cb4d10a),
	.w7(32'h3b91a06d),
	.w8(32'hb9cfd2aa),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44e918),
	.w1(32'h3a29796c),
	.w2(32'hbb61c755),
	.w3(32'h3bf67360),
	.w4(32'h3c7b3f5e),
	.w5(32'hbadd45bb),
	.w6(32'h3b9630c4),
	.w7(32'h3c14d185),
	.w8(32'h39c615aa),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fa9f9),
	.w1(32'h3b6b89cd),
	.w2(32'h3bd25b28),
	.w3(32'h3c2396be),
	.w4(32'h3bda1eae),
	.w5(32'h3c503a59),
	.w6(32'h3c98559b),
	.w7(32'h3c4c1863),
	.w8(32'h3c2f375b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd4c3c),
	.w1(32'h3b305a3e),
	.w2(32'hbd158188),
	.w3(32'h3cabbc30),
	.w4(32'h3c500954),
	.w5(32'hbd0f35bd),
	.w6(32'h3cacb8b7),
	.w7(32'h3c49afea),
	.w8(32'hbcab9338),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd475bec),
	.w1(32'hbcca245a),
	.w2(32'hba973120),
	.w3(32'hbd738f4e),
	.w4(32'hbd1df783),
	.w5(32'h3b1e867f),
	.w6(32'hbd2760c1),
	.w7(32'hbd09093c),
	.w8(32'h39ea4f5c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4dac1),
	.w1(32'h3c0f2ec6),
	.w2(32'h3bbe4528),
	.w3(32'h3c59c9aa),
	.w4(32'h3c78e5e4),
	.w5(32'h3c6b9e7a),
	.w6(32'h3c2ee633),
	.w7(32'h3c3b9fc1),
	.w8(32'h3c137b3b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac55efa),
	.w1(32'hbbbea42b),
	.w2(32'hbc69d03d),
	.w3(32'h3c23bf5b),
	.w4(32'hbc434c31),
	.w5(32'hbc3fe343),
	.w6(32'h3c4e9bb7),
	.w7(32'hbc123355),
	.w8(32'hbb757604),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdd37),
	.w1(32'h3b5854db),
	.w2(32'h3c32a3e2),
	.w3(32'hbb1222fc),
	.w4(32'h3aff2ada),
	.w5(32'h3bf8323e),
	.w6(32'hbb5b2400),
	.w7(32'hb9bd56f6),
	.w8(32'hbb3465b7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc99e56),
	.w1(32'hba9ffd21),
	.w2(32'hbadb73dd),
	.w3(32'h3ce3854f),
	.w4(32'h3c87f5b0),
	.w5(32'hbbc908ac),
	.w6(32'h3c940d00),
	.w7(32'h3c901f61),
	.w8(32'hbc1fd8cb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11afd9),
	.w1(32'h3ba23161),
	.w2(32'hbbd94795),
	.w3(32'h3c65864d),
	.w4(32'h3baf56e9),
	.w5(32'hbb1395c6),
	.w6(32'h3c262bb4),
	.w7(32'hbb3f40cc),
	.w8(32'hbb4dd4c2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa16b19),
	.w1(32'h3adb1eb5),
	.w2(32'hbc0918ae),
	.w3(32'h3bc44f7a),
	.w4(32'h3c081053),
	.w5(32'hba894833),
	.w6(32'h3b0614a6),
	.w7(32'h3bf2cbce),
	.w8(32'hbb197c6e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ed5e6),
	.w1(32'hbaa36dc3),
	.w2(32'hbbfa6c3a),
	.w3(32'hbc457264),
	.w4(32'hbaf1e521),
	.w5(32'hbb0b8409),
	.w6(32'hbbba8521),
	.w7(32'hbbfec802),
	.w8(32'h3b9b15ce),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8829b),
	.w1(32'hba5b919a),
	.w2(32'hba0c43f1),
	.w3(32'hbc0e5cd7),
	.w4(32'hbb863a24),
	.w5(32'h3b4854df),
	.w6(32'hbae7cb05),
	.w7(32'hbb05576a),
	.w8(32'hba8ce612),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d8b0c),
	.w1(32'hbb1f4b04),
	.w2(32'hbb4e5b9c),
	.w3(32'hbb571cc7),
	.w4(32'hbc0d83fe),
	.w5(32'hba9d228d),
	.w6(32'hbabaf277),
	.w7(32'hbb87d250),
	.w8(32'h3b7a9fb4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc539b5a),
	.w1(32'h3b0c82ef),
	.w2(32'h3b91598c),
	.w3(32'hbc554bc2),
	.w4(32'h3b7cdc4c),
	.w5(32'h3c4ad2bf),
	.w6(32'hbb63ff5a),
	.w7(32'h3bcf02bb),
	.w8(32'h3b561fb3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3215db),
	.w1(32'hbb2d3d42),
	.w2(32'h3c30cad3),
	.w3(32'h3b9a3d46),
	.w4(32'h3c197dd0),
	.w5(32'h3c512066),
	.w6(32'h3b1c5eb3),
	.w7(32'h3b77c657),
	.w8(32'h3c0fa9a4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59fe99),
	.w1(32'hba0b8efd),
	.w2(32'hbb8afd17),
	.w3(32'hbaa5892a),
	.w4(32'h39a05967),
	.w5(32'h3b1ac354),
	.w6(32'h3c10c675),
	.w7(32'hbac00672),
	.w8(32'h3b9eb62a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fbc5e),
	.w1(32'h3b6795e6),
	.w2(32'hba86459a),
	.w3(32'h3bbc1171),
	.w4(32'h3bce1bac),
	.w5(32'hba9c1893),
	.w6(32'hbc4e64fe),
	.w7(32'h39d4f6ec),
	.w8(32'hbc017c2e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6117de),
	.w1(32'h3b4b04be),
	.w2(32'hbbc87918),
	.w3(32'hb90e1afc),
	.w4(32'hbab61606),
	.w5(32'hbc0c0fbe),
	.w6(32'hbaa74015),
	.w7(32'hbbf474f4),
	.w8(32'hba0d9ba7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba1cc),
	.w1(32'h3aad2361),
	.w2(32'hba1b2652),
	.w3(32'h3c4d4d04),
	.w4(32'h3bc11664),
	.w5(32'hbae1b2f2),
	.w6(32'h3c5a3738),
	.w7(32'h3c3ce71f),
	.w8(32'h3b93b39e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b18b4),
	.w1(32'h3c52e6a0),
	.w2(32'hbbd33262),
	.w3(32'h3bab8e95),
	.w4(32'h3c87fafc),
	.w5(32'hbbd629e3),
	.w6(32'h3c818bef),
	.w7(32'h3cf94422),
	.w8(32'hbbc0d1c2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3202e),
	.w1(32'hbbaba484),
	.w2(32'hbcb18ec2),
	.w3(32'hbc5d8684),
	.w4(32'hbb8ea696),
	.w5(32'hbcb26fef),
	.w6(32'hbb949746),
	.w7(32'hbb7018ef),
	.w8(32'hbca2a3c6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33185c),
	.w1(32'hbb84862b),
	.w2(32'h3b2944ae),
	.w3(32'hbc2c4b02),
	.w4(32'hbaeb1c4b),
	.w5(32'h3a9eb854),
	.w6(32'hbc29ecde),
	.w7(32'hbb66daf3),
	.w8(32'h37f1d16b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9a471),
	.w1(32'hbaf6f098),
	.w2(32'h3b977b3f),
	.w3(32'h3ace6268),
	.w4(32'hbb5455a9),
	.w5(32'h3bbab2fd),
	.w6(32'h3c094758),
	.w7(32'hbb39c866),
	.w8(32'hbb0ab158),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27da2),
	.w1(32'h3c1e384d),
	.w2(32'hbb79e250),
	.w3(32'hbbb480c5),
	.w4(32'h3be32a98),
	.w5(32'hbab7c1c4),
	.w6(32'h3be9c138),
	.w7(32'h3b86b690),
	.w8(32'h3b1ab326),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e32bd),
	.w1(32'hbb2eba39),
	.w2(32'hbb7b2497),
	.w3(32'h3b5f8a98),
	.w4(32'h3c08029d),
	.w5(32'hbcc2f4f2),
	.w6(32'h3ba193eb),
	.w7(32'h3bbd3dca),
	.w8(32'hbc8c76b4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8231),
	.w1(32'hbbd4c3b7),
	.w2(32'hbad074ca),
	.w3(32'hbd157eb9),
	.w4(32'hbcc0d271),
	.w5(32'hbaebbdf9),
	.w6(32'hbcfbf12d),
	.w7(32'hbc7b1764),
	.w8(32'hbb322034),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db7173),
	.w1(32'hbb5dd86f),
	.w2(32'hbc1cf936),
	.w3(32'h3b554de8),
	.w4(32'hba58c956),
	.w5(32'hbc3af11b),
	.w6(32'h3ad7a8fd),
	.w7(32'hbaaac60a),
	.w8(32'hbc03650c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0d74d),
	.w1(32'hbb9cdc9c),
	.w2(32'h3b92b215),
	.w3(32'h3a6aa9dc),
	.w4(32'hba60791a),
	.w5(32'h3c4aa2a3),
	.w6(32'h3ad390c1),
	.w7(32'h39ef0cbb),
	.w8(32'h3c8f882b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9de64c),
	.w1(32'h3cc091ed),
	.w2(32'h3b910972),
	.w3(32'h3d1c4bdd),
	.w4(32'h3cd24eaf),
	.w5(32'hbb1bff5e),
	.w6(32'h3cc179b2),
	.w7(32'h3c5d918f),
	.w8(32'h3bc9347f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96efe6),
	.w1(32'h3bc060a1),
	.w2(32'h39c91366),
	.w3(32'hbbfa8fab),
	.w4(32'h3963c021),
	.w5(32'h3bddff1d),
	.w6(32'h3a75a905),
	.w7(32'hba0260b8),
	.w8(32'h3bced587),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960010),
	.w1(32'hbaa3c801),
	.w2(32'hbbef0d2b),
	.w3(32'h3c387ca0),
	.w4(32'h3bcd6d4e),
	.w5(32'hbb8d5b92),
	.w6(32'h3c40265c),
	.w7(32'h3bf6ec3e),
	.w8(32'hbbfda0ed),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2863d8),
	.w1(32'h3afebb18),
	.w2(32'h3c2234c2),
	.w3(32'h3c0d384d),
	.w4(32'h3c0fd7e2),
	.w5(32'h3c53cf81),
	.w6(32'h3c315e80),
	.w7(32'h3c254c41),
	.w8(32'h3c272aad),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081fc0),
	.w1(32'hba34fed4),
	.w2(32'h3c9cb216),
	.w3(32'h3c655b89),
	.w4(32'h3b885899),
	.w5(32'h3c92c35b),
	.w6(32'h3c0cca0c),
	.w7(32'h3ba53eb0),
	.w8(32'h3c0f99d2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0324f8),
	.w1(32'h3ca516a7),
	.w2(32'h3aa593fa),
	.w3(32'h3d69f3f8),
	.w4(32'h3d0ddfac),
	.w5(32'hbb37fe40),
	.w6(32'h3ceaf2bd),
	.w7(32'h3cff3ddf),
	.w8(32'h3b021fc2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45c941),
	.w1(32'h3c4fce27),
	.w2(32'hbc4dc130),
	.w3(32'hbcaceac9),
	.w4(32'hbad60349),
	.w5(32'hbc058f30),
	.w6(32'h3b998c0c),
	.w7(32'h3c05cf9d),
	.w8(32'hbc0df3ed),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3d54f),
	.w1(32'hbbace50a),
	.w2(32'hbc4136d4),
	.w3(32'h3b9fc06d),
	.w4(32'h3a0ed638),
	.w5(32'hbbe04b64),
	.w6(32'h3b857bbc),
	.w7(32'hba449d48),
	.w8(32'hbc06c9bc),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba02752),
	.w1(32'h3b4e1c57),
	.w2(32'h3a7a53e2),
	.w3(32'hbb885e2e),
	.w4(32'h3b74e938),
	.w5(32'hbc1cba68),
	.w6(32'hba461dcf),
	.w7(32'h3ad95c30),
	.w8(32'hbc82ba13),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb82a76),
	.w1(32'hbc727ce3),
	.w2(32'hbc8a4455),
	.w3(32'hbd23e2e5),
	.w4(32'hbca16007),
	.w5(32'hbce6644f),
	.w6(32'hbc8f7ab1),
	.w7(32'hbc0894de),
	.w8(32'hbccf7a93),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cea63),
	.w1(32'hbd052be6),
	.w2(32'h3bc291c3),
	.w3(32'hbd61c5f8),
	.w4(32'hbd1c4404),
	.w5(32'h3ba970c6),
	.w6(32'hbd1b011e),
	.w7(32'hbc7f71fc),
	.w8(32'h3b3e5c76),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf545f0),
	.w1(32'h3bada686),
	.w2(32'h3b216db4),
	.w3(32'h3c2cdb3e),
	.w4(32'h3bdd9a98),
	.w5(32'h3c489708),
	.w6(32'h3c3703dc),
	.w7(32'hbb48e0ce),
	.w8(32'h3a51928c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ec080),
	.w1(32'hbac808a0),
	.w2(32'hbb451cda),
	.w3(32'h3ca9e34d),
	.w4(32'h3bc12b91),
	.w5(32'hbb4ffa00),
	.w6(32'h3b43729a),
	.w7(32'hbb4dd893),
	.w8(32'hbbddb314),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07bbed),
	.w1(32'h382af9a2),
	.w2(32'hbb538a3b),
	.w3(32'h3c2ba722),
	.w4(32'h3bbaacd3),
	.w5(32'hbb94e8b1),
	.w6(32'h3b9f25c5),
	.w7(32'h3abdcdfa),
	.w8(32'hbb753c30),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa06abb),
	.w1(32'hbada40dc),
	.w2(32'h3be4a241),
	.w3(32'h3b7e3586),
	.w4(32'h39eb4dbb),
	.w5(32'h3b8ba6f4),
	.w6(32'h3b93f741),
	.w7(32'hbb069b8e),
	.w8(32'h3c0603ab),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90b57c),
	.w1(32'h3c3365de),
	.w2(32'h3c2dd05c),
	.w3(32'h3c7fa488),
	.w4(32'h3cb69125),
	.w5(32'h3c307972),
	.w6(32'h3c93a158),
	.w7(32'h3c77b322),
	.w8(32'hbb3fe605),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c0a0a),
	.w1(32'h3bab7890),
	.w2(32'h3c85b961),
	.w3(32'h3c804da1),
	.w4(32'h3c16e89d),
	.w5(32'h3ca050ee),
	.w6(32'h3bc4ea7e),
	.w7(32'h3c053943),
	.w8(32'h3c286a09),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2cc47),
	.w1(32'h3b99e49e),
	.w2(32'h3b863a8c),
	.w3(32'h3d0498dd),
	.w4(32'h3c98dcf0),
	.w5(32'h3bb8838b),
	.w6(32'h3cc6ab5e),
	.w7(32'h3c905aa8),
	.w8(32'hbac50fbf),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be59655),
	.w1(32'h3b3f0656),
	.w2(32'hbc6d3278),
	.w3(32'h3bc8b804),
	.w4(32'h3c3d3d29),
	.w5(32'hbc7bcf50),
	.w6(32'h3ba95808),
	.w7(32'h3c03875a),
	.w8(32'hbc26745f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43118c),
	.w1(32'hbb42716e),
	.w2(32'h3aae005d),
	.w3(32'hba10858e),
	.w4(32'hbae6e167),
	.w5(32'h3b3cda33),
	.w6(32'hb8391007),
	.w7(32'hba11ca2a),
	.w8(32'h3b65ee6c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b458133),
	.w1(32'h3a2a5a7e),
	.w2(32'hbc0abb9e),
	.w3(32'h3a830a3f),
	.w4(32'h3b0bbcdf),
	.w5(32'hbbe36e7a),
	.w6(32'h3b81b98b),
	.w7(32'h3b6f1a43),
	.w8(32'hbb8aab1c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dedab),
	.w1(32'hbaa4c3d6),
	.w2(32'h3b24f38d),
	.w3(32'hbc7da240),
	.w4(32'h3b6d82b9),
	.w5(32'h3bb6f3c3),
	.w6(32'hb8a75ff4),
	.w7(32'h3a9d758e),
	.w8(32'h3bad87f1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c327b34),
	.w1(32'h3bac6b2e),
	.w2(32'hbb079008),
	.w3(32'h3cc590c7),
	.w4(32'h3c519fd9),
	.w5(32'hbc2f133b),
	.w6(32'h3c6c1231),
	.w7(32'h3c88837a),
	.w8(32'hbc3f2d80),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd015ac),
	.w1(32'h3c1408f4),
	.w2(32'hbcd3de4c),
	.w3(32'hbb06fae1),
	.w4(32'h3bb11786),
	.w5(32'hbcf7bea3),
	.w6(32'hbb370745),
	.w7(32'h3bf7ccb4),
	.w8(32'hbcd7e057),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb497f5),
	.w1(32'hbc5c3c6e),
	.w2(32'h3c563b97),
	.w3(32'hbc629552),
	.w4(32'hbc0efde5),
	.w5(32'h3c9239e9),
	.w6(32'hbc1ae95e),
	.w7(32'hba0aeebe),
	.w8(32'h3c8cd5e8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c8ee4),
	.w1(32'h3bdff3a3),
	.w2(32'hbb5af5b7),
	.w3(32'h3c8ad16c),
	.w4(32'h3c4069b9),
	.w5(32'hbad81c40),
	.w6(32'h3c886d78),
	.w7(32'h3c5e59fe),
	.w8(32'hbb0afcc7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8ac41),
	.w1(32'h3a7ba4a8),
	.w2(32'h3b44ed88),
	.w3(32'h3bd2ec20),
	.w4(32'h3bcc97a8),
	.w5(32'h3b408367),
	.w6(32'h3bc9918e),
	.w7(32'h3bc0277d),
	.w8(32'hb99dba29),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986f107),
	.w1(32'h3b882227),
	.w2(32'h3b2fa265),
	.w3(32'hbc051ad6),
	.w4(32'h3b9665b6),
	.w5(32'h3c4ce94d),
	.w6(32'h3b6e2de0),
	.w7(32'h3bdd2cdf),
	.w8(32'h3b8d2938),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb798c00),
	.w1(32'h3be8f235),
	.w2(32'h3b51fc70),
	.w3(32'h3be08026),
	.w4(32'h3c09ab7f),
	.w5(32'h3c3a0274),
	.w6(32'h3b0404dd),
	.w7(32'h3bda9b58),
	.w8(32'h3c024483),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23d198),
	.w1(32'h3c2124ac),
	.w2(32'hbc1fc350),
	.w3(32'h3c5d1285),
	.w4(32'h3c1bc16f),
	.w5(32'hbc76a4c3),
	.w6(32'h3c4446e4),
	.w7(32'h3bd24be6),
	.w8(32'hbbd90e2d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc559ebb),
	.w1(32'hba46daae),
	.w2(32'hbc86f24f),
	.w3(32'hbcce89c0),
	.w4(32'hbc4fd21c),
	.w5(32'hbc4ba7a5),
	.w6(32'hbc0f3bfe),
	.w7(32'hbb1799da),
	.w8(32'hbc3339b0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcded825),
	.w1(32'hbca532b3),
	.w2(32'hbae52647),
	.w3(32'hbd076f20),
	.w4(32'hbcb64d09),
	.w5(32'h3bc241d3),
	.w6(32'hbce32120),
	.w7(32'hbc9d13a5),
	.w8(32'hbb79e620),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9dfb0),
	.w1(32'hbbb312c5),
	.w2(32'hbceb999a),
	.w3(32'h3c42ac84),
	.w4(32'h3b5bdd49),
	.w5(32'hbd456f88),
	.w6(32'h3b6bb1c5),
	.w7(32'hbad4779a),
	.w8(32'hbcb047ba),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd28eb76),
	.w1(32'hbc9ce55b),
	.w2(32'hbca90e63),
	.w3(32'hbd87e801),
	.w4(32'hbd4648c9),
	.w5(32'hbd16c1e5),
	.w6(32'hbd16fa98),
	.w7(32'hbcc80082),
	.w8(32'hbcde7c01),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd163b08),
	.w1(32'hbcb2135e),
	.w2(32'hbb7e0013),
	.w3(32'hbd71c88c),
	.w4(32'hbd35255b),
	.w5(32'hbb402dac),
	.w6(32'hbd568a48),
	.w7(32'hbcf50757),
	.w8(32'h391f6c3a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb516251),
	.w1(32'hbba1a876),
	.w2(32'h3bc2b83c),
	.w3(32'h3b789687),
	.w4(32'hbb0ff6a5),
	.w5(32'h3b41b064),
	.w6(32'hbaf6da6c),
	.w7(32'hbb40f181),
	.w8(32'h3a26a4bd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d94e),
	.w1(32'hbbc462f1),
	.w2(32'h3cc60921),
	.w3(32'hbacbaa68),
	.w4(32'hbbffed67),
	.w5(32'h3c967d42),
	.w6(32'h3b438fc5),
	.w7(32'hbbcfbe20),
	.w8(32'h3c1c469f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfd7cf),
	.w1(32'h3c8563d7),
	.w2(32'h3a74f774),
	.w3(32'h3d0420bd),
	.w4(32'h3ca14561),
	.w5(32'h3b178674),
	.w6(32'h3ca77f7f),
	.w7(32'h3bf9d546),
	.w8(32'hba86b369),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57858b),
	.w1(32'hbb82b541),
	.w2(32'h3b934a05),
	.w3(32'h3b46da83),
	.w4(32'hba85b3d3),
	.w5(32'h3b826fcc),
	.w6(32'hba998a88),
	.w7(32'h3a9408b9),
	.w8(32'h3b263c91),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ceb53),
	.w1(32'h3bcd8736),
	.w2(32'hbc1b9ca6),
	.w3(32'h3ca5a60d),
	.w4(32'h3c12122f),
	.w5(32'h3af0802d),
	.w6(32'h3c453adc),
	.w7(32'h3b6d0ef2),
	.w8(32'hbb6d6b89),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1202),
	.w1(32'hbc49e169),
	.w2(32'h3c264efd),
	.w3(32'h3a48a50d),
	.w4(32'hbba1d50a),
	.w5(32'h3bd18aff),
	.w6(32'hbba5389b),
	.w7(32'hbc156489),
	.w8(32'h3b8c92a9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8344c1),
	.w1(32'h3ba07502),
	.w2(32'hbcce7a74),
	.w3(32'h3c85d8bd),
	.w4(32'h3c27010f),
	.w5(32'hbcdffc30),
	.w6(32'h3c548e84),
	.w7(32'h3bd28f12),
	.w8(32'hbc8c57ef),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06f2db),
	.w1(32'hbc9ed143),
	.w2(32'hbc812d34),
	.w3(32'hbd3a12f2),
	.w4(32'hbcf0f652),
	.w5(32'hbc7f6512),
	.w6(32'hbce8f619),
	.w7(32'hbc9b033b),
	.w8(32'hbb3b8afc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87624c),
	.w1(32'h3a8765a1),
	.w2(32'h3c0ae46e),
	.w3(32'hbd034c16),
	.w4(32'hbc3d7490),
	.w5(32'h3b7c4cb0),
	.w6(32'hbc30ad18),
	.w7(32'hbc3124b0),
	.w8(32'hba3a02cb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f458f),
	.w1(32'h3b487d2c),
	.w2(32'hbb8baac5),
	.w3(32'h3cb16118),
	.w4(32'h3c17d139),
	.w5(32'h3b831f2b),
	.w6(32'h3bd2040f),
	.w7(32'h39e604a3),
	.w8(32'hb98e9355),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e6eaf),
	.w1(32'h3bd33926),
	.w2(32'hbcd306bc),
	.w3(32'hba6dc025),
	.w4(32'h3bc9497a),
	.w5(32'hbd083fa0),
	.w6(32'h37d51a0f),
	.w7(32'h3bdb7b8a),
	.w8(32'hbc839770),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfd4046),
	.w1(32'hbc9ef8b9),
	.w2(32'h3c0a4eab),
	.w3(32'hbd3393d4),
	.w4(32'hbcd02f52),
	.w5(32'h3bf7cb7b),
	.w6(32'hbd13bf22),
	.w7(32'hbcfda5b1),
	.w8(32'h3be63e5c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3782c),
	.w1(32'h3bd7f33f),
	.w2(32'hbaccbdf7),
	.w3(32'hbae9fca7),
	.w4(32'hbc126325),
	.w5(32'h3b5fa4b4),
	.w6(32'hbb3ba61f),
	.w7(32'hbbee2f38),
	.w8(32'h3b9ae779),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb469c0a),
	.w1(32'h3ad284f2),
	.w2(32'hbc1e9d58),
	.w3(32'h3b0725b4),
	.w4(32'h3bbc8e7a),
	.w5(32'hbbdae3c4),
	.w6(32'h3b325fe8),
	.w7(32'h3b14ddf8),
	.w8(32'hbc107bec),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c33e9),
	.w1(32'hbba88fa6),
	.w2(32'h3aae14ba),
	.w3(32'h3b4b6acd),
	.w4(32'h3baa23fa),
	.w5(32'hb9ca1f40),
	.w6(32'hb95b92cd),
	.w7(32'h3bb041dc),
	.w8(32'h3b4434ce),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0242),
	.w1(32'hbacc7563),
	.w2(32'hbcb3f567),
	.w3(32'h3a87add7),
	.w4(32'h3acfcea2),
	.w5(32'hbd182f46),
	.w6(32'h3ab80423),
	.w7(32'hba1c9341),
	.w8(32'hbcc0a80b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd194896),
	.w1(32'hbcf2c790),
	.w2(32'hbcab7414),
	.w3(32'hbd55ed7e),
	.w4(32'hbd25216e),
	.w5(32'hbd1e78c9),
	.w6(32'hbd0a8a77),
	.w7(32'hbca5c0c9),
	.w8(32'hbcacf1f4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf6c2e0),
	.w1(32'hbc61b2c2),
	.w2(32'h3bdf7bf9),
	.w3(32'hbd66397c),
	.w4(32'hbd1f422c),
	.w5(32'h3b5837d5),
	.w6(32'hbd2d17d4),
	.w7(32'hbcf61386),
	.w8(32'h3b27255a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53a216),
	.w1(32'h3c499810),
	.w2(32'hbb1d66ae),
	.w3(32'hbb59f3ba),
	.w4(32'h3c06302d),
	.w5(32'hbaccf2ca),
	.w6(32'h3b15318e),
	.w7(32'h3be865ea),
	.w8(32'h3acce6c7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55d377),
	.w1(32'hbafa8b9f),
	.w2(32'h3a857ae1),
	.w3(32'hbb38acea),
	.w4(32'hbb0a3afe),
	.w5(32'h3b2d6b9d),
	.w6(32'h3a4bc957),
	.w7(32'h3b1dfc59),
	.w8(32'h3b8a18cd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba862f0),
	.w1(32'h3bebb94e),
	.w2(32'h3a48d851),
	.w3(32'h3baf961b),
	.w4(32'h3bd80fc4),
	.w5(32'h3ba9135c),
	.w6(32'h3bbee3c5),
	.w7(32'h3c1697a1),
	.w8(32'hbaa6778b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc0b4f),
	.w1(32'hba0e12c7),
	.w2(32'hbbd7d89a),
	.w3(32'h3c522c60),
	.w4(32'h3c98318b),
	.w5(32'hbb3ebc40),
	.w6(32'h3c5d65c7),
	.w7(32'h3b8bdf5f),
	.w8(32'hbb95d0bb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293969),
	.w1(32'hbbac88c1),
	.w2(32'hbaf4bbc0),
	.w3(32'h3b4ecb92),
	.w4(32'hbafd9967),
	.w5(32'hbb2c854f),
	.w6(32'hbb353a51),
	.w7(32'hbbc298ad),
	.w8(32'h3b80b363),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f047e),
	.w1(32'hba675289),
	.w2(32'h3c6587d4),
	.w3(32'h3bddf389),
	.w4(32'h3c178826),
	.w5(32'h3c8b578a),
	.w6(32'h3a4a8616),
	.w7(32'h3c19bb29),
	.w8(32'h3c776753),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce85021),
	.w1(32'h3ccd091e),
	.w2(32'h3c9f6202),
	.w3(32'h3d39b44f),
	.w4(32'h3d030d68),
	.w5(32'h3ce4eab6),
	.w6(32'h3d014039),
	.w7(32'h3ca7d685),
	.w8(32'h3ce674dd),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe9214),
	.w1(32'h3c681432),
	.w2(32'h3c66d089),
	.w3(32'h3d5b3ee0),
	.w4(32'h3cdf8c97),
	.w5(32'h3c644eb9),
	.w6(32'h3d1bff80),
	.w7(32'h3ca0f773),
	.w8(32'h3b9ee3a9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule