module layer_6_featuremap_15(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f2332d),
	.w1(32'hb795ee0b),
	.w2(32'hb790aabe),
	.w3(32'hb7a0886b),
	.w4(32'hb73d7952),
	.w5(32'hb70ebdb5),
	.w6(32'hb75bf18d),
	.w7(32'hb71ca87b),
	.w8(32'hb6bcb218),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7989f4f),
	.w1(32'hb5a59428),
	.w2(32'h36df782f),
	.w3(32'hb68b4292),
	.w4(32'h375331bf),
	.w5(32'h37925f7b),
	.w6(32'hb6e4285e),
	.w7(32'h36fd3a68),
	.w8(32'h37455327),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77c4f37),
	.w1(32'hb7aa4444),
	.w2(32'hb728e170),
	.w3(32'hb84a9967),
	.w4(32'hb846a9e0),
	.w5(32'hb8251554),
	.w6(32'hb7a9aa81),
	.w7(32'hb77a6ffb),
	.w8(32'hb2d1d0b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addf9be),
	.w1(32'h3af1de89),
	.w2(32'h3ae849ef),
	.w3(32'h3ac09bd0),
	.w4(32'h3a92c6eb),
	.w5(32'h3a40b5f0),
	.w6(32'h3a4bbf51),
	.w7(32'h3a2b1e3d),
	.w8(32'h39b14234),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c751c),
	.w1(32'hba83cbd4),
	.w2(32'hba4f5ff2),
	.w3(32'hba76f1a9),
	.w4(32'hba750548),
	.w5(32'hba444c7e),
	.w6(32'hba62ebbf),
	.w7(32'hba467e59),
	.w8(32'hba1aad10),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e43393),
	.w1(32'h37eaac39),
	.w2(32'h37b6a423),
	.w3(32'h372a3470),
	.w4(32'h37670485),
	.w5(32'h36458e0a),
	.w6(32'h370ec833),
	.w7(32'h37117533),
	.w8(32'h35545a18),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ac5378),
	.w1(32'h3848af03),
	.w2(32'h38e547dc),
	.w3(32'hb8528967),
	.w4(32'hb7e199fa),
	.w5(32'h379e66f1),
	.w6(32'hb8a87d0d),
	.w7(32'hb723b7f6),
	.w8(32'h37be669f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39451b00),
	.w1(32'h38ec8415),
	.w2(32'h389f06ee),
	.w3(32'h395299b0),
	.w4(32'h38f046a7),
	.w5(32'h384d562b),
	.w6(32'h394cdb43),
	.w7(32'h38f72ef8),
	.w8(32'h382970da),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a008841),
	.w1(32'h39cee522),
	.w2(32'h399b4c5d),
	.w3(32'h39ad4753),
	.w4(32'h39363491),
	.w5(32'h3891e84d),
	.w6(32'h39bf8a89),
	.w7(32'h394d59d8),
	.w8(32'h38e9c3ae),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c6a90),
	.w1(32'hb785892d),
	.w2(32'h37daafad),
	.w3(32'hb825d9c1),
	.w4(32'hb8b7f062),
	.w5(32'hb89c186f),
	.w6(32'hb87d4a1f),
	.w7(32'hb8d5eb33),
	.w8(32'hb90ed490),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0685c),
	.w1(32'h3a82c5ac),
	.w2(32'h3a1c830a),
	.w3(32'h3a8686c9),
	.w4(32'h39e3db6b),
	.w5(32'hb89970f3),
	.w6(32'h3ab9966a),
	.w7(32'h3a7175b9),
	.w8(32'h3a04cf26),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1676d),
	.w1(32'hb7edb77c),
	.w2(32'hb85e47fc),
	.w3(32'h3716cdce),
	.w4(32'h3710ad33),
	.w5(32'hb7b017f0),
	.w6(32'h375f0db0),
	.w7(32'h3789b8b1),
	.w8(32'hb7a42c72),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368d96a0),
	.w1(32'hb6523579),
	.w2(32'h38010081),
	.w3(32'h3725051f),
	.w4(32'h37921f1c),
	.w5(32'h38279f52),
	.w6(32'hb6d2f5e4),
	.w7(32'hb7b5ba20),
	.w8(32'h37f66fae),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f366c9),
	.w1(32'hba34bda1),
	.w2(32'hba40b869),
	.w3(32'hba089c79),
	.w4(32'hba616b05),
	.w5(32'hba62f421),
	.w6(32'h37373323),
	.w7(32'hb8a8d1b5),
	.w8(32'hb95f53a4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3870553a),
	.w1(32'h380a01a7),
	.w2(32'h3840703d),
	.w3(32'h36f4d23c),
	.w4(32'h35b30613),
	.w5(32'hb670c027),
	.w6(32'hb6b9ea57),
	.w7(32'hb797625e),
	.w8(32'hb79e02ac),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31f4b7),
	.w1(32'h3a0ff6c0),
	.w2(32'h39c0c71a),
	.w3(32'h3a32c9ae),
	.w4(32'h39d53034),
	.w5(32'h391902c8),
	.w6(32'h3a360319),
	.w7(32'h39daf998),
	.w8(32'h3914f3d7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3bef8),
	.w1(32'hba393d4e),
	.w2(32'hba14d0f8),
	.w3(32'hbaa2285b),
	.w4(32'hbabab93d),
	.w5(32'hba8c0d93),
	.w6(32'hb9f8841f),
	.w7(32'hba644ca2),
	.w8(32'hb9fcd80b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6893d76),
	.w1(32'h3609ecb9),
	.w2(32'hb2796607),
	.w3(32'h36842dac),
	.w4(32'h37655bd1),
	.w5(32'h36a6ecce),
	.w6(32'h3502b076),
	.w7(32'h374921d1),
	.w8(32'h36960af7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb49e4),
	.w1(32'hb9d2fe7a),
	.w2(32'hb9ad85b3),
	.w3(32'hb9a53785),
	.w4(32'hb9a2b102),
	.w5(32'hb999fda9),
	.w6(32'hb9ed9bb3),
	.w7(32'hba01813a),
	.w8(32'hb9c241e7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9493430),
	.w1(32'hb9b2bcf7),
	.w2(32'hb983652a),
	.w3(32'hb9de4ee5),
	.w4(32'hba1398f0),
	.w5(32'hb9ebe4e0),
	.w6(32'hb9165c39),
	.w7(32'hb9b97be1),
	.w8(32'hb932409a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a426398),
	.w1(32'h3a28bd89),
	.w2(32'h3a2eb02d),
	.w3(32'h3941bf75),
	.w4(32'h38e3ed4d),
	.w5(32'h3918a204),
	.w6(32'h3a23361b),
	.w7(32'h39d48ba1),
	.w8(32'h39f561ff),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba816a8e),
	.w1(32'hba9da0c1),
	.w2(32'hba7b73d5),
	.w3(32'hbaa11fb4),
	.w4(32'hbaa56a29),
	.w5(32'hba57ae48),
	.w6(32'hba39a6a2),
	.w7(32'hba432a3a),
	.w8(32'hb9e1c512),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6cca4),
	.w1(32'hb829fbd9),
	.w2(32'hb91ba588),
	.w3(32'h3940cbd9),
	.w4(32'h38461f79),
	.w5(32'hb8d6452a),
	.w6(32'h398359d1),
	.w7(32'h374ef1c1),
	.w8(32'hb8cab52a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bbac2),
	.w1(32'hba804457),
	.w2(32'hba9b0b17),
	.w3(32'hba30987f),
	.w4(32'hba9bfcbb),
	.w5(32'hbab3b0c3),
	.w6(32'h37ec53c4),
	.w7(32'hb9b797cb),
	.w8(32'hba40cc6e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914417),
	.w1(32'h3b834638),
	.w2(32'h3b645c98),
	.w3(32'h3b109b0a),
	.w4(32'h3a8da7e2),
	.w5(32'h3a04684c),
	.w6(32'h3b5adb5a),
	.w7(32'h3b0b29d1),
	.w8(32'h3afb988e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c9bfa),
	.w1(32'h3b4898dc),
	.w2(32'h3b2843ac),
	.w3(32'h3b3887aa),
	.w4(32'h3af3223e),
	.w5(32'h3aa28d95),
	.w6(32'h3b1e58f8),
	.w7(32'h3ac1eca3),
	.w8(32'h3a84d71b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82ab7b),
	.w1(32'hba41ae3f),
	.w2(32'hba107b7d),
	.w3(32'hba2022e3),
	.w4(32'hba1c17d8),
	.w5(32'hb9d63130),
	.w6(32'hba11e2e4),
	.w7(32'hb9893b1c),
	.w8(32'hb95ce99c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cb3a78),
	.w1(32'h361f1a90),
	.w2(32'h37303ac8),
	.w3(32'h3633abaf),
	.w4(32'h3650541d),
	.w5(32'h354786c2),
	.w6(32'h368b6cea),
	.w7(32'h367e930d),
	.w8(32'h3706916b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2c65d),
	.w1(32'hb878226c),
	.w2(32'hb8881294),
	.w3(32'hb7fef569),
	.w4(32'hb8277512),
	.w5(32'hb7ece970),
	.w6(32'h36807ad0),
	.w7(32'h361ab7e8),
	.w8(32'hb6d5e45e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53b046),
	.w1(32'h3b323a5f),
	.w2(32'h3b172a7e),
	.w3(32'h3b6312a6),
	.w4(32'h3b1eb0ed),
	.w5(32'h3aeea353),
	.w6(32'h3b3cb048),
	.w7(32'h3b00ee8d),
	.w8(32'h3aa02e04),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3639a1a1),
	.w1(32'hbccf787c),
	.w2(32'h3b89deee),
	.w3(32'h374df8be),
	.w4(32'hbc3fb652),
	.w5(32'hbcfb10e8),
	.w6(32'hbb529dfe),
	.w7(32'hbc0f1fd3),
	.w8(32'hbcd2efa0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dcdbf),
	.w1(32'h3b79a978),
	.w2(32'h3b89df37),
	.w3(32'hbcd20df2),
	.w4(32'hbc615062),
	.w5(32'hbc939e2f),
	.w6(32'h3bc7ab3a),
	.w7(32'h3b9ce011),
	.w8(32'h3cbff19f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f14b5),
	.w1(32'hbc4f79d2),
	.w2(32'hbdc5c131),
	.w3(32'hbc8cf789),
	.w4(32'h3d0083f0),
	.w5(32'h3c0d305f),
	.w6(32'hbd3ea216),
	.w7(32'hbdd3a2e6),
	.w8(32'hbd41cf2d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96fdd7),
	.w1(32'hbd0b271d),
	.w2(32'hbc7c2c90),
	.w3(32'h3d348af5),
	.w4(32'h3cce03af),
	.w5(32'h3d289e5a),
	.w6(32'hbc3bcd2b),
	.w7(32'hbc772473),
	.w8(32'hbbb5195c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8a28c),
	.w1(32'h3b52eb59),
	.w2(32'hbc8b3047),
	.w3(32'h3bcd0527),
	.w4(32'hbb4dd9f2),
	.w5(32'hbaf00e89),
	.w6(32'h3caa0615),
	.w7(32'hbc1adf81),
	.w8(32'h3b4efc38),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c714d),
	.w1(32'hbbabdbba),
	.w2(32'h3ca43d8b),
	.w3(32'h3b1ee488),
	.w4(32'h3bd18355),
	.w5(32'h3c66c7a4),
	.w6(32'hbc0ecb08),
	.w7(32'hbd0237c5),
	.w8(32'hbb608310),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45e0b4),
	.w1(32'h3ba5a190),
	.w2(32'h3c548108),
	.w3(32'hbc858a4e),
	.w4(32'h3c023319),
	.w5(32'h3c677961),
	.w6(32'hbc615ede),
	.w7(32'hbc9518a5),
	.w8(32'hbb83a6cd),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5580b9),
	.w1(32'hbc9e03c4),
	.w2(32'hbc9c00cb),
	.w3(32'h3b4dcd34),
	.w4(32'hbc11e9cd),
	.w5(32'hbc221198),
	.w6(32'hbb31976a),
	.w7(32'h3cc01e72),
	.w8(32'hbc0aa474),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0907),
	.w1(32'h3c4e89b0),
	.w2(32'h3bfdcd71),
	.w3(32'hbd14ee8a),
	.w4(32'hbbd4f678),
	.w5(32'hbc149c40),
	.w6(32'h3c83b9db),
	.w7(32'h3c43c731),
	.w8(32'h3b8ae1be),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa13476),
	.w1(32'h3bab10e6),
	.w2(32'hbcbfc239),
	.w3(32'hbc1129f6),
	.w4(32'h3d0a2311),
	.w5(32'h3c90f546),
	.w6(32'hbb415174),
	.w7(32'hbd17b433),
	.w8(32'h3b50f76b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b884e),
	.w1(32'hbb0c0a1f),
	.w2(32'h3bd24d20),
	.w3(32'h3c598800),
	.w4(32'hb7b6244d),
	.w5(32'h3bcde686),
	.w6(32'hb9ecf412),
	.w7(32'hbc95757c),
	.w8(32'hbc09e85e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaef61),
	.w1(32'h3c1e5a4a),
	.w2(32'h3bdc8e49),
	.w3(32'hbad07559),
	.w4(32'hb9c85b4a),
	.w5(32'hbb2474fd),
	.w6(32'h3c3adb2e),
	.w7(32'h3bf22b42),
	.w8(32'h3b925dd5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5142),
	.w1(32'hbb958cee),
	.w2(32'h3c183f68),
	.w3(32'h3a334230),
	.w4(32'hba8a76c6),
	.w5(32'h3b0d4861),
	.w6(32'hbd14569b),
	.w7(32'hbd27575c),
	.w8(32'hbc776268),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc092f),
	.w1(32'h3bb60737),
	.w2(32'h3bc306b2),
	.w3(32'hbbaa93a6),
	.w4(32'h3c422945),
	.w5(32'h3bef7b52),
	.w6(32'hbbaf794a),
	.w7(32'hbbcd6263),
	.w8(32'h3a6fa72f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdca33),
	.w1(32'hbc2ac4a8),
	.w2(32'hbcf999cf),
	.w3(32'hbbf5487b),
	.w4(32'hbc109d9b),
	.w5(32'hbd2e875e),
	.w6(32'h3d0dec45),
	.w7(32'h3d0e0f7f),
	.w8(32'h3c62d9bd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359ab6),
	.w1(32'hbb2cfb98),
	.w2(32'hbcc05038),
	.w3(32'hbc0b0b2a),
	.w4(32'hbcad0f2c),
	.w5(32'hbcbe4973),
	.w6(32'h3b470165),
	.w7(32'hbb007667),
	.w8(32'h3b985ab1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805252),
	.w1(32'hbc9a5071),
	.w2(32'hbcb25584),
	.w3(32'hbb929031),
	.w4(32'hbcf995fc),
	.w5(32'hbcc1dda6),
	.w6(32'h377c313a),
	.w7(32'hbc9e7a05),
	.w8(32'h3c818177),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc39389),
	.w1(32'h3a8e70c6),
	.w2(32'h3d0325fc),
	.w3(32'hbbb0f84c),
	.w4(32'hbd19fa21),
	.w5(32'hbcdc1755),
	.w6(32'hbc8510fb),
	.w7(32'hbc053db5),
	.w8(32'h3b4a1582),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8001b),
	.w1(32'h3c0d7cf8),
	.w2(32'hbcc64141),
	.w3(32'hbd02eca9),
	.w4(32'h3c8a820a),
	.w5(32'h3c6f082c),
	.w6(32'hbc99b430),
	.w7(32'hbc331b08),
	.w8(32'hbc25794d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f02e5),
	.w1(32'hbc4608ec),
	.w2(32'h3c18cb7e),
	.w3(32'hbc0adbc5),
	.w4(32'hbcbea674),
	.w5(32'hbc9287f6),
	.w6(32'h3c6897a0),
	.w7(32'h3c53315a),
	.w8(32'hbbc482f2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c997502),
	.w1(32'h3b0f3126),
	.w2(32'h3c01820f),
	.w3(32'hbc6583ff),
	.w4(32'h3bed2943),
	.w5(32'h3b82361f),
	.w6(32'hbbf4ce1f),
	.w7(32'hbc5126e2),
	.w8(32'hbbae5b15),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5856c3),
	.w1(32'h3c33dac0),
	.w2(32'hbc3182cb),
	.w3(32'h3b261af0),
	.w4(32'h3bdd6875),
	.w5(32'h3c33e7db),
	.w6(32'hbb24b79b),
	.w7(32'hbbc22d60),
	.w8(32'hbbd8acd4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32b984),
	.w1(32'h3bfce526),
	.w2(32'h3afa84b1),
	.w3(32'h3a8a6d1a),
	.w4(32'h3c785a04),
	.w5(32'h3cfd435f),
	.w6(32'h3baba143),
	.w7(32'hbcbff13b),
	.w8(32'hbbb97c0b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aa187),
	.w1(32'h3b912fc5),
	.w2(32'h3a8a4531),
	.w3(32'h3bec3e76),
	.w4(32'h3c04d398),
	.w5(32'hbb37dbea),
	.w6(32'hbb93262b),
	.w7(32'hbca9e446),
	.w8(32'hbc36d0c0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e34d),
	.w1(32'hbc807c9c),
	.w2(32'hbce4bc62),
	.w3(32'hbbb524c7),
	.w4(32'hbc260cea),
	.w5(32'hbc910374),
	.w6(32'h3c21b467),
	.w7(32'hbb8a181d),
	.w8(32'h37f21db9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c862c),
	.w1(32'h3c2b6ecc),
	.w2(32'hbc2147ad),
	.w3(32'hbb2ef8bc),
	.w4(32'h3c663d9b),
	.w5(32'hbc5e289f),
	.w6(32'hbc2b3db0),
	.w7(32'hbca56a09),
	.w8(32'h3cd19c3d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d8e32),
	.w1(32'h3c136e7f),
	.w2(32'hbb34a61f),
	.w3(32'hbca12e35),
	.w4(32'h3b84e499),
	.w5(32'h3cce3afc),
	.w6(32'hbb489c1f),
	.w7(32'h3c102e6f),
	.w8(32'hbc85d606),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055ed9),
	.w1(32'hbbbc0631),
	.w2(32'h3c28ea1b),
	.w3(32'hbca75e84),
	.w4(32'hba9cfb9f),
	.w5(32'h3afbd390),
	.w6(32'h3cae7f4e),
	.w7(32'hbbb984f9),
	.w8(32'h3b990105),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd089),
	.w1(32'hbb7dabc9),
	.w2(32'hbcf0cb9d),
	.w3(32'hbbec637b),
	.w4(32'h3a1e1630),
	.w5(32'h36679cd2),
	.w6(32'h3c879684),
	.w7(32'hbc410fa8),
	.w8(32'hbc40c774),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0f42),
	.w1(32'h3ccd487b),
	.w2(32'h3cc490be),
	.w3(32'hbb0433ad),
	.w4(32'hbd4967b1),
	.w5(32'hbd729132),
	.w6(32'hbaa5565c),
	.w7(32'h3a57466e),
	.w8(32'h3c41b125),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82b8ac),
	.w1(32'hbbebe80c),
	.w2(32'h3ae4603f),
	.w3(32'hbcc80497),
	.w4(32'hbc419743),
	.w5(32'hbd0e6b4f),
	.w6(32'h3c5a54a9),
	.w7(32'h3b86c9ed),
	.w8(32'h3ad6f580),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfa86c),
	.w1(32'h3c1ece19),
	.w2(32'hbb829c3d),
	.w3(32'hbc2cc0a9),
	.w4(32'h3c4a4317),
	.w5(32'h3bc036b9),
	.w6(32'h3c28c3a2),
	.w7(32'hbc4b63a3),
	.w8(32'h3b6ce33a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c297),
	.w1(32'hbc3084c5),
	.w2(32'hbc361b41),
	.w3(32'h3cb9d988),
	.w4(32'hbc74a0d8),
	.w5(32'h3c175e1c),
	.w6(32'h3ce8a226),
	.w7(32'hbb08440a),
	.w8(32'hbcb0b8d6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4749f7),
	.w1(32'h39b6bcfb),
	.w2(32'h3c43a7e6),
	.w3(32'h3a6f382c),
	.w4(32'hbd07af6a),
	.w5(32'h3c4b7193),
	.w6(32'h3d0f5181),
	.w7(32'h3c8c7294),
	.w8(32'h3c2c456d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule