module layer_10_featuremap_326(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f05f38),
	.w1(32'h36e1cff7),
	.w2(32'h36833b3e),
	.w3(32'hb5a22dba),
	.w4(32'hb51071e6),
	.w5(32'hb5087f99),
	.w6(32'hb734d92a),
	.w7(32'hb647addf),
	.w8(32'hb6756a6a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c765ac),
	.w1(32'hb9284914),
	.w2(32'hb8ddfc7c),
	.w3(32'hb8d0c8ca),
	.w4(32'hb8c0d1e6),
	.w5(32'hb8cb4282),
	.w6(32'hb7913bf6),
	.w7(32'hb8450ccb),
	.w8(32'hb8827376),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb642cf2b),
	.w1(32'hb6f21e86),
	.w2(32'hb67802f1),
	.w3(32'hb60eefbe),
	.w4(32'h343a0fb4),
	.w5(32'h367e9672),
	.w6(32'hb5861e09),
	.w7(32'hb59eac91),
	.w8(32'h36ae27b4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6471d8c),
	.w1(32'h37037c04),
	.w2(32'h37a9a263),
	.w3(32'h3493e0bf),
	.w4(32'h3701a898),
	.w5(32'h380c8bc9),
	.w6(32'h36e420e1),
	.w7(32'h3781fea2),
	.w8(32'hb707ec9f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62309df),
	.w1(32'hb7db387c),
	.w2(32'h38095598),
	.w3(32'h373e6381),
	.w4(32'hb7cf2ede),
	.w5(32'hb7866dfd),
	.w6(32'h381606b5),
	.w7(32'hb8126139),
	.w8(32'h36cb5a14),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33a32d25),
	.w1(32'h3506bd0d),
	.w2(32'h35d596a5),
	.w3(32'hb620ee3d),
	.w4(32'hb585c23e),
	.w5(32'hb5ab8c0b),
	.w6(32'hb6b0e4a0),
	.w7(32'hb6a22223),
	.w8(32'h3495e909),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb763e0db),
	.w1(32'h3815760c),
	.w2(32'hb79924db),
	.w3(32'h3842a681),
	.w4(32'h380bf00a),
	.w5(32'h363d99bb),
	.w6(32'hb82f8d0e),
	.w7(32'hb483a5a2),
	.w8(32'hb8209983),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c59ce),
	.w1(32'hb889ba04),
	.w2(32'h383eb712),
	.w3(32'hb98ca15a),
	.w4(32'hb7e51fbb),
	.w5(32'h38c9e4d5),
	.w6(32'hb8363780),
	.w7(32'hb7cb0fc5),
	.w8(32'h37d35ef3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3734835d),
	.w1(32'hb8d6f397),
	.w2(32'hb88366ed),
	.w3(32'hb9281666),
	.w4(32'hb8f461a4),
	.w5(32'hb84abe2d),
	.w6(32'hb9036d42),
	.w7(32'hb78bb4bd),
	.w8(32'hb86fa7a2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b7ad3),
	.w1(32'h39808854),
	.w2(32'hb8b3d34d),
	.w3(32'hb7b4f552),
	.w4(32'hb98def5a),
	.w5(32'hb98a362a),
	.w6(32'hb9df5c9f),
	.w7(32'hb99a7b7c),
	.w8(32'hb913bf21),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899acea),
	.w1(32'hb90c2e3b),
	.w2(32'h383d24d6),
	.w3(32'hb8c23ccc),
	.w4(32'hb7ec3f6b),
	.w5(32'h392e6f9a),
	.w6(32'hb846cc2f),
	.w7(32'h36a2e756),
	.w8(32'h39426926),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8840e00),
	.w1(32'h38f59569),
	.w2(32'h385f5f7a),
	.w3(32'h38ebd228),
	.w4(32'h392010ca),
	.w5(32'h392b5e26),
	.w6(32'h389f99d9),
	.w7(32'h38f07ccc),
	.w8(32'h38cdf15e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39862239),
	.w1(32'h393e598c),
	.w2(32'hb8a362c7),
	.w3(32'hb92014b7),
	.w4(32'hb8b7415b),
	.w5(32'hb9486b43),
	.w6(32'hb94609cd),
	.w7(32'hb84a34ef),
	.w8(32'hb958e658),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2c120),
	.w1(32'hb8da0cb9),
	.w2(32'hb7760554),
	.w3(32'h37a199ca),
	.w4(32'hb8f91eb6),
	.w5(32'hb90a12c9),
	.w6(32'h38387b2d),
	.w7(32'hb8084930),
	.w8(32'h37bd27f6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a669d5),
	.w1(32'hb9548a6a),
	.w2(32'hb97dd4e0),
	.w3(32'hba135ecd),
	.w4(32'hba2d7b36),
	.w5(32'hba12db64),
	.w6(32'hb7524f26),
	.w7(32'hb9344c30),
	.w8(32'hb9d8d035),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c2726),
	.w1(32'hb7a9113e),
	.w2(32'hb9237cd2),
	.w3(32'hb8fab097),
	.w4(32'hb890b2a2),
	.w5(32'h3766122f),
	.w6(32'hb87cac5c),
	.w7(32'h38bc1491),
	.w8(32'h38aac046),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h337dc279),
	.w1(32'h38aeb4ba),
	.w2(32'h38a7a160),
	.w3(32'h38b96a9f),
	.w4(32'h3859ff2b),
	.w5(32'h3920ebef),
	.w6(32'hb82b3356),
	.w7(32'hb804f9f9),
	.w8(32'h3720e079),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bb2de),
	.w1(32'h3989c205),
	.w2(32'h3932ece3),
	.w3(32'hb85c86db),
	.w4(32'h38ccdecd),
	.w5(32'h39401404),
	.w6(32'h38dd41c4),
	.w7(32'h3990edb6),
	.w8(32'h399bae2a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385b243e),
	.w1(32'h3953fcf2),
	.w2(32'h38a98d00),
	.w3(32'h37cd0a80),
	.w4(32'h3981ca82),
	.w5(32'h3946aeac),
	.w6(32'hb836fb18),
	.w7(32'h39303f18),
	.w8(32'h392c992c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb690afb3),
	.w1(32'hb6ebfb2f),
	.w2(32'h35d833ee),
	.w3(32'hb5fa3d17),
	.w4(32'h36f68f71),
	.w5(32'hb6b056d1),
	.w6(32'hb6952078),
	.w7(32'h35c02102),
	.w8(32'hb6c48ce4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62b72c2),
	.w1(32'h36fa986e),
	.w2(32'h3600a77e),
	.w3(32'hb34fcfff),
	.w4(32'h370d8355),
	.w5(32'h36e4afc0),
	.w6(32'hb69edd18),
	.w7(32'hb4562c39),
	.w8(32'h365a65bd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8b9df),
	.w1(32'hb8507d17),
	.w2(32'h386f2b7b),
	.w3(32'hb7aabdfc),
	.w4(32'hb76aec97),
	.w5(32'h385b068d),
	.w6(32'h38973b94),
	.w7(32'hb6a361e3),
	.w8(32'h3867688b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf3f91),
	.w1(32'h396738d5),
	.w2(32'hb90f4cb5),
	.w3(32'hba20cb2c),
	.w4(32'hba179160),
	.w5(32'hb9a3927c),
	.w6(32'hb924df95),
	.w7(32'hb9175fa6),
	.w8(32'h36bee293),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399bffed),
	.w1(32'h39185c71),
	.w2(32'hb869234c),
	.w3(32'hb8b8c823),
	.w4(32'hb92227ff),
	.w5(32'hb90ed580),
	.w6(32'hb72b4c62),
	.w7(32'h38a7fd3e),
	.w8(32'h3832fd82),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a33dd1),
	.w1(32'hb8c33816),
	.w2(32'hb7684d7d),
	.w3(32'hb90ed960),
	.w4(32'hb9199e24),
	.w5(32'hb7f09939),
	.w6(32'hb8cfd8b1),
	.w7(32'hb90532de),
	.w8(32'h378f11e6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888d558),
	.w1(32'hb91ad621),
	.w2(32'hb88919b8),
	.w3(32'hb94cc811),
	.w4(32'hb9936a9f),
	.w5(32'hb9115fd0),
	.w6(32'hb8fa95c4),
	.w7(32'hb943476e),
	.w8(32'hb914d9aa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362628c8),
	.w1(32'h36a5eb44),
	.w2(32'h34b3ffd9),
	.w3(32'h372faa64),
	.w4(32'h36d0292a),
	.w5(32'h367d7837),
	.w6(32'h3784f72a),
	.w7(32'h36989bf7),
	.w8(32'hb713f693),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f60e3),
	.w1(32'h38513a15),
	.w2(32'hb85ffb83),
	.w3(32'h39324c2e),
	.w4(32'h38832759),
	.w5(32'hb8b7c269),
	.w6(32'h39142761),
	.w7(32'h38ffdf5f),
	.w8(32'hb7dcdb1f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0b04f),
	.w1(32'hb7769932),
	.w2(32'hb77f0b79),
	.w3(32'h37f9ef29),
	.w4(32'h37a246ee),
	.w5(32'hb8262d2b),
	.w6(32'h390ac233),
	.w7(32'h388b4dcb),
	.w8(32'h38636b68),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa50fd),
	.w1(32'h346e742a),
	.w2(32'hb9780f24),
	.w3(32'hb97b8cc4),
	.w4(32'hb9e72d81),
	.w5(32'hb9d82b02),
	.w6(32'hb9449ac7),
	.w7(32'hb941876a),
	.w8(32'hb98dda7a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356dbe1e),
	.w1(32'h36743eed),
	.w2(32'h361ad583),
	.w3(32'h37a01dc7),
	.w4(32'h3748612f),
	.w5(32'hb5ec5054),
	.w6(32'hb7832221),
	.w7(32'hb72f41d9),
	.w8(32'h3747baf8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7239193),
	.w1(32'hb6914983),
	.w2(32'hb6ba7483),
	.w3(32'hb56a7096),
	.w4(32'hb5ae2a0a),
	.w5(32'h36c964aa),
	.w6(32'h3705107b),
	.w7(32'h374b3136),
	.w8(32'hb611d69b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39168653),
	.w1(32'h39158a63),
	.w2(32'h3843c9c6),
	.w3(32'hb8c2be7d),
	.w4(32'hb8a66c75),
	.w5(32'hb83686ad),
	.w6(32'hb8c2a686),
	.w7(32'hb860e74d),
	.w8(32'hb7189154),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39655200),
	.w1(32'h390c4318),
	.w2(32'h38b603f5),
	.w3(32'h38d1caeb),
	.w4(32'h3860b3de),
	.w5(32'h38e2a133),
	.w6(32'hb88b6feb),
	.w7(32'h3889da61),
	.w8(32'h38b5849e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fad183),
	.w1(32'h375443f8),
	.w2(32'h3469632f),
	.w3(32'h374b1c8d),
	.w4(32'h37811205),
	.w5(32'h367600c4),
	.w6(32'h36c6d0ba),
	.w7(32'h35d43198),
	.w8(32'hb62290f0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6993007),
	.w1(32'h38081604),
	.w2(32'h36d7bcbc),
	.w3(32'h373300f7),
	.w4(32'h38145c23),
	.w5(32'h382be2dc),
	.w6(32'hb7bbda33),
	.w7(32'h373c420d),
	.w8(32'hb66449d9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63d7e96),
	.w1(32'hb882674c),
	.w2(32'h38d8b1df),
	.w3(32'hb8bb2080),
	.w4(32'hb97621f6),
	.w5(32'h37bc3539),
	.w6(32'hb9b525e5),
	.w7(32'hb9a48a53),
	.w8(32'hb7efef03),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01b6bd),
	.w1(32'hb9b06f02),
	.w2(32'h38f01be2),
	.w3(32'h383389ea),
	.w4(32'hb8b1b013),
	.w5(32'h3955048b),
	.w6(32'h3a0239f5),
	.w7(32'hb55e3643),
	.w8(32'h3994359e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6fe28),
	.w1(32'hb9d7d044),
	.w2(32'hb8d7d9e0),
	.w3(32'h39012cfd),
	.w4(32'hb9132acb),
	.w5(32'hb7a106b8),
	.w6(32'h39c385be),
	.w7(32'hb7dc4668),
	.w8(32'h391011b1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7954bc8),
	.w1(32'hb842fce8),
	.w2(32'hb806c0aa),
	.w3(32'hb817f4ed),
	.w4(32'hb82fc979),
	.w5(32'hb81158f1),
	.w6(32'hb7874c6f),
	.w7(32'hb7998aa8),
	.w8(32'hb7967e4d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e6dfb2),
	.w1(32'hb696396f),
	.w2(32'hb6e885cc),
	.w3(32'hb753dc13),
	.w4(32'hb700c426),
	.w5(32'hb6bf529e),
	.w6(32'hb7af9369),
	.w7(32'hb7979671),
	.w8(32'hb737ae0e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7218a71),
	.w1(32'h36e2544a),
	.w2(32'h379740b2),
	.w3(32'h3725122b),
	.w4(32'h373f0c9d),
	.w5(32'h37c0d6ba),
	.w6(32'h379c741d),
	.w7(32'h373d2a9f),
	.w8(32'h372e2364),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384fd113),
	.w1(32'hb75a1f82),
	.w2(32'hb8506a14),
	.w3(32'h381dc603),
	.w4(32'hb8bd5361),
	.w5(32'h36fc0f90),
	.w6(32'h3855fa33),
	.w7(32'hb7fde153),
	.w8(32'h38979738),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc95ac),
	.w1(32'hb7ff545e),
	.w2(32'hb986b49d),
	.w3(32'hb9e0a8d7),
	.w4(32'hb9867d37),
	.w5(32'hb9a98a0a),
	.w6(32'hb9aad8b1),
	.w7(32'hb8c4b40f),
	.w8(32'hb98b7bf6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987f331),
	.w1(32'h38e03968),
	.w2(32'hb78c5fb3),
	.w3(32'hb984b534),
	.w4(32'hb9a73e43),
	.w5(32'hb962dd33),
	.w6(32'hb976439b),
	.w7(32'hb914b1e9),
	.w8(32'hb899feb5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395472c8),
	.w1(32'h38d1e9a7),
	.w2(32'hb86040e5),
	.w3(32'hb98ca1bd),
	.w4(32'hb98ee397),
	.w5(32'hb955465f),
	.w6(32'hb95236d8),
	.w7(32'hb8c7f2f5),
	.w8(32'hb9034d4d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39063f7e),
	.w1(32'h3900537e),
	.w2(32'h378e4905),
	.w3(32'hb8fd362d),
	.w4(32'hb91fed87),
	.w5(32'hb8f1cb09),
	.w6(32'hb91bcea9),
	.w7(32'hb8a2cb64),
	.w8(32'hb8b1c80a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386078f3),
	.w1(32'hb8f3cb2c),
	.w2(32'hb91dda04),
	.w3(32'h37adf010),
	.w4(32'hb8c03c61),
	.w5(32'hb9d70b7f),
	.w6(32'hb68ca5e0),
	.w7(32'h3782edbe),
	.w8(32'hb9650338),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e0357),
	.w1(32'hb8630b1f),
	.w2(32'hb830ff68),
	.w3(32'hb8bdd166),
	.w4(32'hb89ed8d3),
	.w5(32'hb84af9d8),
	.w6(32'hb78d3e1e),
	.w7(32'hb8785a46),
	.w8(32'hb833ed06),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387588b4),
	.w1(32'h38df64c0),
	.w2(32'h37ba2b91),
	.w3(32'h37c39ccb),
	.w4(32'h38b19aa2),
	.w5(32'hb6ec22ae),
	.w6(32'h38c49f19),
	.w7(32'h39748f67),
	.w8(32'h394256c4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8130f05),
	.w1(32'hb7f56160),
	.w2(32'hb74c7ce9),
	.w3(32'hb7ffda4a),
	.w4(32'hb8206f4a),
	.w5(32'hb72664d2),
	.w6(32'hb887f9b3),
	.w7(32'hb8cbbb97),
	.w8(32'hb858fb35),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38142ecf),
	.w1(32'h3814c4c9),
	.w2(32'h377bf80c),
	.w3(32'h38007fdb),
	.w4(32'h37ec0165),
	.w5(32'h37a91274),
	.w6(32'hb784dac8),
	.w7(32'h3603de48),
	.w8(32'h360d26b3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e7384),
	.w1(32'hb7d3334c),
	.w2(32'h370b3ef5),
	.w3(32'hb8fe4426),
	.w4(32'hb8b20a6c),
	.w5(32'h378df0f7),
	.w6(32'hb92dc005),
	.w7(32'hb8ee543d),
	.w8(32'hb8265a10),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395fc22e),
	.w1(32'hb8b62468),
	.w2(32'hb912d1c7),
	.w3(32'h38c7ecb5),
	.w4(32'hb96bb922),
	.w5(32'hb9b94ea4),
	.w6(32'hb8dee12b),
	.w7(32'h3868aebd),
	.w8(32'h3926a511),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379bbbac),
	.w1(32'h37261800),
	.w2(32'h3747c6bf),
	.w3(32'h37ffe3f7),
	.w4(32'h380e3d46),
	.w5(32'h370b5ec5),
	.w6(32'h3885f2df),
	.w7(32'h384f1966),
	.w8(32'h371a94a0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37067a0e),
	.w1(32'hb632d22b),
	.w2(32'hb69f2b56),
	.w3(32'h36d7d861),
	.w4(32'h34f287e6),
	.w5(32'hb6817e69),
	.w6(32'h368657d5),
	.w7(32'hb61ae3a5),
	.w8(32'hb5d48ff3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cfc732),
	.w1(32'h3556871a),
	.w2(32'h35d678d5),
	.w3(32'h36631d38),
	.w4(32'h36893d7f),
	.w5(32'h35c59454),
	.w6(32'h36614a2f),
	.w7(32'h364446c4),
	.w8(32'h3654a08b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d93dc9),
	.w1(32'hb6b09119),
	.w2(32'hb7058ce3),
	.w3(32'h366257d5),
	.w4(32'h358f183c),
	.w5(32'hb70b31d9),
	.w6(32'h36bb3d1f),
	.w7(32'h36708d0e),
	.w8(32'hb55c29f0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d162f),
	.w1(32'hb731fe66),
	.w2(32'h3730eb00),
	.w3(32'hb631a412),
	.w4(32'hb6112582),
	.w5(32'h379aed56),
	.w6(32'h37b7be82),
	.w7(32'hb72409f0),
	.w8(32'h37bff8b5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c7683),
	.w1(32'hb821013d),
	.w2(32'hb6258bb0),
	.w3(32'hb88f0bc5),
	.w4(32'h3719252b),
	.w5(32'h3600f43f),
	.w6(32'h38858174),
	.w7(32'h38988f7c),
	.w8(32'h385309c3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83fad81),
	.w1(32'h38562b00),
	.w2(32'h374cfacf),
	.w3(32'hb99f967a),
	.w4(32'h390c0c4a),
	.w5(32'hb67d3e19),
	.w6(32'hb91b7967),
	.w7(32'h395ba527),
	.w8(32'h37ea9f30),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e2e0d),
	.w1(32'h390dc9d5),
	.w2(32'h3873f17d),
	.w3(32'h384e2f0f),
	.w4(32'h38386941),
	.w5(32'h38525cd4),
	.w6(32'h37b1aec4),
	.w7(32'h360c9c1d),
	.w8(32'hb813b7f1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3714c66d),
	.w1(32'h37037df6),
	.w2(32'h360d82d8),
	.w3(32'h378f9d42),
	.w4(32'h3732c90a),
	.w5(32'hb5b3fc48),
	.w6(32'hb79c003d),
	.w7(32'hb784a41b),
	.w8(32'hb66a139a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3590d103),
	.w1(32'h364d6c2d),
	.w2(32'hb69d6dc2),
	.w3(32'h33ce93c2),
	.w4(32'h368776a6),
	.w5(32'h36503fb4),
	.w6(32'hb5d20f90),
	.w7(32'hb5c46a73),
	.w8(32'h364ceb3b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f6b9b5),
	.w1(32'h35aaf6ce),
	.w2(32'hb6a44c2c),
	.w3(32'h3637b096),
	.w4(32'h3491c19f),
	.w5(32'h379096c5),
	.w6(32'h36e8ae43),
	.w7(32'h36927aef),
	.w8(32'h36aacb1b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360aa2d3),
	.w1(32'hb6222efd),
	.w2(32'hb69ce404),
	.w3(32'h37815901),
	.w4(32'h37250a8e),
	.w5(32'h35fe5f67),
	.w6(32'hb6395229),
	.w7(32'hb5af3b8e),
	.w8(32'hb6c0ace6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2e063),
	.w1(32'h3908854a),
	.w2(32'h382704ba),
	.w3(32'h392a636a),
	.w4(32'h395e511c),
	.w5(32'h38ca59f2),
	.w6(32'h38aa57ab),
	.w7(32'h38d3a6c4),
	.w8(32'h3830994d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b683cb),
	.w1(32'h37944b66),
	.w2(32'hb882d3c4),
	.w3(32'hb85d7f37),
	.w4(32'hb87caa36),
	.w5(32'hb867830e),
	.w6(32'h384ab576),
	.w7(32'h388f341a),
	.w8(32'h37d093e3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f8644),
	.w1(32'h39032c21),
	.w2(32'h391c62a2),
	.w3(32'h3923fca7),
	.w4(32'h390f4cf7),
	.w5(32'h393a16b3),
	.w6(32'h3985878e),
	.w7(32'h396fc768),
	.w8(32'h39792892),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398702d7),
	.w1(32'hb9121708),
	.w2(32'hb86cc8ce),
	.w3(32'hb949eb49),
	.w4(32'hb9df3d9d),
	.w5(32'hb9aac087),
	.w6(32'hb7b0d6bc),
	.w7(32'hb961bfe5),
	.w8(32'hb9106d1b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3586a76c),
	.w1(32'h366528d2),
	.w2(32'hb5a0268c),
	.w3(32'hb616c016),
	.w4(32'hb63caf6f),
	.w5(32'hb609b574),
	.w6(32'hb7245cb2),
	.w7(32'hb713ea77),
	.w8(32'hb70c3f8b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360f0eaf),
	.w1(32'h35a28670),
	.w2(32'hb6e27aec),
	.w3(32'h36f1176b),
	.w4(32'h36817e71),
	.w5(32'hb48308fa),
	.w6(32'hb614e8de),
	.w7(32'hb6e5376d),
	.w8(32'hb6f0e28a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb754e40f),
	.w1(32'hb6cdab73),
	.w2(32'hb70f5ac1),
	.w3(32'hb19106aa),
	.w4(32'h36296620),
	.w5(32'h3708c2f1),
	.w6(32'h368734d8),
	.w7(32'h36323e64),
	.w8(32'hb4a84f0a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a28a90),
	.w1(32'hb68b6fa4),
	.w2(32'h37b02a45),
	.w3(32'h37622014),
	.w4(32'h38232340),
	.w5(32'h384e17d6),
	.w6(32'h380d9dc2),
	.w7(32'h375148be),
	.w8(32'h374cc097),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37123e43),
	.w1(32'h3531c9af),
	.w2(32'hb6330bb1),
	.w3(32'h3669e474),
	.w4(32'hb5024eba),
	.w5(32'hb668165a),
	.w6(32'hb5a0515b),
	.w7(32'hb6c7ea1e),
	.w8(32'hb7779741),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8377156),
	.w1(32'h3867eba2),
	.w2(32'h3831246f),
	.w3(32'hb6eeebc1),
	.w4(32'h38c3eaa6),
	.w5(32'h38744068),
	.w6(32'h37d1fe45),
	.w7(32'h383437c6),
	.w8(32'h37ad3f93),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db680e),
	.w1(32'hb917b78a),
	.w2(32'hb98c842a),
	.w3(32'hb9e29a6f),
	.w4(32'h397b0284),
	.w5(32'hb8c4c267),
	.w6(32'h38989065),
	.w7(32'h39511817),
	.w8(32'hb8cba6d7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79b0528),
	.w1(32'h38261551),
	.w2(32'h38791285),
	.w3(32'hb86794e5),
	.w4(32'h35f81ab1),
	.w5(32'h37612320),
	.w6(32'hb7f2ba08),
	.w7(32'h385a150d),
	.w8(32'h37f764f0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3854c053),
	.w1(32'hb8fb1030),
	.w2(32'hb8ab5dea),
	.w3(32'hb8fd7f23),
	.w4(32'hb8b034da),
	.w5(32'h37a6cdf3),
	.w6(32'h39158043),
	.w7(32'h38940842),
	.w8(32'h393759ff),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866a187),
	.w1(32'h387d205d),
	.w2(32'hb6982eb2),
	.w3(32'h38976c6d),
	.w4(32'h389520b6),
	.w5(32'hb7b93218),
	.w6(32'h37c8accf),
	.w7(32'h3801a670),
	.w8(32'h376ec17c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39189dcc),
	.w1(32'h3760233a),
	.w2(32'hb8eb2abf),
	.w3(32'hb8c299c7),
	.w4(32'hb93f47b5),
	.w5(32'hb931a43f),
	.w6(32'h37ce9f35),
	.w7(32'h3843a107),
	.w8(32'hb8501753),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb843483b),
	.w1(32'h3884045b),
	.w2(32'h37d86f7b),
	.w3(32'h364b5c55),
	.w4(32'h38a9c63f),
	.w5(32'h3857da1e),
	.w6(32'hb888a9f8),
	.w7(32'h38369309),
	.w8(32'h37ec9335),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35262c48),
	.w1(32'hb4be2862),
	.w2(32'h3634ac30),
	.w3(32'hb6323e0b),
	.w4(32'hb6096c5b),
	.w5(32'hb5d721d9),
	.w6(32'hb6f632fa),
	.w7(32'hb71d4709),
	.w8(32'h3546fe8d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ca24ab),
	.w1(32'hb71b19b7),
	.w2(32'hb70ade41),
	.w3(32'hb649004d),
	.w4(32'hb7a92256),
	.w5(32'hb7acbb38),
	.w6(32'hb7a70204),
	.w7(32'hb7f153b6),
	.w8(32'hb7c19238),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h32e052ec),
	.w1(32'hb60878ab),
	.w2(32'hb5f34c49),
	.w3(32'hb5ad7c82),
	.w4(32'h34f7fd80),
	.w5(32'h36ae94b2),
	.w6(32'hb6a29fd8),
	.w7(32'hb6b5e421),
	.w8(32'hb66a6b9e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb620334d),
	.w1(32'hb6d9f091),
	.w2(32'hb691bc79),
	.w3(32'hb58e16eb),
	.w4(32'hb744a0dd),
	.w5(32'hb7d15328),
	.w6(32'hb584b58e),
	.w7(32'hb6e17723),
	.w8(32'hb582ca17),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8040181),
	.w1(32'hb880267d),
	.w2(32'hb8399713),
	.w3(32'hb7dd5f07),
	.w4(32'hb82f1e06),
	.w5(32'hb79baf51),
	.w6(32'hb72e507e),
	.w7(32'hb7e869ec),
	.w8(32'hb7dcfea4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82dfc86),
	.w1(32'h37b1042f),
	.w2(32'h37f5d8c4),
	.w3(32'h3716cb76),
	.w4(32'h377c7c46),
	.w5(32'h370f7e88),
	.w6(32'hb5c2df69),
	.w7(32'hb7b5c2d4),
	.w8(32'hb7b36d2b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984320c),
	.w1(32'h3932cf99),
	.w2(32'hb8b13517),
	.w3(32'h375feb0f),
	.w4(32'hb89bf70d),
	.w5(32'hb88fba71),
	.w6(32'hb8db56b2),
	.w7(32'h3890634d),
	.w8(32'hb8519150),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378991bd),
	.w1(32'h39127229),
	.w2(32'h39150013),
	.w3(32'h385a7f14),
	.w4(32'h393d42f2),
	.w5(32'h3936c92c),
	.w6(32'h377b3234),
	.w7(32'h38e310d6),
	.w8(32'h38cf2e3f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85354f9),
	.w1(32'hb900996e),
	.w2(32'h36f614ff),
	.w3(32'h38991a8b),
	.w4(32'hb81b05ea),
	.w5(32'hb52c0cda),
	.w6(32'h392fd9d6),
	.w7(32'hb80f8474),
	.w8(32'h370f5ffd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39400a27),
	.w1(32'hb9f762ea),
	.w2(32'hb992999b),
	.w3(32'hb98b4a80),
	.w4(32'hba9a0931),
	.w5(32'hba307b32),
	.w6(32'hb94101b5),
	.w7(32'hba01b5e2),
	.w8(32'hba102b46),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4d663),
	.w1(32'hb73596f8),
	.w2(32'h37c939b0),
	.w3(32'h388c683d),
	.w4(32'hb887d78a),
	.w5(32'hb7954582),
	.w6(32'h38ee1b9c),
	.w7(32'hb76b55dc),
	.w8(32'h388ea3e8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc4c50),
	.w1(32'hb70afca3),
	.w2(32'hba077f17),
	.w3(32'hb95e0771),
	.w4(32'hb842c06b),
	.w5(32'hb9a289c6),
	.w6(32'hb8e24eef),
	.w7(32'h38ce0956),
	.w8(32'hb9603ccc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974bcbc),
	.w1(32'h38621976),
	.w2(32'hb98e8678),
	.w3(32'hb9e26f82),
	.w4(32'hb7cd82e6),
	.w5(32'hb9be41bf),
	.w6(32'hb9133766),
	.w7(32'h388c9d7e),
	.w8(32'hb90573b9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949d31b),
	.w1(32'h37d63e13),
	.w2(32'hb844f9b4),
	.w3(32'h382bf38b),
	.w4(32'hb881a4a3),
	.w5(32'hb83cc101),
	.w6(32'h389f93e1),
	.w7(32'h3785e767),
	.w8(32'hb8275d6d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8132140),
	.w1(32'hb71ba340),
	.w2(32'hb86d83df),
	.w3(32'h37f6ba6e),
	.w4(32'hb80cc2d9),
	.w5(32'hb8651cb9),
	.w6(32'h3890c2f2),
	.w7(32'hb7e929a3),
	.w8(32'hb85d8163),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939c942),
	.w1(32'h38658216),
	.w2(32'hb9401145),
	.w3(32'hb9f0c150),
	.w4(32'hb9cf4760),
	.w5(32'hb9abe65c),
	.w6(32'hb9d6a43e),
	.w7(32'hb983afad),
	.w8(32'hb991bf82),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d520cc),
	.w1(32'h38a54b7e),
	.w2(32'h3832e15b),
	.w3(32'h39a69698),
	.w4(32'h3902e454),
	.w5(32'h394fb7c4),
	.w6(32'h3924800a),
	.w7(32'h392e7c8f),
	.w8(32'h399ec4ee),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e0006),
	.w1(32'hb8daac23),
	.w2(32'h395372f0),
	.w3(32'hb91c1b1b),
	.w4(32'h389a7f4b),
	.w5(32'h3965d5c6),
	.w6(32'hb8f83b03),
	.w7(32'h38c3a57d),
	.w8(32'h393cc121),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b883bc),
	.w1(32'hba0d5ace),
	.w2(32'h391e60b5),
	.w3(32'h389010b6),
	.w4(32'hba82d4f0),
	.w5(32'hb9f7715a),
	.w6(32'h3a5d7d09),
	.w7(32'hb9882192),
	.w8(32'hb7fc0bd1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394337e0),
	.w1(32'hb792eaee),
	.w2(32'hb8da5ef4),
	.w3(32'hb9b7516a),
	.w4(32'hb9d24b69),
	.w5(32'hb9288c55),
	.w6(32'hb9d3c115),
	.w7(32'hb93f1feb),
	.w8(32'hb780b026),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39747e45),
	.w1(32'h39625dd7),
	.w2(32'h39031877),
	.w3(32'h39316b26),
	.w4(32'hb7a85d71),
	.w5(32'h38e916f2),
	.w6(32'hb9b7a0fe),
	.w7(32'hb9db87f4),
	.w8(32'hb9d3ac75),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84117bf),
	.w1(32'h37a2edb4),
	.w2(32'h384d242d),
	.w3(32'hb90b0ba8),
	.w4(32'hb80fbe14),
	.w5(32'hb6788358),
	.w6(32'hb9115cbf),
	.w7(32'hb89799b1),
	.w8(32'hb814fd40),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed91f8),
	.w1(32'h39960d2a),
	.w2(32'h39b77785),
	.w3(32'hb8d0f55f),
	.w4(32'h395d2e04),
	.w5(32'h39178e51),
	.w6(32'hb9abda53),
	.w7(32'hb9a51083),
	.w8(32'h37c015d6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ac80b),
	.w1(32'h38f43519),
	.w2(32'h384f913d),
	.w3(32'hb966f81b),
	.w4(32'h37e2348d),
	.w5(32'hb8b597d9),
	.w6(32'hb926af02),
	.w7(32'hb92360fe),
	.w8(32'hb9419b8d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b02126),
	.w1(32'hb6fa4cb8),
	.w2(32'h384ca7ee),
	.w3(32'h382170d0),
	.w4(32'h379358dd),
	.w5(32'h385e254f),
	.w6(32'hb7585178),
	.w7(32'hb78cbe0a),
	.w8(32'h37db0d30),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ba3ab0),
	.w1(32'hb895fee8),
	.w2(32'hb8285f51),
	.w3(32'hb821c16c),
	.w4(32'hb7096b2a),
	.w5(32'h37c87a3b),
	.w6(32'hb8ed0f4e),
	.w7(32'hb896933c),
	.w8(32'hb6ca3362),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39419aa4),
	.w1(32'h384ff23f),
	.w2(32'hb8b50c5d),
	.w3(32'hb9a8b0c7),
	.w4(32'hb98f5cca),
	.w5(32'hb941a298),
	.w6(32'hb9ace80c),
	.w7(32'hb94b09da),
	.w8(32'hb9758319),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ecd9f),
	.w1(32'hb6f307eb),
	.w2(32'hb949610d),
	.w3(32'hb9aac0c4),
	.w4(32'hb9970241),
	.w5(32'hb9b1303c),
	.w6(32'hb9c8ba6c),
	.w7(32'hb99d5ba9),
	.w8(32'hb9909fc0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b6f1b),
	.w1(32'hb94a4d95),
	.w2(32'hb92e3c2c),
	.w3(32'hb990d633),
	.w4(32'hba16f5eb),
	.w5(32'hb9ec6de2),
	.w6(32'hb905b7b4),
	.w7(32'hb912f086),
	.w8(32'hb99fa980),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b94c5),
	.w1(32'h3805f584),
	.w2(32'hb887fd19),
	.w3(32'h38283410),
	.w4(32'hb8a9a76b),
	.w5(32'hb88eca37),
	.w6(32'hb952af1e),
	.w7(32'hb94903cf),
	.w8(32'hb92e31d5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0c462),
	.w1(32'hb73a4682),
	.w2(32'hb824c790),
	.w3(32'h379202cb),
	.w4(32'hb666b565),
	.w5(32'hb7adb6cd),
	.w6(32'h38da9c8a),
	.w7(32'h3856c08b),
	.w8(32'h380f1306),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dfc81e),
	.w1(32'h389578d3),
	.w2(32'hb6b243ec),
	.w3(32'hb8053b78),
	.w4(32'h38a3755e),
	.w5(32'h36c7f58f),
	.w6(32'h390a98ea),
	.w7(32'h392c90ff),
	.w8(32'hb924101a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b45619),
	.w1(32'h37e64cc2),
	.w2(32'h3829a238),
	.w3(32'hb839306e),
	.w4(32'h37dd8e0a),
	.w5(32'h37f5ea0d),
	.w6(32'hb8abee61),
	.w7(32'h37f9659f),
	.w8(32'h37d1aa23),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79a2311),
	.w1(32'hb7c17aaa),
	.w2(32'h37defa70),
	.w3(32'hb7e7f863),
	.w4(32'hb79218c9),
	.w5(32'hb7986f7d),
	.w6(32'hb86ee7ef),
	.w7(32'hb805851c),
	.w8(32'hb7888456),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72874e7),
	.w1(32'hb70f8d1f),
	.w2(32'hb59672c3),
	.w3(32'hb7bda087),
	.w4(32'hb7975d92),
	.w5(32'h3823384f),
	.w6(32'hb69aa92e),
	.w7(32'hb685bd51),
	.w8(32'hb7a11445),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb1848),
	.w1(32'h37fb99d2),
	.w2(32'h36c24d9f),
	.w3(32'h3799327e),
	.w4(32'h382d0d14),
	.w5(32'h3875c9c4),
	.w6(32'hb83348d2),
	.w7(32'hb816c361),
	.w8(32'h3795e92f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94797db),
	.w1(32'hb9799852),
	.w2(32'hb897dc21),
	.w3(32'hb955cf16),
	.w4(32'hb98fff0c),
	.w5(32'hb9844d1a),
	.w6(32'hb906d8d5),
	.w7(32'hb920ccb8),
	.w8(32'hb7b97866),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e9069),
	.w1(32'hb95f19b7),
	.w2(32'hb98f3ac8),
	.w3(32'hb9b4d382),
	.w4(32'hb9c61fe5),
	.w5(32'hb9dc20b0),
	.w6(32'h3737dade),
	.w7(32'h392596cd),
	.w8(32'hb983316f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96821f8),
	.w1(32'hb967da9f),
	.w2(32'hb93b0aa8),
	.w3(32'hb9585c60),
	.w4(32'hb9908fae),
	.w5(32'hb93eaa0f),
	.w6(32'h39057fee),
	.w7(32'hb8c4085d),
	.w8(32'hb8adc191),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38819a28),
	.w1(32'hb6cd1e9f),
	.w2(32'hb864c3f0),
	.w3(32'hb7d70c95),
	.w4(32'hb8a328c3),
	.w5(32'hb8244223),
	.w6(32'hb912b3f1),
	.w7(32'hb91c1a4f),
	.w8(32'hb8974cdc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805f7d6),
	.w1(32'hb8aaa60e),
	.w2(32'hb8ac6271),
	.w3(32'h35827168),
	.w4(32'hb900587b),
	.w5(32'hb8f59d01),
	.w6(32'h384acded),
	.w7(32'hb832a758),
	.w8(32'hb83b6090),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37454199),
	.w1(32'hb582497b),
	.w2(32'hb7a9ee3d),
	.w3(32'h3605b3f5),
	.w4(32'hb6286c8a),
	.w5(32'hb77eeabe),
	.w6(32'h364bc884),
	.w7(32'hb72235a6),
	.w8(32'hb76caa07),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a8cccf),
	.w1(32'hb7a64a51),
	.w2(32'hb8576e75),
	.w3(32'h356e8bdc),
	.w4(32'hb56ade7d),
	.w5(32'h37447269),
	.w6(32'h369748cd),
	.w7(32'h3677fc96),
	.w8(32'hb79c987f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375bd08d),
	.w1(32'h37b87951),
	.w2(32'hb5121f9f),
	.w3(32'h37edb589),
	.w4(32'h37b70778),
	.w5(32'h370e75da),
	.w6(32'hb7047118),
	.w7(32'hb7906bd6),
	.w8(32'hb708481e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8433532),
	.w1(32'hb8cff732),
	.w2(32'hb85362b3),
	.w3(32'hb7b46203),
	.w4(32'hb8cf5090),
	.w5(32'hb8471d78),
	.w6(32'hb76ea289),
	.w7(32'hb89984b4),
	.w8(32'hb7e1409b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39734bb4),
	.w1(32'h39d8d860),
	.w2(32'hb7ffe741),
	.w3(32'h3937312b),
	.w4(32'hb887b7f2),
	.w5(32'h3925a446),
	.w6(32'hb9036371),
	.w7(32'h39380da7),
	.w8(32'h397c99e9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a110c52),
	.w1(32'h38fe491d),
	.w2(32'h3805de13),
	.w3(32'h399a19e8),
	.w4(32'h3878cb39),
	.w5(32'hb96cd09c),
	.w6(32'hb9b65883),
	.w7(32'hb7bfa0c0),
	.w8(32'hb9b8c9db),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66a3a37),
	.w1(32'h36e10342),
	.w2(32'hb604c1da),
	.w3(32'h36a3539d),
	.w4(32'h37f7f036),
	.w5(32'h3650cb9b),
	.w6(32'h36d5588f),
	.w7(32'h37993c0a),
	.w8(32'h37b44ed2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863944a),
	.w1(32'hb8900ae1),
	.w2(32'hb7f9fd79),
	.w3(32'hb792a563),
	.w4(32'h379c785b),
	.w5(32'hb5a77b37),
	.w6(32'h382d7951),
	.w7(32'hb883a5ed),
	.w8(32'hb856a68f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3634b05e),
	.w1(32'hb7134ddd),
	.w2(32'hb7a4cfc5),
	.w3(32'h368ca2da),
	.w4(32'hb6982a41),
	.w5(32'h38ad8c49),
	.w6(32'h3706adfe),
	.w7(32'hb63ebc8a),
	.w8(32'hb83d0067),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39224acf),
	.w1(32'h38620fb6),
	.w2(32'h37d99a8c),
	.w3(32'hb7ea6c5e),
	.w4(32'h38391a87),
	.w5(32'hb8956d12),
	.w6(32'hb91a8d34),
	.w7(32'hb88577d0),
	.w8(32'hb8839c06),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb764967a),
	.w1(32'h3824539d),
	.w2(32'h35d7f9ba),
	.w3(32'hb912b024),
	.w4(32'h39218be2),
	.w5(32'h38c3e923),
	.w6(32'h38bc975e),
	.w7(32'h39df9024),
	.w8(32'h398044e1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ea6e3),
	.w1(32'h39396257),
	.w2(32'h37e28ecb),
	.w3(32'h38a9c218),
	.w4(32'h38a35505),
	.w5(32'h37da6ac7),
	.w6(32'h38dc6254),
	.w7(32'h39038d4f),
	.w8(32'h388039d4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964bbde),
	.w1(32'h38d87421),
	.w2(32'h38b3ea79),
	.w3(32'h38961c3c),
	.w4(32'h36538ca2),
	.w5(32'hb6acb6db),
	.w6(32'hb7e31f82),
	.w7(32'hb7ac0a5c),
	.w8(32'hb7cd5324),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390fb695),
	.w1(32'h382b38b5),
	.w2(32'h38cebd58),
	.w3(32'hb89f301d),
	.w4(32'hb9800001),
	.w5(32'hb95a4182),
	.w6(32'hb88cdd47),
	.w7(32'hb8e3ff25),
	.w8(32'hb951440f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907d706),
	.w1(32'hb7015fb3),
	.w2(32'hb89fa0f5),
	.w3(32'hb831dcad),
	.w4(32'hb8bd1705),
	.w5(32'hb89f0afb),
	.w6(32'h3701493e),
	.w7(32'h37ea1a11),
	.w8(32'hb8eec093),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88de503),
	.w1(32'hb8885a42),
	.w2(32'h38b86ee7),
	.w3(32'h38504927),
	.w4(32'hb8fd6924),
	.w5(32'hb8996472),
	.w6(32'h3892c439),
	.w7(32'hb7bef18e),
	.w8(32'h380fb662),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39015558),
	.w1(32'h391298c4),
	.w2(32'hb8687ae4),
	.w3(32'hb9bec03d),
	.w4(32'hb9929026),
	.w5(32'hb9219587),
	.w6(32'hb94db048),
	.w7(32'hb8aa4e88),
	.w8(32'h35e51a9f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384de145),
	.w1(32'hb78782b0),
	.w2(32'hb72705af),
	.w3(32'hb8a63285),
	.w4(32'hb85a735c),
	.w5(32'hb82c921b),
	.w6(32'hb8b7b8fc),
	.w7(32'hb8281dee),
	.w8(32'hb6f2bcfa),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39907ab6),
	.w1(32'h369d8003),
	.w2(32'hb8ce9c8d),
	.w3(32'h380f99fb),
	.w4(32'hb9891045),
	.w5(32'hb932b38e),
	.w6(32'h37334d0c),
	.w7(32'hb7b9037b),
	.w8(32'hb8919f70),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f5bfe),
	.w1(32'hb95b6c63),
	.w2(32'hb954f294),
	.w3(32'hb98b25ba),
	.w4(32'hb9ce69aa),
	.w5(32'hb9976d81),
	.w6(32'hb920ce90),
	.w7(32'hb969a007),
	.w8(32'hb8ff5bac),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370274c1),
	.w1(32'hb78e17a4),
	.w2(32'h36fac421),
	.w3(32'hb79814b4),
	.w4(32'h373abc4f),
	.w5(32'h345885d9),
	.w6(32'hb7c48efb),
	.w7(32'h372fa2cd),
	.w8(32'h3734fd44),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bec23b),
	.w1(32'hb7781282),
	.w2(32'hb5b1c770),
	.w3(32'hb7a3eecd),
	.w4(32'hb61356dc),
	.w5(32'h37424557),
	.w6(32'hb74d0880),
	.w7(32'h365430c9),
	.w8(32'h3685a8bb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e2e713),
	.w1(32'h35a4bc48),
	.w2(32'h37dd94f5),
	.w3(32'hb49ef8f2),
	.w4(32'h382f7fd2),
	.w5(32'h381c2079),
	.w6(32'hb80de6c9),
	.w7(32'hb57a1114),
	.w8(32'hb818b818),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c31fb6),
	.w1(32'h39615f69),
	.w2(32'h39938057),
	.w3(32'h394618ae),
	.w4(32'h37789022),
	.w5(32'h38dcc907),
	.w6(32'h38ddf88d),
	.w7(32'h378dc1fa),
	.w8(32'hb8ab01ee),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db0fee),
	.w1(32'hb9837910),
	.w2(32'hb9a277d2),
	.w3(32'hb9733dbd),
	.w4(32'hb978a2e0),
	.w5(32'hb99be77f),
	.w6(32'hb929ae6c),
	.w7(32'hb9cb2db2),
	.w8(32'hba0641ab),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ee3fd5),
	.w1(32'hb74f2b79),
	.w2(32'h364f658c),
	.w3(32'hb7a51987),
	.w4(32'hb5b29d08),
	.w5(32'hb76db8ae),
	.w6(32'hb7cf939d),
	.w7(32'h36133cb7),
	.w8(32'hb68ce05d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ea8ec),
	.w1(32'h3904e0a2),
	.w2(32'hb73907af),
	.w3(32'hb9a6869d),
	.w4(32'hb9314ff8),
	.w5(32'hb941e0c2),
	.w6(32'hb88f0e6d),
	.w7(32'h38e03032),
	.w8(32'hb7976542),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe7f93),
	.w1(32'h39de2b58),
	.w2(32'h391daf9d),
	.w3(32'h39ed7ac5),
	.w4(32'h39b6e84a),
	.w5(32'h393ddee9),
	.w6(32'hb99ccdcb),
	.w7(32'h38d7ab7d),
	.w8(32'h3a1c4622),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934e600),
	.w1(32'h39548a36),
	.w2(32'h39136abb),
	.w3(32'h39c8bf6a),
	.w4(32'h397e8772),
	.w5(32'h3916b00e),
	.w6(32'h396745e3),
	.w7(32'h395f7be5),
	.w8(32'h398655ad),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885310e),
	.w1(32'h3780b688),
	.w2(32'hb9132cef),
	.w3(32'hb83df860),
	.w4(32'hb93ca27e),
	.w5(32'hb95621c3),
	.w6(32'h38def7a7),
	.w7(32'hb79f69a6),
	.w8(32'hb88623a7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae74cf),
	.w1(32'h376a8c7c),
	.w2(32'hb8daac2a),
	.w3(32'hb88f7e22),
	.w4(32'hb83972d9),
	.w5(32'hb859064c),
	.w6(32'h3849930a),
	.w7(32'h389054a7),
	.w8(32'h363ccad1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fa5eda),
	.w1(32'h37cb6c2d),
	.w2(32'h3761c9e7),
	.w3(32'h384f7e13),
	.w4(32'h384f8c22),
	.w5(32'h3890765e),
	.w6(32'h38ba6182),
	.w7(32'h3863b80e),
	.w8(32'h382b7cdc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3951ca30),
	.w1(32'h386c2535),
	.w2(32'h37d3bf48),
	.w3(32'hb91a0833),
	.w4(32'hb946aadd),
	.w5(32'hb8aa5884),
	.w6(32'hb983ad30),
	.w7(32'hb96e6f82),
	.w8(32'hb88a6311),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb720636a),
	.w1(32'hb8b5bf3e),
	.w2(32'hb7bdd4a1),
	.w3(32'h39a1b659),
	.w4(32'hb9169b7a),
	.w5(32'hb91924d1),
	.w6(32'h398ba01a),
	.w7(32'h39afafe5),
	.w8(32'h39d2327b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e6b1d),
	.w1(32'hb8d81afc),
	.w2(32'hb801f0ad),
	.w3(32'hb887bd93),
	.w4(32'hb8346187),
	.w5(32'h386c6840),
	.w6(32'h380e6af4),
	.w7(32'hb6ea7d02),
	.w8(32'hb80f889d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c276d),
	.w1(32'h385e2f0f),
	.w2(32'h385611e0),
	.w3(32'h3734bfbb),
	.w4(32'h381ba607),
	.w5(32'hb5c9db19),
	.w6(32'hb88185d0),
	.w7(32'hb796ff4d),
	.w8(32'h38143ada),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d143a5),
	.w1(32'hb841e6fe),
	.w2(32'hb7cee412),
	.w3(32'h351c4a11),
	.w4(32'hb6bc81ad),
	.w5(32'h3789b550),
	.w6(32'h37ca2e9c),
	.w7(32'h380a957c),
	.w8(32'hb81fee2f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39104074),
	.w1(32'h38d77a00),
	.w2(32'h37f42936),
	.w3(32'hb8267566),
	.w4(32'hb88e6710),
	.w5(32'hb8b57944),
	.w6(32'h397ea681),
	.w7(32'h38bfe2c3),
	.w8(32'hb639add2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb43616e4),
	.w1(32'hb7fbf83c),
	.w2(32'hb7708a9a),
	.w3(32'hb8147f34),
	.w4(32'h37a99257),
	.w5(32'hb5ab3e36),
	.w6(32'hb850093a),
	.w7(32'hb623203e),
	.w8(32'hb734ea3c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39214e82),
	.w1(32'h38053915),
	.w2(32'hb8ae5bba),
	.w3(32'hb8de4e2f),
	.w4(32'hb9a2875e),
	.w5(32'hb9016bfa),
	.w6(32'hb9692486),
	.w7(32'hb986de50),
	.w8(32'hb91cbea8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3732b233),
	.w1(32'hb835f471),
	.w2(32'hb6630a51),
	.w3(32'h381d7498),
	.w4(32'h385cd9a2),
	.w5(32'h3896d98f),
	.w6(32'h36385f89),
	.w7(32'h37532f63),
	.w8(32'h37799425),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c3648),
	.w1(32'hb7b88171),
	.w2(32'hb817b2f0),
	.w3(32'h38a666c5),
	.w4(32'h3910d0d5),
	.w5(32'h37b15b20),
	.w6(32'h39225662),
	.w7(32'h38a7c107),
	.w8(32'hb8154fe6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad90c1),
	.w1(32'h3837e2e8),
	.w2(32'h37091ffb),
	.w3(32'h380e64ef),
	.w4(32'h3619c438),
	.w5(32'hb6ef55bc),
	.w6(32'h35beacc3),
	.w7(32'hb8718fa8),
	.w8(32'hb8253f34),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3727472d),
	.w1(32'hb8268f9d),
	.w2(32'hb8277974),
	.w3(32'h380d475e),
	.w4(32'hb7598e58),
	.w5(32'h35453016),
	.w6(32'h38037ce7),
	.w7(32'hb817d809),
	.w8(32'hb783ee2e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a58335),
	.w1(32'hb94492a5),
	.w2(32'hb91845ae),
	.w3(32'hb9b32240),
	.w4(32'hba27be6c),
	.w5(32'hb9d51b70),
	.w6(32'h38ef547c),
	.w7(32'hb92d781d),
	.w8(32'hb99707d4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39736189),
	.w1(32'h3934e7f3),
	.w2(32'hb8262dbe),
	.w3(32'hb9661b65),
	.w4(32'hb974cdbb),
	.w5(32'hb9b0637b),
	.w6(32'hb8b8b9e5),
	.w7(32'h39ae5220),
	.w8(32'hb913cb99),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fd860),
	.w1(32'hb8d695af),
	.w2(32'h37790d71),
	.w3(32'hb73d85b0),
	.w4(32'hb7e8b97b),
	.w5(32'h38fdaa84),
	.w6(32'h390e58ba),
	.w7(32'hb64ec6fe),
	.w8(32'h38479e69),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e99df),
	.w1(32'h3925f854),
	.w2(32'h3994fe11),
	.w3(32'hb939b12b),
	.w4(32'hb8babacf),
	.w5(32'h39bcb5e3),
	.w6(32'hb9efa3ed),
	.w7(32'hb9712522),
	.w8(32'h3988cfab),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba05a3),
	.w1(32'h376df715),
	.w2(32'h379073cf),
	.w3(32'h387ddef4),
	.w4(32'h38b59d69),
	.w5(32'h35d69b8c),
	.w6(32'h375fcb79),
	.w7(32'h387ddd4b),
	.w8(32'h369512ea),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398173ac),
	.w1(32'h37a95eba),
	.w2(32'hb84fbbe6),
	.w3(32'h3901c789),
	.w4(32'hb99176e1),
	.w5(32'hb897fb6b),
	.w6(32'h3780a9b6),
	.w7(32'hb99836a3),
	.w8(32'h38de7852),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381836f8),
	.w1(32'hb6d01c48),
	.w2(32'hb78fd39d),
	.w3(32'hb70e4023),
	.w4(32'h37e106fe),
	.w5(32'h36720883),
	.w6(32'h3852cb01),
	.w7(32'h38cb0a45),
	.w8(32'h390420e2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913507e),
	.w1(32'h390849ff),
	.w2(32'h385e7692),
	.w3(32'hb993dbaa),
	.w4(32'hb8be644f),
	.w5(32'hb9837801),
	.w6(32'hb9e6b8b3),
	.w7(32'hb84225ae),
	.w8(32'h39263a92),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382aec65),
	.w1(32'h375ee6f5),
	.w2(32'h379c6077),
	.w3(32'hb79f648a),
	.w4(32'hb8b28fa3),
	.w5(32'hb8326013),
	.w6(32'h377e4439),
	.w7(32'hb8f6a1da),
	.w8(32'hb8f93c63),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39302cd9),
	.w1(32'hb89fdabd),
	.w2(32'hb8bb48de),
	.w3(32'hb8bc6634),
	.w4(32'hb9306ce5),
	.w5(32'hb8f940f4),
	.w6(32'hb7ba3da0),
	.w7(32'hb7f4d9cc),
	.w8(32'hb8b8dc08),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5bce706),
	.w1(32'h376a2a79),
	.w2(32'h367deb66),
	.w3(32'hb527fe2b),
	.w4(32'hb6e59baf),
	.w5(32'h389bdbc3),
	.w6(32'h37ad2ff7),
	.w7(32'h371c9066),
	.w8(32'h382f13d0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3834cc94),
	.w1(32'hb8c3d067),
	.w2(32'h379e8e7f),
	.w3(32'hb6a5e26c),
	.w4(32'h373a5d53),
	.w5(32'h3883f865),
	.w6(32'hb71d6e1d),
	.w7(32'hb8313131),
	.w8(32'h37b3f1b6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b1f59),
	.w1(32'hb78b900c),
	.w2(32'hb6200ba9),
	.w3(32'h3617c494),
	.w4(32'h37b03679),
	.w5(32'hb78db6bf),
	.w6(32'hb81f369b),
	.w7(32'hb74c4c5f),
	.w8(32'hb5341f9d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d7b235),
	.w1(32'hb8247f86),
	.w2(32'h37dba5a5),
	.w3(32'h3724eab6),
	.w4(32'hb69b63ee),
	.w5(32'hb855c190),
	.w6(32'h3891990b),
	.w7(32'hb757359c),
	.w8(32'hb7b946ce),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a0b24f),
	.w1(32'h3801cf7b),
	.w2(32'hb8356aad),
	.w3(32'h37cedaa9),
	.w4(32'hb81a46e3),
	.w5(32'hb7b92fdb),
	.w6(32'h387c62c9),
	.w7(32'hb83c718a),
	.w8(32'hb7374c25),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37db239b),
	.w1(32'hb61496d2),
	.w2(32'hb793af4e),
	.w3(32'hb7906c3d),
	.w4(32'h3796cbfb),
	.w5(32'h385fb6a4),
	.w6(32'hb66ae712),
	.w7(32'hb7bab945),
	.w8(32'h3740dc3a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386cbe0d),
	.w1(32'hb80c96e3),
	.w2(32'h379ac0e4),
	.w3(32'h369d5257),
	.w4(32'h388436d1),
	.w5(32'hb7112420),
	.w6(32'hb825edf3),
	.w7(32'h37cb7ec2),
	.w8(32'h363db347),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bffaba),
	.w1(32'hb80d1582),
	.w2(32'h381ee1e2),
	.w3(32'h384ead44),
	.w4(32'h38b0b2bc),
	.w5(32'h36da82e0),
	.w6(32'h3940ba08),
	.w7(32'h386dc3d9),
	.w8(32'h386396d4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8617caa),
	.w1(32'h37ffc429),
	.w2(32'h38d519dc),
	.w3(32'hb715986a),
	.w4(32'h387fdabf),
	.w5(32'h382540d8),
	.w6(32'hb79b6195),
	.w7(32'hb6d10764),
	.w8(32'h381656f7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937fbba),
	.w1(32'hb8f8f17f),
	.w2(32'hb8549d62),
	.w3(32'hb92007b9),
	.w4(32'hb8b1eed0),
	.w5(32'hb8afdeb8),
	.w6(32'hb8bd304d),
	.w7(32'hb742d251),
	.w8(32'hb78bbca5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791dbdd),
	.w1(32'hb99aa597),
	.w2(32'hba12e87d),
	.w3(32'hba1623a2),
	.w4(32'hb9ba4b65),
	.w5(32'hba127d07),
	.w6(32'hb9a5292f),
	.w7(32'h37addbba),
	.w8(32'hba0c01bb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88767d0),
	.w1(32'hb91729ea),
	.w2(32'hb85e2c0d),
	.w3(32'hb9e47fd1),
	.w4(32'hb9a6d973),
	.w5(32'hb98c83a7),
	.w6(32'hb9b9742f),
	.w7(32'hb9d92f16),
	.w8(32'hb9cba4e6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7247ede),
	.w1(32'h3719ecf7),
	.w2(32'h37809d8c),
	.w3(32'hb76ae85f),
	.w4(32'h382304ff),
	.w5(32'h38548809),
	.w6(32'hb782cb28),
	.w7(32'h36cdc339),
	.w8(32'hb847cd4f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374c51c3),
	.w1(32'h37a63d18),
	.w2(32'h37e9c040),
	.w3(32'h37a49e61),
	.w4(32'h37c10c6d),
	.w5(32'h37f13dbe),
	.w6(32'hb866b537),
	.w7(32'hb855eadc),
	.w8(32'h37c81e58),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7924212),
	.w1(32'hb865f9a0),
	.w2(32'hb74c38e4),
	.w3(32'hb8b01d99),
	.w4(32'hb86de1d1),
	.w5(32'hb7a52a08),
	.w6(32'hb8cf5178),
	.w7(32'hb8ac1724),
	.w8(32'hb7f7e419),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37949af9),
	.w1(32'hb80a2c60),
	.w2(32'h362b2097),
	.w3(32'hb8371401),
	.w4(32'hb67d2fa1),
	.w5(32'hb78d6c78),
	.w6(32'hb80f481a),
	.w7(32'h36b62be7),
	.w8(32'hb838b7b7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db3ddc),
	.w1(32'h38e1abaa),
	.w2(32'h3838bafd),
	.w3(32'h37837269),
	.w4(32'h36950817),
	.w5(32'h374122d4),
	.w6(32'hb8fc6ed0),
	.w7(32'hb8d0ea91),
	.w8(32'hb82d7aa8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c44d3),
	.w1(32'h381c2ab1),
	.w2(32'hb8d6ffbd),
	.w3(32'h397ceb2c),
	.w4(32'h3905edea),
	.w5(32'hb89fff6f),
	.w6(32'h38eb498c),
	.w7(32'h393bfd33),
	.w8(32'h376fc92d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b6670),
	.w1(32'hb9ded724),
	.w2(32'hb98bb80e),
	.w3(32'hb9a6c69d),
	.w4(32'hb9afa9a7),
	.w5(32'hb965b4e6),
	.w6(32'hb8f0e028),
	.w7(32'hb9807884),
	.w8(32'hb9388766),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bf845),
	.w1(32'hb762c0a6),
	.w2(32'hb7baed52),
	.w3(32'h376dc993),
	.w4(32'h374e6caf),
	.w5(32'hb83d4cc0),
	.w6(32'hb74e5037),
	.w7(32'h38aa6b1f),
	.w8(32'hb7aa2c8e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909c145),
	.w1(32'hb980a078),
	.w2(32'hb87375e5),
	.w3(32'hb9d6cfcc),
	.w4(32'hb9b8fea6),
	.w5(32'hb8da5f3e),
	.w6(32'hb966d32e),
	.w7(32'hb9c69877),
	.w8(32'hb5021a20),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842bac4),
	.w1(32'h37b8d661),
	.w2(32'h3787af18),
	.w3(32'h37f3e1d7),
	.w4(32'h3813b1b4),
	.w5(32'h380c8ce2),
	.w6(32'h38617d87),
	.w7(32'h36fe8a6b),
	.w8(32'h37accaef),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bfc943),
	.w1(32'hb78ba45e),
	.w2(32'h37009318),
	.w3(32'hb658a087),
	.w4(32'hb356d02e),
	.w5(32'hb507e1b8),
	.w6(32'hb790ff57),
	.w7(32'hb620e439),
	.w8(32'hb65eb13b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8320330),
	.w1(32'hb6d7dec5),
	.w2(32'h380f365a),
	.w3(32'hb82cae47),
	.w4(32'hb6032340),
	.w5(32'h389a7ef3),
	.w6(32'hb8040c43),
	.w7(32'hb6a286aa),
	.w8(32'h3831e71e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374af8ac),
	.w1(32'h373c8941),
	.w2(32'hb6efb6c0),
	.w3(32'h3577a3b3),
	.w4(32'h37971b57),
	.w5(32'h37689f79),
	.w6(32'hb7b581f2),
	.w7(32'hb7bc5e53),
	.w8(32'h374a8e9e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3864b796),
	.w1(32'hb86a4f3a),
	.w2(32'hb884dcdd),
	.w3(32'hb896a8e1),
	.w4(32'hb8862dcd),
	.w5(32'hb8d0f3bc),
	.w6(32'hb7f0cb34),
	.w7(32'hb8b2228c),
	.w8(32'hb81bd6fa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987b2ae),
	.w1(32'h39983333),
	.w2(32'h39461616),
	.w3(32'hb79a3a87),
	.w4(32'h39a3205a),
	.w5(32'h3951c076),
	.w6(32'hb91d5282),
	.w7(32'h394f8e87),
	.w8(32'h391c4dde),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b0545),
	.w1(32'hb678cd34),
	.w2(32'h389fe9d9),
	.w3(32'hb81558c2),
	.w4(32'hb8a29407),
	.w5(32'hb798597e),
	.w6(32'h37628a56),
	.w7(32'hb6d12415),
	.w8(32'h385edc56),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c63548),
	.w1(32'hb78cb19e),
	.w2(32'h39237c5e),
	.w3(32'h37ae6c75),
	.w4(32'h37d4b019),
	.w5(32'h38c263d6),
	.w6(32'h388ba666),
	.w7(32'h3737e5ba),
	.w8(32'h38456a2e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e74f6),
	.w1(32'h38cd299e),
	.w2(32'hb667a136),
	.w3(32'hb93efd9a),
	.w4(32'hb8823514),
	.w5(32'hb89f3811),
	.w6(32'hb8d21031),
	.w7(32'hb745e0c8),
	.w8(32'h37567cfa),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383b28e3),
	.w1(32'h3898127b),
	.w2(32'h37228a60),
	.w3(32'hb99d6fed),
	.w4(32'hb9855c6b),
	.w5(32'hb982e404),
	.w6(32'hb9e74a20),
	.w7(32'hb9aa663b),
	.w8(32'hb97da7e9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b54d47),
	.w1(32'h39b65818),
	.w2(32'hb841164a),
	.w3(32'hb9587f19),
	.w4(32'h39b81d1f),
	.w5(32'h38f8d848),
	.w6(32'hb9db6864),
	.w7(32'h39bd6132),
	.w8(32'h38582349),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372805ed),
	.w1(32'h3520622f),
	.w2(32'h36828445),
	.w3(32'h3701ac74),
	.w4(32'h37148e8d),
	.w5(32'hb5799a09),
	.w6(32'hb824d0c1),
	.w7(32'hb8027cba),
	.w8(32'hb60957e4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb642d629),
	.w1(32'hb8370e51),
	.w2(32'h377caa7e),
	.w3(32'hb855ad15),
	.w4(32'hb7026e86),
	.w5(32'hb7d72205),
	.w6(32'hb8781802),
	.w7(32'hb714a1f1),
	.w8(32'hb7327ecb),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fb83e),
	.w1(32'h3891cfa0),
	.w2(32'hb4a41626),
	.w3(32'h385a01c8),
	.w4(32'h38b228c6),
	.w5(32'h38249b9b),
	.w6(32'h395b4644),
	.w7(32'h3915b2fc),
	.w8(32'h388e3ea7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c379e),
	.w1(32'h3a10021c),
	.w2(32'h3992a1ea),
	.w3(32'hb73cede0),
	.w4(32'h370fc380),
	.w5(32'h3904ba4a),
	.w6(32'h38c3155c),
	.w7(32'h3a25432f),
	.w8(32'h399c0ea6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d7992),
	.w1(32'hb8e0ff70),
	.w2(32'hb90cf121),
	.w3(32'hb9916165),
	.w4(32'hb932f851),
	.w5(32'hb976b32d),
	.w6(32'hb95f4ea5),
	.w7(32'hb8d96a56),
	.w8(32'hb94c37d3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eaef3c),
	.w1(32'h38aaf1c4),
	.w2(32'h37453225),
	.w3(32'h38ed258e),
	.w4(32'h38e11116),
	.w5(32'h38896d3a),
	.w6(32'h37c8cdf1),
	.w7(32'hb6acca12),
	.w8(32'hb81df9a7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aebd2d),
	.w1(32'h3801979c),
	.w2(32'h37bf7b2e),
	.w3(32'h3792aa60),
	.w4(32'h3705e6c6),
	.w5(32'hb5fd3c96),
	.w6(32'hb7e2295b),
	.w7(32'hb80b249d),
	.w8(32'hb7a0a746),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d373d),
	.w1(32'h39257f25),
	.w2(32'h393c5526),
	.w3(32'h369f0111),
	.w4(32'h3936ed2c),
	.w5(32'h3936c6fd),
	.w6(32'hb74b7f90),
	.w7(32'h380a337d),
	.w8(32'h38912ab2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f11896),
	.w1(32'h37a0b489),
	.w2(32'h37f66d94),
	.w3(32'hb819cca7),
	.w4(32'h384b59b4),
	.w5(32'h38c60201),
	.w6(32'hb90d1d08),
	.w7(32'h380736b8),
	.w8(32'h38599326),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c5ca4),
	.w1(32'h395524a7),
	.w2(32'hb8ba8976),
	.w3(32'h3937ebf2),
	.w4(32'hb6af7282),
	.w5(32'hb88d29b0),
	.w6(32'h3887608d),
	.w7(32'h386900da),
	.w8(32'hb822d56e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872aa76),
	.w1(32'h37d86b5b),
	.w2(32'h38404f86),
	.w3(32'hb8720eea),
	.w4(32'h38aacfd0),
	.w5(32'h38944d27),
	.w6(32'hb8ca8e07),
	.w7(32'h3802b5fc),
	.w8(32'h38429aa3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3743c621),
	.w1(32'hb8b8cb8a),
	.w2(32'h375e0eaf),
	.w3(32'hb7874548),
	.w4(32'h3712583d),
	.w5(32'h386e76d9),
	.w6(32'h38a7d946),
	.w7(32'h3900aaf1),
	.w8(32'h38b7952c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974d14d),
	.w1(32'hb8fd8582),
	.w2(32'hb8b048df),
	.w3(32'hb9251003),
	.w4(32'hb9641f97),
	.w5(32'hb945957d),
	.w6(32'hb9426375),
	.w7(32'hb9138494),
	.w8(32'hb8b35f07),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375b879a),
	.w1(32'h35feba37),
	.w2(32'h36fdd700),
	.w3(32'hb73f69bf),
	.w4(32'hb6ae2f4a),
	.w5(32'hb706f7e4),
	.w6(32'hb709e4fb),
	.w7(32'hb624249a),
	.w8(32'h358f54ed),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74d5719),
	.w1(32'hb7eaf1b0),
	.w2(32'hb7ec7f45),
	.w3(32'h37ac4a43),
	.w4(32'h36f243c2),
	.w5(32'hb7c1ebc3),
	.w6(32'h36c01357),
	.w7(32'hb5f1d105),
	.w8(32'hb7ac2b58),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3581c86d),
	.w1(32'h37815b6b),
	.w2(32'h36bc58d2),
	.w3(32'h379ecd3b),
	.w4(32'h37b1b153),
	.w5(32'h37d06868),
	.w6(32'h35c747f7),
	.w7(32'hb70c07e7),
	.w8(32'hb7c186f3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e7d3b3),
	.w1(32'hb78f9cd7),
	.w2(32'h385e9c0d),
	.w3(32'hb8477a65),
	.w4(32'h37d561f1),
	.w5(32'hb9f5323d),
	.w6(32'hb88337ea),
	.w7(32'h381a14c9),
	.w8(32'hba6d638e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d1160),
	.w1(32'hbac56114),
	.w2(32'hb9c3e6a5),
	.w3(32'hba97f20c),
	.w4(32'hb98c97d7),
	.w5(32'hba848ac1),
	.w6(32'hbafdbba7),
	.w7(32'hba330081),
	.w8(32'hba23b385),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06d968),
	.w1(32'hb97ef109),
	.w2(32'h3a132820),
	.w3(32'hb962920f),
	.w4(32'h393c1a59),
	.w5(32'h38d44c95),
	.w6(32'hba913bf1),
	.w7(32'h39c21785),
	.w8(32'hba301e1b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a265e7),
	.w1(32'hba053cb5),
	.w2(32'hba3b0dba),
	.w3(32'hb90aa25c),
	.w4(32'hb825f18e),
	.w5(32'hb91ff9ff),
	.w6(32'hba8a0a78),
	.w7(32'hba946821),
	.w8(32'hba5bdadd),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3817281b),
	.w1(32'h3986a3e9),
	.w2(32'h39bf0b16),
	.w3(32'hb9b2c1bd),
	.w4(32'hb9f808d2),
	.w5(32'h39d8b6b2),
	.w6(32'hba113711),
	.w7(32'hb8877cf4),
	.w8(32'h38ff20c9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dfbc6),
	.w1(32'h3919c7ef),
	.w2(32'h3a360ad0),
	.w3(32'hb7bf8ea4),
	.w4(32'h3a3cc45b),
	.w5(32'hba6147c2),
	.w6(32'hb95a5e11),
	.w7(32'h39efa174),
	.w8(32'hba9902c6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba487c15),
	.w1(32'hb9dd3e60),
	.w2(32'hbaa74fa6),
	.w3(32'hba74d52f),
	.w4(32'hbaabc455),
	.w5(32'hba23f918),
	.w6(32'hbac26e81),
	.w7(32'hba937f9b),
	.w8(32'hb9fd5158),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31fcb2),
	.w1(32'hbad12ce1),
	.w2(32'hbac1a613),
	.w3(32'hb9fe1f30),
	.w4(32'hba90f662),
	.w5(32'h3a0cbab7),
	.w6(32'hba24642b),
	.w7(32'hba9b1d06),
	.w8(32'h39a3f071),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398853aa),
	.w1(32'hb9954634),
	.w2(32'h394ddfc6),
	.w3(32'hb90097bd),
	.w4(32'h39f48bbb),
	.w5(32'hba6fe21d),
	.w6(32'hb9611c60),
	.w7(32'hb881834d),
	.w8(32'hb96db4e5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30e0f9),
	.w1(32'hb9834529),
	.w2(32'hbaf542ba),
	.w3(32'hbacaa4e9),
	.w4(32'hbaed601d),
	.w5(32'hb87aca32),
	.w6(32'hba8fe4cf),
	.w7(32'hbb007ea1),
	.w8(32'hba45d14e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b9bc8),
	.w1(32'hb9ccc6eb),
	.w2(32'h3a2f51ee),
	.w3(32'h37ee12ac),
	.w4(32'h3a4efd14),
	.w5(32'hbaa3e349),
	.w6(32'hba0fb68c),
	.w7(32'h3a16d236),
	.w8(32'hbaeb6ba6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee63d7),
	.w1(32'hbb23d951),
	.w2(32'hbac061f4),
	.w3(32'hbaeede85),
	.w4(32'hba868203),
	.w5(32'h3a303b78),
	.w6(32'hbb32d65a),
	.w7(32'hbadefc5f),
	.w8(32'h3a0bed1a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b849f),
	.w1(32'h38d43396),
	.w2(32'h3ab31e9d),
	.w3(32'h388b6144),
	.w4(32'h3ad24756),
	.w5(32'hb94b6c33),
	.w6(32'hb889fcb2),
	.w7(32'h3a98744d),
	.w8(32'hb8f504a2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d34db),
	.w1(32'hb85d4aa3),
	.w2(32'h3989bdd8),
	.w3(32'hb98f4fb9),
	.w4(32'h3a7dea3c),
	.w5(32'hba34218d),
	.w6(32'hb62f2673),
	.w7(32'h3a6fbb50),
	.w8(32'hb9c69123),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6de25),
	.w1(32'h3964a045),
	.w2(32'hb935b708),
	.w3(32'hba442393),
	.w4(32'hba2fda22),
	.w5(32'h3a1fe0f6),
	.w6(32'hba061ed8),
	.w7(32'hb9f61d48),
	.w8(32'h3a0f1a94),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9888a4),
	.w1(32'h39bd4953),
	.w2(32'h3ab41c7b),
	.w3(32'h3a3088be),
	.w4(32'h3b058996),
	.w5(32'h3a75fc84),
	.w6(32'h39aa733b),
	.w7(32'h3aa6c3eb),
	.w8(32'h3a7ef4d2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de02c5),
	.w1(32'h39b568dd),
	.w2(32'h3936aafd),
	.w3(32'h3a165711),
	.w4(32'h393346f0),
	.w5(32'hbb158e04),
	.w6(32'h3970a378),
	.w7(32'h3a4f317b),
	.w8(32'hbb040cb1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135ec7),
	.w1(32'hbaf74d95),
	.w2(32'h3a5b5f5f),
	.w3(32'hba795932),
	.w4(32'hb9f4d712),
	.w5(32'hb9fa6dfc),
	.w6(32'hba799863),
	.w7(32'h396d35a4),
	.w8(32'hba5a660d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2272e),
	.w1(32'h39cf6170),
	.w2(32'h39e08f74),
	.w3(32'hb9b16cf3),
	.w4(32'h392f780c),
	.w5(32'h3a84a75b),
	.w6(32'hb993eea2),
	.w7(32'h39e1a4be),
	.w8(32'h3a8d9efd),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadba68),
	.w1(32'h3a971708),
	.w2(32'h3a633ce7),
	.w3(32'h3a282ae9),
	.w4(32'h3a6546fd),
	.w5(32'hb9eea5fa),
	.w6(32'h3a254af0),
	.w7(32'h3a3dd465),
	.w8(32'h3a502ff3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06363b),
	.w1(32'hba7a2514),
	.w2(32'hbac0c7d1),
	.w3(32'hba611e73),
	.w4(32'hbaf61aca),
	.w5(32'hb7c5ea9e),
	.w6(32'hba0ee8de),
	.w7(32'hba05822c),
	.w8(32'hba18a480),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aee54),
	.w1(32'hbb0040c0),
	.w2(32'hb91dd726),
	.w3(32'hbab47b1e),
	.w4(32'h3916c663),
	.w5(32'hb9a4d840),
	.w6(32'hbb0ec53f),
	.w7(32'hb97026f4),
	.w8(32'hbaa24db5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba226d55),
	.w1(32'hbaa60e79),
	.w2(32'hba755212),
	.w3(32'hba8d772a),
	.w4(32'hba51d303),
	.w5(32'h39de4b47),
	.w6(32'hbb14374a),
	.w7(32'hbaf0de52),
	.w8(32'h39b4151c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ac885),
	.w1(32'h39dee42c),
	.w2(32'h3a3ab4d2),
	.w3(32'h3a4f59b1),
	.w4(32'h39b98fb7),
	.w5(32'hba3a863c),
	.w6(32'hb838084c),
	.w7(32'h3a179dfe),
	.w8(32'hba7f9f05),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc54b),
	.w1(32'hbaae3027),
	.w2(32'hb7a62752),
	.w3(32'hba58c5c9),
	.w4(32'h37961464),
	.w5(32'hb93a5458),
	.w6(32'hb9d4c017),
	.w7(32'hb9a7bba7),
	.w8(32'hb8f762f4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e997c),
	.w1(32'hb7f18912),
	.w2(32'h380f85c6),
	.w3(32'hb993d1fb),
	.w4(32'h394a7669),
	.w5(32'h3a2c32bc),
	.w6(32'hb991556d),
	.w7(32'hb9db8e2b),
	.w8(32'h38e09b89),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39890468),
	.w1(32'h3a86322c),
	.w2(32'h3a376318),
	.w3(32'h3a38eedb),
	.w4(32'h3a807e07),
	.w5(32'h398070f1),
	.w6(32'h3a97f833),
	.w7(32'h39d32219),
	.w8(32'hb8eb8858),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38906363),
	.w1(32'h3848bda6),
	.w2(32'h3940044f),
	.w3(32'hb8fb9651),
	.w4(32'h39a20f38),
	.w5(32'h398c8a5a),
	.w6(32'hb993a78b),
	.w7(32'hb973cf5a),
	.w8(32'h398a47ef),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25b7d1),
	.w1(32'h3a16642d),
	.w2(32'h39a7f8c8),
	.w3(32'h3947e386),
	.w4(32'hb9900fe6),
	.w5(32'h3a3ab2e5),
	.w6(32'h38b2ae12),
	.w7(32'h38ff6359),
	.w8(32'h3a1ce482),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09f8c9),
	.w1(32'h39a707f6),
	.w2(32'h39cb603d),
	.w3(32'h38d7b149),
	.w4(32'h3a382911),
	.w5(32'h39ea89a8),
	.w6(32'h3950a24a),
	.w7(32'h3a1fe3d5),
	.w8(32'h39fcd6fa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e51a99),
	.w1(32'h3a653406),
	.w2(32'h3a802b34),
	.w3(32'h3a88193e),
	.w4(32'h3a3573fe),
	.w5(32'h3aa2bc6e),
	.w6(32'h3af50004),
	.w7(32'h3a8d2969),
	.w8(32'h3a5b6ace),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule