module layer_10_featuremap_405(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47e744),
	.w1(32'hbb0a9f3e),
	.w2(32'hba5309da),
	.w3(32'h3b91eed4),
	.w4(32'hba9025b9),
	.w5(32'h3a8b7780),
	.w6(32'h3b89b402),
	.w7(32'hbb41d10a),
	.w8(32'hba82a019),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980be05),
	.w1(32'hb9149c25),
	.w2(32'hbbb2ee47),
	.w3(32'h3a247689),
	.w4(32'h3baae1de),
	.w5(32'h3bbc6e33),
	.w6(32'hbb73dd61),
	.w7(32'hbb92b96d),
	.w8(32'h3a7929b0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb5fb4),
	.w1(32'hba8c7ef5),
	.w2(32'hbb815a74),
	.w3(32'h3a9aabfc),
	.w4(32'h3b88a0a7),
	.w5(32'hbbd51501),
	.w6(32'h3b88404e),
	.w7(32'h3c0f483d),
	.w8(32'h3bc0a0d1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2bd0f),
	.w1(32'hbbe67566),
	.w2(32'hb8c4e37c),
	.w3(32'hbb0cf45e),
	.w4(32'hbc13a9f3),
	.w5(32'h3b48f4e3),
	.w6(32'h3a9daf7e),
	.w7(32'hbbff5147),
	.w8(32'h3b304470),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6807c),
	.w1(32'hba9a84f3),
	.w2(32'hb9af893a),
	.w3(32'h3b39028f),
	.w4(32'hbb8e45a8),
	.w5(32'hbb7639d4),
	.w6(32'h3b01afb6),
	.w7(32'h3ad99f9d),
	.w8(32'h3919042c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6aec1),
	.w1(32'h3b118460),
	.w2(32'hbaac0387),
	.w3(32'hbaaf8649),
	.w4(32'h3a63aa99),
	.w5(32'hbb8cfc6f),
	.w6(32'hbb3d1def),
	.w7(32'hba304541),
	.w8(32'hbb3a2d5e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1848cc),
	.w1(32'hbb58487d),
	.w2(32'h39e0797f),
	.w3(32'hbb2eeb1d),
	.w4(32'h3ba46069),
	.w5(32'h3b731ca7),
	.w6(32'hbc0fbdfb),
	.w7(32'hbb588b45),
	.w8(32'hbb0303b3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58a32),
	.w1(32'h3bc400c8),
	.w2(32'h3c23f756),
	.w3(32'hbbd9cab2),
	.w4(32'h3aad2d6d),
	.w5(32'hbb7d84f4),
	.w6(32'h3d1a54a7),
	.w7(32'h3ce6aa1b),
	.w8(32'h3ab7378b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb533e29),
	.w1(32'hbb8a81a0),
	.w2(32'hbb487391),
	.w3(32'hbbe8c92e),
	.w4(32'hbb916fe1),
	.w5(32'hbabeb087),
	.w6(32'h3ad44fb8),
	.w7(32'h3a012b5b),
	.w8(32'h3a578f94),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccf487),
	.w1(32'hbb411539),
	.w2(32'h3b509df8),
	.w3(32'hbb580999),
	.w4(32'hbb3b822b),
	.w5(32'h3aadfc09),
	.w6(32'hba3208e5),
	.w7(32'h3a01a90a),
	.w8(32'hbac51b1a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b501062),
	.w1(32'h3b7ecd9f),
	.w2(32'h3bccdd73),
	.w3(32'hbb14929a),
	.w4(32'h3a998c39),
	.w5(32'h3bb66e48),
	.w6(32'hbba9e45d),
	.w7(32'h3b87effc),
	.w8(32'h3ba9e033),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9855),
	.w1(32'hbbdf8dd8),
	.w2(32'hb8b452c9),
	.w3(32'h3b7773b4),
	.w4(32'hbc4adc90),
	.w5(32'h3a451477),
	.w6(32'h3be4925f),
	.w7(32'hbaa0aa3e),
	.w8(32'hbb8dbab5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0f687),
	.w1(32'hbbd1e7b1),
	.w2(32'hbc28d201),
	.w3(32'h3b5715a7),
	.w4(32'hbbef82ae),
	.w5(32'hbb29729f),
	.w6(32'h3b71958a),
	.w7(32'hbaac60fe),
	.w8(32'hba8994fa),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacb4ac),
	.w1(32'hbb04f5f7),
	.w2(32'h3bdc65b5),
	.w3(32'hbc5adea3),
	.w4(32'hbbcf55f0),
	.w5(32'hbaccacfe),
	.w6(32'hbb44163e),
	.w7(32'hbb438b1b),
	.w8(32'hbb046823),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e85314),
	.w1(32'hba30ae59),
	.w2(32'h3a3a4319),
	.w3(32'h3bb4d607),
	.w4(32'hbad9cdd8),
	.w5(32'h3b1a6b53),
	.w6(32'h39ba621d),
	.w7(32'hbb7c43ae),
	.w8(32'hbb1d4fd7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab713ac),
	.w1(32'hb942b9ba),
	.w2(32'hbbcf718e),
	.w3(32'hbb38743b),
	.w4(32'h39dafacb),
	.w5(32'h3a1ba068),
	.w6(32'hbb7c572d),
	.w7(32'hbbc3a6bd),
	.w8(32'hbbc17ec4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7e07),
	.w1(32'h3b003638),
	.w2(32'h3348e14e),
	.w3(32'hbbb7f079),
	.w4(32'h3a55f5b2),
	.w5(32'h3b828a59),
	.w6(32'h39f831ed),
	.w7(32'hbb99cc7e),
	.w8(32'hbb900d6b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45731f),
	.w1(32'h3a2eec1d),
	.w2(32'hbb33605f),
	.w3(32'h3ae0ba87),
	.w4(32'hbb9dba88),
	.w5(32'hbabf30fc),
	.w6(32'h3c6ac828),
	.w7(32'h3c3afb62),
	.w8(32'h3bcc6fba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64cd82),
	.w1(32'h3b42f854),
	.w2(32'h3b4d4a75),
	.w3(32'h3b7c21d6),
	.w4(32'hbb9130e1),
	.w5(32'h3a983efe),
	.w6(32'h3c3ae569),
	.w7(32'h3b864f78),
	.w8(32'h3665cbce),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a716a91),
	.w1(32'hbb0c8516),
	.w2(32'h3b25abd7),
	.w3(32'h3b6b7d03),
	.w4(32'hbb48e0e9),
	.w5(32'h3bef04dc),
	.w6(32'h396519b1),
	.w7(32'hbbe31398),
	.w8(32'hb9c47886),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dfe3e),
	.w1(32'h3ac9d678),
	.w2(32'hba341b7a),
	.w3(32'hbb8b7fb2),
	.w4(32'hbb8c5716),
	.w5(32'hbb634aec),
	.w6(32'hbb546db8),
	.w7(32'hba6c556f),
	.w8(32'hbba3d419),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c26c17),
	.w1(32'h3abd70a1),
	.w2(32'hbb5b09e0),
	.w3(32'hb9a3de0e),
	.w4(32'hba38eae8),
	.w5(32'h3ae171f1),
	.w6(32'hbbadecbd),
	.w7(32'hbbdda493),
	.w8(32'h3b95b98c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cbf70),
	.w1(32'hb9e61e77),
	.w2(32'hbb35258a),
	.w3(32'hbaaddf2c),
	.w4(32'h3bcd0bb7),
	.w5(32'hbb8b45a3),
	.w6(32'h3ae94460),
	.w7(32'h3b8e5d2a),
	.w8(32'h3c353331),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fed8d9),
	.w1(32'h3b221684),
	.w2(32'h3a832a5b),
	.w3(32'h3b53bbfb),
	.w4(32'h3aac74b8),
	.w5(32'h3b93e467),
	.w6(32'hbb2cd4f8),
	.w7(32'hba9618e9),
	.w8(32'h3a4301e0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a317cd8),
	.w1(32'h3b21b538),
	.w2(32'h3bc8f485),
	.w3(32'hbad55951),
	.w4(32'h3be24921),
	.w5(32'h3b9df0b0),
	.w6(32'hbc32b210),
	.w7(32'hbb62381e),
	.w8(32'h3b9ee4a9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c23cc),
	.w1(32'h3b50bff3),
	.w2(32'hb9a64cae),
	.w3(32'h3a8920af),
	.w4(32'h3abf4d20),
	.w5(32'hbb493623),
	.w6(32'h3ba675e2),
	.w7(32'hb9c92087),
	.w8(32'h3b62f671),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3bafa),
	.w1(32'hbb1ffcae),
	.w2(32'hbb14ca5b),
	.w3(32'h3ab04211),
	.w4(32'hb8f516d2),
	.w5(32'hbbff594b),
	.w6(32'h3b35c250),
	.w7(32'h3b436e9d),
	.w8(32'hbae526e8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1365c),
	.w1(32'hba99b0a4),
	.w2(32'hbc7333eb),
	.w3(32'hbb79a159),
	.w4(32'h3c07546f),
	.w5(32'h3b2010f8),
	.w6(32'hbc2fafca),
	.w7(32'hbc2026ca),
	.w8(32'hbbaf8a15),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51d61f),
	.w1(32'hba488d0a),
	.w2(32'hbb33f98f),
	.w3(32'hb83d5015),
	.w4(32'h3b2e252c),
	.w5(32'h39dbae61),
	.w6(32'h3aee41bb),
	.w7(32'hbad7dd0b),
	.w8(32'hbb4ae605),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18d564),
	.w1(32'h3bcbc54e),
	.w2(32'h3b28abf0),
	.w3(32'hbbb29dec),
	.w4(32'hbac6e100),
	.w5(32'h3ba47e8e),
	.w6(32'hbc6744f3),
	.w7(32'hbc48da11),
	.w8(32'hbc33cf32),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d2e6c),
	.w1(32'hbb7e9785),
	.w2(32'hba2c3079),
	.w3(32'hb81e2064),
	.w4(32'h3be0e03a),
	.w5(32'h3c4ff5c4),
	.w6(32'hbbbbd25c),
	.w7(32'hbbbe5c7e),
	.w8(32'hbb3265fc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43290d),
	.w1(32'hbb01fac1),
	.w2(32'hbacc71be),
	.w3(32'h3c1599fd),
	.w4(32'h3bc7357f),
	.w5(32'h3bb8acf0),
	.w6(32'h3b7e19f6),
	.w7(32'h3b404141),
	.w8(32'h3a35b30c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd4975),
	.w1(32'h3b09f65a),
	.w2(32'h39db7f8f),
	.w3(32'hba845fa8),
	.w4(32'h3c0d4451),
	.w5(32'h3baf7415),
	.w6(32'h3bcd182b),
	.w7(32'h3b92e01e),
	.w8(32'h3c51e519),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed4b9c),
	.w1(32'h3a9302a1),
	.w2(32'h3b11a76d),
	.w3(32'hbb448861),
	.w4(32'h3ba3527a),
	.w5(32'hba6447bc),
	.w6(32'h3ba4de10),
	.w7(32'hb9fcc6dc),
	.w8(32'h3b392c73),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02fceb),
	.w1(32'hbb72eecc),
	.w2(32'h3abd96e1),
	.w3(32'hbaa37eb1),
	.w4(32'hbb728eb9),
	.w5(32'hbb2434b0),
	.w6(32'h3bfe8692),
	.w7(32'h3b20a194),
	.w8(32'hbbc6dd65),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af67ff4),
	.w1(32'hbb7cfa14),
	.w2(32'h3a8ddd60),
	.w3(32'h3af6ee72),
	.w4(32'hbbcbb7b3),
	.w5(32'h3b092408),
	.w6(32'h3b07d274),
	.w7(32'h3add6d5d),
	.w8(32'h3bb436a3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba894828),
	.w1(32'hbb906a52),
	.w2(32'h3c0acbd5),
	.w3(32'h3b335bff),
	.w4(32'hbc4550a7),
	.w5(32'h3b80234b),
	.w6(32'h3bc36efd),
	.w7(32'hbc109d15),
	.w8(32'hb8b7aacc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d698),
	.w1(32'hba333f82),
	.w2(32'hbbbfaf3e),
	.w3(32'h3b8423ff),
	.w4(32'h3c58d078),
	.w5(32'h3c9549d1),
	.w6(32'h3ad115a2),
	.w7(32'hbc648659),
	.w8(32'h3a3c5133),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1afa47),
	.w1(32'hba1ca3ba),
	.w2(32'h3c11a371),
	.w3(32'hbab05c34),
	.w4(32'hbbe1ab90),
	.w5(32'hbb93f59c),
	.w6(32'hbc3b1781),
	.w7(32'hbc0ac095),
	.w8(32'hbbd4584e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3216f2),
	.w1(32'hbb4217f8),
	.w2(32'hbb877c2b),
	.w3(32'h38ebb28a),
	.w4(32'h3b9916a5),
	.w5(32'h3c329486),
	.w6(32'hbbd2dc7c),
	.w7(32'hbaf47033),
	.w8(32'h3be336e3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a946116),
	.w1(32'hbb0e4c2f),
	.w2(32'hb9cef8f0),
	.w3(32'h3ac498c3),
	.w4(32'hbb0f6c62),
	.w5(32'h3a00df33),
	.w6(32'h3b4a2f3e),
	.w7(32'h3b830a56),
	.w8(32'h3b42c590),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fffa0),
	.w1(32'h3a807a58),
	.w2(32'h3b2a3375),
	.w3(32'h36397b10),
	.w4(32'hbb1b3b70),
	.w5(32'hbba3bc63),
	.w6(32'hbb087281),
	.w7(32'h3a539e07),
	.w8(32'h3b070a76),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0844),
	.w1(32'hbb795ccd),
	.w2(32'hbba6d131),
	.w3(32'hba995a8f),
	.w4(32'hbb437e7d),
	.w5(32'hbaf97667),
	.w6(32'hbaf25a4d),
	.w7(32'hbbb79e52),
	.w8(32'hbb738ce5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb169d7e),
	.w1(32'hba73d849),
	.w2(32'hbbf12200),
	.w3(32'hbb9e271a),
	.w4(32'hbb9d738d),
	.w5(32'hbb70feb5),
	.w6(32'h3af9e4fa),
	.w7(32'hbb512071),
	.w8(32'h3b403b9c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf2b6e),
	.w1(32'h3b5070a0),
	.w2(32'h3901f363),
	.w3(32'h3ad4b26a),
	.w4(32'hbb1c72da),
	.w5(32'hbb98b305),
	.w6(32'h39ccd315),
	.w7(32'hbb4ab225),
	.w8(32'h3a5ee58e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b156ea5),
	.w1(32'hbb671d35),
	.w2(32'h3bdc96ea),
	.w3(32'h3b420731),
	.w4(32'hbb09f18f),
	.w5(32'hbb101bed),
	.w6(32'h3adfdd8f),
	.w7(32'h3acd9b49),
	.w8(32'h3b0699a6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee909b),
	.w1(32'h3af230bf),
	.w2(32'h3c075bd2),
	.w3(32'hbb8b0c5f),
	.w4(32'hbbbd2603),
	.w5(32'hbabe7aeb),
	.w6(32'h3a0f7b0d),
	.w7(32'hbb880967),
	.w8(32'hbbd1319a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dfdae),
	.w1(32'hbb5103be),
	.w2(32'hbba2681e),
	.w3(32'hbb1b8b5f),
	.w4(32'hbbf4a2ae),
	.w5(32'hbb427f9d),
	.w6(32'h3c41dbee),
	.w7(32'h3c1445a8),
	.w8(32'h3bf3423b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040875),
	.w1(32'h3b8a8768),
	.w2(32'h3ba582e3),
	.w3(32'hbba70fe4),
	.w4(32'hbb8c12e3),
	.w5(32'hbafd45bd),
	.w6(32'hbb8fcc0b),
	.w7(32'h3b605cc8),
	.w8(32'h38d2f3e2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06d8db),
	.w1(32'h3b92c41b),
	.w2(32'h3b8a5537),
	.w3(32'hbaa85870),
	.w4(32'h3bec9071),
	.w5(32'h3b85ae60),
	.w6(32'hbc07f858),
	.w7(32'h3be8a866),
	.w8(32'h3b161afd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87c88),
	.w1(32'h3b51b3c0),
	.w2(32'h3b592d28),
	.w3(32'h3b839087),
	.w4(32'h3a8582cf),
	.w5(32'hba6ebcf7),
	.w6(32'h3a8a6c41),
	.w7(32'hb9c74c32),
	.w8(32'h39ef5b4d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989f779),
	.w1(32'hb8b7cc99),
	.w2(32'hbaf9a0c4),
	.w3(32'h3b64c572),
	.w4(32'h3b42837d),
	.w5(32'h39fe7195),
	.w6(32'hbb6d85c5),
	.w7(32'hbb0bc340),
	.w8(32'h3b5087d2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86197),
	.w1(32'h3b6a0214),
	.w2(32'h3ab59b82),
	.w3(32'hbadfb93e),
	.w4(32'h3b698873),
	.w5(32'h395e2db3),
	.w6(32'h399f34a6),
	.w7(32'h3b290e0f),
	.w8(32'hba33dad8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91600d),
	.w1(32'hbb74dba8),
	.w2(32'hbc1f749d),
	.w3(32'hbc49a4df),
	.w4(32'hba0fe298),
	.w5(32'hba93e6f7),
	.w6(32'h3c690827),
	.w7(32'h3bf037b2),
	.w8(32'h3ae9740b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3308f),
	.w1(32'hbbb4a3ad),
	.w2(32'hbc1b8b3e),
	.w3(32'hbbb99621),
	.w4(32'h3b6c1a30),
	.w5(32'h3bfd0e3c),
	.w6(32'h3ba8ab71),
	.w7(32'hba84f0ba),
	.w8(32'h3af40315),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9feb0),
	.w1(32'hbbb344fd),
	.w2(32'hbc381990),
	.w3(32'hbb77d1d5),
	.w4(32'h3c12e45a),
	.w5(32'h3c26d916),
	.w6(32'h3a8e6a16),
	.w7(32'hbb6f7839),
	.w8(32'h3bc2889a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0a1dc),
	.w1(32'hba3b897a),
	.w2(32'hb888dad0),
	.w3(32'hbb919075),
	.w4(32'hbba114d8),
	.w5(32'h3aefb3b8),
	.w6(32'h3a8c9d54),
	.w7(32'hbb7db299),
	.w8(32'hbafe78df),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad45569),
	.w1(32'hba53eb7c),
	.w2(32'hba5080b8),
	.w3(32'h3b610bc2),
	.w4(32'h39197df8),
	.w5(32'hbb7eb097),
	.w6(32'h3b12d3a4),
	.w7(32'h39811344),
	.w8(32'h3a16b0a3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9947cc7),
	.w1(32'hbaff7d3c),
	.w2(32'hbbb4cdfb),
	.w3(32'hbae01f78),
	.w4(32'h3984ff2c),
	.w5(32'hba9f3ade),
	.w6(32'hbc0325fc),
	.w7(32'hbb1be605),
	.w8(32'hba15f4a7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6387ef),
	.w1(32'hbba2acbc),
	.w2(32'h3a4c3baf),
	.w3(32'h3a5e4d83),
	.w4(32'hbb721b38),
	.w5(32'hbb50b993),
	.w6(32'h3aeb8004),
	.w7(32'hbbbbf322),
	.w8(32'hbc3bb83c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8555a),
	.w1(32'h3a17402d),
	.w2(32'hba36f4d8),
	.w3(32'h37f32ad7),
	.w4(32'hbafee03e),
	.w5(32'hbba94c60),
	.w6(32'hbaba5af8),
	.w7(32'h3b832fe1),
	.w8(32'h3add4492),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70d868),
	.w1(32'h3b949f16),
	.w2(32'hbb20072f),
	.w3(32'hbc0ae896),
	.w4(32'hbbaa84f0),
	.w5(32'hbbfaf2e4),
	.w6(32'hb98fd427),
	.w7(32'hbb040ea2),
	.w8(32'hbb08f2fe),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93dc4fe),
	.w1(32'hbbb17314),
	.w2(32'hbbe179c1),
	.w3(32'hb9d22e24),
	.w4(32'hbab6da7d),
	.w5(32'h3bbcf3bc),
	.w6(32'hbb250faa),
	.w7(32'h3b60aefd),
	.w8(32'h3b818b97),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be099),
	.w1(32'h3af7937a),
	.w2(32'h3b770cbf),
	.w3(32'hb911c2df),
	.w4(32'hbac5435f),
	.w5(32'h3b128209),
	.w6(32'hbabf59e5),
	.w7(32'hbbae43d5),
	.w8(32'hbb6bcee2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68fa6e),
	.w1(32'h3b81bb24),
	.w2(32'h39a6cd8a),
	.w3(32'h3bba8aa4),
	.w4(32'h3b39780c),
	.w5(32'h3b90f685),
	.w6(32'hbae46b3f),
	.w7(32'hbaaa8bfd),
	.w8(32'hba48ee64),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f654c),
	.w1(32'hba33becb),
	.w2(32'h3bc7fe1d),
	.w3(32'h3b98d9ba),
	.w4(32'hbc083c68),
	.w5(32'hbc3b4e4e),
	.w6(32'hb789006e),
	.w7(32'h3b203420),
	.w8(32'hbb6f048b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd5fde),
	.w1(32'h3c03c6c5),
	.w2(32'hbb575823),
	.w3(32'hbbb8eadc),
	.w4(32'h3c2360df),
	.w5(32'h3c32f47a),
	.w6(32'h3bd183ce),
	.w7(32'hbb636db9),
	.w8(32'hbc085129),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d49e5),
	.w1(32'h3bd2846c),
	.w2(32'h3bbca4b5),
	.w3(32'h3c1d4a18),
	.w4(32'h3b144e7a),
	.w5(32'hbaf08c05),
	.w6(32'h3c9abf2b),
	.w7(32'h3cabbdae),
	.w8(32'h3c820ed8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2bb95),
	.w1(32'hbb8a6041),
	.w2(32'hb9f2d4ea),
	.w3(32'hba8bc1d5),
	.w4(32'hbb44c826),
	.w5(32'h38696a92),
	.w6(32'h3938659d),
	.w7(32'hb98be410),
	.w8(32'h3c25f658),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd83a4),
	.w1(32'h3ac74cef),
	.w2(32'h3991198e),
	.w3(32'hbb98079f),
	.w4(32'hbbb3e0f0),
	.w5(32'hbb2f3781),
	.w6(32'hbba278ba),
	.w7(32'hbbd72b05),
	.w8(32'hbbd4c07f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed85bc),
	.w1(32'hba423a98),
	.w2(32'h3c099e04),
	.w3(32'hbbe01678),
	.w4(32'hbae7fcb0),
	.w5(32'h3c398ab3),
	.w6(32'hbb4f610f),
	.w7(32'hbb98f308),
	.w8(32'hbbafa703),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85dc2b),
	.w1(32'hbab658bd),
	.w2(32'h3be206ae),
	.w3(32'hbb8df9d0),
	.w4(32'h3b84c58e),
	.w5(32'hbc1aa762),
	.w6(32'hbc1debd1),
	.w7(32'h3b299ea9),
	.w8(32'h3b20a9e8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badaaa7),
	.w1(32'h3c08b641),
	.w2(32'h3c0541cb),
	.w3(32'h3c1c4c3a),
	.w4(32'hbb0df185),
	.w5(32'h3c3a4042),
	.w6(32'h3ba28502),
	.w7(32'h3b66d9e4),
	.w8(32'h3c2ea526),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57b591),
	.w1(32'hbb95ab5e),
	.w2(32'hbc16e42c),
	.w3(32'h3b229a2d),
	.w4(32'hbc20c6bf),
	.w5(32'h3b7e6bd5),
	.w6(32'h3c0b24fb),
	.w7(32'hbc01c1de),
	.w8(32'hba5ebe5a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11332d),
	.w1(32'h3bc1a4b3),
	.w2(32'h3c456d7e),
	.w3(32'hbb7966c7),
	.w4(32'h3c4e62e4),
	.w5(32'hbb08f1fe),
	.w6(32'hbb28df01),
	.w7(32'h3c4b18fd),
	.w8(32'h3c7d7392),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee85d2),
	.w1(32'h3b42b6ed),
	.w2(32'hbab88ec5),
	.w3(32'h3bb4c54e),
	.w4(32'hbc5b4be3),
	.w5(32'hbc681d89),
	.w6(32'h3c9c6998),
	.w7(32'hbc8777b4),
	.w8(32'hbbc9a24e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f742),
	.w1(32'h3c1a3c1a),
	.w2(32'hb9edee4e),
	.w3(32'hbc0d02a0),
	.w4(32'hbb5e2a27),
	.w5(32'hbc8a2eca),
	.w6(32'h3c482b06),
	.w7(32'h3c3a5b03),
	.w8(32'h3b8dce3e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af77e4a),
	.w1(32'hbb86f58c),
	.w2(32'hbb98ab8d),
	.w3(32'h3bc5e3a5),
	.w4(32'hbb9e6dc1),
	.w5(32'hbcd530ce),
	.w6(32'hbb838006),
	.w7(32'hbbad2161),
	.w8(32'hbac59fec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22a28d),
	.w1(32'h3af255a5),
	.w2(32'hbcb4aae3),
	.w3(32'hbb20d2e7),
	.w4(32'hbbaba885),
	.w5(32'hbd3f7ffe),
	.w6(32'h3c63235d),
	.w7(32'hbb1689b2),
	.w8(32'hbca91326),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92146c),
	.w1(32'h3b1481f7),
	.w2(32'hbbab28e9),
	.w3(32'h3bd4fa57),
	.w4(32'h3baeeff4),
	.w5(32'hbba42c8a),
	.w6(32'h3c488094),
	.w7(32'h3a7f5f37),
	.w8(32'hbb1c6998),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27fa3),
	.w1(32'h3c85b39d),
	.w2(32'h3be85b03),
	.w3(32'h3a5c903f),
	.w4(32'h3c2d2b5e),
	.w5(32'hbbb84cae),
	.w6(32'hbabefe0b),
	.w7(32'h3c4fdbf1),
	.w8(32'h3b9f3b67),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6423fb),
	.w1(32'h394dfb16),
	.w2(32'h3b23f6cd),
	.w3(32'h3bb42674),
	.w4(32'hbb8e849c),
	.w5(32'hbb0d5765),
	.w6(32'h3c70d94f),
	.w7(32'h3b75d0c8),
	.w8(32'h3af41599),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b3096),
	.w1(32'hbbab4894),
	.w2(32'h3abca103),
	.w3(32'h3a2e2d38),
	.w4(32'hb9ca998d),
	.w5(32'hbc20734f),
	.w6(32'hbb99def0),
	.w7(32'hbb5e66b1),
	.w8(32'hbb3da74e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1efcc0),
	.w1(32'hbb47f028),
	.w2(32'h3c2923a8),
	.w3(32'hb860b312),
	.w4(32'h398339cc),
	.w5(32'h3c37260a),
	.w6(32'hb8d34ac4),
	.w7(32'hbaceec5f),
	.w8(32'hbae7f475),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96a8d7),
	.w1(32'hbb04e16f),
	.w2(32'h3aa80b21),
	.w3(32'h3b52f495),
	.w4(32'hbc02430b),
	.w5(32'h3c8330c5),
	.w6(32'hba8dde38),
	.w7(32'h39a112dd),
	.w8(32'hb9a6f031),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077ae7),
	.w1(32'hbbda5f70),
	.w2(32'hbbda849a),
	.w3(32'h3bba479f),
	.w4(32'h3b039dcb),
	.w5(32'hbb5f44aa),
	.w6(32'hba57cfee),
	.w7(32'hbc21354f),
	.w8(32'h3b02ec30),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3cf78),
	.w1(32'h3bf66f4b),
	.w2(32'h3a169bfd),
	.w3(32'h3b2a5129),
	.w4(32'h3c24eafd),
	.w5(32'hbc89f0fc),
	.w6(32'hbb8027db),
	.w7(32'hbb89db1a),
	.w8(32'hbbf22a1d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2c8bd),
	.w1(32'h3b3a3586),
	.w2(32'hbc3dcac8),
	.w3(32'h3c87bedf),
	.w4(32'hbc3ffb46),
	.w5(32'hbc574788),
	.w6(32'h3b49c9e0),
	.w7(32'hbbf5e8ca),
	.w8(32'h3ba6195d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5659c9),
	.w1(32'h3b9c1891),
	.w2(32'h3b412ccf),
	.w3(32'h3c129e43),
	.w4(32'h3b7de18f),
	.w5(32'h3b8a3cd0),
	.w6(32'h3b862786),
	.w7(32'h3b4ef985),
	.w8(32'hbb0b9e6d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c30ea),
	.w1(32'h3acb9c94),
	.w2(32'hbbfc415d),
	.w3(32'hbb9da856),
	.w4(32'h3c0e405a),
	.w5(32'hbc1ecd09),
	.w6(32'h3c2353db),
	.w7(32'h3c093a23),
	.w8(32'hbb64ef1b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc605fe),
	.w1(32'hbb985ea5),
	.w2(32'h3b0d8c36),
	.w3(32'hba3360bf),
	.w4(32'h3a9b45c9),
	.w5(32'h3c7abe0f),
	.w6(32'hbc3ac781),
	.w7(32'hbbee6215),
	.w8(32'hba95effd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865231),
	.w1(32'hba90f383),
	.w2(32'h3baca38b),
	.w3(32'hbbeeadd9),
	.w4(32'h3c28a2a5),
	.w5(32'h3c651063),
	.w6(32'h3c186b0a),
	.w7(32'hbbf86733),
	.w8(32'h3bb2076e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac28c07),
	.w1(32'hbb809390),
	.w2(32'h3c49433c),
	.w3(32'h3bab0113),
	.w4(32'hbbbfd3d7),
	.w5(32'hbb8afb8e),
	.w6(32'hbb23c28b),
	.w7(32'hbb44f967),
	.w8(32'h3ae9ab1e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafd0b0),
	.w1(32'hbb1d06e5),
	.w2(32'hbb9f66c0),
	.w3(32'h3b05d85e),
	.w4(32'hbb0e9a85),
	.w5(32'h3c5cb051),
	.w6(32'h3c3d852a),
	.w7(32'hbbde6b5f),
	.w8(32'h3b994d96),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bbd26),
	.w1(32'h3ba7f0c1),
	.w2(32'hbb79c309),
	.w3(32'hbb325150),
	.w4(32'h3b94c50a),
	.w5(32'hba1b9cda),
	.w6(32'h3bcef91e),
	.w7(32'hbbac7970),
	.w8(32'h3b95a2a5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f2020),
	.w1(32'h3a3e11de),
	.w2(32'hbc11527d),
	.w3(32'hb948d0ac),
	.w4(32'hbb152e29),
	.w5(32'h3d75182a),
	.w6(32'hbbf77e3f),
	.w7(32'hbc26eb6e),
	.w8(32'hbba4c616),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc69df),
	.w1(32'hba6b4f51),
	.w2(32'hbc892120),
	.w3(32'hbc0c0a3f),
	.w4(32'hbc3cc7cf),
	.w5(32'h3cce6cfa),
	.w6(32'hbc269424),
	.w7(32'hbc20354b),
	.w8(32'h3be04b0d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add2632),
	.w1(32'hbb25cfc3),
	.w2(32'h3bf40f95),
	.w3(32'h3be22805),
	.w4(32'hbb0aea51),
	.w5(32'h3c06a963),
	.w6(32'h3bd35bab),
	.w7(32'h3c63cee3),
	.w8(32'h3c392646),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9965c8b),
	.w1(32'hbb0fe205),
	.w2(32'hbc115650),
	.w3(32'h3b21cf03),
	.w4(32'hbc15a18e),
	.w5(32'h3c03857d),
	.w6(32'h3c2b1904),
	.w7(32'hba946d5e),
	.w8(32'hbb1c669f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4b212),
	.w1(32'hbb7b6fc7),
	.w2(32'h3c11a4cb),
	.w3(32'h3aacec08),
	.w4(32'hbbaaa9dc),
	.w5(32'hbc139ed6),
	.w6(32'h3c132f0c),
	.w7(32'h3c39fe76),
	.w8(32'h3c238348),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af31ea),
	.w1(32'h3b18d0e0),
	.w2(32'hb97b954a),
	.w3(32'h3b144a3c),
	.w4(32'hbb51172f),
	.w5(32'hbbd034ef),
	.w6(32'hbbf37bb7),
	.w7(32'hbca49c5a),
	.w8(32'hbb77ec64),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c088b99),
	.w1(32'hbc54ad36),
	.w2(32'hbb9ee0bd),
	.w3(32'h3b479546),
	.w4(32'hbb0b2e26),
	.w5(32'h3c878b96),
	.w6(32'h3ab1d362),
	.w7(32'hbbc341f4),
	.w8(32'hbc57aaea),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29938a),
	.w1(32'h3a1dfd68),
	.w2(32'hbbd7fb07),
	.w3(32'h3ac06373),
	.w4(32'hbc843a74),
	.w5(32'h3cdfe9c4),
	.w6(32'h3bcfe39d),
	.w7(32'hbb8eeba2),
	.w8(32'hbb8e363e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5365a),
	.w1(32'h38698420),
	.w2(32'hba5c4033),
	.w3(32'hbc175ad4),
	.w4(32'h3c12a51d),
	.w5(32'h3ada8ede),
	.w6(32'hbc629ac6),
	.w7(32'h3a7aa624),
	.w8(32'hbbc4f483),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db386),
	.w1(32'hbc4184de),
	.w2(32'h3c3cd342),
	.w3(32'h3c22d942),
	.w4(32'hbc723ec9),
	.w5(32'hbca25d6a),
	.w6(32'h3c2858d5),
	.w7(32'hba8660c8),
	.w8(32'h3aad4e27),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d9f60),
	.w1(32'hba482268),
	.w2(32'hbbffec89),
	.w3(32'h3be0d690),
	.w4(32'hbc167486),
	.w5(32'hbbe0288f),
	.w6(32'hba70f456),
	.w7(32'hbbcc4569),
	.w8(32'h3b35197d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1fae),
	.w1(32'h3c376381),
	.w2(32'hbb87ac1c),
	.w3(32'h385ae747),
	.w4(32'h3c9cec9e),
	.w5(32'hbcbd3384),
	.w6(32'h3a712b70),
	.w7(32'h3bdca842),
	.w8(32'hbbde70d2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ed9cb),
	.w1(32'h3aa8a1aa),
	.w2(32'h3ba7de85),
	.w3(32'h3c37bbc4),
	.w4(32'hba113a88),
	.w5(32'h3d0aeda8),
	.w6(32'hbb83eb60),
	.w7(32'h3b338a3a),
	.w8(32'h3c1e1216),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb012aae),
	.w1(32'hbc3aaf82),
	.w2(32'h3a005952),
	.w3(32'hbc2d5f70),
	.w4(32'hbc9f320f),
	.w5(32'h3af4c341),
	.w6(32'h39ad4ac6),
	.w7(32'hbc8b1630),
	.w8(32'hb8822f44),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb81091),
	.w1(32'h3a649eac),
	.w2(32'h3a752a86),
	.w3(32'hbb9e9b53),
	.w4(32'hbac4452b),
	.w5(32'h3cad62d7),
	.w6(32'hbaab7a62),
	.w7(32'hbbabf49f),
	.w8(32'hbbf72632),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d06f6),
	.w1(32'h3c157ca8),
	.w2(32'hba921510),
	.w3(32'hbc956216),
	.w4(32'h3b8170a6),
	.w5(32'h3b31cfa8),
	.w6(32'hbc0cfc4a),
	.w7(32'hbc0671ce),
	.w8(32'hbc1c19ad),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1dc9a),
	.w1(32'hba299ed3),
	.w2(32'hbb766cae),
	.w3(32'hbc1b9f56),
	.w4(32'hbb933fbd),
	.w5(32'h3b814ce7),
	.w6(32'hbb2611b5),
	.w7(32'h3bb52e6c),
	.w8(32'hbad799c7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b807f1a),
	.w1(32'hbbc361b5),
	.w2(32'h3baffd73),
	.w3(32'h3b5cdae6),
	.w4(32'hbcb6a7bc),
	.w5(32'h3d311bd9),
	.w6(32'h3c28f09b),
	.w7(32'h3c68a65d),
	.w8(32'h3cabaf49),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38f082),
	.w1(32'hba220eab),
	.w2(32'hbb779b3d),
	.w3(32'hbc711e91),
	.w4(32'h3cbeb135),
	.w5(32'hbcb584d9),
	.w6(32'hbc5b0437),
	.w7(32'hbc333db6),
	.w8(32'hbb97ddfc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ea5b0),
	.w1(32'hbb6bf400),
	.w2(32'h3a980a65),
	.w3(32'h3bb98543),
	.w4(32'h3bc4e19b),
	.w5(32'hbc1e174b),
	.w6(32'h3bbbfe67),
	.w7(32'h3b97d407),
	.w8(32'hba7e20cf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c0bc),
	.w1(32'hbb372f2f),
	.w2(32'hbb9e610b),
	.w3(32'h3c8263c3),
	.w4(32'hbc0de1ba),
	.w5(32'hbc283f8d),
	.w6(32'h3c001619),
	.w7(32'hbb87eddd),
	.w8(32'hbb91976d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad31258),
	.w1(32'h3afda4a8),
	.w2(32'hbb60de9e),
	.w3(32'hbb6e2f20),
	.w4(32'hbb9af04e),
	.w5(32'h3cda3121),
	.w6(32'hbb5fa723),
	.w7(32'hbc0879c1),
	.w8(32'h394d2c04),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc376016),
	.w1(32'h3c055056),
	.w2(32'hbb11c727),
	.w3(32'hbc389f4d),
	.w4(32'h3bb79e58),
	.w5(32'hbc95d38e),
	.w6(32'hbc03b8d3),
	.w7(32'h3b0a67da),
	.w8(32'h3af76494),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe13bae),
	.w1(32'hbc0a5ea5),
	.w2(32'hbc0d6a3f),
	.w3(32'h3b437b1c),
	.w4(32'hbc83bb8d),
	.w5(32'hbbdfadca),
	.w6(32'h3bd6a99e),
	.w7(32'hbcb3ed41),
	.w8(32'hbb2cbdb8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc166a38),
	.w1(32'hbb406c7c),
	.w2(32'h3c0ee95c),
	.w3(32'hbbb59dcc),
	.w4(32'hbc274f14),
	.w5(32'h3d839f67),
	.w6(32'hbb6b83d0),
	.w7(32'hbbdb3010),
	.w8(32'h3c8872ff),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39703b),
	.w1(32'h3a2509ac),
	.w2(32'h39c5135f),
	.w3(32'hbad877d3),
	.w4(32'h3b72b370),
	.w5(32'h3ae5351e),
	.w6(32'hbad28789),
	.w7(32'h3a702f54),
	.w8(32'hbb2d07d4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6d0a7),
	.w1(32'h3b1a6117),
	.w2(32'h3a0bbbdd),
	.w3(32'h3bfc371d),
	.w4(32'hbbab0172),
	.w5(32'h3c6d7fc3),
	.w6(32'h3c1843ab),
	.w7(32'h3bccbee3),
	.w8(32'h3b590f7f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a126137),
	.w1(32'h3c2bc9fa),
	.w2(32'h3b6fafb0),
	.w3(32'hbbdd3755),
	.w4(32'h3aed3273),
	.w5(32'h3d17c52d),
	.w6(32'h3a692434),
	.w7(32'hba02086e),
	.w8(32'h3c4db608),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a933),
	.w1(32'hbbe9c15b),
	.w2(32'h3b3ca0cd),
	.w3(32'h3be90458),
	.w4(32'hbc1ce237),
	.w5(32'h3d722572),
	.w6(32'hbb48db0b),
	.w7(32'hbb35b014),
	.w8(32'h3c8be1b4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014b64),
	.w1(32'h3c1425a2),
	.w2(32'h3c52e7fb),
	.w3(32'hbc19eddd),
	.w4(32'h3bacbd62),
	.w5(32'h3b726bca),
	.w6(32'hbbec2d57),
	.w7(32'h3ba61cd4),
	.w8(32'h3b92a5a0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43c37e),
	.w1(32'hbc3afade),
	.w2(32'h3b87b0d5),
	.w3(32'h3ad86c41),
	.w4(32'h39e8cb09),
	.w5(32'hbc81aaae),
	.w6(32'h3ad52fca),
	.w7(32'h3a82b74e),
	.w8(32'h3c1e24d9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20ee3a),
	.w1(32'hbc489085),
	.w2(32'hbc17ce3c),
	.w3(32'h3c01572f),
	.w4(32'hbc7f62ae),
	.w5(32'hbc93ecb6),
	.w6(32'h3c15982c),
	.w7(32'hbbd42495),
	.w8(32'hbc27d970),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2de9),
	.w1(32'hba5439b4),
	.w2(32'h3c1e2be2),
	.w3(32'hbc64b8cb),
	.w4(32'hbc387dad),
	.w5(32'hbc119648),
	.w6(32'h3be9a989),
	.w7(32'h3c805f65),
	.w8(32'h3c84ba60),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801033),
	.w1(32'h3b986b34),
	.w2(32'hbb7ee0b6),
	.w3(32'h3b59b3d3),
	.w4(32'h3bb8b458),
	.w5(32'hbc46977a),
	.w6(32'h3c751047),
	.w7(32'h3b9f57c6),
	.w8(32'h3a334752),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36b12a),
	.w1(32'hbc1b395e),
	.w2(32'hbc4235c6),
	.w3(32'h38f234d2),
	.w4(32'h3b018589),
	.w5(32'hbb5eba55),
	.w6(32'h3bf662ff),
	.w7(32'hbc413f91),
	.w8(32'hbc25c886),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff1822),
	.w1(32'h3b052c4a),
	.w2(32'h3a650213),
	.w3(32'h3b300473),
	.w4(32'h3ba2c49b),
	.w5(32'h39e05aeb),
	.w6(32'h3b9cd444),
	.w7(32'hb96fea69),
	.w8(32'h3bd63b60),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45bec6),
	.w1(32'hb926e263),
	.w2(32'hbbc40476),
	.w3(32'hbc91ece3),
	.w4(32'h3c3c0f64),
	.w5(32'hbca390c3),
	.w6(32'hbc2edeaa),
	.w7(32'h3b18ee11),
	.w8(32'hbbf277d5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c086983),
	.w1(32'hbbf9a2b7),
	.w2(32'h3c1f679d),
	.w3(32'h3bf9253d),
	.w4(32'hbc05ef93),
	.w5(32'h3cee1ac0),
	.w6(32'h3c9704b3),
	.w7(32'hbb8db20f),
	.w8(32'h3c153dff),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8b9fd),
	.w1(32'hbb273740),
	.w2(32'hbb80a833),
	.w3(32'hbbccec46),
	.w4(32'h3bf2b6f6),
	.w5(32'hbc2292e7),
	.w6(32'hbb8f675c),
	.w7(32'h3b080bae),
	.w8(32'hbb0cb0ef),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44c063),
	.w1(32'h3ba6f508),
	.w2(32'hbba80ee5),
	.w3(32'h3b702203),
	.w4(32'hbc4bb921),
	.w5(32'h3c0a7916),
	.w6(32'h3c6e9210),
	.w7(32'hb795bce4),
	.w8(32'h3a9cb96e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbac33a),
	.w1(32'hbb9d88b8),
	.w2(32'hbbee2d74),
	.w3(32'hba965e6f),
	.w4(32'hba203032),
	.w5(32'h3ae13635),
	.w6(32'hbc1c4ae2),
	.w7(32'hbbd5e332),
	.w8(32'h3aacd8c7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44e736),
	.w1(32'h3ac284d0),
	.w2(32'hbae858d2),
	.w3(32'hbba17d91),
	.w4(32'h3b895727),
	.w5(32'h3bcd9ff9),
	.w6(32'h3b470004),
	.w7(32'hb92b7f66),
	.w8(32'h3bc2169f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38fb29),
	.w1(32'h3b15a1e1),
	.w2(32'hbb0c6546),
	.w3(32'h3c0ee222),
	.w4(32'hbbcfdb79),
	.w5(32'hbc63b6d1),
	.w6(32'h3c64bb40),
	.w7(32'hbba6eff6),
	.w8(32'h39c38754),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befa56f),
	.w1(32'hbb8a6f3f),
	.w2(32'h3b0c9d07),
	.w3(32'h3c0309c8),
	.w4(32'hbc36cec0),
	.w5(32'h3b0f7390),
	.w6(32'h3c1c3369),
	.w7(32'h3af671dd),
	.w8(32'h3b60e3fc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e8dd8),
	.w1(32'hbafd84b9),
	.w2(32'hbb3da6c2),
	.w3(32'h3ba5f7a7),
	.w4(32'h378f0cd8),
	.w5(32'h39bcb7ea),
	.w6(32'h3b898a14),
	.w7(32'h3a38ab90),
	.w8(32'h3b5c7d67),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e9799),
	.w1(32'hbb85c5d4),
	.w2(32'hbb721e7c),
	.w3(32'h3bf2375b),
	.w4(32'h3b47c0c4),
	.w5(32'hbcadfd2d),
	.w6(32'hb82ba91a),
	.w7(32'hbbaf2151),
	.w8(32'hbbe5d242),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8045ac),
	.w1(32'hbb041975),
	.w2(32'h3c5ab466),
	.w3(32'h3c589ecf),
	.w4(32'hbc3ede4f),
	.w5(32'h3b7d70da),
	.w6(32'hbc72829f),
	.w7(32'hbbf8e0c8),
	.w8(32'hbb86f8ff),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59fa8d),
	.w1(32'h3b3c5807),
	.w2(32'hb9d7adb8),
	.w3(32'hbb8132bd),
	.w4(32'hbb212c0b),
	.w5(32'h3d0d2420),
	.w6(32'hbbc40911),
	.w7(32'hb9ca4501),
	.w8(32'hbb48ea65),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc30da9),
	.w1(32'h3b17d6f3),
	.w2(32'h3bd0a47d),
	.w3(32'hbb8e50cd),
	.w4(32'h3c250337),
	.w5(32'h3c414785),
	.w6(32'hbb2b1458),
	.w7(32'h3c0fbd83),
	.w8(32'h3b8d1edc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfae21a),
	.w1(32'hbb1c2d11),
	.w2(32'hbb747446),
	.w3(32'hbbc62ac5),
	.w4(32'hba0d98ba),
	.w5(32'hbbd09b8a),
	.w6(32'hbc0dae07),
	.w7(32'h3c1fecc0),
	.w8(32'h3bde75ca),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95f004),
	.w1(32'hbb45d9bf),
	.w2(32'hba5b3db9),
	.w3(32'h3a48ce31),
	.w4(32'h3b61bf2d),
	.w5(32'hbb84d57b),
	.w6(32'h3b8fd510),
	.w7(32'h39bf81b7),
	.w8(32'hbb5952bf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1580b0),
	.w1(32'hbbb734df),
	.w2(32'hba306974),
	.w3(32'hbc02961c),
	.w4(32'hb9cb1cff),
	.w5(32'h3ca13c0b),
	.w6(32'hbbf49862),
	.w7(32'hbb4b4bc7),
	.w8(32'hbb24292f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b46d6),
	.w1(32'hbb230f07),
	.w2(32'hb84c1ba2),
	.w3(32'h3ab7a8ec),
	.w4(32'h3b96d543),
	.w5(32'hbbdb8527),
	.w6(32'hbac86fe8),
	.w7(32'h3b79861e),
	.w8(32'hbb76dc3a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb26e8d),
	.w1(32'h3bc42e74),
	.w2(32'h3aa2570e),
	.w3(32'h3b2833d0),
	.w4(32'h3c997273),
	.w5(32'h3b140a3c),
	.w6(32'h3b9480ef),
	.w7(32'h3c0eda52),
	.w8(32'h3b4fc8c6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69fade),
	.w1(32'hbbc1faf0),
	.w2(32'hbc5bfc4c),
	.w3(32'h3c38ef69),
	.w4(32'h3a327099),
	.w5(32'hbc977b90),
	.w6(32'h3c0d808f),
	.w7(32'hbbed0789),
	.w8(32'hbc6ab974),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78883),
	.w1(32'hbaca439b),
	.w2(32'hbb3df009),
	.w3(32'hbbefc16a),
	.w4(32'hbbd00a5b),
	.w5(32'hbbe3affb),
	.w6(32'hbb81171f),
	.w7(32'hbbb6f8c8),
	.w8(32'hbb90317b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b238),
	.w1(32'hbb7f985c),
	.w2(32'hbbaba78b),
	.w3(32'hb80a6252),
	.w4(32'h3bb37a5a),
	.w5(32'h39f41a72),
	.w6(32'h3b911aff),
	.w7(32'h395da9cf),
	.w8(32'hbbef3259),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf298e),
	.w1(32'h3c0a4604),
	.w2(32'hbbe5880e),
	.w3(32'hbc00d269),
	.w4(32'h3c33305b),
	.w5(32'h3bd998f1),
	.w6(32'hbc4c8538),
	.w7(32'h39e5ced3),
	.w8(32'h3b22fab0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6661a),
	.w1(32'h3b4969be),
	.w2(32'hbb40bee7),
	.w3(32'h3aa82c6d),
	.w4(32'h3bff7bfc),
	.w5(32'hbbefba70),
	.w6(32'h3a3af509),
	.w7(32'hbb1250f5),
	.w8(32'hba5329c2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928180),
	.w1(32'h3bd5cc97),
	.w2(32'h3a1231c6),
	.w3(32'h3c24fd35),
	.w4(32'hbb2e416d),
	.w5(32'hbab8d95c),
	.w6(32'h3b395c88),
	.w7(32'hbb95c5ac),
	.w8(32'hbb710bac),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fde73),
	.w1(32'h3b85dfab),
	.w2(32'h3b88ffdc),
	.w3(32'hbb4ba01c),
	.w4(32'h3ad7295d),
	.w5(32'h3c951220),
	.w6(32'h3bcca5bc),
	.w7(32'h3aad6152),
	.w8(32'hba7510e8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dfa93),
	.w1(32'h3bab1215),
	.w2(32'hbac92a02),
	.w3(32'hbb5f843c),
	.w4(32'h39339d09),
	.w5(32'hbc60a5b3),
	.w6(32'hbb741bd9),
	.w7(32'hbb448a70),
	.w8(32'h3b04aad1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b767655),
	.w1(32'h3b658a31),
	.w2(32'h3b2e40dc),
	.w3(32'h3b89ac07),
	.w4(32'h3b5afae6),
	.w5(32'hbc814982),
	.w6(32'h3b419310),
	.w7(32'hba82f0b3),
	.w8(32'hbb03d8dd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba379b32),
	.w1(32'h3b848a58),
	.w2(32'h3b732ddb),
	.w3(32'h3be1546a),
	.w4(32'h3ba517ae),
	.w5(32'hbb2145b9),
	.w6(32'h3b8227c1),
	.w7(32'h3af67d04),
	.w8(32'hbb29b195),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f05af),
	.w1(32'h3ac5b6e7),
	.w2(32'h3bb37253),
	.w3(32'hb9a20ff9),
	.w4(32'hba825195),
	.w5(32'h3cb8e264),
	.w6(32'hba75873e),
	.w7(32'hbae47cc1),
	.w8(32'h3bd53b88),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b456938),
	.w1(32'h3c34679b),
	.w2(32'h3bbcb253),
	.w3(32'h3ad694b4),
	.w4(32'h38580b9c),
	.w5(32'hbc121088),
	.w6(32'hba52d791),
	.w7(32'h3c8a3f8b),
	.w8(32'h3aceeb5d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6fea9),
	.w1(32'hbb744f62),
	.w2(32'hbb8f2adb),
	.w3(32'hba98768d),
	.w4(32'hba0ae75c),
	.w5(32'h3c9f37a6),
	.w6(32'hbbab238c),
	.w7(32'h3bc1e5f3),
	.w8(32'h3be7da97),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb8db4),
	.w1(32'hbb06d294),
	.w2(32'h3b4405d4),
	.w3(32'hbc0c3eae),
	.w4(32'h3c10895c),
	.w5(32'hbba5c429),
	.w6(32'hbbb4c14e),
	.w7(32'h3bc562e2),
	.w8(32'hbb237bb2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a3612),
	.w1(32'h3c28038f),
	.w2(32'hbc653ed8),
	.w3(32'hbb26771e),
	.w4(32'h3c70d1e1),
	.w5(32'hbd32484f),
	.w6(32'hbb6b0fde),
	.w7(32'h3bdec24a),
	.w8(32'hbc67daba),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b755951),
	.w1(32'h3a7aa572),
	.w2(32'h3bd677bb),
	.w3(32'h3c1dd409),
	.w4(32'hbbdf2e0a),
	.w5(32'h3b0d5807),
	.w6(32'h3c6435d9),
	.w7(32'h3c1966b0),
	.w8(32'h3c587e98),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53f233),
	.w1(32'h3c35ffeb),
	.w2(32'hbc03fc7f),
	.w3(32'h3b2c48c7),
	.w4(32'h3c39583c),
	.w5(32'hbcb79aa5),
	.w6(32'hbb689a37),
	.w7(32'h3bc96ff4),
	.w8(32'hbbf79d8e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004a7b),
	.w1(32'hbc041d3e),
	.w2(32'hbb42e4e9),
	.w3(32'h3c555369),
	.w4(32'hbcc3a061),
	.w5(32'h3d4ff19e),
	.w6(32'h3c26d2c7),
	.w7(32'hbc24f401),
	.w8(32'hbaef0b67),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d02cf),
	.w1(32'hbc15a9d6),
	.w2(32'hbc5489af),
	.w3(32'hbc330b69),
	.w4(32'hbb8183a4),
	.w5(32'hbcc38112),
	.w6(32'hbb9e7079),
	.w7(32'hb8186fbe),
	.w8(32'hbc501db7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86c321),
	.w1(32'hbca0bdd2),
	.w2(32'h3c59f125),
	.w3(32'h3cc1ab39),
	.w4(32'hbce82732),
	.w5(32'h3c072e1d),
	.w6(32'h3c54bb9b),
	.w7(32'h39b89e7e),
	.w8(32'h3c367ba8),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e461),
	.w1(32'hbc0f33e3),
	.w2(32'hbc4823cd),
	.w3(32'h3b844817),
	.w4(32'hbc0387f6),
	.w5(32'h3cf8d459),
	.w6(32'hbb653cd1),
	.w7(32'hbc22ccdc),
	.w8(32'hbb6dbea2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24080),
	.w1(32'hbb292763),
	.w2(32'hbb7744df),
	.w3(32'h3b46af42),
	.w4(32'h3c302f68),
	.w5(32'hbbe6e75e),
	.w6(32'hbc22c732),
	.w7(32'h3b11fbf8),
	.w8(32'hba53c02d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc073d03),
	.w1(32'h3b699c9c),
	.w2(32'hbc3994de),
	.w3(32'h3ad6e11c),
	.w4(32'h3c0054fa),
	.w5(32'hbc8295cb),
	.w6(32'h3b4830b2),
	.w7(32'h3bae25f5),
	.w8(32'hbc529178),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd21195),
	.w1(32'h3bea367a),
	.w2(32'h3a2d6e12),
	.w3(32'hbb92596f),
	.w4(32'h3b9fda52),
	.w5(32'h3cd3be05),
	.w6(32'hb9b7a744),
	.w7(32'hbb3eb6eb),
	.w8(32'h3ac65e1f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7eed1),
	.w1(32'h3b2f3db8),
	.w2(32'h3c3c1e15),
	.w3(32'hba40b5be),
	.w4(32'h3c08c889),
	.w5(32'h3c87b0fe),
	.w6(32'h3bfe0990),
	.w7(32'h3ba993a4),
	.w8(32'h3a8da7e3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f82e6a),
	.w1(32'hba045481),
	.w2(32'hbb171cc6),
	.w3(32'hbc4037ff),
	.w4(32'h388ecdff),
	.w5(32'hbc477f9a),
	.w6(32'h399f696f),
	.w7(32'h3bba4ea3),
	.w8(32'hbbfb36d8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00f248),
	.w1(32'hbba51029),
	.w2(32'hbbacb06f),
	.w3(32'hba881264),
	.w4(32'hbcab317d),
	.w5(32'hba8abe95),
	.w6(32'hbbf02289),
	.w7(32'hbc3b4907),
	.w8(32'hbbb01e67),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72b018),
	.w1(32'h3b529ce3),
	.w2(32'hbac6a16e),
	.w3(32'h3b10be3a),
	.w4(32'h3b80875a),
	.w5(32'h3bd2f7ef),
	.w6(32'h3be156e5),
	.w7(32'h3a7c74b7),
	.w8(32'hbbd816c8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaae23a),
	.w1(32'hbba05d08),
	.w2(32'h3bb51a92),
	.w3(32'hba8f566f),
	.w4(32'hbbaec31e),
	.w5(32'h3cac3408),
	.w6(32'hbb3166f1),
	.w7(32'hbb1b8d49),
	.w8(32'h3b9e4212),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac11880),
	.w1(32'h3af2af72),
	.w2(32'hbaaf5f5a),
	.w3(32'h3bbc1558),
	.w4(32'hba1fa0ff),
	.w5(32'hbb9275f4),
	.w6(32'hbb98ef34),
	.w7(32'hb9d73caf),
	.w8(32'hbbaa41fb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f025),
	.w1(32'h3b8603cb),
	.w2(32'hbb871679),
	.w3(32'h3be6e9ab),
	.w4(32'h3c05ca26),
	.w5(32'hbc0b8594),
	.w6(32'h38b57cd8),
	.w7(32'h3c30f860),
	.w8(32'hbb1db84f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a754024),
	.w1(32'hbb95194f),
	.w2(32'h3b7d03b4),
	.w3(32'h3aafd701),
	.w4(32'hbb9d371c),
	.w5(32'h3c54b9ae),
	.w6(32'h3a53d0c6),
	.w7(32'hbba398f4),
	.w8(32'h3bb9d22a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6823),
	.w1(32'h3c2bbc2f),
	.w2(32'h378ff5f4),
	.w3(32'h3bb6e138),
	.w4(32'h3ba2f23f),
	.w5(32'hbd06b665),
	.w6(32'h3b176a1c),
	.w7(32'h3b8e65d0),
	.w8(32'hbb5573ac),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafddc3),
	.w1(32'hbc18a706),
	.w2(32'hbb9d6f23),
	.w3(32'h3ab0f647),
	.w4(32'hbb3271e6),
	.w5(32'hbc147887),
	.w6(32'h3b2106c4),
	.w7(32'h3a950fd6),
	.w8(32'hba83387a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d1316),
	.w1(32'hba1c902b),
	.w2(32'hba8185e5),
	.w3(32'h3c089b61),
	.w4(32'h3c974953),
	.w5(32'hbc35beed),
	.w6(32'hba53c2f7),
	.w7(32'hbc2a26fa),
	.w8(32'hbaca9506),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46a16f),
	.w1(32'h3c27c99a),
	.w2(32'h3afb20a4),
	.w3(32'h3c207c32),
	.w4(32'h3c96a7f5),
	.w5(32'hbc72a498),
	.w6(32'hbbd596f8),
	.w7(32'h3b478887),
	.w8(32'hbb969295),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b322a),
	.w1(32'hbb7fb7d4),
	.w2(32'h3a2f4979),
	.w3(32'hbac2ba58),
	.w4(32'hbc17d72d),
	.w5(32'hbb97d4ed),
	.w6(32'h3b3b58b8),
	.w7(32'hba0bc291),
	.w8(32'h3b6bfc4a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc42a),
	.w1(32'hbc0141ea),
	.w2(32'hbc12ac2c),
	.w3(32'h3ab113ed),
	.w4(32'hbb0838be),
	.w5(32'hbc472893),
	.w6(32'hba0bd00b),
	.w7(32'hba95e732),
	.w8(32'hbb8dc22c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ef06a),
	.w1(32'hbbce902c),
	.w2(32'hbbe543ba),
	.w3(32'h3c1daa0a),
	.w4(32'hbbd610a7),
	.w5(32'hb849200b),
	.w6(32'h3c7d5dd2),
	.w7(32'h3c732938),
	.w8(32'h3b6215a9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4ebfe),
	.w1(32'h3b53047f),
	.w2(32'hbc92048a),
	.w3(32'hbc148cde),
	.w4(32'h3c37cec4),
	.w5(32'hbabedc72),
	.w6(32'hbc097d79),
	.w7(32'hbc380b00),
	.w8(32'hbc6776b2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5ff6),
	.w1(32'hbb0e57a6),
	.w2(32'h3a56bb32),
	.w3(32'hbb926283),
	.w4(32'hbc66204c),
	.w5(32'h3d824941),
	.w6(32'h3b4bb7ff),
	.w7(32'hbb626c85),
	.w8(32'h3c26b74d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef8ef6),
	.w1(32'hbc0a29a8),
	.w2(32'hbbb6db67),
	.w3(32'hbcb07e8c),
	.w4(32'h3c53d0e5),
	.w5(32'h3aa8991e),
	.w6(32'hbc08e066),
	.w7(32'hbb39e7bf),
	.w8(32'hbbb3c0f7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b3967),
	.w1(32'h3c090dd7),
	.w2(32'hbb05a12e),
	.w3(32'hb9fdbd9e),
	.w4(32'h3ba713a4),
	.w5(32'hbc3f9059),
	.w6(32'hbbd73dbf),
	.w7(32'h3ba5263e),
	.w8(32'h3adacdf5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84d388),
	.w1(32'h3c8b95c4),
	.w2(32'h3b8d6af6),
	.w3(32'hbae5abb5),
	.w4(32'h3cb048ae),
	.w5(32'hbca3004b),
	.w6(32'hba38ae99),
	.w7(32'h3cad8994),
	.w8(32'h3b06fd82),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee822),
	.w1(32'hbc69c885),
	.w2(32'h3b6d1199),
	.w3(32'h3bcdc1a1),
	.w4(32'hbc6de889),
	.w5(32'h3d64b3ab),
	.w6(32'h3c0a96a5),
	.w7(32'hbb971807),
	.w8(32'h3c5a1d5a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc073283),
	.w1(32'h3c4de850),
	.w2(32'hbba7acaf),
	.w3(32'h3b512530),
	.w4(32'h3c054405),
	.w5(32'hba0fb78f),
	.w6(32'hbb8080e5),
	.w7(32'h3c2a0728),
	.w8(32'h3bb36618),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc27e91),
	.w1(32'h3b432ebc),
	.w2(32'hbb4535fa),
	.w3(32'hbb6ab4bc),
	.w4(32'hbaeb15f0),
	.w5(32'h3bd53a4e),
	.w6(32'hbaa198fc),
	.w7(32'h3b08b93c),
	.w8(32'hb9f522af),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc558494),
	.w1(32'hba1ac60f),
	.w2(32'h3b4e2daf),
	.w3(32'hbce976b0),
	.w4(32'hba639ec7),
	.w5(32'h3c459568),
	.w6(32'hbc46a83b),
	.w7(32'h3b30b62a),
	.w8(32'h3b8222d9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef750c),
	.w1(32'hba67e3bc),
	.w2(32'hbc647ac8),
	.w3(32'h3b1fb97d),
	.w4(32'h39d530ee),
	.w5(32'hbc6a47ab),
	.w6(32'h3b6dde9b),
	.w7(32'h3ac2cda8),
	.w8(32'hbc350018),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc8a9),
	.w1(32'h38f13ef1),
	.w2(32'h3ba23b21),
	.w3(32'hbb754e8d),
	.w4(32'h3b3f4938),
	.w5(32'h3884d9f5),
	.w6(32'hbb570d11),
	.w7(32'h3b921738),
	.w8(32'hbb03cc5a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41c538),
	.w1(32'h3be5bd45),
	.w2(32'h3bdb5bf0),
	.w3(32'hbb7aa9e5),
	.w4(32'hba8bd5f1),
	.w5(32'hbb46b560),
	.w6(32'hbb535c3d),
	.w7(32'h3bc6dcf2),
	.w8(32'h3babab62),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955343a),
	.w1(32'h394a31f0),
	.w2(32'h3b576fb9),
	.w3(32'h3b0d6797),
	.w4(32'hbb91a246),
	.w5(32'hbb3d3a59),
	.w6(32'h3c05ec77),
	.w7(32'h3c1d72f4),
	.w8(32'h3b044a2a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c016a79),
	.w1(32'hbbeb3421),
	.w2(32'hbad7e0fc),
	.w3(32'h3bc5988a),
	.w4(32'hbb74f580),
	.w5(32'h39e4a15a),
	.w6(32'h3b78f074),
	.w7(32'h39bd70cb),
	.w8(32'hbaaa73d7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f17706),
	.w1(32'hbb4f8416),
	.w2(32'hbb8bf314),
	.w3(32'hbb391256),
	.w4(32'hbbba4ca3),
	.w5(32'hbb0e5267),
	.w6(32'h3b149dd8),
	.w7(32'hbb28ce03),
	.w8(32'h3a2258b8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58cd8),
	.w1(32'hbb3674f1),
	.w2(32'hbbad798a),
	.w3(32'hbc5c56c2),
	.w4(32'hbb3ae0ce),
	.w5(32'hbb75ce86),
	.w6(32'hbb43840c),
	.w7(32'hbbbccc8d),
	.w8(32'hbb3a32d4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e76c4),
	.w1(32'h3b1ea558),
	.w2(32'h3bad6e3c),
	.w3(32'hbc049791),
	.w4(32'hbad823a8),
	.w5(32'h3c61a5f0),
	.w6(32'hbabf83e6),
	.w7(32'hbb2308c5),
	.w8(32'h3c4d4802),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee7d3),
	.w1(32'hb93ac4f8),
	.w2(32'h3b6b0870),
	.w3(32'h3c3fe12f),
	.w4(32'h3b1f6a89),
	.w5(32'hbbdaaaf1),
	.w6(32'h3c2c6125),
	.w7(32'h3b733be4),
	.w8(32'h3c09060d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7bb15),
	.w1(32'h3b9217ea),
	.w2(32'h3c184acb),
	.w3(32'hbb79b8f7),
	.w4(32'h3ba7ff93),
	.w5(32'hbad48445),
	.w6(32'hbb0002cb),
	.w7(32'hbaa7a34b),
	.w8(32'h39363bf4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02e1ad),
	.w1(32'h3a5cf538),
	.w2(32'h3afd4b09),
	.w3(32'h3add4474),
	.w4(32'hbc27135c),
	.w5(32'h3b7be72d),
	.w6(32'h3b0ee196),
	.w7(32'hbb2d0f3c),
	.w8(32'hbbc32f0d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d6c52),
	.w1(32'h3c7adb6a),
	.w2(32'h3ca4b4a4),
	.w3(32'h3baec25e),
	.w4(32'hbb5d3647),
	.w5(32'h3c21f6b5),
	.w6(32'hb983007d),
	.w7(32'h3b7d81f8),
	.w8(32'h3bb5646c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c643966),
	.w1(32'h3c0d0e24),
	.w2(32'h3c852809),
	.w3(32'h3c59cfda),
	.w4(32'hbb515563),
	.w5(32'hbbbff705),
	.w6(32'h3ad9fd2d),
	.w7(32'h3b861709),
	.w8(32'h3b8ad932),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c064c11),
	.w1(32'hba966db0),
	.w2(32'hbb14c6a5),
	.w3(32'h3bae1b09),
	.w4(32'hba8bea81),
	.w5(32'hbae5310f),
	.w6(32'h3bc922c7),
	.w7(32'hbbc46154),
	.w8(32'hbbcf8a99),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5f85),
	.w1(32'h39dd9d59),
	.w2(32'hbb4e1c2c),
	.w3(32'h3bc674c5),
	.w4(32'hbc80ca7a),
	.w5(32'hbb817834),
	.w6(32'h3b7e726e),
	.w7(32'h3c84eb88),
	.w8(32'h3a5b9044),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab75fb),
	.w1(32'h3ac32171),
	.w2(32'h3bffeb4f),
	.w3(32'h3bceb0cf),
	.w4(32'hbb4acdcf),
	.w5(32'h3a85a97d),
	.w6(32'h3aa4c2c2),
	.w7(32'h3bb4b203),
	.w8(32'h3c74e60a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaba40),
	.w1(32'hbbedc580),
	.w2(32'hba635e08),
	.w3(32'h3b362d97),
	.w4(32'h3b244aea),
	.w5(32'hbb93bf7a),
	.w6(32'h3bbda81e),
	.w7(32'hbb807c66),
	.w8(32'hbc0f9f41),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacfeeb),
	.w1(32'hbbcfd382),
	.w2(32'hbc3fc4ca),
	.w3(32'h3ab0d3b7),
	.w4(32'h3ac8ac3b),
	.w5(32'h3c866cd3),
	.w6(32'hbbf64218),
	.w7(32'hbc633897),
	.w8(32'hbc9ad2d2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc6311),
	.w1(32'hbac4ceec),
	.w2(32'h3be06907),
	.w3(32'hbbc22de9),
	.w4(32'h3bb8619b),
	.w5(32'h3b9bc199),
	.w6(32'hbb3033ea),
	.w7(32'hbb1285ca),
	.w8(32'hbb376c3e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc95f2),
	.w1(32'h3a34d9a8),
	.w2(32'h39abe2e0),
	.w3(32'hbc271e87),
	.w4(32'h3b03a746),
	.w5(32'h3add8122),
	.w6(32'hba2e1f6c),
	.w7(32'hbb02248e),
	.w8(32'h3953823b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69e6eb),
	.w1(32'hbbdfbe71),
	.w2(32'hbbe27f59),
	.w3(32'hbb29dfe9),
	.w4(32'hbc608b34),
	.w5(32'hbcc38a0c),
	.w6(32'h39b73845),
	.w7(32'h3c8937cd),
	.w8(32'h3be9bd9c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db8b74),
	.w1(32'hbc14e3b0),
	.w2(32'hbbe53e82),
	.w3(32'hba4fe53f),
	.w4(32'hbc00989a),
	.w5(32'h3c258343),
	.w6(32'h3c30fc33),
	.w7(32'h3a90f7f1),
	.w8(32'h3b8bd764),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba13066),
	.w1(32'hbb24ed2d),
	.w2(32'hbba42b18),
	.w3(32'hba1e4562),
	.w4(32'h3c4898dc),
	.w5(32'h3a11108f),
	.w6(32'hba6f14cd),
	.w7(32'h3c06fb75),
	.w8(32'h3baa3c15),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59fd0a),
	.w1(32'hbb4eac34),
	.w2(32'h3c13592b),
	.w3(32'hbb925c64),
	.w4(32'h3a7235b4),
	.w5(32'h3b13be4d),
	.w6(32'hba676314),
	.w7(32'hbb5c0886),
	.w8(32'h3bcf3a73),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce4b0),
	.w1(32'hbb19b1ca),
	.w2(32'h3b5a6d6e),
	.w3(32'hba82fcc0),
	.w4(32'hba6d4437),
	.w5(32'h3b4db7f8),
	.w6(32'h3950a7b7),
	.w7(32'hbb4b84c6),
	.w8(32'h39e1c7ae),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ef7e6),
	.w1(32'h3bc0cfdd),
	.w2(32'hbaa8af86),
	.w3(32'hbb8905dc),
	.w4(32'h3b7121a7),
	.w5(32'hbb09a5d9),
	.w6(32'h3b8b23bc),
	.w7(32'hbb8fdfd8),
	.w8(32'hbbb10251),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c027d),
	.w1(32'hbac50130),
	.w2(32'hbc3628d1),
	.w3(32'hbc429a52),
	.w4(32'hbbb01ab2),
	.w5(32'h3a60c692),
	.w6(32'hb8f0cfee),
	.w7(32'h3a79efc5),
	.w8(32'hba78e8dc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07eff8),
	.w1(32'h3b743a23),
	.w2(32'h3c3b112b),
	.w3(32'hbbf4358d),
	.w4(32'h3c0bffb3),
	.w5(32'h3aacbcd9),
	.w6(32'h3a15ad8d),
	.w7(32'h3c10c953),
	.w8(32'h3ae69f9e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0d9da),
	.w1(32'h3bead5f0),
	.w2(32'hbb47a67d),
	.w3(32'hbaf7c84f),
	.w4(32'h3b9991eb),
	.w5(32'hbab967ca),
	.w6(32'h3ae0bc45),
	.w7(32'h3bcd2aa9),
	.w8(32'h3bdb8c26),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a43b5),
	.w1(32'h3bf3f378),
	.w2(32'hbb3fe204),
	.w3(32'h3b2eb874),
	.w4(32'h3b7cafd8),
	.w5(32'hbc067802),
	.w6(32'h3b6df214),
	.w7(32'h3c4ce1b9),
	.w8(32'h3b9912f0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa77ac),
	.w1(32'hbc2397a3),
	.w2(32'hbc40165d),
	.w3(32'h3c008f51),
	.w4(32'h3b57cbad),
	.w5(32'hbb825871),
	.w6(32'h3c2ffba1),
	.w7(32'h3b38cf40),
	.w8(32'hba17b4e4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c9e75),
	.w1(32'hbb9790a7),
	.w2(32'h3b770b5e),
	.w3(32'hbc53b532),
	.w4(32'hbb45dc85),
	.w5(32'h3b486c64),
	.w6(32'hbbb21556),
	.w7(32'h39f1971e),
	.w8(32'hba504f58),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e4679),
	.w1(32'hbbf2f68c),
	.w2(32'hbbd6fe44),
	.w3(32'hbaef2897),
	.w4(32'hbb375957),
	.w5(32'hbb8b6eb8),
	.w6(32'h3b9eed80),
	.w7(32'hbb6e8cf9),
	.w8(32'h39f99141),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1994),
	.w1(32'hbb670d24),
	.w2(32'hbc05aa3e),
	.w3(32'hbb28f7db),
	.w4(32'hbc27b27b),
	.w5(32'hbbc816c8),
	.w6(32'h3c03d697),
	.w7(32'h3c5bb298),
	.w8(32'h3bd7d986),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb117),
	.w1(32'hbb884b26),
	.w2(32'hbb31817a),
	.w3(32'hbbbd8f56),
	.w4(32'hba753078),
	.w5(32'hbc6419c3),
	.w6(32'h3b8171d8),
	.w7(32'h3c3e89eb),
	.w8(32'h3bcd0ef1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c078d),
	.w1(32'hbbfdf967),
	.w2(32'hba863970),
	.w3(32'h3b79656b),
	.w4(32'h3b52d54e),
	.w5(32'h3b6c04d6),
	.w6(32'hba84a442),
	.w7(32'h3b07b65a),
	.w8(32'hbb8422a7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c186f),
	.w1(32'h3ab55d5a),
	.w2(32'hbb231ed4),
	.w3(32'hbac84f09),
	.w4(32'h3b959ef6),
	.w5(32'hbb0f2dae),
	.w6(32'h3bcdf791),
	.w7(32'h3ba30b26),
	.w8(32'h3bf2d2f1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f357),
	.w1(32'h3b43065f),
	.w2(32'h3c15ea8e),
	.w3(32'hbb90d79c),
	.w4(32'h3b0288c3),
	.w5(32'hbc0f439f),
	.w6(32'hbab680ad),
	.w7(32'hbb20e622),
	.w8(32'hbb20c03d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98cc88),
	.w1(32'hbbc74553),
	.w2(32'hbb9365ca),
	.w3(32'h3b8a32c6),
	.w4(32'hbb0a727f),
	.w5(32'h3c08b433),
	.w6(32'hb98d6599),
	.w7(32'h3b513f68),
	.w8(32'hbb3a84e0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1572c2),
	.w1(32'h3b7b8cb3),
	.w2(32'h3b615d2c),
	.w3(32'hbc1d8233),
	.w4(32'h3b3d974a),
	.w5(32'h3b4d18f9),
	.w6(32'hbb8f1dd6),
	.w7(32'h3bd21f47),
	.w8(32'h3b373fef),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06353c),
	.w1(32'hbb89631e),
	.w2(32'hbc04781b),
	.w3(32'h3b098a8e),
	.w4(32'h3b46c784),
	.w5(32'h3aea3b6a),
	.w6(32'h3ae732b4),
	.w7(32'h3b592c2f),
	.w8(32'hbb78a983),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3b416),
	.w1(32'h3b7c559b),
	.w2(32'hbae5197d),
	.w3(32'hbba1f7a8),
	.w4(32'hbb845fa5),
	.w5(32'hbc1c7eb5),
	.w6(32'hbb93abe7),
	.w7(32'hbbee350a),
	.w8(32'h3ae9f1b6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6683),
	.w1(32'h39899a2d),
	.w2(32'hbbf7ab7d),
	.w3(32'h3b6f9933),
	.w4(32'h3c86eee0),
	.w5(32'hbc27a761),
	.w6(32'h3c82b002),
	.w7(32'h3adb2202),
	.w8(32'hbb79caf1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba165352),
	.w1(32'hba31cbc6),
	.w2(32'h3ab0fe2c),
	.w3(32'hbb009161),
	.w4(32'hb993aa1c),
	.w5(32'hba8c15bc),
	.w6(32'h3c126240),
	.w7(32'h3bd98ddb),
	.w8(32'hba94aa46),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da454),
	.w1(32'hbc06675b),
	.w2(32'hbc06c24d),
	.w3(32'hba67a467),
	.w4(32'hbb3c379f),
	.w5(32'h3b46c431),
	.w6(32'h3b35f6e2),
	.w7(32'h3a79b95e),
	.w8(32'hbc21feeb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba296a2),
	.w1(32'hbc3b9863),
	.w2(32'hbbcd87a6),
	.w3(32'h3b81043a),
	.w4(32'h3b6b8272),
	.w5(32'h3bd02365),
	.w6(32'hbb1c1abb),
	.w7(32'hbb6c2236),
	.w8(32'hbaae6200),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae72ba),
	.w1(32'h3b7cd589),
	.w2(32'h3b6488a1),
	.w3(32'hbbf9f90e),
	.w4(32'h3c15cbad),
	.w5(32'hbb84babd),
	.w6(32'h3a87825f),
	.w7(32'h3be091a7),
	.w8(32'h3a262658),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14284e),
	.w1(32'hbc096afb),
	.w2(32'hbc84bff8),
	.w3(32'hb9146c43),
	.w4(32'hbb564997),
	.w5(32'h3b924c8a),
	.w6(32'hbb225179),
	.w7(32'hbbe6ff7f),
	.w8(32'h3b215a49),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0df9),
	.w1(32'hb9dd89e9),
	.w2(32'h3b9924ba),
	.w3(32'hbbc6711f),
	.w4(32'hbb0c7a14),
	.w5(32'hbb119c63),
	.w6(32'hbc057985),
	.w7(32'hba3576c3),
	.w8(32'h3b15181b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f79a3),
	.w1(32'hbb9bdb87),
	.w2(32'hbbdb0094),
	.w3(32'hbba3ef18),
	.w4(32'hbc0908e6),
	.w5(32'hbc454613),
	.w6(32'h3a84d3f9),
	.w7(32'hbbb344ce),
	.w8(32'hbb2353f9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34a50),
	.w1(32'hbb08d910),
	.w2(32'hbbea8371),
	.w3(32'hbae4f730),
	.w4(32'hbbbfa696),
	.w5(32'h3b430f4e),
	.w6(32'h3a5dcb89),
	.w7(32'hba2035a6),
	.w8(32'h3b233ac6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6087f9),
	.w1(32'h3b9fec63),
	.w2(32'h3b9fb1fa),
	.w3(32'h3a922b01),
	.w4(32'hbadc4231),
	.w5(32'h3bbc52e9),
	.w6(32'h3b833c1b),
	.w7(32'hbaf7c120),
	.w8(32'h3ac43eba),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149aff),
	.w1(32'h39e734a5),
	.w2(32'hb9a1ee89),
	.w3(32'hb9c48b3f),
	.w4(32'hba3bc30a),
	.w5(32'hbb567a16),
	.w6(32'hba6df7fa),
	.w7(32'h3a6460bb),
	.w8(32'hbbaf2fff),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb218ca3),
	.w1(32'hba632ba3),
	.w2(32'h3bd1c53d),
	.w3(32'hbc2f4010),
	.w4(32'h3afa8583),
	.w5(32'h3acf5513),
	.w6(32'hbbb920fc),
	.w7(32'h398396b0),
	.w8(32'h3a96a30c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b547eb8),
	.w1(32'hbbb55201),
	.w2(32'h3b9ec52e),
	.w3(32'hbac86d9d),
	.w4(32'hba030b9b),
	.w5(32'hbbd7e5d0),
	.w6(32'h3a284f17),
	.w7(32'hbb9b0ce0),
	.w8(32'h3b887f65),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cd171),
	.w1(32'h3bb9e9ae),
	.w2(32'h3a0d3653),
	.w3(32'hbaadb8b3),
	.w4(32'h3b3ff873),
	.w5(32'hbc4d5bb9),
	.w6(32'hba5a9f91),
	.w7(32'h39f1d9c6),
	.w8(32'h3ae78f78),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f964ec),
	.w1(32'hbb7f978c),
	.w2(32'hbabafd36),
	.w3(32'hbbb3eb39),
	.w4(32'h3ba94c44),
	.w5(32'h3be2a7cb),
	.w6(32'hbbda99e6),
	.w7(32'hbc2b2f46),
	.w8(32'hbbde5081),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad969a0),
	.w1(32'hbad98ac8),
	.w2(32'hbb5db392),
	.w3(32'hbafca89d),
	.w4(32'hb8f5246d),
	.w5(32'h3aa14afd),
	.w6(32'h3b9d4d6e),
	.w7(32'hbb52d3b9),
	.w8(32'h3aa1e820),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cab3b),
	.w1(32'h3bfcd63f),
	.w2(32'hbb1e5be9),
	.w3(32'hbc17a01e),
	.w4(32'h3b5c4091),
	.w5(32'hbb701787),
	.w6(32'hbbb4c681),
	.w7(32'h3c4d8562),
	.w8(32'h3b59397c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule