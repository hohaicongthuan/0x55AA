module layer_6_featuremap_91(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d222c51),
	.w1(32'hbc23cd18),
	.w2(32'hbc3da716),
	.w3(32'h3b7c0637),
	.w4(32'h3c48091f),
	.w5(32'h3bd52804),
	.w6(32'h3b80e9f2),
	.w7(32'h3bd7fb8c),
	.w8(32'h3b54c969),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11f335),
	.w1(32'h3abc9d46),
	.w2(32'h3bc099aa),
	.w3(32'hbb18561d),
	.w4(32'hbc1c62ad),
	.w5(32'hbbde2bf4),
	.w6(32'h3bc48504),
	.w7(32'hbb133870),
	.w8(32'h3b1ce4af),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3c807),
	.w1(32'hbc859acf),
	.w2(32'hbd19787d),
	.w3(32'h3c2ffd78),
	.w4(32'h3cb76043),
	.w5(32'h3b9c5fdf),
	.w6(32'h3c672da8),
	.w7(32'h3afdd6a5),
	.w8(32'hbc83a299),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37ee6c),
	.w1(32'h3b592c9e),
	.w2(32'h3c4f939e),
	.w3(32'hbb7d23cf),
	.w4(32'hbb8ed5f7),
	.w5(32'hbb6e17f0),
	.w6(32'h3b051650),
	.w7(32'h3be9e44c),
	.w8(32'h3bd57b58),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ccfec),
	.w1(32'hbcd68d03),
	.w2(32'hbd60322a),
	.w3(32'hbb2890fa),
	.w4(32'h3c3a47ee),
	.w5(32'h3a3edd59),
	.w6(32'hbcd1ed41),
	.w7(32'hbc9109cf),
	.w8(32'hbc800eae),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1afe0a),
	.w1(32'hbc4ce00c),
	.w2(32'hbc31628a),
	.w3(32'h3b41ec63),
	.w4(32'h3c80d745),
	.w5(32'h3c831914),
	.w6(32'hb9ba2d20),
	.w7(32'h3c08a65c),
	.w8(32'h3c2770ed),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e926),
	.w1(32'h3c060666),
	.w2(32'h3cb6a73e),
	.w3(32'hbcdfe697),
	.w4(32'hbd0583c9),
	.w5(32'hbcf4b7d9),
	.w6(32'hbbd07632),
	.w7(32'hbbbdb305),
	.w8(32'hbc10b7da),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1eec0),
	.w1(32'h3cb16d61),
	.w2(32'h3d0c661c),
	.w3(32'hbcff9b08),
	.w4(32'hbcabbc8c),
	.w5(32'h3bc56647),
	.w6(32'h3a98b79e),
	.w7(32'h3c0c6367),
	.w8(32'h3c46a39b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca43e7e),
	.w1(32'hbc4011b0),
	.w2(32'hbccbd138),
	.w3(32'hbc4ec34d),
	.w4(32'hbc31c0f6),
	.w5(32'h3b73156d),
	.w6(32'hbcdf8424),
	.w7(32'hbd302c2e),
	.w8(32'hbc2de257),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44c021),
	.w1(32'hbcabac5d),
	.w2(32'hbcc0accb),
	.w3(32'h3a22f5fa),
	.w4(32'h3bd1a874),
	.w5(32'h3b8673e1),
	.w6(32'hbc1eeded),
	.w7(32'hbc3a6db8),
	.w8(32'hbc3f90ae),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5cfb9),
	.w1(32'h3a012964),
	.w2(32'h3be38fce),
	.w3(32'h3c2fa4f3),
	.w4(32'h3c9ce670),
	.w5(32'h3bac6f1e),
	.w6(32'h3c9aa725),
	.w7(32'h3cf9bf9e),
	.w8(32'hbb3fc950),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0adf2d),
	.w1(32'h3b984c35),
	.w2(32'hbc9a939f),
	.w3(32'h3b859640),
	.w4(32'h3c5f656c),
	.w5(32'h3c664c2e),
	.w6(32'hbb8daacc),
	.w7(32'hbc0ce5df),
	.w8(32'hbc2ce996),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc800d1d),
	.w1(32'hbbde55c1),
	.w2(32'h3c330086),
	.w3(32'hbbec9143),
	.w4(32'h3bdd7e42),
	.w5(32'hbc1a376e),
	.w6(32'h3b0841c3),
	.w7(32'h3c75c351),
	.w8(32'h3aefb12c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37bcc9),
	.w1(32'h3b0c68a2),
	.w2(32'hbc0deb6d),
	.w3(32'hbbb043d9),
	.w4(32'hbc8c1a0c),
	.w5(32'hbbb4a633),
	.w6(32'hbcb2c19e),
	.w7(32'hbcd5d0d3),
	.w8(32'hbc08e6f3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dfa63),
	.w1(32'hbbc742e9),
	.w2(32'hbbd56100),
	.w3(32'h3bb0efba),
	.w4(32'h3c133748),
	.w5(32'h3bb45927),
	.w6(32'h3a973853),
	.w7(32'h3c1605a5),
	.w8(32'h3beee621),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba39ae1),
	.w1(32'h39d0bc90),
	.w2(32'h3b71c892),
	.w3(32'h381ee8f1),
	.w4(32'h3ba8ac0e),
	.w5(32'h3c120037),
	.w6(32'h3bc5de18),
	.w7(32'h3c42c16b),
	.w8(32'h3c38eb1d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936dd5e),
	.w1(32'h3cc8b449),
	.w2(32'h3cdae706),
	.w3(32'h3c84376e),
	.w4(32'h3ca65ba3),
	.w5(32'h3c86d52f),
	.w6(32'h3ce9568a),
	.w7(32'h3cf18eeb),
	.w8(32'h3cb2d5e2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbfcd2d),
	.w1(32'hbc04163b),
	.w2(32'hbc197e65),
	.w3(32'h3ba227e3),
	.w4(32'h3beac479),
	.w5(32'h3bb57d51),
	.w6(32'h3b30413b),
	.w7(32'hba08c03a),
	.w8(32'hbb88ef56),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48b176),
	.w1(32'h3ace0006),
	.w2(32'h3bd8841a),
	.w3(32'hbb83f83b),
	.w4(32'hbb5b7dcc),
	.w5(32'hbb2ddfe8),
	.w6(32'h3addf036),
	.w7(32'h3bc7907c),
	.w8(32'h3b921891),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c282),
	.w1(32'h3ca44ce7),
	.w2(32'h3c7aadd1),
	.w3(32'hbada133f),
	.w4(32'h3c929831),
	.w5(32'h3bcdb91e),
	.w6(32'h3c3aa0c4),
	.w7(32'h3c40706b),
	.w8(32'h3bddc002),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8443b8),
	.w1(32'h3bc2a201),
	.w2(32'h3bd5a55d),
	.w3(32'h3ac860fe),
	.w4(32'hbb13ff8f),
	.w5(32'hba065b2a),
	.w6(32'h3b4b2748),
	.w7(32'h3b1b230c),
	.w8(32'h3af75e9e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969376),
	.w1(32'h3bee06ea),
	.w2(32'h3c029ef7),
	.w3(32'h3b164bd9),
	.w4(32'h3bdf5c7f),
	.w5(32'h3b8180fb),
	.w6(32'h3bc2d7e2),
	.w7(32'h3bb52a47),
	.w8(32'h3b9ffb74),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c666198),
	.w1(32'hbcb6b1c4),
	.w2(32'hbb0d9520),
	.w3(32'h3b5fd394),
	.w4(32'h3c124268),
	.w5(32'h39e020cf),
	.w6(32'hbc32beb3),
	.w7(32'hbc300c8c),
	.w8(32'hbc048179),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badcd26),
	.w1(32'hbc1ee9f4),
	.w2(32'h3c599c45),
	.w3(32'hbc3c22eb),
	.w4(32'hbd1e36f4),
	.w5(32'hbca5263d),
	.w6(32'hbd018385),
	.w7(32'hbccd05bf),
	.w8(32'hbc3f6863),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5927cd),
	.w1(32'hbc201420),
	.w2(32'hbcc4ba79),
	.w3(32'hbb1cb56c),
	.w4(32'hbab61d10),
	.w5(32'h3c0fd2f3),
	.w6(32'hbc86cb5a),
	.w7(32'hbd0d0697),
	.w8(32'hbc6b12e6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc071a),
	.w1(32'h3b23e02c),
	.w2(32'h3c0e73fe),
	.w3(32'h3bdac332),
	.w4(32'h3c8526d4),
	.w5(32'h3b605eb1),
	.w6(32'hbbcddb48),
	.w7(32'h3c02f8a3),
	.w8(32'h387b2acb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bd94c),
	.w1(32'hbb8af4fa),
	.w2(32'hbbda3a9b),
	.w3(32'hbaadca56),
	.w4(32'h3c017958),
	.w5(32'h3ade9e6e),
	.w6(32'h3cb2a724),
	.w7(32'h3c8b7f3a),
	.w8(32'hbaa2f388),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf51eb),
	.w1(32'h3c38143d),
	.w2(32'h3cb90a24),
	.w3(32'hbca29005),
	.w4(32'hbca76c52),
	.w5(32'hbc5351f3),
	.w6(32'hbaf38cf3),
	.w7(32'h3b8f63a9),
	.w8(32'h3b54c085),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c800a99),
	.w1(32'h3afb8d30),
	.w2(32'h3b092702),
	.w3(32'hbb7ae8fe),
	.w4(32'hbbadba26),
	.w5(32'hbb19a005),
	.w6(32'hba9c315e),
	.w7(32'hbaffa266),
	.w8(32'hb9a2cb5f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8637ec),
	.w1(32'hbbaa9d3d),
	.w2(32'hbbc70b87),
	.w3(32'hbcbd2405),
	.w4(32'hbc16e52c),
	.w5(32'h3bf506e8),
	.w6(32'hbcfc6d9b),
	.w7(32'hbcfe3dc6),
	.w8(32'hbc850d06),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb24e7a),
	.w1(32'hbc847586),
	.w2(32'h3c6c34ef),
	.w3(32'hbd0d8cb7),
	.w4(32'hbbf04852),
	.w5(32'h3b04047b),
	.w6(32'h39c2c0d0),
	.w7(32'h3d521ead),
	.w8(32'h3d47b55f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2c242),
	.w1(32'hbce3e10a),
	.w2(32'hbcef1021),
	.w3(32'h3c0f94c1),
	.w4(32'h3cb3a481),
	.w5(32'h3c8db913),
	.w6(32'h3c414806),
	.w7(32'h3cc73280),
	.w8(32'h3c345c76),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb8293),
	.w1(32'h3c2e6c4c),
	.w2(32'h3bb6dc9d),
	.w3(32'hb98e08d7),
	.w4(32'h3c22fa2a),
	.w5(32'h3a27d542),
	.w6(32'hbbb1b4af),
	.w7(32'hbba6b7cf),
	.w8(32'h3b68e9c8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5d0b),
	.w1(32'h3c36fb62),
	.w2(32'h3cabc008),
	.w3(32'h3c6820c8),
	.w4(32'h3c91dd21),
	.w5(32'h3c2264d0),
	.w6(32'h3c8234ad),
	.w7(32'h3c473145),
	.w8(32'h3c422bfe),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86736d),
	.w1(32'hbc5494d7),
	.w2(32'hbc7065bc),
	.w3(32'h3c51c581),
	.w4(32'h3c7fbb58),
	.w5(32'h3c67cc44),
	.w6(32'hbba0c8ac),
	.w7(32'hbb96b37a),
	.w8(32'h3a6fbbc3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd87828),
	.w1(32'hba83a931),
	.w2(32'hba5ba30f),
	.w3(32'h3c0e70a2),
	.w4(32'h3ba5b8e6),
	.w5(32'hbbc0757c),
	.w6(32'h3bf3abb7),
	.w7(32'h3c357d82),
	.w8(32'h3c11af0c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941641),
	.w1(32'hbbde841c),
	.w2(32'hbbba4d59),
	.w3(32'h3c0aaf1e),
	.w4(32'h3c99e9b0),
	.w5(32'h3b978e67),
	.w6(32'h3be742c2),
	.w7(32'h3cac63d6),
	.w8(32'h3c286b03),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb832423),
	.w1(32'h3bd23df4),
	.w2(32'h3c0ba6f1),
	.w3(32'h3ad48858),
	.w4(32'hbb07afff),
	.w5(32'hbb3b5ba2),
	.w6(32'h3b864bf1),
	.w7(32'h3b042ae0),
	.w8(32'h39f8935c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d7ac3),
	.w1(32'hbc683e59),
	.w2(32'hbcdfe1a7),
	.w3(32'h3c448e76),
	.w4(32'hbbf3f5f5),
	.w5(32'hbc9e8b6e),
	.w6(32'hbbe29a15),
	.w7(32'hbccccbb7),
	.w8(32'hbcfa096f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc751bed),
	.w1(32'hbc1bbf4f),
	.w2(32'hbc6c60c4),
	.w3(32'h3c4c9f40),
	.w4(32'h3c1f95e3),
	.w5(32'h3c1fa43e),
	.w6(32'h3adaa16a),
	.w7(32'h3bbe69da),
	.w8(32'h3b88437c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fca33),
	.w1(32'hbc85ce11),
	.w2(32'h3bf5b495),
	.w3(32'hbb8f4221),
	.w4(32'h3b9b8f6a),
	.w5(32'hbb703399),
	.w6(32'hbc8f7dde),
	.w7(32'hbbbb126b),
	.w8(32'hbae7ecc3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb34173),
	.w1(32'h3c1cd721),
	.w2(32'h3c8e3168),
	.w3(32'hb9bb1e27),
	.w4(32'h3810ebe6),
	.w5(32'hba8306e0),
	.w6(32'h3bbb8d57),
	.w7(32'h3c24bef6),
	.w8(32'h3bc528e9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f27b4),
	.w1(32'hbb6ebc03),
	.w2(32'hbc205cd7),
	.w3(32'h3c24725c),
	.w4(32'h3c8ee6bd),
	.w5(32'h3c7f4223),
	.w6(32'h3bb29f1d),
	.w7(32'h3b59d5c0),
	.w8(32'hbb46c589),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5d39),
	.w1(32'h3b357d16),
	.w2(32'h3c24902b),
	.w3(32'h3a82dcba),
	.w4(32'h3b8935a0),
	.w5(32'hbb90844d),
	.w6(32'h3b31e78d),
	.w7(32'h3c1690d8),
	.w8(32'hbb27f100),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68a120),
	.w1(32'hba8b7bd8),
	.w2(32'hbaf8eb79),
	.w3(32'h3ba75833),
	.w4(32'h3ad2a908),
	.w5(32'h3a9c988d),
	.w6(32'h3ae70cd1),
	.w7(32'hbb73a964),
	.w8(32'hb91610d1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe158d),
	.w1(32'hbc485a2c),
	.w2(32'hbcbcdafc),
	.w3(32'h3cd15f00),
	.w4(32'h3cdbb3d1),
	.w5(32'hbb34aa7f),
	.w6(32'h3ca7a15d),
	.w7(32'hbc3f9974),
	.w8(32'hbc7d877d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d151f),
	.w1(32'hbba06ee9),
	.w2(32'h3d160aed),
	.w3(32'hbb9158cf),
	.w4(32'hbbf8316b),
	.w5(32'hbc888299),
	.w6(32'h3baab0ce),
	.w7(32'h3c0a74ed),
	.w8(32'h3c6b2e93),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28bd9c),
	.w1(32'h3cb8292d),
	.w2(32'h3cfef00e),
	.w3(32'h3cb12790),
	.w4(32'h3cb5172b),
	.w5(32'h3c2c5fcb),
	.w6(32'h3c2743b6),
	.w7(32'h3c5cbdbf),
	.w8(32'h3c86f115),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9849e5),
	.w1(32'hb95f2e49),
	.w2(32'h3bc8f27b),
	.w3(32'hbb8fbc55),
	.w4(32'hbadb1ed1),
	.w5(32'h3b7e5472),
	.w6(32'hbb8a9183),
	.w7(32'h3a098a66),
	.w8(32'h3baf2901),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f2cac),
	.w1(32'h3c1a56b5),
	.w2(32'h3c60bc5b),
	.w3(32'h3c3a38f6),
	.w4(32'h3c9d9763),
	.w5(32'hba53469b),
	.w6(32'h3c82ba5d),
	.w7(32'h3c7b0efc),
	.w8(32'h3bbb1c65),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48cfb3),
	.w1(32'hba206932),
	.w2(32'h3c8b6a5e),
	.w3(32'hbb43b4c8),
	.w4(32'hbbd6a033),
	.w5(32'hbc13cafe),
	.w6(32'h3998a731),
	.w7(32'h3bc63752),
	.w8(32'hbb7f3bc1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c4ea8),
	.w1(32'h3b1d608e),
	.w2(32'h3c19df37),
	.w3(32'hbb6c406b),
	.w4(32'hbb96d3eb),
	.w5(32'hbb64cb25),
	.w6(32'h3afd8e8e),
	.w7(32'h3a957518),
	.w8(32'h3bb19c78),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e1f5),
	.w1(32'h3c0e1c91),
	.w2(32'h3cb60176),
	.w3(32'hbca7543a),
	.w4(32'hbcd001ae),
	.w5(32'hbc8d538f),
	.w6(32'hbb9eee2b),
	.w7(32'hbb0fdc5e),
	.w8(32'h3ba89f0c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf70b56),
	.w1(32'h3cbc7721),
	.w2(32'h3d024008),
	.w3(32'hbccee58e),
	.w4(32'hbce24a23),
	.w5(32'hbcb76645),
	.w6(32'hbbf8159c),
	.w7(32'hbb43bb95),
	.w8(32'h3b5b35f5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc44f7),
	.w1(32'hbb3f3065),
	.w2(32'h3c4488eb),
	.w3(32'hbc4d069f),
	.w4(32'hbc71d36f),
	.w5(32'hbc7db5ee),
	.w6(32'hbc345098),
	.w7(32'hbc23a311),
	.w8(32'hbc55b84a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c5b21),
	.w1(32'hbc10d886),
	.w2(32'hba1ef12b),
	.w3(32'h3bb3a233),
	.w4(32'h3bbb9047),
	.w5(32'h3aacac95),
	.w6(32'hbbb2715d),
	.w7(32'hbba27015),
	.w8(32'h39d03b46),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd985a),
	.w1(32'hbc7e3509),
	.w2(32'hbccf33a0),
	.w3(32'hbb1971bb),
	.w4(32'hbc00cc14),
	.w5(32'hbb8361e1),
	.w6(32'hbc3e208b),
	.w7(32'hbca68f60),
	.w8(32'hbc63a8ef),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b1df3),
	.w1(32'hba99bd5f),
	.w2(32'h3b0bc7b1),
	.w3(32'h3c012bdb),
	.w4(32'h3c47c9a7),
	.w5(32'h3c5bc249),
	.w6(32'h3b622595),
	.w7(32'h3bff9094),
	.w8(32'h3b589827),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96907b),
	.w1(32'h3c0a0df7),
	.w2(32'h3c6abd5f),
	.w3(32'hbb454f2f),
	.w4(32'h3a044c77),
	.w5(32'h3a83cb69),
	.w6(32'h3b88a7c4),
	.w7(32'h3c183319),
	.w8(32'h3c12a61e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58335b),
	.w1(32'hbc0c08fc),
	.w2(32'hbbb70faf),
	.w3(32'h3c359b46),
	.w4(32'hbb9ee6d2),
	.w5(32'hbb5a16a4),
	.w6(32'hbbb4aaa5),
	.w7(32'hbc225f96),
	.w8(32'h3bd767a1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf9a3e),
	.w1(32'h3b9ff012),
	.w2(32'h3c3327b8),
	.w3(32'hbb5be9bb),
	.w4(32'hbb98ea41),
	.w5(32'hbb764066),
	.w6(32'hbb13b9e7),
	.w7(32'hbb9ccd87),
	.w8(32'hbb1dbcec),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1af163),
	.w1(32'hbc06181e),
	.w2(32'hbb81c304),
	.w3(32'hbb480945),
	.w4(32'h3ba70253),
	.w5(32'h3bc9f448),
	.w6(32'hbb8022d7),
	.w7(32'h3ba0bf00),
	.w8(32'h3b97dfb2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc695302),
	.w1(32'h3c818e22),
	.w2(32'h3c543e57),
	.w3(32'hbb9dd3e5),
	.w4(32'h3a48e2cc),
	.w5(32'h3c2eccf3),
	.w6(32'h3bb95c38),
	.w7(32'h3b96a101),
	.w8(32'h3c3a8d47),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4e38b),
	.w1(32'h3d38577f),
	.w2(32'h3da3cb77),
	.w3(32'hbc814857),
	.w4(32'h3a5b552c),
	.w5(32'hbb7bfed7),
	.w6(32'h3cd2c875),
	.w7(32'h3d71d15d),
	.w8(32'h3d564c3b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule