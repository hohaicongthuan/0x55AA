module layer_10_featuremap_137(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65bd5c),
	.w1(32'h3b42bdfe),
	.w2(32'h3b9dbafa),
	.w3(32'hbc016b07),
	.w4(32'h3c086d3a),
	.w5(32'h3c45801e),
	.w6(32'h3b7b5614),
	.w7(32'h3ba0f198),
	.w8(32'h3c1773aa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d12d0),
	.w1(32'hbc9c9bc5),
	.w2(32'h3c334281),
	.w3(32'h3c27e24f),
	.w4(32'hbbebdb7e),
	.w5(32'h3ba32f90),
	.w6(32'hbc850766),
	.w7(32'hbb3f721d),
	.w8(32'h3b2798cf),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5961b5),
	.w1(32'hbc4df166),
	.w2(32'h3baed4d3),
	.w3(32'h3b72a307),
	.w4(32'hbbb9e2df),
	.w5(32'h3af68cc2),
	.w6(32'hbba988d9),
	.w7(32'h3b89e10b),
	.w8(32'h3bcb9dc4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5463e),
	.w1(32'hbb717c13),
	.w2(32'hbb38d0fb),
	.w3(32'h3ba6aebf),
	.w4(32'h3c0efc14),
	.w5(32'h3b8b652f),
	.w6(32'hba1f74fd),
	.w7(32'h3b82c0b5),
	.w8(32'h3c7a962c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c518c24),
	.w1(32'hbbb9412e),
	.w2(32'hbb95840a),
	.w3(32'h3c6ebffb),
	.w4(32'hbaf8b772),
	.w5(32'hbb9ab4bf),
	.w6(32'hbc0753ee),
	.w7(32'hbb0cbd9b),
	.w8(32'hba33d806),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f941),
	.w1(32'h3c18b9b2),
	.w2(32'hbabacc41),
	.w3(32'hb7c99a99),
	.w4(32'hba5944d7),
	.w5(32'hbb2b16a8),
	.w6(32'h39ad4eba),
	.w7(32'h3a3d3084),
	.w8(32'hbb917bcf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed2bb),
	.w1(32'hbcdbc6ff),
	.w2(32'hbb85f917),
	.w3(32'hbb3f7d01),
	.w4(32'hbc59f05b),
	.w5(32'hbc2e64da),
	.w6(32'hbc8cc663),
	.w7(32'hbc3aaf88),
	.w8(32'hbc032b27),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4167cb),
	.w1(32'h3cf79002),
	.w2(32'hbc159520),
	.w3(32'hbb96f845),
	.w4(32'h3bf786b2),
	.w5(32'hbc395942),
	.w6(32'h3cab5928),
	.w7(32'hbbe5b6b5),
	.w8(32'hbcc3199b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff27ce),
	.w1(32'h3c3dc821),
	.w2(32'hbc2a0c35),
	.w3(32'hbcb82951),
	.w4(32'h3b61de3e),
	.w5(32'hbbfc731d),
	.w6(32'h3b274656),
	.w7(32'hbba6daa4),
	.w8(32'hbbdc2af1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124283),
	.w1(32'hbd3ce1f3),
	.w2(32'h3b39a9c6),
	.w3(32'hbb196804),
	.w4(32'hbcaa846a),
	.w5(32'h39c6c35c),
	.w6(32'hbd074028),
	.w7(32'hbc15dcea),
	.w8(32'h3c961da7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d41967a),
	.w1(32'h3bafb571),
	.w2(32'h3b70f3df),
	.w3(32'h3cf1ab46),
	.w4(32'hba832b44),
	.w5(32'hbabf6cb5),
	.w6(32'h3c618e03),
	.w7(32'h3c24427d),
	.w8(32'h3adb1124),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902623d),
	.w1(32'h3c2c53ae),
	.w2(32'hbbfaf127),
	.w3(32'hb9f903ba),
	.w4(32'h3bd665d0),
	.w5(32'hbc1eb14c),
	.w6(32'h3c42e0ea),
	.w7(32'h3b893d2e),
	.w8(32'hbbf6873d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf01521),
	.w1(32'h3c864140),
	.w2(32'hbb98201a),
	.w3(32'hbc0c90fa),
	.w4(32'h3b189649),
	.w5(32'hbc2c2481),
	.w6(32'h3c8f9b7c),
	.w7(32'h3a57aaff),
	.w8(32'hbc57eff1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6228eb),
	.w1(32'h3d8b8a60),
	.w2(32'hbac5433f),
	.w3(32'hbc47dd41),
	.w4(32'h3d1aa070),
	.w5(32'hbc0e2c8f),
	.w6(32'h3d6453ab),
	.w7(32'h3c2ecb89),
	.w8(32'hbcf35b20),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd63ef56),
	.w1(32'h3c0ee5e0),
	.w2(32'h3c3956a3),
	.w3(32'hbd45408e),
	.w4(32'h3c882f8f),
	.w5(32'h3bfb1689),
	.w6(32'h3be2ca47),
	.w7(32'h3c5cd7e7),
	.w8(32'h3c312282),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3ba66),
	.w1(32'h3c6b1649),
	.w2(32'hba6e287c),
	.w3(32'hbc22edb2),
	.w4(32'h3b69972b),
	.w5(32'hba4e6f54),
	.w6(32'hb997bf1b),
	.w7(32'hbba2a813),
	.w8(32'hbc02e01b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe61126),
	.w1(32'h3acb312c),
	.w2(32'h3990edf5),
	.w3(32'hba6e919d),
	.w4(32'h3abc3d10),
	.w5(32'h3b097af8),
	.w6(32'h3aca61ff),
	.w7(32'h3b3d93fa),
	.w8(32'hbb806cc1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38124d),
	.w1(32'hbd1d0fda),
	.w2(32'h3bcb6430),
	.w3(32'hbc0f60ff),
	.w4(32'hbcd8b385),
	.w5(32'hbb19c67a),
	.w6(32'hbd179fdf),
	.w7(32'hbcc0771b),
	.w8(32'h3b7d2434),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0979df),
	.w1(32'hbbfaa79e),
	.w2(32'hbb957be6),
	.w3(32'h3c8776d6),
	.w4(32'hbba1512f),
	.w5(32'hbbd6eab5),
	.w6(32'hbc079647),
	.w7(32'hbc742604),
	.w8(32'hbc30816e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf4068),
	.w1(32'h3c1f31a4),
	.w2(32'hbc38a527),
	.w3(32'hba9e6629),
	.w4(32'h3b48475b),
	.w5(32'hbc0da77c),
	.w6(32'h3ba8d0bd),
	.w7(32'hbbb298c0),
	.w8(32'hbbc930c7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bd945),
	.w1(32'h3cc4f74a),
	.w2(32'hbc42a288),
	.w3(32'hbbcdd484),
	.w4(32'h3c21442e),
	.w5(32'hbc336e56),
	.w6(32'h3c647b44),
	.w7(32'hbb94cb87),
	.w8(32'hbc0bc254),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92ed8b),
	.w1(32'h3c4cc96d),
	.w2(32'h3c257c51),
	.w3(32'hbc103096),
	.w4(32'h3bb4bfb7),
	.w5(32'h3c46484a),
	.w6(32'h3cbf80f9),
	.w7(32'h3be5b871),
	.w8(32'h3afcd4ac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb556),
	.w1(32'hbacf4d28),
	.w2(32'hbbd7e989),
	.w3(32'hb9f97242),
	.w4(32'hbb222198),
	.w5(32'hbbe048a4),
	.w6(32'hbc44a3eb),
	.w7(32'hbc679485),
	.w8(32'hbc8e3f62),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e80fb),
	.w1(32'h3d03cce0),
	.w2(32'hbbd87fd0),
	.w3(32'h3c101991),
	.w4(32'h3c56e1bb),
	.w5(32'hbc1057e9),
	.w6(32'h3cbd2899),
	.w7(32'h3aebf881),
	.w8(32'hbca19e8c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3a3fb),
	.w1(32'h3b506617),
	.w2(32'h3b67dc89),
	.w3(32'hbca2737b),
	.w4(32'h3b571b2e),
	.w5(32'hbad0a302),
	.w6(32'h3aa781e0),
	.w7(32'h3bcbdd55),
	.w8(32'h3c37daee),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b848c37),
	.w1(32'h3c4e20d9),
	.w2(32'h3ad45593),
	.w3(32'hb999c160),
	.w4(32'h3c05319f),
	.w5(32'h3b58d88a),
	.w6(32'h3c2c6e88),
	.w7(32'h3c010424),
	.w8(32'hbb22af60),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093a40),
	.w1(32'h3c300c7f),
	.w2(32'hbbd89623),
	.w3(32'hba17a31f),
	.w4(32'h3b11f78a),
	.w5(32'hbbd66442),
	.w6(32'h3bf45236),
	.w7(32'hbafb44c3),
	.w8(32'hbbd27974),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c2c98),
	.w1(32'hbc2d7536),
	.w2(32'hbb07125f),
	.w3(32'hbc394c9f),
	.w4(32'hbc2796b1),
	.w5(32'hbb7e19fe),
	.w6(32'hbc04b4db),
	.w7(32'hb8d28dda),
	.w8(32'h3b8fa616),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd449a3),
	.w1(32'h3be0fc72),
	.w2(32'hbba122a1),
	.w3(32'h3bf94642),
	.w4(32'hb8f5707e),
	.w5(32'hbba326aa),
	.w6(32'h3b461c61),
	.w7(32'hbacb13d2),
	.w8(32'h3bbda805),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4411d2),
	.w1(32'h3ba90013),
	.w2(32'hb973c557),
	.w3(32'hba86b237),
	.w4(32'h3b660576),
	.w5(32'h3a34a672),
	.w6(32'h3bc8ee80),
	.w7(32'h3ae53cb3),
	.w8(32'h3aa89c23),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526a14),
	.w1(32'h3c528197),
	.w2(32'hbc04ba65),
	.w3(32'h3baa097b),
	.w4(32'h3b42b0d9),
	.w5(32'hbc03a257),
	.w6(32'h3c0c80a5),
	.w7(32'hbb5d8859),
	.w8(32'hbc0a9f00),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60bc86),
	.w1(32'h3c94aec0),
	.w2(32'h3a7e7437),
	.w3(32'hbc0feb37),
	.w4(32'h3bda1041),
	.w5(32'hbaba53db),
	.w6(32'h3c6c9d9d),
	.w7(32'h3bb07df0),
	.w8(32'hbb8befd8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc191256),
	.w1(32'h3c1e7892),
	.w2(32'hbcd44cc6),
	.w3(32'hbb84b2f8),
	.w4(32'h3b4951ab),
	.w5(32'hbca21b9b),
	.w6(32'h3c528660),
	.w7(32'hbc46499d),
	.w8(32'hbc342cf2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc689852),
	.w1(32'hbc05ac5f),
	.w2(32'hbb12ca4a),
	.w3(32'hbc2c5cd8),
	.w4(32'hbb1a040d),
	.w5(32'hbb5281e1),
	.w6(32'hbb3aa428),
	.w7(32'hbbfbb4f6),
	.w8(32'hbae43883),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ba69),
	.w1(32'hbd34571f),
	.w2(32'h3c113eba),
	.w3(32'h39e0e221),
	.w4(32'hbcd045e4),
	.w5(32'h3bd4f338),
	.w6(32'hbd163ad9),
	.w7(32'hbbbb9d0f),
	.w8(32'h3ccf63d5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d408a07),
	.w1(32'h3c1fb82f),
	.w2(32'hbbd435ee),
	.w3(32'h3d016df9),
	.w4(32'hba049546),
	.w5(32'hbbeb233a),
	.w6(32'h3c2613cf),
	.w7(32'h3a810ccd),
	.w8(32'hbc1cdab8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc637efb),
	.w1(32'hbc77a2fa),
	.w2(32'h3c890c96),
	.w3(32'h3c2f8adb),
	.w4(32'h3a6b237b),
	.w5(32'h3a714e21),
	.w6(32'hbbedd5eb),
	.w7(32'h3c093eb6),
	.w8(32'h3b07eeab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb65883),
	.w1(32'hbcd41d3d),
	.w2(32'h3be90b5a),
	.w3(32'h3bb39e7a),
	.w4(32'hbbd00aee),
	.w5(32'h3bede395),
	.w6(32'hbcdc9809),
	.w7(32'hbb099fb4),
	.w8(32'h3c08d9de),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21651e),
	.w1(32'h3c888dbb),
	.w2(32'hbc0fcf27),
	.w3(32'hbadb0341),
	.w4(32'h3a8153e4),
	.w5(32'hbc3f11be),
	.w6(32'h3c3faf66),
	.w7(32'hbb3fcc34),
	.w8(32'hbc34ac82),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc922b6a),
	.w1(32'hbc4edc0f),
	.w2(32'h3b886dbd),
	.w3(32'hbc3bd428),
	.w4(32'hbb4f3577),
	.w5(32'h39ebe7f3),
	.w6(32'hbc37bb3c),
	.w7(32'hbb4828da),
	.w8(32'h3b171145),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21a501),
	.w1(32'h3b33b83b),
	.w2(32'h3b5aefd4),
	.w3(32'h3b111519),
	.w4(32'h3abe9d16),
	.w5(32'h3baad7ea),
	.w6(32'h3b43f73b),
	.w7(32'h3af4854d),
	.w8(32'h392a66d1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb0186),
	.w1(32'hbafa1312),
	.w2(32'h3b66ed90),
	.w3(32'h3b44cbb9),
	.w4(32'hba32090f),
	.w5(32'hbad220f5),
	.w6(32'h3a6e17a8),
	.w7(32'h3b97c556),
	.w8(32'h3b674e14),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90de60),
	.w1(32'h3c9c8edc),
	.w2(32'h3b189240),
	.w3(32'hbb3d5fe8),
	.w4(32'h3c0f410e),
	.w5(32'hbb0e9577),
	.w6(32'h3c6b0e96),
	.w7(32'h3bc650ca),
	.w8(32'hbb89a0d9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc741e73),
	.w1(32'hbd5c0eae),
	.w2(32'h3c05e2d8),
	.w3(32'hbc7549ca),
	.w4(32'hbced17bf),
	.w5(32'hbaba7661),
	.w6(32'hbd38152b),
	.w7(32'hbc9a065f),
	.w8(32'h3c5e1503),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3ef7e0),
	.w1(32'h3b2c105b),
	.w2(32'h3c2dc304),
	.w3(32'h3cdcb743),
	.w4(32'h3c2b967f),
	.w5(32'h3bfa24a3),
	.w6(32'h3c2e3282),
	.w7(32'h3bfd6abe),
	.w8(32'hbb0c6bfd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06582d),
	.w1(32'hbc51275f),
	.w2(32'hbbf0cdc1),
	.w3(32'h3b8cf4e2),
	.w4(32'hbb8d8f9f),
	.w5(32'hbb97759a),
	.w6(32'hbaa21632),
	.w7(32'hbbc89dcb),
	.w8(32'hbb91d663),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b076410),
	.w1(32'hbb958cbb),
	.w2(32'hbc174903),
	.w3(32'h3bba9067),
	.w4(32'h3bdff96c),
	.w5(32'h3b6a86ca),
	.w6(32'hbb8e52c0),
	.w7(32'h3b0f67b4),
	.w8(32'hbb08f269),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34e0b),
	.w1(32'h3bad7edf),
	.w2(32'hbc3ce771),
	.w3(32'h3b3e1a83),
	.w4(32'hbb7f11ea),
	.w5(32'hbc9d99ea),
	.w6(32'h3af00a58),
	.w7(32'hbcab9dbc),
	.w8(32'hbc823786),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af27432),
	.w1(32'h3c44aa00),
	.w2(32'hbb24a732),
	.w3(32'h3ac18692),
	.w4(32'h3b9df4d5),
	.w5(32'hbb6bafef),
	.w6(32'h3c36f9fd),
	.w7(32'h3b494138),
	.w8(32'hbb91df53),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42d3b0),
	.w1(32'h3d1f8f5a),
	.w2(32'hbab1f28a),
	.w3(32'hbc0dcf67),
	.w4(32'h3c9fc109),
	.w5(32'hbba73bf5),
	.w6(32'h3ce56d32),
	.w7(32'h3b970b9b),
	.w8(32'hbc994ad5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceba383),
	.w1(32'hbb35ba7e),
	.w2(32'h3bab27aa),
	.w3(32'hbcb6327f),
	.w4(32'h3bed31e2),
	.w5(32'h3b5902fc),
	.w6(32'h3aa7c4dc),
	.w7(32'hb9539386),
	.w8(32'hb9a1a4ef),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fa250),
	.w1(32'h3b9e862c),
	.w2(32'hbc259475),
	.w3(32'hbbd32299),
	.w4(32'hbb56f8ad),
	.w5(32'h39c9f2b7),
	.w6(32'hba47c3cc),
	.w7(32'hbbdf986d),
	.w8(32'h3b5756b5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16319a),
	.w1(32'h3bedd0fa),
	.w2(32'hba2cb2d2),
	.w3(32'h3c41039e),
	.w4(32'h3a1819c2),
	.w5(32'hbab22ae1),
	.w6(32'hba5f5388),
	.w7(32'hb9a4186c),
	.w8(32'hbba72a9d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc655af0),
	.w1(32'hbc9d04b1),
	.w2(32'hbc42e672),
	.w3(32'hbbe14cbd),
	.w4(32'hbc7e7157),
	.w5(32'hbc252735),
	.w6(32'hbc9f2015),
	.w7(32'hbc9b563d),
	.w8(32'hbc3e26c3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5adc5),
	.w1(32'hbc6d9c93),
	.w2(32'hbb1ead59),
	.w3(32'h3b5d453e),
	.w4(32'hbbec9726),
	.w5(32'hb994a01c),
	.w6(32'hbc6b2632),
	.w7(32'hbba54ab4),
	.w8(32'hbb78a034),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d31c4),
	.w1(32'h3bbfd77e),
	.w2(32'hbb78f856),
	.w3(32'h3a360dde),
	.w4(32'h3b220b4b),
	.w5(32'h3aab2919),
	.w6(32'h3b7e584f),
	.w7(32'hbb39f94c),
	.w8(32'hb8b3e3ef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba392ccb),
	.w1(32'h3bb84e16),
	.w2(32'h3b9c71b2),
	.w3(32'h3a590cb1),
	.w4(32'h3c1960e8),
	.w5(32'h3b3e99a9),
	.w6(32'h3c1b8fe4),
	.w7(32'h3a0ab508),
	.w8(32'hbbfc08a9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaf21e),
	.w1(32'h3b5fa617),
	.w2(32'hbc0e7519),
	.w3(32'hbc09aad0),
	.w4(32'h3c241bb8),
	.w5(32'hbbff49fa),
	.w6(32'h3b439d59),
	.w7(32'hbbd29567),
	.w8(32'hbc0cb922),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eea97),
	.w1(32'hbc8f2cb5),
	.w2(32'h3c641e68),
	.w3(32'hbbe03596),
	.w4(32'hbbd8257e),
	.w5(32'h3c09cf2b),
	.w6(32'hbc988b11),
	.w7(32'hbb2e8555),
	.w8(32'h3b8fe08f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c837f4e),
	.w1(32'h3cec843a),
	.w2(32'hbb7f9908),
	.w3(32'h3c10757f),
	.w4(32'h3c29a3fd),
	.w5(32'hbbc171fb),
	.w6(32'h3c995ab0),
	.w7(32'h3ab169e5),
	.w8(32'hbc3f6351),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5f3ce),
	.w1(32'hbc76788b),
	.w2(32'h3ac9e80c),
	.w3(32'hbc632512),
	.w4(32'hbc409e77),
	.w5(32'hbb9a5529),
	.w6(32'hbc5f4c9b),
	.w7(32'hbc29f868),
	.w8(32'hbbe2a4dc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ea3d7),
	.w1(32'h3cd7d33f),
	.w2(32'hbada0ab7),
	.w3(32'hbbefe4cf),
	.w4(32'h3bfe85fd),
	.w5(32'hbb49ce14),
	.w6(32'h3c51e1d2),
	.w7(32'hbb068813),
	.w8(32'hbc236944),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97b76b),
	.w1(32'h3b806a0a),
	.w2(32'hbc989f57),
	.w3(32'hbc5b36f5),
	.w4(32'h3b0baf48),
	.w5(32'hbc173b38),
	.w6(32'hba949b2a),
	.w7(32'hbc16b720),
	.w8(32'h39dc29b0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5aff5),
	.w1(32'hbd299dd9),
	.w2(32'h3bfecca2),
	.w3(32'h3ba4adc3),
	.w4(32'hbc98c016),
	.w5(32'h3b86d20f),
	.w6(32'hbcf7dc94),
	.w7(32'hbbddf9f8),
	.w8(32'h3ca2e95d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d19ee2c),
	.w1(32'hbc172ad6),
	.w2(32'hba8d537f),
	.w3(32'h3cb93260),
	.w4(32'hbba1a545),
	.w5(32'hba32e3e4),
	.w6(32'hbc1d036e),
	.w7(32'hbb951b6c),
	.w8(32'h3b996663),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27764d),
	.w1(32'h3b98d0f5),
	.w2(32'hbc492589),
	.w3(32'h3b4f76f9),
	.w4(32'h3b880d74),
	.w5(32'hbc0f94ef),
	.w6(32'h3ba99498),
	.w7(32'hbc14ba44),
	.w8(32'hbbd3018b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31bdd9),
	.w1(32'h3aa258d8),
	.w2(32'h3aade034),
	.w3(32'hbb0a1862),
	.w4(32'h3b5ae883),
	.w5(32'h3c24f8a4),
	.w6(32'h3a6b625b),
	.w7(32'hbbef3e4f),
	.w8(32'hbbd8b088),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1920a),
	.w1(32'hbc24bda6),
	.w2(32'hbb5b89f2),
	.w3(32'h3b104e6e),
	.w4(32'hbb1f4da3),
	.w5(32'hb8a3e9ac),
	.w6(32'hbb2dd1ec),
	.w7(32'hba1e9a5c),
	.w8(32'hbc106421),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab6407),
	.w1(32'h3c674210),
	.w2(32'hbb870bda),
	.w3(32'h3b99dc14),
	.w4(32'hbb0b0e8c),
	.w5(32'hbb688a7e),
	.w6(32'h3b05a7d7),
	.w7(32'hbb5b63a4),
	.w8(32'hbc1a0d71),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf33430),
	.w1(32'h3b8f39d5),
	.w2(32'hbc67d51a),
	.w3(32'hba9a035b),
	.w4(32'h3bfaca35),
	.w5(32'hbc995507),
	.w6(32'h3c49a0dc),
	.w7(32'hbbd93ef4),
	.w8(32'hbc4386a1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf935b6),
	.w1(32'hbcc30fd3),
	.w2(32'h3c310bf3),
	.w3(32'hbc722e44),
	.w4(32'hbc369e6c),
	.w5(32'h3bd10f0e),
	.w6(32'hbca838d7),
	.w7(32'hbabb0384),
	.w8(32'h3c2d2380),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1c900),
	.w1(32'h3c907dd3),
	.w2(32'hbbd433d1),
	.w3(32'h3c717270),
	.w4(32'h3b7e3f1b),
	.w5(32'hbc00ca66),
	.w6(32'h3c176e68),
	.w7(32'hbb0342ea),
	.w8(32'hbc48e6f4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa0ae3),
	.w1(32'h3cbc1412),
	.w2(32'hbb537cf6),
	.w3(32'hbc66fb08),
	.w4(32'h3c078152),
	.w5(32'hbb837ba1),
	.w6(32'h3c55f724),
	.w7(32'h3a35eab9),
	.w8(32'hbc06519e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84c4e8),
	.w1(32'h3ca3d25f),
	.w2(32'hba9c35bf),
	.w3(32'hbc1ea281),
	.w4(32'h3b5be514),
	.w5(32'hbb6ce936),
	.w6(32'h3c703eda),
	.w7(32'h3abfafa7),
	.w8(32'hbbf0b472),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc497714),
	.w1(32'hbc56c1f5),
	.w2(32'h3c1bb75c),
	.w3(32'hbbae74aa),
	.w4(32'hbc0f2d51),
	.w5(32'h3ab80034),
	.w6(32'hbc8221ac),
	.w7(32'hbb699980),
	.w8(32'h3b45bcb3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb7ce),
	.w1(32'h3c512671),
	.w2(32'hbc499338),
	.w3(32'h3ab67a81),
	.w4(32'h3bea8785),
	.w5(32'hbb8aec3f),
	.w6(32'h3c9174b5),
	.w7(32'h3b61aaae),
	.w8(32'hbbeb64fb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc467e1d),
	.w1(32'h3d3aca26),
	.w2(32'hbc206352),
	.w3(32'hbb59ee2c),
	.w4(32'h3c555028),
	.w5(32'hbc9221f7),
	.w6(32'h3d0e56a1),
	.w7(32'hbbacbc2a),
	.w8(32'hbce4e602),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd23c00f),
	.w1(32'hbb7fd3bb),
	.w2(32'h3b2a82b8),
	.w3(32'hbce6bdc8),
	.w4(32'h3b848198),
	.w5(32'h3b00986e),
	.w6(32'hbb8aaa79),
	.w7(32'hbb801935),
	.w8(32'hbbf5bf45),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8cc8),
	.w1(32'hbaefbcca),
	.w2(32'hbbddfeac),
	.w3(32'h3aba59c9),
	.w4(32'hbab10622),
	.w5(32'hbb857175),
	.w6(32'hbb96edb0),
	.w7(32'hbbe79360),
	.w8(32'hbbda2f19),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3af8),
	.w1(32'h3caa6260),
	.w2(32'hbc8e3a70),
	.w3(32'h3af7fb98),
	.w4(32'h3bcbdc76),
	.w5(32'hbc724c76),
	.w6(32'h3c9e36ff),
	.w7(32'hbbe8ef01),
	.w8(32'hbc593e23),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91e924),
	.w1(32'hbb38e506),
	.w2(32'h3b28467c),
	.w3(32'hbc2873e7),
	.w4(32'hba09ffcf),
	.w5(32'h3b899285),
	.w6(32'hba13daee),
	.w7(32'h3983d833),
	.w8(32'h398eea8d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01b214),
	.w1(32'hbb36f63c),
	.w2(32'h3c1d5cd7),
	.w3(32'h3b6e04b0),
	.w4(32'h3aee049a),
	.w5(32'h3bc18361),
	.w6(32'hbb0416c0),
	.w7(32'hbb14c01e),
	.w8(32'hbb5cebe5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c339bc0),
	.w1(32'h3bdae86d),
	.w2(32'hbab2d476),
	.w3(32'h3b4eff68),
	.w4(32'h3b7a0d9c),
	.w5(32'hbbadf4e6),
	.w6(32'h3b8d55d6),
	.w7(32'h3adb5e28),
	.w8(32'h3b6b96ea),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079e07),
	.w1(32'hbc539a39),
	.w2(32'h3c071427),
	.w3(32'hbb99ecc5),
	.w4(32'hbb889fea),
	.w5(32'h3bd09ee4),
	.w6(32'hbc564618),
	.w7(32'hbb9ec925),
	.w8(32'hba2e87b4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2671b8),
	.w1(32'hbc137791),
	.w2(32'h3ab7b9dc),
	.w3(32'h3b833bc2),
	.w4(32'hbbe10fec),
	.w5(32'hb992e978),
	.w6(32'hbc1e0af6),
	.w7(32'h39f2e779),
	.w8(32'hb8c2b285),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96e88d),
	.w1(32'h3b100206),
	.w2(32'h3bc8e4f8),
	.w3(32'hbb216209),
	.w4(32'h3be26686),
	.w5(32'h3bb207ef),
	.w6(32'h3b7b4ac6),
	.w7(32'h3a7e2dfd),
	.w8(32'hbbd3c8ff),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c6030),
	.w1(32'h3c2d651a),
	.w2(32'h3be43518),
	.w3(32'hbbf999bf),
	.w4(32'h3c9f2c08),
	.w5(32'h3b93a3cd),
	.w6(32'h3c35b3f9),
	.w7(32'h3baa99f8),
	.w8(32'hbc2bd5ff),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc529599),
	.w1(32'h3c6a0214),
	.w2(32'hbb7a1216),
	.w3(32'hbc13678c),
	.w4(32'h3b97f86f),
	.w5(32'hbb83d9d7),
	.w6(32'h3c16cef0),
	.w7(32'hb9a12097),
	.w8(32'hbb86b620),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bdbd5),
	.w1(32'hbc545f29),
	.w2(32'h399e6750),
	.w3(32'hbb9464bc),
	.w4(32'hbaec901b),
	.w5(32'h3abf8668),
	.w6(32'hbc2eaf4b),
	.w7(32'hbb315682),
	.w8(32'hbba24bdc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c698),
	.w1(32'h3ca1663a),
	.w2(32'hbc505715),
	.w3(32'hbba6021d),
	.w4(32'hbad26fe8),
	.w5(32'hbc71d1d4),
	.w6(32'h3bd2354c),
	.w7(32'hbc82cd36),
	.w8(32'hbcadeb9e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92bb59),
	.w1(32'h3c91077a),
	.w2(32'h3a455003),
	.w3(32'hbc374b4c),
	.w4(32'h3bf14539),
	.w5(32'h39e71a81),
	.w6(32'h3c768338),
	.w7(32'h3bbd264d),
	.w8(32'hbb0e02d0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd39f6),
	.w1(32'hbcd4d335),
	.w2(32'hbafcf078),
	.w3(32'h3b0001a4),
	.w4(32'hbc244a3e),
	.w5(32'hbbf48a36),
	.w6(32'hbc831d52),
	.w7(32'hbc238aae),
	.w8(32'hbbe60196),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a3bba),
	.w1(32'hbc834a6a),
	.w2(32'h3bc3bc40),
	.w3(32'h3bafb8a3),
	.w4(32'hbc04f010),
	.w5(32'h3baae042),
	.w6(32'hbc896cde),
	.w7(32'hbb57acf0),
	.w8(32'h3c120759),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f9828),
	.w1(32'h3c16d1c9),
	.w2(32'hbb31cf59),
	.w3(32'h3c639967),
	.w4(32'h3bc417cb),
	.w5(32'h3a416588),
	.w6(32'h3bbad8f3),
	.w7(32'hbbf3a010),
	.w8(32'hbb36731c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20cc26),
	.w1(32'hbc857292),
	.w2(32'h3aae0310),
	.w3(32'h3b88d686),
	.w4(32'hbbd0bc12),
	.w5(32'h39fb8be2),
	.w6(32'hbbb61025),
	.w7(32'h39d19987),
	.w8(32'h3b02c279),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853188),
	.w1(32'hbc02d920),
	.w2(32'hbbdd44a8),
	.w3(32'h3b427e8b),
	.w4(32'hbba47612),
	.w5(32'h3bb530a5),
	.w6(32'hbb6a1a2d),
	.w7(32'hba8003d6),
	.w8(32'h3a994a80),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78da8),
	.w1(32'hbc20fbde),
	.w2(32'hb9944591),
	.w3(32'h3b215c64),
	.w4(32'hba808ae1),
	.w5(32'h3adf49fb),
	.w6(32'hbbbe7a21),
	.w7(32'hbb81b348),
	.w8(32'h3b20ee09),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ca833),
	.w1(32'h3a7ed97d),
	.w2(32'hbcbf53a0),
	.w3(32'h3c3ea414),
	.w4(32'hbb7bfdf5),
	.w5(32'hbc9b9d68),
	.w6(32'hbbc41c25),
	.w7(32'hbcde3f2b),
	.w8(32'h3a27b866),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85cc25),
	.w1(32'hbc497502),
	.w2(32'h3b3ec14c),
	.w3(32'h3cd084f9),
	.w4(32'hb9e83586),
	.w5(32'h3b5dee06),
	.w6(32'hbbc1f278),
	.w7(32'hbbcec34f),
	.w8(32'hbbf1e63e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cda98),
	.w1(32'h3c09aa4f),
	.w2(32'h3c228dd9),
	.w3(32'h3b306892),
	.w4(32'h3c098daa),
	.w5(32'h3b806800),
	.w6(32'h39cd39a0),
	.w7(32'h3b89e7cb),
	.w8(32'h3b3e9844),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f6f12),
	.w1(32'h3a7dd1df),
	.w2(32'hbbab555b),
	.w3(32'h3bd6c6e7),
	.w4(32'h3cab184f),
	.w5(32'h3bba7fb7),
	.w6(32'h38bcd3f7),
	.w7(32'h3b4df344),
	.w8(32'h3c8153e2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52eaa6),
	.w1(32'hbbcc9421),
	.w2(32'hbc80a089),
	.w3(32'h3bd2984e),
	.w4(32'hbbff8162),
	.w5(32'hbbe20a50),
	.w6(32'hbb383c6d),
	.w7(32'hbbf5f16a),
	.w8(32'hbc7ed90d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919444),
	.w1(32'h3d9107c7),
	.w2(32'hbc93cc55),
	.w3(32'h3c2fd1d5),
	.w4(32'h3d03ffbe),
	.w5(32'hbccf9905),
	.w6(32'h3d69e334),
	.w7(32'h3b58dc03),
	.w8(32'hbd1f6897),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd64a7b3),
	.w1(32'h3c9836a1),
	.w2(32'hbb446cca),
	.w3(32'hbd1f805c),
	.w4(32'h3bcd3ab1),
	.w5(32'hbb8a7110),
	.w6(32'h3c0d7d25),
	.w7(32'h3ab35c62),
	.w8(32'hbc2e7504),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf6c2f3),
	.w1(32'h3d16fe8c),
	.w2(32'hbc1aea3c),
	.w3(32'hbc8dda8f),
	.w4(32'h3c99a264),
	.w5(32'hbc3df184),
	.w6(32'h3cdf1de8),
	.w7(32'hbac1d39f),
	.w8(32'hbcc74a2a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6557f),
	.w1(32'h3c0d6d78),
	.w2(32'hbca19c24),
	.w3(32'hbc7f5654),
	.w4(32'h3b652c15),
	.w5(32'hbc966f59),
	.w6(32'h3c35fac2),
	.w7(32'hbb5d9717),
	.w8(32'hbc427ebc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55484b),
	.w1(32'hbc591350),
	.w2(32'h3bde408a),
	.w3(32'hbc0605bc),
	.w4(32'hbba4e572),
	.w5(32'h3bd25243),
	.w6(32'hbc113198),
	.w7(32'h3ac5c8bf),
	.w8(32'h3bedd7df),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c197605),
	.w1(32'h3c94ac11),
	.w2(32'hbb98dd51),
	.w3(32'h3bc6dec2),
	.w4(32'h3c047dbc),
	.w5(32'hbb6daff2),
	.w6(32'h3c2690be),
	.w7(32'hbac1578c),
	.w8(32'hbc170282),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25f33a),
	.w1(32'h3d1eb768),
	.w2(32'hbc0f72c0),
	.w3(32'hbb9de63c),
	.w4(32'h3c690784),
	.w5(32'hbc6e6658),
	.w6(32'h3ce5b632),
	.w7(32'hbb074034),
	.w8(32'hbcbe26b9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec080f),
	.w1(32'hbb920215),
	.w2(32'h3c5e6c41),
	.w3(32'hbca7bf50),
	.w4(32'h3b949ab5),
	.w5(32'h3bf95ab6),
	.w6(32'h3b0b24dc),
	.w7(32'h3befc96f),
	.w8(32'hb9ea2bec),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5363c),
	.w1(32'h3c85b7ee),
	.w2(32'hbba4f3c1),
	.w3(32'hba63a089),
	.w4(32'h3b91962a),
	.w5(32'hbb4e6032),
	.w6(32'h3c3105c7),
	.w7(32'hbb3370f5),
	.w8(32'hbafe729a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb81830),
	.w1(32'h3c976b36),
	.w2(32'h3b62bcb6),
	.w3(32'h3acd83bc),
	.w4(32'h3c687f11),
	.w5(32'h3bff1db9),
	.w6(32'h3c38c046),
	.w7(32'h3be7c92a),
	.w8(32'hbb25c40d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0c79),
	.w1(32'h3c9662bb),
	.w2(32'h3bd94aa2),
	.w3(32'h3aa86a65),
	.w4(32'h3c037cb2),
	.w5(32'h3b6ca47b),
	.w6(32'h3be39d18),
	.w7(32'h3c1a9183),
	.w8(32'h3b2f0b9b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc284cd3),
	.w1(32'hbc3f1b98),
	.w2(32'h3c38af45),
	.w3(32'hba694252),
	.w4(32'hbba8711c),
	.w5(32'h3b9ddee4),
	.w6(32'hbc23fd05),
	.w7(32'h3a81fc99),
	.w8(32'h3b53eaba),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c274ddb),
	.w1(32'h3d0fd38b),
	.w2(32'h3b8e690f),
	.w3(32'hba374941),
	.w4(32'h3cc19b15),
	.w5(32'h3a753495),
	.w6(32'h3ce0b454),
	.w7(32'h3c3c128f),
	.w8(32'hbc32e720),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf6581),
	.w1(32'h3d4aeeed),
	.w2(32'hbc484c5f),
	.w3(32'hbc9a27f1),
	.w4(32'h3ca74161),
	.w5(32'hbc63776d),
	.w6(32'h3d14c7f5),
	.w7(32'h3ad06264),
	.w8(32'hbcbb1a5d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2c4788),
	.w1(32'h3ccb8990),
	.w2(32'hbbd4d0f3),
	.w3(32'hbcf2fcab),
	.w4(32'h3c012c25),
	.w5(32'hbc097edd),
	.w6(32'h3c8290c6),
	.w7(32'h39c699c5),
	.w8(32'hbc756382),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcbade),
	.w1(32'h3ccfff32),
	.w2(32'hbbae2d5a),
	.w3(32'hbc85d8ee),
	.w4(32'h3becf701),
	.w5(32'hbbd49011),
	.w6(32'h3c842f64),
	.w7(32'h3af65081),
	.w8(32'hbc2b7ed2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca08e7e),
	.w1(32'h3c62eaed),
	.w2(32'h3aa8d0f6),
	.w3(32'hbc42e044),
	.w4(32'h3b0057fb),
	.w5(32'hbab94663),
	.w6(32'h3c8d853d),
	.w7(32'h3b6df10f),
	.w8(32'hbbd7ed65),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22e5f0),
	.w1(32'hbc2d6f15),
	.w2(32'hbc6a4cc1),
	.w3(32'hbb9fa347),
	.w4(32'h3a98fae1),
	.w5(32'hbc4aec38),
	.w6(32'hbb36a454),
	.w7(32'hbc5f9cf1),
	.w8(32'hbbb9f67b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a790f),
	.w1(32'h3c3f27ad),
	.w2(32'hba34e400),
	.w3(32'hbaf46bf9),
	.w4(32'h3b2dbb6c),
	.w5(32'hbb2c3f38),
	.w6(32'h3c078b02),
	.w7(32'h3b19ecc5),
	.w8(32'hbbf44e8b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc266cb3),
	.w1(32'h3c264529),
	.w2(32'hbbd7d1ea),
	.w3(32'hbbd2f84d),
	.w4(32'h3b790706),
	.w5(32'hbbf663e8),
	.w6(32'h3bea0376),
	.w7(32'hbbbc655e),
	.w8(32'hbc1c704e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2186a8),
	.w1(32'h3d093ac6),
	.w2(32'hbaeeda20),
	.w3(32'hbc1d1735),
	.w4(32'h3c45e93d),
	.w5(32'hbbb3f1f4),
	.w6(32'h3ca9e572),
	.w7(32'h3b0bc488),
	.w8(32'hbc80bd5e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcfe76),
	.w1(32'hba164de6),
	.w2(32'hbb7f04fb),
	.w3(32'hbc9aa553),
	.w4(32'hb8d80373),
	.w5(32'h3bc09562),
	.w6(32'h3b02f4ed),
	.w7(32'hbb239037),
	.w8(32'h39cbbf52),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2da2ed),
	.w1(32'h3b5ed730),
	.w2(32'h3bd90507),
	.w3(32'h3ba9793c),
	.w4(32'hbac7642f),
	.w5(32'h3be8fd69),
	.w6(32'hbb8bdb8f),
	.w7(32'h3b86320d),
	.w8(32'h3aee82ae),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28692),
	.w1(32'h3ca29566),
	.w2(32'hbc12cfbe),
	.w3(32'hb916e095),
	.w4(32'h3bb94a5e),
	.w5(32'hbc0a2bf2),
	.w6(32'h3c62c493),
	.w7(32'hbb1a2ee5),
	.w8(32'hbbe0c642),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61130b),
	.w1(32'h3976e7fe),
	.w2(32'h395b2c56),
	.w3(32'hbbdd75d5),
	.w4(32'h37da37bb),
	.w5(32'hb989efb1),
	.w6(32'hb6a3e2d4),
	.w7(32'hb8eb5363),
	.w8(32'hb9357d7f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1311a1),
	.w1(32'hbb69390d),
	.w2(32'hbb879006),
	.w3(32'h3a27270b),
	.w4(32'hbb61e593),
	.w5(32'hbc09d070),
	.w6(32'h3b0fd800),
	.w7(32'hb9afc953),
	.w8(32'hbc061db4),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8472c6),
	.w1(32'h39a46922),
	.w2(32'hbb85d9ad),
	.w3(32'hb9dd4938),
	.w4(32'hbb9249e5),
	.w5(32'hbbb06654),
	.w6(32'hbaf33852),
	.w7(32'hbbfd95dd),
	.w8(32'hbc09b433),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a213e92),
	.w1(32'h3a1349a0),
	.w2(32'hb9c4ae29),
	.w3(32'h3ab1ec7c),
	.w4(32'h39c2b493),
	.w5(32'hba26c2e8),
	.w6(32'h3a3b62a7),
	.w7(32'hba2e36b2),
	.w8(32'hbaa947e0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011bb9),
	.w1(32'hbb2099df),
	.w2(32'hb953d557),
	.w3(32'hbadde55d),
	.w4(32'hbb03737b),
	.w5(32'hba9eb3ba),
	.w6(32'hba5c508e),
	.w7(32'hbad78ca9),
	.w8(32'hbb0fa79d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2acd35),
	.w1(32'hb9219fb7),
	.w2(32'hb98d6353),
	.w3(32'h38df7a3b),
	.w4(32'h39a4936d),
	.w5(32'h38522f85),
	.w6(32'h3a13d454),
	.w7(32'h39838a5e),
	.w8(32'hb9aca09f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01db8e),
	.w1(32'h3a806d96),
	.w2(32'h39afc91f),
	.w3(32'h39de0bf7),
	.w4(32'hb7ec0d71),
	.w5(32'h3884b3d7),
	.w6(32'hb8ee99e3),
	.w7(32'hba960d4b),
	.w8(32'hbafa076b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbff695),
	.w1(32'hbaaa6262),
	.w2(32'hba0072e6),
	.w3(32'hbad6b6ef),
	.w4(32'h3b550259),
	.w5(32'h3aef1dbb),
	.w6(32'h3af9652b),
	.w7(32'h3aac80cf),
	.w8(32'hba5111bd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eba32),
	.w1(32'hba2028ba),
	.w2(32'hbbafe13f),
	.w3(32'h3a75119c),
	.w4(32'hbb7fbf49),
	.w5(32'hbbaaaadb),
	.w6(32'hbb07c024),
	.w7(32'hbc38fd3a),
	.w8(32'hbc4b39be),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9999373),
	.w1(32'hb95d4370),
	.w2(32'h3a97007e),
	.w3(32'hb98ccb42),
	.w4(32'h3a9cbd91),
	.w5(32'h3a76590f),
	.w6(32'h3a651d3c),
	.w7(32'h3b0f877e),
	.w8(32'h3aebbbfb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16299e),
	.w1(32'h3aafa365),
	.w2(32'hbac65c70),
	.w3(32'h3accfffd),
	.w4(32'h3b19a7e8),
	.w5(32'hbaf392e5),
	.w6(32'hbaa54df3),
	.w7(32'hb83f88f2),
	.w8(32'hbb881b73),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ee44e),
	.w1(32'hba981d39),
	.w2(32'hbb8c70ee),
	.w3(32'h3adf545c),
	.w4(32'hbb397dec),
	.w5(32'hbbc39798),
	.w6(32'hba064665),
	.w7(32'hbbbbd9c0),
	.w8(32'hbc123e90),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26020e),
	.w1(32'h3ad356c7),
	.w2(32'h3b0bf316),
	.w3(32'hba2902bb),
	.w4(32'h3b33dae6),
	.w5(32'h3b018a38),
	.w6(32'h39a8b611),
	.w7(32'h3b71385c),
	.w8(32'h3b0e7caa),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0e974),
	.w1(32'h3aa9e35b),
	.w2(32'hb835ab5c),
	.w3(32'h3b6a146e),
	.w4(32'h39d142f7),
	.w5(32'hbb1f061a),
	.w6(32'h3a7746ce),
	.w7(32'hbb3eb2a8),
	.w8(32'hbbd839ea),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed2909),
	.w1(32'h39e3117a),
	.w2(32'hb92500a5),
	.w3(32'h399cb000),
	.w4(32'h39dd1402),
	.w5(32'hb93d01fc),
	.w6(32'h3998d930),
	.w7(32'h38561d0a),
	.w8(32'hba3698dc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18056c),
	.w1(32'hbb0a3014),
	.w2(32'h3ad877a4),
	.w3(32'h3b2c549f),
	.w4(32'hbb165098),
	.w5(32'hbb4d7dce),
	.w6(32'h3b78ec56),
	.w7(32'h398f27e8),
	.w8(32'hbaaaa8c3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b71d42),
	.w1(32'h39e17c88),
	.w2(32'hba6a3af6),
	.w3(32'hb9d3f37b),
	.w4(32'h398b3aae),
	.w5(32'hba162c20),
	.w6(32'hba8d6dc5),
	.w7(32'hbae43c33),
	.w8(32'hbb09c6e7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8182510),
	.w1(32'hb8ebec4c),
	.w2(32'hb8ae3ce0),
	.w3(32'hb7930fb4),
	.w4(32'hb83dabb3),
	.w5(32'hb887fd79),
	.w6(32'h38a60226),
	.w7(32'hb772faa3),
	.w8(32'hb8b40c5c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79174ae),
	.w1(32'hb8a663cf),
	.w2(32'hb89b500b),
	.w3(32'h37a954b0),
	.w4(32'hb5d97c02),
	.w5(32'hb87e028f),
	.w6(32'h3752139b),
	.w7(32'h379e0cdd),
	.w8(32'hb7ac050a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e79a88),
	.w1(32'h39dc8e9a),
	.w2(32'hb9344bdd),
	.w3(32'h3a910ca3),
	.w4(32'h3a120b73),
	.w5(32'hba4459e6),
	.w6(32'h3aa3adce),
	.w7(32'h3a33ddb9),
	.w8(32'h3988d4fe),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2e4b),
	.w1(32'h38846535),
	.w2(32'hb9a54a9e),
	.w3(32'hb9b05b20),
	.w4(32'h3b39acd0),
	.w5(32'h3a3415d8),
	.w6(32'h39d80ef8),
	.w7(32'h3ad871bc),
	.w8(32'hba8d22c3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc7e57),
	.w1(32'hba46fc1f),
	.w2(32'hbb22c00e),
	.w3(32'h39634b5d),
	.w4(32'hbb42e483),
	.w5(32'hbb70f7dd),
	.w6(32'h3b0453fb),
	.w7(32'hbb15f60a),
	.w8(32'hbb3be51c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b042db),
	.w1(32'hb82a8f14),
	.w2(32'h375f7e55),
	.w3(32'hb8049bc5),
	.w4(32'hb733ff73),
	.w5(32'h37e9f677),
	.w6(32'hb7679a89),
	.w7(32'h37667f9d),
	.w8(32'h37f215bf),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7529816),
	.w1(32'hba4f42b2),
	.w2(32'hbb481b3c),
	.w3(32'h3b0299b3),
	.w4(32'hbb096d2e),
	.w5(32'hbb67d0a7),
	.w6(32'hba3d760e),
	.w7(32'hbba5dc8e),
	.w8(32'hbbda1935),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac68e99),
	.w1(32'hb9b879bd),
	.w2(32'hba958360),
	.w3(32'h3aad6552),
	.w4(32'hba7166a7),
	.w5(32'hbb361da4),
	.w6(32'h3a030930),
	.w7(32'hbae2a0dc),
	.w8(32'hbb618333),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39458a1b),
	.w1(32'hb8e232b2),
	.w2(32'hbafd8a2d),
	.w3(32'h3b9070bb),
	.w4(32'h3a313345),
	.w5(32'hbb351364),
	.w6(32'h3b16b14e),
	.w7(32'hbb82094a),
	.w8(32'hbbb57e67),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed9342),
	.w1(32'hbbe94bfd),
	.w2(32'hbbc7ddf4),
	.w3(32'h3abdf258),
	.w4(32'hbb3bbb80),
	.w5(32'hbbf43a5f),
	.w6(32'h3a91db01),
	.w7(32'hbb7bf0d6),
	.w8(32'hbb3da4b9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b6ea0),
	.w1(32'h39d6dc96),
	.w2(32'h3a59a819),
	.w3(32'h3919dcb9),
	.w4(32'h3a887f51),
	.w5(32'h39b54b15),
	.w6(32'h39823085),
	.w7(32'h3945462b),
	.w8(32'hb69f5c0b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b015cd3),
	.w1(32'h3af39b5c),
	.w2(32'h3b0dd20f),
	.w3(32'h3b16b3a2),
	.w4(32'h3b22a312),
	.w5(32'h3afbfd20),
	.w6(32'h3b26445a),
	.w7(32'h3af0c667),
	.w8(32'h3aa845e7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c34ce),
	.w1(32'hb9edccfd),
	.w2(32'hba224ab6),
	.w3(32'hba992b06),
	.w4(32'h3a3c3f1f),
	.w5(32'hb8afbbbb),
	.w6(32'hb9b112a8),
	.w7(32'h3af525e3),
	.w8(32'h3a146215),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4009c9),
	.w1(32'hba6bae47),
	.w2(32'h39bfd901),
	.w3(32'hbab37c12),
	.w4(32'h3b164812),
	.w5(32'h3ad58c59),
	.w6(32'hbaf10af3),
	.w7(32'h37d3a05f),
	.w8(32'h3a87a733),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a145c5),
	.w1(32'h39d9efdd),
	.w2(32'h3ae66860),
	.w3(32'hb8daa918),
	.w4(32'h3ad92b2b),
	.w5(32'h3b384b1e),
	.w6(32'h3a14a6b4),
	.w7(32'h3b0ed23c),
	.w8(32'h3b3ecb6d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3552cdc4),
	.w1(32'hb9e3e385),
	.w2(32'hb9d8c71d),
	.w3(32'h39e9f8d8),
	.w4(32'hba4f36a8),
	.w5(32'hba8c7714),
	.w6(32'hb95d81a9),
	.w7(32'hbaf5cba1),
	.w8(32'hbb2217aa),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93354f6),
	.w1(32'hb880efec),
	.w2(32'h370db1ea),
	.w3(32'h3900c124),
	.w4(32'h390c5ecc),
	.w5(32'h389c0e91),
	.w6(32'hb904ccb4),
	.w7(32'hb862d8bb),
	.w8(32'hb921e06a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa108d),
	.w1(32'hb955f1de),
	.w2(32'hbb1c4049),
	.w3(32'h3b560922),
	.w4(32'hb9c0623a),
	.w5(32'hbb3e847c),
	.w6(32'h3aede982),
	.w7(32'hbb39a7fc),
	.w8(32'hbbadc3e5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bce7f),
	.w1(32'hbab86472),
	.w2(32'hbaf9d402),
	.w3(32'h3a3ff96e),
	.w4(32'hba9af542),
	.w5(32'hbb0361d3),
	.w6(32'h3a847c10),
	.w7(32'hb983e32b),
	.w8(32'hb9237f9c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba844ff6),
	.w1(32'hba636f49),
	.w2(32'hba28dd1c),
	.w3(32'hbacb35f6),
	.w4(32'hba907e0e),
	.w5(32'h3900e47f),
	.w6(32'hbaa1f998),
	.w7(32'h38e7bebb),
	.w8(32'hb9c0bc4d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39907e85),
	.w1(32'h390525fb),
	.w2(32'h36974b40),
	.w3(32'h390203fd),
	.w4(32'h38ac1224),
	.w5(32'h38f2064d),
	.w6(32'h394dfa48),
	.w7(32'h39ed8eac),
	.w8(32'h39770436),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10e220),
	.w1(32'h3a968569),
	.w2(32'hb9b9bd6e),
	.w3(32'h3bfec9ca),
	.w4(32'h3946907d),
	.w5(32'hba90a37e),
	.w6(32'h3bc9de2e),
	.w7(32'hbaafa01f),
	.w8(32'hbb8e4ca3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d6177),
	.w1(32'h39839f64),
	.w2(32'h39e73518),
	.w3(32'h397a20de),
	.w4(32'h39d6365a),
	.w5(32'h3a3e7dc0),
	.w6(32'h39eb0f0d),
	.w7(32'h3a04b01a),
	.w8(32'h3a15084f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39515b80),
	.w1(32'hb99a3cbb),
	.w2(32'hba03f6f9),
	.w3(32'h3917f112),
	.w4(32'hb9933894),
	.w5(32'hb9ecc5f3),
	.w6(32'h38128cfc),
	.w7(32'hba0fedac),
	.w8(32'hba0ae955),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22f525),
	.w1(32'hb75d7973),
	.w2(32'hb90823d6),
	.w3(32'h39bf608b),
	.w4(32'h3b139e75),
	.w5(32'h3acd5e1e),
	.w6(32'h39b794d1),
	.w7(32'h3b053946),
	.w8(32'h3afa40d3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36471),
	.w1(32'hbacf7ce8),
	.w2(32'hbb4b78de),
	.w3(32'h3b65ddf9),
	.w4(32'hbb081d93),
	.w5(32'hbbb98bcd),
	.w6(32'hba6ede4c),
	.w7(32'hbbaec8db),
	.w8(32'hbc1a3d58),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926cd84),
	.w1(32'h39d350b9),
	.w2(32'h3a03de0a),
	.w3(32'h395b6b25),
	.w4(32'h3a05ded3),
	.w5(32'hb80cfaa0),
	.w6(32'h39c879e8),
	.w7(32'h3a134694),
	.w8(32'hb8e0e550),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bc800),
	.w1(32'h3a0401f2),
	.w2(32'h3a7be7f1),
	.w3(32'h3a5e59b2),
	.w4(32'h3a94838a),
	.w5(32'hb89179eb),
	.w6(32'h3b310c3b),
	.w7(32'h3afa2103),
	.w8(32'h39ac5442),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f8b3a),
	.w1(32'h39b8a8dd),
	.w2(32'hbabbeb49),
	.w3(32'hbaa082df),
	.w4(32'hba067e3a),
	.w5(32'hbaa8fffb),
	.w6(32'hba90e9a9),
	.w7(32'hba3bd9b6),
	.w8(32'hba2f6fa2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb776c99),
	.w1(32'hbb4349e0),
	.w2(32'hbb5b8566),
	.w3(32'hbbc576d9),
	.w4(32'hbc111cfe),
	.w5(32'hbbad4d72),
	.w6(32'hbbc4c1c4),
	.w7(32'hbc05b710),
	.w8(32'hbb99a644),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f3f31),
	.w1(32'hbab15b4f),
	.w2(32'hbb41bbe0),
	.w3(32'h3a8cfb31),
	.w4(32'h38a0e039),
	.w5(32'hba7fe320),
	.w6(32'h3a3d7fbf),
	.w7(32'hbaa5b4dc),
	.w8(32'hbb141495),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27172e),
	.w1(32'hb9bd64a4),
	.w2(32'hbb4098ab),
	.w3(32'hba227fb2),
	.w4(32'hbb3ef165),
	.w5(32'hbb6b591e),
	.w6(32'hbb2dcb28),
	.w7(32'hbbf440a9),
	.w8(32'hbc038706),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f200f7),
	.w1(32'h3a4012ca),
	.w2(32'h3a3172d7),
	.w3(32'h3a806c7f),
	.w4(32'h3a729294),
	.w5(32'h3a85df68),
	.w6(32'h3a509444),
	.w7(32'h3a7e06bd),
	.w8(32'h3a6ab9b2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ac608),
	.w1(32'h37d94ef4),
	.w2(32'hbaa25f72),
	.w3(32'h3aa37c4c),
	.w4(32'h3ac51c34),
	.w5(32'h39ade68e),
	.w6(32'h3a58b8e7),
	.w7(32'h38df84d4),
	.w8(32'hba98d0ff),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7647012),
	.w1(32'hb7d3d535),
	.w2(32'hb76b43c9),
	.w3(32'h352f7ddf),
	.w4(32'hb8092378),
	.w5(32'hb71ef94a),
	.w6(32'h382921f9),
	.w7(32'h368f8d9e),
	.w8(32'h3823f6ea),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a166e),
	.w1(32'h39c17b2c),
	.w2(32'h393645c4),
	.w3(32'h3941c050),
	.w4(32'hb9b6f155),
	.w5(32'hb4fb3658),
	.w6(32'hb7c38147),
	.w7(32'hba49cc23),
	.w8(32'hb98c7dd3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e5f16),
	.w1(32'h39ce01bb),
	.w2(32'h3a418318),
	.w3(32'h39849e92),
	.w4(32'h39d89fa1),
	.w5(32'h3a302685),
	.w6(32'hb8c4430d),
	.w7(32'h3982f46b),
	.w8(32'h3a2fe19e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39484b),
	.w1(32'hba645147),
	.w2(32'hba12e74b),
	.w3(32'hbb251b36),
	.w4(32'hbabd73a8),
	.w5(32'hba37480f),
	.w6(32'hbb2073f3),
	.w7(32'hbb73a18d),
	.w8(32'hbb3bac9d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7830813),
	.w1(32'h3630ba6f),
	.w2(32'h37749082),
	.w3(32'hb7932a18),
	.w4(32'h370bb20c),
	.w5(32'h37c51c14),
	.w6(32'hb751823c),
	.w7(32'h374fbd11),
	.w8(32'h37a5d8d8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7376142),
	.w1(32'hb80ec675),
	.w2(32'hb80f776b),
	.w3(32'h3809af77),
	.w4(32'h38df26e2),
	.w5(32'hb7ed753b),
	.w6(32'h38579c05),
	.w7(32'h3715fc7b),
	.w8(32'hb91841e7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930ffe1),
	.w1(32'hb983f757),
	.w2(32'h39f72cb4),
	.w3(32'hba2cc980),
	.w4(32'h398d7085),
	.w5(32'h39efe3ff),
	.w6(32'hbaa2ebd4),
	.w7(32'hba9f28da),
	.w8(32'hbab4fb98),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c664b9),
	.w1(32'hbb0506cb),
	.w2(32'hbbe4fa97),
	.w3(32'hb943f116),
	.w4(32'h392bd61e),
	.w5(32'hbbf47cca),
	.w6(32'h3aa66a69),
	.w7(32'hbadc4ef1),
	.w8(32'hbbfd3edc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb613ff6),
	.w1(32'h39e5b548),
	.w2(32'h3a81483e),
	.w3(32'h3b51038c),
	.w4(32'h3b49066a),
	.w5(32'hba89ec55),
	.w6(32'h3b14585f),
	.w7(32'h39bd7647),
	.w8(32'hbba456b5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e65208),
	.w1(32'hba7ab2a8),
	.w2(32'hba50424e),
	.w3(32'hb9b9ed98),
	.w4(32'hba2161cb),
	.w5(32'hb945b666),
	.w6(32'hb9ff7e7c),
	.w7(32'hba616e9a),
	.w8(32'hb967907d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4543fb),
	.w1(32'hbb88d858),
	.w2(32'hbbc813ff),
	.w3(32'hbab9b3a9),
	.w4(32'hbc028f1f),
	.w5(32'hbc2e6cad),
	.w6(32'h3b3552d2),
	.w7(32'hbbaeaed2),
	.w8(32'hbbd7e899),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb420834),
	.w1(32'hbb15fcfb),
	.w2(32'h3a72068e),
	.w3(32'hb792db78),
	.w4(32'h3b71a2ea),
	.w5(32'h3b4c1b02),
	.w6(32'hb91f952c),
	.w7(32'hb9d19ae2),
	.w8(32'h39eacbdf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab53bdd),
	.w1(32'hba2b7459),
	.w2(32'hbb1a7a93),
	.w3(32'h3b1a9f45),
	.w4(32'hba868b99),
	.w5(32'hbb220a46),
	.w6(32'h3b138ea1),
	.w7(32'hba868050),
	.w8(32'hbb57d5e6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eee099),
	.w1(32'hb8bbd18d),
	.w2(32'hb7dc21b2),
	.w3(32'hb8e1336e),
	.w4(32'hb8bfff84),
	.w5(32'hb88966f6),
	.w6(32'hb830208f),
	.w7(32'hb8ae2f3b),
	.w8(32'hb84ec956),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e80da8),
	.w1(32'hb8e572f6),
	.w2(32'hb8d63ae6),
	.w3(32'hb8e7e29b),
	.w4(32'hb8eb46a4),
	.w5(32'hb98e9b9d),
	.w6(32'hb91ce36e),
	.w7(32'hb981baea),
	.w8(32'hb9cb4fa5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c85b84),
	.w1(32'h35ac41ba),
	.w2(32'h3725a725),
	.w3(32'h37f0bea1),
	.w4(32'hb7a0614b),
	.w5(32'hb7cad340),
	.w6(32'hb7d18fdd),
	.w7(32'hb8177584),
	.w8(32'h36995613),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46de1c),
	.w1(32'h3a262c3b),
	.w2(32'hbb057b82),
	.w3(32'h3b803b62),
	.w4(32'hb96d3be6),
	.w5(32'hbb907f83),
	.w6(32'h3b388477),
	.w7(32'hb981f471),
	.w8(32'hbbba329a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ebab9d),
	.w1(32'hbb1220b9),
	.w2(32'hbad26f37),
	.w3(32'h3acaec08),
	.w4(32'hba7aeb6e),
	.w5(32'hbac512d9),
	.w6(32'hba67e97b),
	.w7(32'hbba280d5),
	.w8(32'hbbbc2168),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae66062),
	.w1(32'h393b3cd9),
	.w2(32'hb99d51e4),
	.w3(32'hb9ff33bd),
	.w4(32'h3b0c8913),
	.w5(32'h392d8db4),
	.w6(32'h3a927437),
	.w7(32'h3b0202ce),
	.w8(32'h3a2781f2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea265b),
	.w1(32'hba2ff171),
	.w2(32'h37855ffb),
	.w3(32'h380864f7),
	.w4(32'hb9c4d8f1),
	.w5(32'h391e8e02),
	.w6(32'hb9e91502),
	.w7(32'hb9d850df),
	.w8(32'hb82d95f8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56868c),
	.w1(32'h3ae62aea),
	.w2(32'hbb015ea9),
	.w3(32'h3b4e648e),
	.w4(32'hbaa66589),
	.w5(32'hbbc42bf7),
	.w6(32'h3b1544ab),
	.w7(32'hbb5bc835),
	.w8(32'hbc0066dd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba942181),
	.w1(32'hba92e975),
	.w2(32'hbb0f0e45),
	.w3(32'hba24db07),
	.w4(32'h3a0509ec),
	.w5(32'hbb36ec62),
	.w6(32'hba56a934),
	.w7(32'h3b16dc24),
	.w8(32'hbaa2d8b3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77d2b89),
	.w1(32'h378e5bd7),
	.w2(32'h385a088c),
	.w3(32'hb703d453),
	.w4(32'h37f43150),
	.w5(32'h3882cd1d),
	.w6(32'h36170274),
	.w7(32'h38185723),
	.w8(32'h3880acbe),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a8c26),
	.w1(32'h397de65c),
	.w2(32'hbab449ed),
	.w3(32'hbb6a5cad),
	.w4(32'hba93e007),
	.w5(32'hbaffefab),
	.w6(32'hbaf53144),
	.w7(32'h3a0a3f9d),
	.w8(32'hbaaf47f1),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81faf03),
	.w1(32'hb86a9c88),
	.w2(32'h380a1b23),
	.w3(32'hb7e9e7e8),
	.w4(32'hb7a3b00b),
	.w5(32'h387c2a62),
	.w6(32'h37f15171),
	.w7(32'h379a2530),
	.w8(32'h38bdc7cf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ef463),
	.w1(32'h3b4f0e8c),
	.w2(32'hba97d052),
	.w3(32'hb99d049b),
	.w4(32'h3a0f77bb),
	.w5(32'hbb28e1fb),
	.w6(32'h3af977da),
	.w7(32'h3a8c7306),
	.w8(32'hbb96236f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb019b),
	.w1(32'hbae65d5c),
	.w2(32'hb9d1c602),
	.w3(32'hba8f4e62),
	.w4(32'h3af9261f),
	.w5(32'h3b2382af),
	.w6(32'hbb2ef089),
	.w7(32'hba4d187e),
	.w8(32'h39e10d02),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53eeda),
	.w1(32'h37a11f43),
	.w2(32'hba1ad32e),
	.w3(32'h3a97f960),
	.w4(32'h3a989ddc),
	.w5(32'hba6519ec),
	.w6(32'h3a44fa92),
	.w7(32'h3a2e612d),
	.w8(32'hba93adb7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a0c8a),
	.w1(32'h3923777c),
	.w2(32'h397daeae),
	.w3(32'hba2eadd6),
	.w4(32'h399b13f6),
	.w5(32'h38acdc2a),
	.w6(32'hba8a206a),
	.w7(32'hb920f945),
	.w8(32'hb8769ea8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a511ba),
	.w1(32'h3912583f),
	.w2(32'h3ab75c73),
	.w3(32'hb9c474a2),
	.w4(32'h3b44db4c),
	.w5(32'h3aafab77),
	.w6(32'h3a58cb48),
	.w7(32'h3b16f855),
	.w8(32'hb92aa39e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20042),
	.w1(32'h3977e245),
	.w2(32'hba3faa46),
	.w3(32'h3a093c36),
	.w4(32'hba4a9bc5),
	.w5(32'hbabe09b1),
	.w6(32'h3799bf77),
	.w7(32'hbb0a9ab7),
	.w8(32'hbb77c963),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0614),
	.w1(32'hbb29203e),
	.w2(32'hbb83f6b2),
	.w3(32'hba3089b0),
	.w4(32'hbb57ae36),
	.w5(32'hbba3c6cc),
	.w6(32'h3ab6de77),
	.w7(32'hbb315dd1),
	.w8(32'hbb4cdb18),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a67881),
	.w1(32'h37ba9c9b),
	.w2(32'h376cb6d5),
	.w3(32'h38828313),
	.w4(32'h37b63723),
	.w5(32'hb84ed459),
	.w6(32'h389df88c),
	.w7(32'hb7f55d04),
	.w8(32'hb8c860c1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394479c5),
	.w1(32'hb954f760),
	.w2(32'h37df3bb0),
	.w3(32'hb7c375f1),
	.w4(32'hb92bbba7),
	.w5(32'hb9087d0c),
	.w6(32'hb838bec0),
	.w7(32'hb9c62e3c),
	.w8(32'hb808143d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c16a),
	.w1(32'hbb88566b),
	.w2(32'hbb9a7b25),
	.w3(32'h3bad67d6),
	.w4(32'hbaeff4fe),
	.w5(32'hbbe22135),
	.w6(32'h3b951b1d),
	.w7(32'hba86102c),
	.w8(32'hbc00f8b1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26f542),
	.w1(32'hbb89b399),
	.w2(32'hbbaafaf1),
	.w3(32'h3ac629da),
	.w4(32'hbb90f899),
	.w5(32'hbbcb754d),
	.w6(32'hbaa79002),
	.w7(32'hbbdf8ecf),
	.w8(32'hbc3b58cd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f3c5c),
	.w1(32'h390dacfa),
	.w2(32'hba47b638),
	.w3(32'h3a69f3de),
	.w4(32'h3aec3aad),
	.w5(32'hba80d725),
	.w6(32'h3a1226d6),
	.w7(32'h37b6bf66),
	.w8(32'hbb43704d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cedb6b),
	.w1(32'h3a30ef04),
	.w2(32'hbb588bd4),
	.w3(32'h3baeb6fe),
	.w4(32'h3b06f537),
	.w5(32'hba7d1cd5),
	.w6(32'h3bf84f0e),
	.w7(32'h3a0bd971),
	.w8(32'hbb1776cd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33b2a4),
	.w1(32'hb9ed6d18),
	.w2(32'hb866599e),
	.w3(32'hb993aef2),
	.w4(32'hba3da75c),
	.w5(32'hb9aa0b95),
	.w6(32'hba22d69a),
	.w7(32'hba2c0b25),
	.w8(32'hba0f5fa6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a8a0c),
	.w1(32'hbad48d31),
	.w2(32'hbab3e51b),
	.w3(32'hba075f48),
	.w4(32'hba6f8aec),
	.w5(32'hba1f55a2),
	.w6(32'hb904c137),
	.w7(32'h37faa448),
	.w8(32'h38858c84),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6e30),
	.w1(32'h3a3d7362),
	.w2(32'hbbd75039),
	.w3(32'h3b4c4b7d),
	.w4(32'hbb47c00c),
	.w5(32'hbc5b5b27),
	.w6(32'h398330dd),
	.w7(32'hb93e86a7),
	.w8(32'hbc63e7d3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67f25),
	.w1(32'hbb17ef3d),
	.w2(32'hbbbe22ca),
	.w3(32'hbb64ad44),
	.w4(32'hbbe0180a),
	.w5(32'hbbeae633),
	.w6(32'hba89addc),
	.w7(32'hbc1316b9),
	.w8(32'hbc04d278),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c3dbd),
	.w1(32'h3ba688e2),
	.w2(32'h3b11fed9),
	.w3(32'h3bc3f605),
	.w4(32'h3b17a22a),
	.w5(32'hbb68b0ee),
	.w6(32'h3b43324b),
	.w7(32'hba6e7ab8),
	.w8(32'hbc05571c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66d5a7),
	.w1(32'hbaad7473),
	.w2(32'hb9c2c653),
	.w3(32'hbb2df846),
	.w4(32'hbaa59a4c),
	.w5(32'h3a6f713f),
	.w6(32'hbb0d4077),
	.w7(32'h395df30e),
	.w8(32'h3b011810),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac497a),
	.w1(32'hbb6c7f5a),
	.w2(32'hba6a7c09),
	.w3(32'hbb8ef74e),
	.w4(32'h38ed8d6b),
	.w5(32'h3a80563d),
	.w6(32'hbb05a39b),
	.w7(32'hbaadda47),
	.w8(32'h38d5c7be),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367943be),
	.w1(32'h36e652aa),
	.w2(32'h37ec842a),
	.w3(32'h35d84635),
	.w4(32'h3781e65e),
	.w5(32'h38049ae8),
	.w6(32'h37c807f6),
	.w7(32'h37d4d0b4),
	.w8(32'h380537cc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64efeff),
	.w1(32'hb6237c6f),
	.w2(32'h37a20451),
	.w3(32'h3686ed3a),
	.w4(32'h362b177c),
	.w5(32'h379b0d05),
	.w6(32'h37a5a427),
	.w7(32'h378f9a7c),
	.w8(32'h3821352b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89e6f2),
	.w1(32'h390f972b),
	.w2(32'hb90886f1),
	.w3(32'h3aab653c),
	.w4(32'hb9d0693b),
	.w5(32'hba145cac),
	.w6(32'h3a48d16c),
	.w7(32'hba3b7058),
	.w8(32'hba9ca94a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813326d),
	.w1(32'hb823d143),
	.w2(32'h365eff5a),
	.w3(32'hb7e48f08),
	.w4(32'hb7b252bb),
	.w5(32'h3785ec68),
	.w6(32'hb618036d),
	.w7(32'h35a6e5fc),
	.w8(32'h38275eeb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac24d28),
	.w1(32'hbab19a07),
	.w2(32'hbb267e38),
	.w3(32'h3a90e9c3),
	.w4(32'hbad3236d),
	.w5(32'hbb6311bd),
	.w6(32'h3ad477bc),
	.w7(32'hb9e3e9b0),
	.w8(32'hbb481a61),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f715e),
	.w1(32'hbb076c77),
	.w2(32'hbb800bc7),
	.w3(32'h3afb8de1),
	.w4(32'hbadbdaf4),
	.w5(32'hbb8f91ae),
	.w6(32'hb927ec08),
	.w7(32'hbb6cfb91),
	.w8(32'hbbd71b9c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41fa36),
	.w1(32'h389c7ab2),
	.w2(32'hba3b1c04),
	.w3(32'h398ccb53),
	.w4(32'hb90e413e),
	.w5(32'hbaa7d919),
	.w6(32'h38d47c0e),
	.w7(32'hb952b072),
	.w8(32'hbb08e37f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6df60ce),
	.w1(32'h389e1090),
	.w2(32'h38a50813),
	.w3(32'h37807fae),
	.w4(32'h38c8de82),
	.w5(32'h38f0d48b),
	.w6(32'h388010ae),
	.w7(32'h38cccd51),
	.w8(32'h38d24d3c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac89ce2),
	.w1(32'hb9ced99c),
	.w2(32'hbb046057),
	.w3(32'h3bbc87e2),
	.w4(32'hba482561),
	.w5(32'hbbde3643),
	.w6(32'h3aaceb61),
	.w7(32'hbbdabfff),
	.w8(32'hbc36045f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfc458),
	.w1(32'h39913072),
	.w2(32'hb9a4711c),
	.w3(32'h3b00ff4d),
	.w4(32'hba519adc),
	.w5(32'hbae54ee2),
	.w6(32'h3a08c2f0),
	.w7(32'hbb6ce97f),
	.w8(32'hbb81d900),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb838e116),
	.w1(32'hb8049c9f),
	.w2(32'h36ef195c),
	.w3(32'hb78134ec),
	.w4(32'hb6b7ace5),
	.w5(32'hb6d0e661),
	.w6(32'h36f84b7e),
	.w7(32'h38175875),
	.w8(32'h381e2044),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a15077),
	.w1(32'hbab960d6),
	.w2(32'hbb0be9fe),
	.w3(32'h3a55d9d5),
	.w4(32'hbb2c4e20),
	.w5(32'hbb563a3f),
	.w6(32'h3993b0bc),
	.w7(32'hbb67df30),
	.w8(32'hbb810775),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccb9df),
	.w1(32'h39998a56),
	.w2(32'h3961da84),
	.w3(32'h39beea8e),
	.w4(32'h3988d9f3),
	.w5(32'h393b6509),
	.w6(32'h39671b4a),
	.w7(32'h3932bc11),
	.w8(32'h38e6466a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38747861),
	.w1(32'hb8304371),
	.w2(32'hb978b3e4),
	.w3(32'h37511a0a),
	.w4(32'h38e290e1),
	.w5(32'hb863791f),
	.w6(32'h37b2cfcb),
	.w7(32'h38a4756a),
	.w8(32'h387ae8e7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371dbc90),
	.w1(32'hb6a89840),
	.w2(32'h36a89cc6),
	.w3(32'h370c36cc),
	.w4(32'h37b67839),
	.w5(32'h375b72a9),
	.w6(32'hb5f4136c),
	.w7(32'h3806165c),
	.w8(32'h37ff128f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807af32),
	.w1(32'h3816f4d5),
	.w2(32'h3905f0c3),
	.w3(32'h37f31c26),
	.w4(32'hb6fb1679),
	.w5(32'h38658739),
	.w6(32'h38b41d02),
	.w7(32'hb8a6be58),
	.w8(32'hb76a98da),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44684c),
	.w1(32'hb995d23e),
	.w2(32'h39702205),
	.w3(32'hbadf0fab),
	.w4(32'hb94f81cb),
	.w5(32'h39ae516f),
	.w6(32'hba540e91),
	.w7(32'h39d631ee),
	.w8(32'h3a818da2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02622c),
	.w1(32'hbab33ef8),
	.w2(32'hbbaf617e),
	.w3(32'h3a1eb555),
	.w4(32'hba9a592d),
	.w5(32'hbb99668d),
	.w6(32'hba3eafb2),
	.w7(32'hbb9d166f),
	.w8(32'hbc096470),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce3d3d),
	.w1(32'hba8c1e95),
	.w2(32'hbb2ae78a),
	.w3(32'h3acb1c9b),
	.w4(32'hba98b80b),
	.w5(32'hbb299e76),
	.w6(32'h3a0c73e5),
	.w7(32'hbb65e56f),
	.w8(32'hbba53cc3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba326015),
	.w1(32'hba1388f2),
	.w2(32'hbb66734f),
	.w3(32'hba529e72),
	.w4(32'hbb22d455),
	.w5(32'hbb4904ac),
	.w6(32'hba99cdd1),
	.w7(32'hbb7e7d38),
	.w8(32'hbb866add),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bdbb1),
	.w1(32'h39168bb8),
	.w2(32'h39959fca),
	.w3(32'hb7598cec),
	.w4(32'h393e31e9),
	.w5(32'h398f0669),
	.w6(32'h381968b5),
	.w7(32'h396c17f8),
	.w8(32'h39a56cb6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6ea6f),
	.w1(32'hb90d104d),
	.w2(32'hb99f640b),
	.w3(32'h3a02108e),
	.w4(32'h39a56833),
	.w5(32'hb839e22e),
	.w6(32'h39fc4a50),
	.w7(32'h39c56617),
	.w8(32'hb89065af),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70940b6),
	.w1(32'hb71bb21d),
	.w2(32'hb4a31aaf),
	.w3(32'hb6da43cb),
	.w4(32'hb7468bec),
	.w5(32'h3581c98d),
	.w6(32'h368d5bc9),
	.w7(32'hb4f01b3b),
	.w8(32'h377fcc9e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb743aec2),
	.w1(32'hb7dc571a),
	.w2(32'hb80798af),
	.w3(32'h37fa7ded),
	.w4(32'h3797e53d),
	.w5(32'hb5584c3f),
	.w6(32'h381b9c29),
	.w7(32'h383b0adb),
	.w8(32'h38201721),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac86d5f),
	.w1(32'h39d825ab),
	.w2(32'hba4b0942),
	.w3(32'hb9db0b77),
	.w4(32'hba8bc00a),
	.w5(32'hbaed251c),
	.w6(32'hb9e6f22c),
	.w7(32'hbb87b6a2),
	.w8(32'hbb85d8c1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd99b0),
	.w1(32'hba166e8c),
	.w2(32'hba10d7b1),
	.w3(32'hb9ea9c60),
	.w4(32'hb9bae964),
	.w5(32'hba0d8c60),
	.w6(32'hb9f19912),
	.w7(32'hba14daf1),
	.w8(32'hba34ac02),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908f729),
	.w1(32'h390fa25b),
	.w2(32'h3a021b1b),
	.w3(32'h39abf09b),
	.w4(32'h39f7a968),
	.w5(32'h3a2abe65),
	.w6(32'h36873748),
	.w7(32'h38e992f0),
	.w8(32'h39c25a40),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147539),
	.w1(32'hba0de501),
	.w2(32'hba21ae0d),
	.w3(32'hbb08f123),
	.w4(32'hba59cdeb),
	.w5(32'hba0070dd),
	.w6(32'hbaff5955),
	.w7(32'h39674578),
	.w8(32'h37c0ca50),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8384416),
	.w1(32'hb7efa0d5),
	.w2(32'hb4a4f85c),
	.w3(32'hb7ac1f8d),
	.w4(32'hb6123368),
	.w5(32'h36fa612c),
	.w6(32'h37b3b530),
	.w7(32'h37f616cc),
	.w8(32'h3811f2ff),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3a308),
	.w1(32'h3a3045f9),
	.w2(32'hba9b0eca),
	.w3(32'h3ac620a9),
	.w4(32'hb9e6db69),
	.w5(32'hbb0b9216),
	.w6(32'h39e955fc),
	.w7(32'hbac62a22),
	.w8(32'hbb128979),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ca0d8),
	.w1(32'hb90d4439),
	.w2(32'hb98759b5),
	.w3(32'hb9692d72),
	.w4(32'hb9639b55),
	.w5(32'hb94aecd5),
	.w6(32'h37eb1252),
	.w7(32'hb9850c2d),
	.w8(32'hba307e04),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd7de1),
	.w1(32'h3b2df6ce),
	.w2(32'h3b6bde56),
	.w3(32'hbb4925f6),
	.w4(32'h3b56e5d4),
	.w5(32'h3bb8c40e),
	.w6(32'hbb94e1ef),
	.w7(32'hbb9a8fea),
	.w8(32'hba8570ec),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec8d17),
	.w1(32'h381b6a96),
	.w2(32'hb900965f),
	.w3(32'h3904894e),
	.w4(32'h38674398),
	.w5(32'hb828efa6),
	.w6(32'h391e1b31),
	.w7(32'hb79e2488),
	.w8(32'hb901f0dc),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a641f),
	.w1(32'hb90bc389),
	.w2(32'h3a239c1d),
	.w3(32'hbb02dcb1),
	.w4(32'h3ae2f266),
	.w5(32'h3a854163),
	.w6(32'hbaf5c99a),
	.w7(32'hb92e10ad),
	.w8(32'hba088b6f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule