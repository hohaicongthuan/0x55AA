module layer_10_featuremap_387(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00d92c),
	.w1(32'h3778da2a),
	.w2(32'hbb0a5bb8),
	.w3(32'hbadc32fe),
	.w4(32'hbb873c47),
	.w5(32'hbad4f4e6),
	.w6(32'hbc16a4ad),
	.w7(32'hbb881ab4),
	.w8(32'h3bba5870),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a6aa),
	.w1(32'hbb14c678),
	.w2(32'h3ad07098),
	.w3(32'hbbb79e5c),
	.w4(32'h3ac589eb),
	.w5(32'h3bdcfef6),
	.w6(32'h3bf2d65a),
	.w7(32'h3bcc0143),
	.w8(32'h3c0c998e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b8747),
	.w1(32'hba55e3e7),
	.w2(32'h38f6dace),
	.w3(32'hbae83035),
	.w4(32'h3b264369),
	.w5(32'hbc36daa0),
	.w6(32'h38cb1289),
	.w7(32'h3aa37095),
	.w8(32'h3c149d18),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbac371),
	.w1(32'hbb7bdb51),
	.w2(32'hbbe0e8a6),
	.w3(32'hbc4a1824),
	.w4(32'hbb8e3fc3),
	.w5(32'hbc8a2306),
	.w6(32'hb9de0641),
	.w7(32'hba3a3484),
	.w8(32'h3b529e70),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d08cf),
	.w1(32'h3afd95ca),
	.w2(32'hbb5fbacc),
	.w3(32'h3b49a4d0),
	.w4(32'h3b94b920),
	.w5(32'hbbf331fb),
	.w6(32'h3bd5077a),
	.w7(32'hbabfbcb2),
	.w8(32'h3b1c0e61),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d31eb),
	.w1(32'hbb146eaa),
	.w2(32'h3b0b2e87),
	.w3(32'hbb6555d2),
	.w4(32'h3c1a874e),
	.w5(32'h3c6d06d8),
	.w6(32'h3ae0b6ff),
	.w7(32'hbbc5c6e7),
	.w8(32'hbb880c28),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09e6c7),
	.w1(32'h3ae300a5),
	.w2(32'h3be3ecfa),
	.w3(32'h3beac11b),
	.w4(32'h3b6835c1),
	.w5(32'hbbcc2125),
	.w6(32'h39cf0d59),
	.w7(32'h3bebbba8),
	.w8(32'h3bf46fc4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040fa7),
	.w1(32'hbb34aa36),
	.w2(32'h3b89d708),
	.w3(32'hbba18c86),
	.w4(32'hbc2b5675),
	.w5(32'hbc2af189),
	.w6(32'h3c1b53fb),
	.w7(32'hbbcc7233),
	.w8(32'hbc4bcd9e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae236c),
	.w1(32'hbac1de79),
	.w2(32'hb9c5a149),
	.w3(32'hbbd4a814),
	.w4(32'hbad59f85),
	.w5(32'hbb475021),
	.w6(32'hbc1680b9),
	.w7(32'hbab38e9f),
	.w8(32'hbbd47779),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc11b4a),
	.w1(32'hbad32ee0),
	.w2(32'hbaa7f1ab),
	.w3(32'hbb24c408),
	.w4(32'hbaf54bd5),
	.w5(32'hbb87b717),
	.w6(32'h3b7b3c65),
	.w7(32'h3a511537),
	.w8(32'h3b9961d3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05bd22),
	.w1(32'hbb651856),
	.w2(32'hbb157a5b),
	.w3(32'h3adc4949),
	.w4(32'h3c2bcfda),
	.w5(32'h3cadad04),
	.w6(32'hba115097),
	.w7(32'hb9e85897),
	.w8(32'h3c386d98),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc24060),
	.w1(32'hbc002a00),
	.w2(32'hbbb643ed),
	.w3(32'h3be0bf14),
	.w4(32'h3a060a87),
	.w5(32'h3afa17e1),
	.w6(32'h3bab4eab),
	.w7(32'hb982e42c),
	.w8(32'hbadd8758),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb5c27),
	.w1(32'h3b634f16),
	.w2(32'hbb4c7ba4),
	.w3(32'hbb434af1),
	.w4(32'h3b8d76aa),
	.w5(32'hbb89d554),
	.w6(32'hbb989a5d),
	.w7(32'h3b59922c),
	.w8(32'h3b5220bf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24f20),
	.w1(32'h3be52ef6),
	.w2(32'h3b95af77),
	.w3(32'h3c3a8c17),
	.w4(32'h3bff1420),
	.w5(32'hbb363e5d),
	.w6(32'h39cd2182),
	.w7(32'h3b89e78a),
	.w8(32'h3c09b72a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf78a0d),
	.w1(32'hbb53963c),
	.w2(32'hbb652bba),
	.w3(32'hbaeff759),
	.w4(32'h3c9444bb),
	.w5(32'hbb79d6f4),
	.w6(32'h3c08b809),
	.w7(32'h3bee63e7),
	.w8(32'h3c5e1811),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e1e4e),
	.w1(32'hbb62d7a6),
	.w2(32'hbb509142),
	.w3(32'hb9c48f2b),
	.w4(32'hba775276),
	.w5(32'hbba305e4),
	.w6(32'h3bb7ecef),
	.w7(32'hbb178214),
	.w8(32'h3b0e1953),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda6f73),
	.w1(32'hbaae084c),
	.w2(32'hbb9052aa),
	.w3(32'hbb45aab4),
	.w4(32'h39933537),
	.w5(32'hbbabbbd1),
	.w6(32'hba59fa23),
	.w7(32'h3bbc067e),
	.w8(32'h3b16a169),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107d57),
	.w1(32'hbb734b72),
	.w2(32'hbbbd0179),
	.w3(32'hbbe643fe),
	.w4(32'hbb1a994b),
	.w5(32'h3b9ebc41),
	.w6(32'h3b342253),
	.w7(32'hbaee2074),
	.w8(32'hbb26918d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc089a3),
	.w1(32'h3afdbc94),
	.w2(32'hbb477ebb),
	.w3(32'hb989419b),
	.w4(32'h3c3fa85f),
	.w5(32'h3b78eed9),
	.w6(32'h39a354c5),
	.w7(32'hbaf21551),
	.w8(32'h3b63256a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6da480),
	.w1(32'hbb68a0b3),
	.w2(32'h3aea0622),
	.w3(32'h3b58ca32),
	.w4(32'h3c208a8e),
	.w5(32'hbad247d8),
	.w6(32'h3bb99413),
	.w7(32'h3c17af54),
	.w8(32'h3c933474),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15c206),
	.w1(32'h3ad4ba0f),
	.w2(32'h3bebd170),
	.w3(32'hbb024c7e),
	.w4(32'hbae081e5),
	.w5(32'h3b65d77e),
	.w6(32'h3b062b33),
	.w7(32'hbc022f10),
	.w8(32'hbb6ee23d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fea849),
	.w1(32'hbb2818b4),
	.w2(32'hba78a7cb),
	.w3(32'h392fe63f),
	.w4(32'hbb8179a3),
	.w5(32'hbabd414c),
	.w6(32'hbbc21d84),
	.w7(32'hbb934142),
	.w8(32'hbc18c2a6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ed84f),
	.w1(32'h3bf96b39),
	.w2(32'h3bf475b4),
	.w3(32'h3b9f295e),
	.w4(32'hbb9f9908),
	.w5(32'h3b865950),
	.w6(32'hbc13913c),
	.w7(32'hbb8b726c),
	.w8(32'h39869ed1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc414a),
	.w1(32'hbb1979ad),
	.w2(32'hbb8c9789),
	.w3(32'h3bac613c),
	.w4(32'h3c07bb66),
	.w5(32'h3b49551d),
	.w6(32'hbb011cbe),
	.w7(32'h3c2a9e61),
	.w8(32'h3bd12d89),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed26d5),
	.w1(32'hbac0ee23),
	.w2(32'h3b166f64),
	.w3(32'h3aa04de0),
	.w4(32'h3b905016),
	.w5(32'hba95f3d2),
	.w6(32'h3a8a702d),
	.w7(32'h3aa65116),
	.w8(32'hbbc677db),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819a8e),
	.w1(32'h3b80b26f),
	.w2(32'h3c059ec3),
	.w3(32'h3b84d586),
	.w4(32'hbbb69038),
	.w5(32'h3bd24c24),
	.w6(32'h3a03d4d6),
	.w7(32'hbc362605),
	.w8(32'hbc5a884f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35b897),
	.w1(32'h3b836604),
	.w2(32'h3b0da83a),
	.w3(32'h3c140762),
	.w4(32'hbbd0b39d),
	.w5(32'hbb584435),
	.w6(32'hbb638886),
	.w7(32'h3b99d5c9),
	.w8(32'h3b83e034),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862ae3),
	.w1(32'hbb812a86),
	.w2(32'hba8e3f55),
	.w3(32'hbb806733),
	.w4(32'h39d88203),
	.w5(32'hbbb16857),
	.w6(32'hba0c1dd1),
	.w7(32'h3b416d3a),
	.w8(32'hba8a2099),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86e4af),
	.w1(32'hbae1b1a5),
	.w2(32'h3c057c0e),
	.w3(32'h3acbbdc8),
	.w4(32'hbbddb8d7),
	.w5(32'h3c6942b8),
	.w6(32'h3abfba12),
	.w7(32'h3badbd87),
	.w8(32'h3ba977a5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aa2fb),
	.w1(32'h3b061e98),
	.w2(32'h392b0c1d),
	.w3(32'h3c8df45c),
	.w4(32'h3bcd9410),
	.w5(32'h3bb85e78),
	.w6(32'h3b21255f),
	.w7(32'h38f778f9),
	.w8(32'h39031114),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893025),
	.w1(32'hbbe4988d),
	.w2(32'hbaf2ad15),
	.w3(32'h3b9cffbc),
	.w4(32'h3b986fcb),
	.w5(32'hb92fd1b8),
	.w6(32'hbb1600ab),
	.w7(32'h3bf68acf),
	.w8(32'h3c08389b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8d613),
	.w1(32'hbb3ef9c0),
	.w2(32'hbb4e629a),
	.w3(32'h3a736a32),
	.w4(32'h3bde3c6c),
	.w5(32'hbb7069a8),
	.w6(32'h3b49cdfa),
	.w7(32'h3c367333),
	.w8(32'h3b6b203c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28e3d7),
	.w1(32'h3a6cad7a),
	.w2(32'h3ae80cc5),
	.w3(32'hbb8351a4),
	.w4(32'hbb165512),
	.w5(32'h3b296f0c),
	.w6(32'h3b846a5e),
	.w7(32'hbb540a58),
	.w8(32'hbbd8aa18),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe845d5),
	.w1(32'h3b4ab28e),
	.w2(32'h3c0ee10d),
	.w3(32'hbb4499b9),
	.w4(32'hba46b787),
	.w5(32'hb94ffc9f),
	.w6(32'hbb158f46),
	.w7(32'hbb92069f),
	.w8(32'hbbcda81a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074933),
	.w1(32'h3bf195d8),
	.w2(32'h3c5bd8bc),
	.w3(32'hbb3e6eb5),
	.w4(32'h3ab9d3b5),
	.w5(32'h3bda82ab),
	.w6(32'h39051f3e),
	.w7(32'hbc09dd9b),
	.w8(32'hbc1db172),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1abb77),
	.w1(32'hbb18e96d),
	.w2(32'hbb1e9375),
	.w3(32'h3b315ea9),
	.w4(32'hb9c02f00),
	.w5(32'hbaee0e09),
	.w6(32'hbb8c5d86),
	.w7(32'hbae3e1dd),
	.w8(32'hbb55a508),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a5338),
	.w1(32'h3b8cf354),
	.w2(32'hbab7755b),
	.w3(32'hbb6eac88),
	.w4(32'h3b26ed39),
	.w5(32'h3c0c08b3),
	.w6(32'hba5115f0),
	.w7(32'hbb920fc4),
	.w8(32'h3bdbf913),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb678eac),
	.w1(32'h3aabdad8),
	.w2(32'h3b39e133),
	.w3(32'hbb44154f),
	.w4(32'h3bc8664a),
	.w5(32'h3c195f6b),
	.w6(32'h3b454fdb),
	.w7(32'h3c05e8ec),
	.w8(32'h3b7beb3f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba671a7),
	.w1(32'hbb88339b),
	.w2(32'hba66c501),
	.w3(32'hb9ac7088),
	.w4(32'h3a7c8e51),
	.w5(32'h3973237b),
	.w6(32'h3aa4ded5),
	.w7(32'hbbe72ad8),
	.w8(32'h3a4eeda9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6117),
	.w1(32'hbb8470b4),
	.w2(32'hbbe9804b),
	.w3(32'hbb8300b8),
	.w4(32'hba7c29a1),
	.w5(32'hbb6bcc19),
	.w6(32'hbb099940),
	.w7(32'hbb3280e9),
	.w8(32'hba86d3dc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2624),
	.w1(32'h3ac81815),
	.w2(32'h3ad75eb6),
	.w3(32'h3ba31569),
	.w4(32'h3c3b0878),
	.w5(32'hba21df53),
	.w6(32'h3b9fe8f6),
	.w7(32'h3c9445d8),
	.w8(32'h3bf46d5a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ef242),
	.w1(32'hbb055604),
	.w2(32'h3b05e816),
	.w3(32'hbaa07ad2),
	.w4(32'h3bbe54d5),
	.w5(32'h3b8e1379),
	.w6(32'h3bb67af3),
	.w7(32'hb7891433),
	.w8(32'h3a7f0afc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb157d1),
	.w1(32'hbbd21afb),
	.w2(32'hbc4059bf),
	.w3(32'hbb4c5ece),
	.w4(32'hbb72c66c),
	.w5(32'hbbda7538),
	.w6(32'hbaa6616a),
	.w7(32'h3b249287),
	.w8(32'h3b82067d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ea1c),
	.w1(32'hba09febe),
	.w2(32'hbb393f34),
	.w3(32'h38ed6b5c),
	.w4(32'hb91625cc),
	.w5(32'hba8d9939),
	.w6(32'h3b6120e3),
	.w7(32'h3aa30ce9),
	.w8(32'hba8350df),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bcbda),
	.w1(32'h3b074f5a),
	.w2(32'hbb99a262),
	.w3(32'h39f42282),
	.w4(32'h3b622b85),
	.w5(32'hbb579e5b),
	.w6(32'hba9aff38),
	.w7(32'hba517da5),
	.w8(32'h3a80b77a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb1a57),
	.w1(32'hbbad10b7),
	.w2(32'hbbd0f93d),
	.w3(32'h3a3c05a9),
	.w4(32'hbb7af43f),
	.w5(32'hbbabbea9),
	.w6(32'h3b4bbc88),
	.w7(32'h3bc945f4),
	.w8(32'h3b8177cf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4816ab),
	.w1(32'hb9874847),
	.w2(32'hb9e921ce),
	.w3(32'hbbde802d),
	.w4(32'h3b74828f),
	.w5(32'hbb8e54f2),
	.w6(32'h3a59c63a),
	.w7(32'hbb9ca644),
	.w8(32'hb9237799),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f60cf),
	.w1(32'hb9d5c709),
	.w2(32'h384955ad),
	.w3(32'h3950e18e),
	.w4(32'hbab2f0fd),
	.w5(32'hb856c01b),
	.w6(32'hb93adafa),
	.w7(32'h3b270fbf),
	.w8(32'h3b865545),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4a739),
	.w1(32'h3bbebcff),
	.w2(32'h3c25a111),
	.w3(32'h3bdb1028),
	.w4(32'hbaad2ec5),
	.w5(32'h3aef724c),
	.w6(32'h3c128582),
	.w7(32'h3a361ead),
	.w8(32'hbb735933),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85551a),
	.w1(32'hbbcb9d9c),
	.w2(32'hba89d4e3),
	.w3(32'h3bd64336),
	.w4(32'h39113208),
	.w5(32'hbb9c4fc9),
	.w6(32'h3b89c32c),
	.w7(32'h3b992411),
	.w8(32'hbb046fb7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1424a6),
	.w1(32'h3aa7a892),
	.w2(32'h3b2f8184),
	.w3(32'h3bbe6b40),
	.w4(32'h3b3ae049),
	.w5(32'h3b4f628c),
	.w6(32'h3a089659),
	.w7(32'h3b157528),
	.w8(32'h3b1fb7cd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba579576),
	.w1(32'hba3061a8),
	.w2(32'h3b27a2bf),
	.w3(32'hbb744a20),
	.w4(32'h3af59dc1),
	.w5(32'hba718cd8),
	.w6(32'h3ba5ebb3),
	.w7(32'h3b4777da),
	.w8(32'h3b10b040),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc070584),
	.w1(32'h3b912495),
	.w2(32'h3c05919b),
	.w3(32'hbb206250),
	.w4(32'h39664d03),
	.w5(32'h3b237d0f),
	.w6(32'hbb83c315),
	.w7(32'hbb8bed41),
	.w8(32'hbbb44f3c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253ff7),
	.w1(32'hba94a4ae),
	.w2(32'h3bbbc3f0),
	.w3(32'h3bb9047a),
	.w4(32'hbc0f6565),
	.w5(32'hbbddcd2f),
	.w6(32'hbb561d99),
	.w7(32'hbc1682ac),
	.w8(32'hbc562526),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba70acc),
	.w1(32'hbb84e7e6),
	.w2(32'hbbd911aa),
	.w3(32'hbbc982fb),
	.w4(32'h3b86cdd9),
	.w5(32'h3aa96c53),
	.w6(32'hbbcf4561),
	.w7(32'h3c13db5d),
	.w8(32'h3c2c79ea),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e471bc),
	.w1(32'hbb6421bd),
	.w2(32'hbc09e5a3),
	.w3(32'hbaad0c35),
	.w4(32'h39e3b6b7),
	.w5(32'hbba98130),
	.w6(32'h3b806b14),
	.w7(32'h3bf009f8),
	.w8(32'h3b97500f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a75d3),
	.w1(32'h3b1fa34d),
	.w2(32'hba6df575),
	.w3(32'hbc01570b),
	.w4(32'h3ba384ab),
	.w5(32'h38088aab),
	.w6(32'hbb24a9da),
	.w7(32'h3b00aeae),
	.w8(32'h3c014ae1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b78f8),
	.w1(32'h39b9e26d),
	.w2(32'hbb2e02c0),
	.w3(32'hb9ac6e8a),
	.w4(32'h3b0b470f),
	.w5(32'hbb892715),
	.w6(32'h3ba4d6fe),
	.w7(32'hbaf7f0f6),
	.w8(32'hbc09faaf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81bf42),
	.w1(32'hb9045721),
	.w2(32'h3b737b8b),
	.w3(32'hbada95f7),
	.w4(32'h3bd7dc67),
	.w5(32'h3c332eda),
	.w6(32'hbbc09ab5),
	.w7(32'hbac56024),
	.w8(32'h3b9d64f0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b3f56),
	.w1(32'h3b119135),
	.w2(32'h3a47407f),
	.w3(32'h3bc37587),
	.w4(32'h3bedbbf0),
	.w5(32'hbc31c9ed),
	.w6(32'h3a4407e4),
	.w7(32'h3bd8e40d),
	.w8(32'h3be3cf3a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb82840),
	.w1(32'hbb89f8e7),
	.w2(32'hbb2e5621),
	.w3(32'h3a548c6a),
	.w4(32'hbb600dd6),
	.w5(32'h3b2c723c),
	.w6(32'h3aeed72f),
	.w7(32'h3acd97d7),
	.w8(32'hb975a732),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fcdf7),
	.w1(32'hbb3f2e8f),
	.w2(32'hbbf257db),
	.w3(32'h3a254f1f),
	.w4(32'h3bd55fdd),
	.w5(32'h39198d72),
	.w6(32'hbaf38189),
	.w7(32'hbba22ee5),
	.w8(32'h3bbbdc19),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fe4b1),
	.w1(32'hbbacb4a6),
	.w2(32'hbbc39fd8),
	.w3(32'hbbfc6296),
	.w4(32'hbb9c0ec4),
	.w5(32'hbc24b854),
	.w6(32'h3aa45fc9),
	.w7(32'h3ba51398),
	.w8(32'h3b7940fd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccdd9a),
	.w1(32'hbbb05e56),
	.w2(32'hbbd4d81b),
	.w3(32'h3b340cb0),
	.w4(32'hbb873b1a),
	.w5(32'hbbc1f456),
	.w6(32'hb9daf7a1),
	.w7(32'h3b35479d),
	.w8(32'h3b5d8f45),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a95b7),
	.w1(32'h3bcf4ea8),
	.w2(32'h3beafaa6),
	.w3(32'hbb7389d7),
	.w4(32'hbb2e5914),
	.w5(32'hb9e25092),
	.w6(32'h3b77a863),
	.w7(32'hbc073608),
	.w8(32'hbba3c714),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38ad0c),
	.w1(32'hbb508673),
	.w2(32'h3ba5f797),
	.w3(32'h3bf2b799),
	.w4(32'h3b16a3b1),
	.w5(32'h3bebe859),
	.w6(32'h3b035b13),
	.w7(32'hbb8477dc),
	.w8(32'hbb9704fa),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab06e5),
	.w1(32'hbb808126),
	.w2(32'hbbe0cdf0),
	.w3(32'hba40b738),
	.w4(32'hbb8c7553),
	.w5(32'hbacf7019),
	.w6(32'h3a45ba1f),
	.w7(32'hbb42dc47),
	.w8(32'hbbe2e234),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76f052),
	.w1(32'hbbbc016f),
	.w2(32'hbbc2d2d1),
	.w3(32'hbb8657bb),
	.w4(32'hbbb1c6fc),
	.w5(32'hbc47dc3e),
	.w6(32'hba4561b4),
	.w7(32'h3bbd065f),
	.w8(32'hbba12ec0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4d9b),
	.w1(32'hbb52ef04),
	.w2(32'h3b262157),
	.w3(32'hbbfd3f0d),
	.w4(32'hbc01deee),
	.w5(32'h3be1f9a7),
	.w6(32'h3b951417),
	.w7(32'hb9f6b92b),
	.w8(32'h3bbf2cc5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7dc8d),
	.w1(32'hbb069b90),
	.w2(32'h3ac57906),
	.w3(32'h3bb15700),
	.w4(32'hbac8c1ad),
	.w5(32'hbb99584d),
	.w6(32'hbb70a780),
	.w7(32'h3b66aec4),
	.w8(32'hbb2ad62d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1960e9),
	.w1(32'hbaa6b5fc),
	.w2(32'hbb8cfcff),
	.w3(32'hbb267ed6),
	.w4(32'hbb686ffe),
	.w5(32'hbb23831b),
	.w6(32'h3bacbdba),
	.w7(32'hbc0c3cc6),
	.w8(32'hbba81226),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a3b1),
	.w1(32'hbc6c893a),
	.w2(32'hbcd45135),
	.w3(32'hbb1e0350),
	.w4(32'hbcc5d0e6),
	.w5(32'h3d5c3a1e),
	.w6(32'hbbfc2a18),
	.w7(32'h3c1e801c),
	.w8(32'h3c572e6c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb3392),
	.w1(32'h3b730b36),
	.w2(32'h3bb2ad9e),
	.w3(32'h3c58c237),
	.w4(32'hba5853be),
	.w5(32'hbb7d224c),
	.w6(32'hbc573bd8),
	.w7(32'hbb5a5362),
	.w8(32'h3ba8d01a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7dcb),
	.w1(32'h3bebf991),
	.w2(32'h3c056196),
	.w3(32'h3adf3350),
	.w4(32'h3c6abbed),
	.w5(32'hbc6926f1),
	.w6(32'h3bb4a029),
	.w7(32'hbbd27562),
	.w8(32'hbc1f272c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04a27e),
	.w1(32'h3bc96c9b),
	.w2(32'hbb06d6b7),
	.w3(32'hbc08f0fa),
	.w4(32'h3c0bbcf4),
	.w5(32'h3aea7d0e),
	.w6(32'h3c0d6563),
	.w7(32'hbaa51a2e),
	.w8(32'hba0a5185),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bb88b),
	.w1(32'hbb9603c1),
	.w2(32'hb99b01a9),
	.w3(32'h3b773357),
	.w4(32'hbb25e252),
	.w5(32'h3bc22de3),
	.w6(32'h3afdeb7c),
	.w7(32'hbb873aed),
	.w8(32'hbb3a85e4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d7692),
	.w1(32'hbb7bba18),
	.w2(32'h3ba725b1),
	.w3(32'h3b16b083),
	.w4(32'h3b49d56a),
	.w5(32'h3acd6506),
	.w6(32'h37a8a717),
	.w7(32'hbb445254),
	.w8(32'hbbe8e78b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a8b75),
	.w1(32'h3b57d2e7),
	.w2(32'h3bac8285),
	.w3(32'hbbce3b05),
	.w4(32'h3be83b00),
	.w5(32'hbc140302),
	.w6(32'h3a1681bc),
	.w7(32'hbae8c723),
	.w8(32'hbbeb235d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac729c6),
	.w1(32'hbc853138),
	.w2(32'hbc82748b),
	.w3(32'h392ef5e7),
	.w4(32'hbc1012f3),
	.w5(32'h3c763f63),
	.w6(32'h3b2bdcd6),
	.w7(32'h3bf409e0),
	.w8(32'h3bd0b41b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69c202),
	.w1(32'hbb9bc34d),
	.w2(32'h3b5b8ee7),
	.w3(32'h3b3ecb9e),
	.w4(32'hbbc3ff35),
	.w5(32'h3ba7eab3),
	.w6(32'hbbdec541),
	.w7(32'hbb5bc37d),
	.w8(32'h3b839f03),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2744eb),
	.w1(32'h3c322485),
	.w2(32'h3be6f6da),
	.w3(32'h3a6f9e6e),
	.w4(32'h3c1695d4),
	.w5(32'h3bc249fe),
	.w6(32'hbb034a0f),
	.w7(32'h3c4e1954),
	.w8(32'h3b80b38a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3697c6),
	.w1(32'h3aa36ebc),
	.w2(32'h3bbe1252),
	.w3(32'h3bfb3a18),
	.w4(32'h3bc34fd3),
	.w5(32'h3a9c7d30),
	.w6(32'hba4e996a),
	.w7(32'hba0c1ede),
	.w8(32'h3ae0dc6d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a8c54),
	.w1(32'hbc45f0b5),
	.w2(32'hbc4ebc9d),
	.w3(32'h3ba51c89),
	.w4(32'hbc7e16ce),
	.w5(32'h3cdf19b1),
	.w6(32'h3b67b061),
	.w7(32'h3c1c4e94),
	.w8(32'h3b02625e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ae8e9),
	.w1(32'hbb012c0f),
	.w2(32'h3b21c350),
	.w3(32'h3bf23e9a),
	.w4(32'h3b52e23b),
	.w5(32'hbbe1e11f),
	.w6(32'hbc954a0a),
	.w7(32'h3b31b158),
	.w8(32'hbb1d1f2d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec4315),
	.w1(32'h3a96b044),
	.w2(32'hbb0bf654),
	.w3(32'hbbf4fa1a),
	.w4(32'h3a58bd31),
	.w5(32'hbb38358a),
	.w6(32'h3b1bc194),
	.w7(32'hb9d8beed),
	.w8(32'h3ba494ca),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e5a07),
	.w1(32'h3ae23255),
	.w2(32'h3ab2444c),
	.w3(32'h3c654649),
	.w4(32'hbb50a24b),
	.w5(32'hbc064a4b),
	.w6(32'h3bf4ae68),
	.w7(32'hbb82261c),
	.w8(32'hbc0e933f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0edc1),
	.w1(32'hbbc3144e),
	.w2(32'hbc16c526),
	.w3(32'hbad32795),
	.w4(32'hbb65f564),
	.w5(32'hbaba33b5),
	.w6(32'hbbe11a9d),
	.w7(32'h3b90211d),
	.w8(32'h3ba36e85),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ceec3),
	.w1(32'hbb093394),
	.w2(32'h3be97c20),
	.w3(32'h39b28f09),
	.w4(32'h3ba502f3),
	.w5(32'hbb828ce6),
	.w6(32'h3760d1b0),
	.w7(32'hbb8bcef2),
	.w8(32'h3b0f8290),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf41c2d),
	.w1(32'hbb1ddebe),
	.w2(32'hbc029477),
	.w3(32'hbb12ca0e),
	.w4(32'hbb4d7603),
	.w5(32'hbbb53b49),
	.w6(32'h3b9bd803),
	.w7(32'hbba45be2),
	.w8(32'hbc49eeb0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00392f),
	.w1(32'hbb606c29),
	.w2(32'hbb6755b4),
	.w3(32'hbc564a51),
	.w4(32'h3a46f3d8),
	.w5(32'h3b223f1c),
	.w6(32'hbbd58ff3),
	.w7(32'hbb3577be),
	.w8(32'hbb37e24f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd830),
	.w1(32'h3adaf7fa),
	.w2(32'h3b9e7e47),
	.w3(32'h3b408844),
	.w4(32'h3b0bd702),
	.w5(32'hb9acfe66),
	.w6(32'hbac769cf),
	.w7(32'h3b257ff2),
	.w8(32'hbbfc2372),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc323362),
	.w1(32'hbbdf39b8),
	.w2(32'hb9ecce87),
	.w3(32'hbc1fed75),
	.w4(32'h3c07eaf0),
	.w5(32'hb9b949dc),
	.w6(32'hba95d757),
	.w7(32'hba561827),
	.w8(32'h3bb31e36),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951e63a),
	.w1(32'hbc23add7),
	.w2(32'h3996352f),
	.w3(32'h3baededb),
	.w4(32'hbc78891d),
	.w5(32'h3cbedb77),
	.w6(32'hbb8578fb),
	.w7(32'h3be16e71),
	.w8(32'h3c10aef2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8aa27),
	.w1(32'hba8ea771),
	.w2(32'h3b2b7c7b),
	.w3(32'h3b33f9b0),
	.w4(32'h3ac847eb),
	.w5(32'hbc52530f),
	.w6(32'hbc6cdbe1),
	.w7(32'h3be2d1cb),
	.w8(32'hbb0d1eab),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba30180),
	.w1(32'h3a87d340),
	.w2(32'h3a85ee39),
	.w3(32'hbb0c609a),
	.w4(32'h3bc71a4e),
	.w5(32'h3a2c2630),
	.w6(32'hb9ef1c7f),
	.w7(32'hbb32093a),
	.w8(32'hbb9a7e16),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1455b8),
	.w1(32'hbb457d3f),
	.w2(32'h3c583fd2),
	.w3(32'hbbc9c98f),
	.w4(32'h3c3fab42),
	.w5(32'hbc83b0a0),
	.w6(32'h3b556199),
	.w7(32'hbc4b5b39),
	.w8(32'hbc2a25c5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15f1ec),
	.w1(32'hbbb1b034),
	.w2(32'h3c39593f),
	.w3(32'hb9b4f5e0),
	.w4(32'h3c5105b7),
	.w5(32'hbbc00c5a),
	.w6(32'h3be03c6d),
	.w7(32'hbc0ff724),
	.w8(32'hbb0d0ea1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1539c4),
	.w1(32'hbb2399a9),
	.w2(32'h3b23234d),
	.w3(32'h3b20d24d),
	.w4(32'hbb0a8069),
	.w5(32'h3bed1ae3),
	.w6(32'h3c92676c),
	.w7(32'h3a3cb92c),
	.w8(32'h3b90fc2c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2382a0),
	.w1(32'h3bb63c61),
	.w2(32'h3bcf58cb),
	.w3(32'h3a96b05b),
	.w4(32'h3bea0484),
	.w5(32'h3c0eb801),
	.w6(32'hba86c6cc),
	.w7(32'h3b963e53),
	.w8(32'h3b0c9fa2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6a122),
	.w1(32'hb8478c72),
	.w2(32'hbb9035d0),
	.w3(32'h3ae8ddf8),
	.w4(32'hba0d5fe9),
	.w5(32'hba11be8b),
	.w6(32'h3c12de66),
	.w7(32'hba33b609),
	.w8(32'h3b0c4a44),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d66af),
	.w1(32'hbb91a7c9),
	.w2(32'h3bba824a),
	.w3(32'hbb7576ab),
	.w4(32'h3c1449ff),
	.w5(32'h3a66ead5),
	.w6(32'hbb10e4d9),
	.w7(32'hbb75f940),
	.w8(32'hbafa6847),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe08e7f),
	.w1(32'hbb1d9714),
	.w2(32'h3a0beaa9),
	.w3(32'hbb4c65bc),
	.w4(32'hbc339c15),
	.w5(32'hbbfbb490),
	.w6(32'h3bb5cd90),
	.w7(32'hbc0af737),
	.w8(32'hb9b287af),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69862a),
	.w1(32'h3b503072),
	.w2(32'h3ba44ac1),
	.w3(32'h3a16c82a),
	.w4(32'h3afcc4fc),
	.w5(32'h3c7d7913),
	.w6(32'h3af2cb8d),
	.w7(32'hbb8a8066),
	.w8(32'hbbc7a9a0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820972),
	.w1(32'hbb06f4b6),
	.w2(32'h3b11fc98),
	.w3(32'hbb5b90b1),
	.w4(32'h3b37e11c),
	.w5(32'hbbd06d5d),
	.w6(32'hbbbb56d1),
	.w7(32'hbbaac18d),
	.w8(32'hba4b3784),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc1286),
	.w1(32'hbbf71758),
	.w2(32'hbc0646d2),
	.w3(32'h37c4fd3a),
	.w4(32'hbc914481),
	.w5(32'h3cd58e2f),
	.w6(32'h3afcc922),
	.w7(32'h3b45b005),
	.w8(32'hb957baab),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e8051),
	.w1(32'hb9d2eb2d),
	.w2(32'h3aabdf96),
	.w3(32'hba761c12),
	.w4(32'hba61469e),
	.w5(32'h3b0487b0),
	.w6(32'hbbd5b02d),
	.w7(32'h3b740084),
	.w8(32'h3b253ded),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78cb0e),
	.w1(32'hbb74a658),
	.w2(32'hbb93c183),
	.w3(32'h3bc78d1c),
	.w4(32'h381d3874),
	.w5(32'h3bc85fd2),
	.w6(32'hbb52326a),
	.w7(32'h38cc8fdf),
	.w8(32'hba2bab52),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1429),
	.w1(32'hbb0cb3d8),
	.w2(32'hba79ece3),
	.w3(32'h3bc927ea),
	.w4(32'h3b94b89d),
	.w5(32'hbb8b588b),
	.w6(32'hbb97b2f5),
	.w7(32'hbabf2d38),
	.w8(32'hbbaf222a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb41af2),
	.w1(32'h3b1780bb),
	.w2(32'h3b47a972),
	.w3(32'hbc09fb18),
	.w4(32'hbc6092c0),
	.w5(32'h3c763c56),
	.w6(32'hb9ac4308),
	.w7(32'hbae19a8a),
	.w8(32'hbbd248c2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddfa53),
	.w1(32'h3ac904e8),
	.w2(32'h3ba58b54),
	.w3(32'h3bc42674),
	.w4(32'hbb8999f4),
	.w5(32'hbc2cb43e),
	.w6(32'hbb6ef398),
	.w7(32'h3ac31b29),
	.w8(32'hbbbdb640),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70efde),
	.w1(32'h3beddbbe),
	.w2(32'hbb602eb9),
	.w3(32'hbbb5ff5c),
	.w4(32'h3ae9080b),
	.w5(32'hba4c2ded),
	.w6(32'hbb949683),
	.w7(32'hba853ed9),
	.w8(32'hba358f0d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6b57c),
	.w1(32'h3b829087),
	.w2(32'hb9bd107c),
	.w3(32'h39eb6fde),
	.w4(32'h3b66600c),
	.w5(32'h3ba5f093),
	.w6(32'hbbb43df9),
	.w7(32'h3b502023),
	.w8(32'hbb19e95c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b679003),
	.w1(32'h3c09e803),
	.w2(32'h3cb337e6),
	.w3(32'h3b0e31ed),
	.w4(32'h3ca19830),
	.w5(32'hbca2afb0),
	.w6(32'h3b288747),
	.w7(32'hbbfd3a8e),
	.w8(32'hbc0fc9b7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc480069),
	.w1(32'h3c17a616),
	.w2(32'h3a82407b),
	.w3(32'hbc2f3892),
	.w4(32'h3c252884),
	.w5(32'h3b580eda),
	.w6(32'h3c87f337),
	.w7(32'h37db3a81),
	.w8(32'hbc3717f6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38d75b),
	.w1(32'hbb39a2de),
	.w2(32'hbc3a78da),
	.w3(32'h3b4ca87b),
	.w4(32'hbbab7b2e),
	.w5(32'h3cc8a0e8),
	.w6(32'hbb6786e3),
	.w7(32'h3c65479c),
	.w8(32'h3c2af838),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c057afb),
	.w1(32'hba9c19df),
	.w2(32'hbb922fd2),
	.w3(32'h3b7f1101),
	.w4(32'hbb7c260d),
	.w5(32'hbb4553f7),
	.w6(32'hbbd3faa7),
	.w7(32'hbbbb3642),
	.w8(32'hbbc63f2f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb326c0),
	.w1(32'hba1312c3),
	.w2(32'h38f872fe),
	.w3(32'hbc417f45),
	.w4(32'h3b6f2ff6),
	.w5(32'hbc6e59c5),
	.w6(32'hbc26f4c5),
	.w7(32'h3b406f63),
	.w8(32'hbbb1945f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aa2ba),
	.w1(32'hbc06be30),
	.w2(32'hbbc20632),
	.w3(32'hbb7aa748),
	.w4(32'hbbc66f9a),
	.w5(32'h3c887e85),
	.w6(32'h3b524c32),
	.w7(32'h3c052c43),
	.w8(32'h3ac7cf97),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a14f4),
	.w1(32'hbb9de0bb),
	.w2(32'h3b42f946),
	.w3(32'h3bec5fcc),
	.w4(32'h3becfb63),
	.w5(32'hbc1939ea),
	.w6(32'hbbf27a8d),
	.w7(32'hbc6b291b),
	.w8(32'hbc83ff63),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc299972),
	.w1(32'hbb86c44c),
	.w2(32'hbbbea67f),
	.w3(32'hbc457047),
	.w4(32'hbc05adcf),
	.w5(32'h3cb252c9),
	.w6(32'hbb53f640),
	.w7(32'h3a3fc5d6),
	.w8(32'h3c1c88dd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169c94),
	.w1(32'hbb85ac75),
	.w2(32'hbb7c4326),
	.w3(32'h3b73fbac),
	.w4(32'h3a3a9e50),
	.w5(32'hbba6ec75),
	.w6(32'hbb26ca35),
	.w7(32'h3b4d7177),
	.w8(32'hbb511f40),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15683a),
	.w1(32'hbaa0fc87),
	.w2(32'hbc100458),
	.w3(32'hbb95a978),
	.w4(32'hbb0cf71d),
	.w5(32'h3b38c2da),
	.w6(32'hbab8bc2d),
	.w7(32'h39b2d30d),
	.w8(32'hbb0f52d5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba917c81),
	.w1(32'h3bce8db9),
	.w2(32'h3c0c048b),
	.w3(32'hbc247522),
	.w4(32'h3b8dc488),
	.w5(32'hb9a03a0e),
	.w6(32'hbb6be0d6),
	.w7(32'hbc06d92c),
	.w8(32'h3aa0d6da),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02d00),
	.w1(32'h3b7e2252),
	.w2(32'h3bfc9228),
	.w3(32'hbb2ba7e6),
	.w4(32'h3c0a0174),
	.w5(32'hbca6ea15),
	.w6(32'h3bcb2398),
	.w7(32'hbc0c4df6),
	.w8(32'hbbd2df79),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f202c),
	.w1(32'hbc2daa02),
	.w2(32'hbc669753),
	.w3(32'hbb3274a5),
	.w4(32'hbc812b19),
	.w5(32'h3cb8d859),
	.w6(32'h3bdc7ef3),
	.w7(32'hba885493),
	.w8(32'h3bca8ff8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf88f96),
	.w1(32'hbb6c22d8),
	.w2(32'hbc3866a4),
	.w3(32'h3bb0aed6),
	.w4(32'hbc05f0cc),
	.w5(32'h3d17e459),
	.w6(32'hbbad19e2),
	.w7(32'h3a8fa046),
	.w8(32'h3b71d0ce),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5f90d),
	.w1(32'hba856ec4),
	.w2(32'hbc3420e0),
	.w3(32'h3b40750e),
	.w4(32'hbbf39813),
	.w5(32'hbb8efd32),
	.w6(32'hbbc13aa9),
	.w7(32'hbbf2345d),
	.w8(32'hbb9fafe9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e02f0),
	.w1(32'hbb09e1f9),
	.w2(32'hbc33ef62),
	.w3(32'hbc02eb68),
	.w4(32'hbbdcdb4b),
	.w5(32'hbc032a48),
	.w6(32'hbc27f274),
	.w7(32'hbb875137),
	.w8(32'hb831d794),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574db9),
	.w1(32'hbaf36d41),
	.w2(32'hbb836de8),
	.w3(32'h38102bf9),
	.w4(32'h3b2fb1bb),
	.w5(32'h3c008736),
	.w6(32'hba8af5c2),
	.w7(32'h3abe6667),
	.w8(32'hbb11203e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b11cd),
	.w1(32'hbb9ab35c),
	.w2(32'hbc0d44eb),
	.w3(32'h3b5776bf),
	.w4(32'hbc19ef07),
	.w5(32'h3c13f4c8),
	.w6(32'h3ac2afd5),
	.w7(32'h3bc766b7),
	.w8(32'h3b2a9629),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa83f7b),
	.w1(32'hbc4224e4),
	.w2(32'h3947e1e8),
	.w3(32'hbb4b1981),
	.w4(32'hbc06154f),
	.w5(32'hbc340189),
	.w6(32'hbb2c6154),
	.w7(32'hbbd83126),
	.w8(32'hbc155317),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65a575),
	.w1(32'hbb2a62d7),
	.w2(32'hbcb7d0ee),
	.w3(32'hbb4ed517),
	.w4(32'hbc302cdf),
	.w5(32'h3d3d2012),
	.w6(32'hbb17b8b0),
	.w7(32'h3bc45e31),
	.w8(32'h3caf8606),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ed32e),
	.w1(32'h3bafd027),
	.w2(32'h3af27d75),
	.w3(32'h3c770716),
	.w4(32'h3baec7d7),
	.w5(32'hbbfe22ee),
	.w6(32'hbbb402c9),
	.w7(32'hbac7d673),
	.w8(32'hbbd13744),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947270),
	.w1(32'h3b5c4b7d),
	.w2(32'h3a7b1e3e),
	.w3(32'hba9fc322),
	.w4(32'hbbadb78d),
	.w5(32'h3a688bf5),
	.w6(32'h3a03f483),
	.w7(32'h39ba9f7f),
	.w8(32'h3b3ba83a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3891c7),
	.w1(32'hbc1ea721),
	.w2(32'h3c4a9eef),
	.w3(32'hba7d097f),
	.w4(32'h3c775630),
	.w5(32'hbc1f3d89),
	.w6(32'h3b90060e),
	.w7(32'hbbbe2730),
	.w8(32'hbb32a706),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43337),
	.w1(32'h3c82eabe),
	.w2(32'h3b033fb5),
	.w3(32'h3b727300),
	.w4(32'h3c427ecf),
	.w5(32'hbcd176db),
	.w6(32'h3c54dc42),
	.w7(32'h39b8b7f6),
	.w8(32'hbae51b4f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc7c8a),
	.w1(32'h3bbece1c),
	.w2(32'h3bf6c16c),
	.w3(32'hbbead1b7),
	.w4(32'h3c5b975c),
	.w5(32'h3ba7e99f),
	.w6(32'h3b9e7147),
	.w7(32'hbb6c5db3),
	.w8(32'hbaa9c4f2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba46d9),
	.w1(32'h3aeae512),
	.w2(32'hbbe2d06e),
	.w3(32'h3a4bc09b),
	.w4(32'hb9df1d0a),
	.w5(32'h3cbecdb0),
	.w6(32'h3c072014),
	.w7(32'h3a81b046),
	.w8(32'h3b4c6371),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4c86),
	.w1(32'hbc2bc669),
	.w2(32'hbb4fe394),
	.w3(32'h3b236ff1),
	.w4(32'h3bb5c7c1),
	.w5(32'h3c1918f0),
	.w6(32'hbbe10bc2),
	.w7(32'h3bc4cf46),
	.w8(32'hbb39ed72),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5054e),
	.w1(32'hba3cfe11),
	.w2(32'h3b28b009),
	.w3(32'hba97ce33),
	.w4(32'h3bb94f7a),
	.w5(32'hbbfd0f4c),
	.w6(32'h3a24405a),
	.w7(32'hbb8347d8),
	.w8(32'hbc27c15e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc66c75),
	.w1(32'hbb8f5e27),
	.w2(32'hbc8f5097),
	.w3(32'hbbbdd8a9),
	.w4(32'hbc2e20a8),
	.w5(32'h3caa66a6),
	.w6(32'hbb231380),
	.w7(32'h39d5a254),
	.w8(32'hba632010),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391dc5b4),
	.w1(32'h3b0da3aa),
	.w2(32'hbb9fb51e),
	.w3(32'h3b50280e),
	.w4(32'hbc4815fc),
	.w5(32'h39872e82),
	.w6(32'hbc3ecfa7),
	.w7(32'hba739e3c),
	.w8(32'hbbcc72e0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5e43f),
	.w1(32'h3ae89231),
	.w2(32'h3c08d203),
	.w3(32'h3aefbc9a),
	.w4(32'h3aba8772),
	.w5(32'hba9614f5),
	.w6(32'hbbf52588),
	.w7(32'hba97c972),
	.w8(32'h3b96b6d4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a3445),
	.w1(32'h3ab01083),
	.w2(32'h3bfa2ad2),
	.w3(32'h3b18031d),
	.w4(32'h3b09e934),
	.w5(32'hbb91b9fd),
	.w6(32'h3ba7ebff),
	.w7(32'hbbb32a21),
	.w8(32'h3918efd0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4d943),
	.w1(32'hbbc371d4),
	.w2(32'hbc258fb1),
	.w3(32'hb93a83fb),
	.w4(32'hbadcbeb4),
	.w5(32'h3ba377dd),
	.w6(32'h3b6127b7),
	.w7(32'h3bb67e1c),
	.w8(32'h3c328d83),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d25ee),
	.w1(32'hbc18bb96),
	.w2(32'hba643e17),
	.w3(32'hbb50ce71),
	.w4(32'h3a215f8a),
	.w5(32'h3c80c866),
	.w6(32'h3b85c1b2),
	.w7(32'hba3a508a),
	.w8(32'hbaa5c936),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d1cc),
	.w1(32'h3acae5d1),
	.w2(32'h3bf6487f),
	.w3(32'h3b7c6c09),
	.w4(32'h3bc6b351),
	.w5(32'hbbc7ec0d),
	.w6(32'h3a8eb3ef),
	.w7(32'hbc05d416),
	.w8(32'hbb75735f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae82f0),
	.w1(32'hba8a9508),
	.w2(32'h3bf199e3),
	.w3(32'h3bfdb2d6),
	.w4(32'h3c469821),
	.w5(32'h3ac84f83),
	.w6(32'h3c60c1af),
	.w7(32'h3a9a61c5),
	.w8(32'h3a6b7356),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb271),
	.w1(32'h3b8c1571),
	.w2(32'h3bd0f7cd),
	.w3(32'h3ad47938),
	.w4(32'h3b5416bd),
	.w5(32'hbc5a92b9),
	.w6(32'hbac90667),
	.w7(32'hbbdd1d22),
	.w8(32'hbc165edb),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8ffde),
	.w1(32'h3b821780),
	.w2(32'h3bb3c9b8),
	.w3(32'hbb774be8),
	.w4(32'h3be16d71),
	.w5(32'hbb2f24c5),
	.w6(32'h3b489b22),
	.w7(32'hbaa1a29e),
	.w8(32'hbba07b4a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa48b),
	.w1(32'hbc005b48),
	.w2(32'hbbba7da5),
	.w3(32'hbb459a2a),
	.w4(32'hbb211fbb),
	.w5(32'hbc489864),
	.w6(32'hba9132bd),
	.w7(32'hbbb70386),
	.w8(32'hbbc4f583),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4afa8),
	.w1(32'h3bc42d0c),
	.w2(32'h3b68eccd),
	.w3(32'hbc1d235b),
	.w4(32'h3a6506c1),
	.w5(32'h3bb68327),
	.w6(32'h3a35b45b),
	.w7(32'hbb844ab1),
	.w8(32'hbb0f182f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26fdce),
	.w1(32'hbbb7d855),
	.w2(32'hbb9636f1),
	.w3(32'hb9dad948),
	.w4(32'hbbc02d3d),
	.w5(32'hbbaac882),
	.w6(32'hbc1e4b5f),
	.w7(32'hbbd254b4),
	.w8(32'hbb1b0d94),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4053),
	.w1(32'h3b44e62a),
	.w2(32'hbc013609),
	.w3(32'h3873405d),
	.w4(32'h3a950396),
	.w5(32'hbc0fd27c),
	.w6(32'h3bc96caf),
	.w7(32'h3bba9a14),
	.w8(32'h3a7422e8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb94f),
	.w1(32'h3b12ef9e),
	.w2(32'h3c1c5b11),
	.w3(32'hbbbb5cc3),
	.w4(32'h3bbb6c1b),
	.w5(32'hbb266e7a),
	.w6(32'hbb0e4c95),
	.w7(32'h3a7a54aa),
	.w8(32'h3b9d1be3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac02fd3),
	.w1(32'h3a89e56f),
	.w2(32'hbb5f311c),
	.w3(32'h3b433e79),
	.w4(32'h3b2735f1),
	.w5(32'h3adbe17c),
	.w6(32'h3c8feb13),
	.w7(32'h3a185a4c),
	.w8(32'hbaa2de67),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25fa52),
	.w1(32'hba94a313),
	.w2(32'hbc06e115),
	.w3(32'hbb3b72a8),
	.w4(32'hbc51dbd3),
	.w5(32'hbc0689b9),
	.w6(32'hbaaa67a2),
	.w7(32'hbbd434c0),
	.w8(32'hbafa658e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80c77c),
	.w1(32'hbba3b86e),
	.w2(32'hbb16b8b3),
	.w3(32'hbb4e8319),
	.w4(32'h3aeac040),
	.w5(32'hbaa4bddf),
	.w6(32'h3bd911aa),
	.w7(32'hbb8148d5),
	.w8(32'hbb827696),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932cca6),
	.w1(32'hbbe1b00c),
	.w2(32'hbb83086f),
	.w3(32'h3bafc97d),
	.w4(32'hbbb3f636),
	.w5(32'h3b28e958),
	.w6(32'h3b02d5f4),
	.w7(32'hbafd616a),
	.w8(32'hbad172a7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8301b9),
	.w1(32'hbc405808),
	.w2(32'hbc4efddc),
	.w3(32'h3b8947e3),
	.w4(32'hbc00d7bc),
	.w5(32'h3ba45d53),
	.w6(32'hbbc7cd5d),
	.w7(32'hba5d540f),
	.w8(32'h3b901991),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbac4f),
	.w1(32'h3b8a97ff),
	.w2(32'h3ba5c1a3),
	.w3(32'hbba89237),
	.w4(32'h3bbdbcd4),
	.w5(32'hbbbfec0f),
	.w6(32'hbbe3bbe1),
	.w7(32'hbc0786a8),
	.w8(32'hbbc9ae66),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba42bd9),
	.w1(32'h3a432d11),
	.w2(32'h3b9b1340),
	.w3(32'hbb43960f),
	.w4(32'h3c3388ec),
	.w5(32'hbb63f218),
	.w6(32'h3b9701a3),
	.w7(32'hbbd1b742),
	.w8(32'hbb1cc94c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94468d),
	.w1(32'hb9c65726),
	.w2(32'h3b9b6330),
	.w3(32'hbb98f830),
	.w4(32'hbc24353c),
	.w5(32'h3c93eee1),
	.w6(32'h3bb716b8),
	.w7(32'h3bc7149c),
	.w8(32'h3aca1048),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed6fab),
	.w1(32'hbc89eabe),
	.w2(32'hbc8de514),
	.w3(32'h3bca56ab),
	.w4(32'hbc5f2f56),
	.w5(32'h3ce27864),
	.w6(32'hbc24f517),
	.w7(32'h3c18c024),
	.w8(32'h3be779c9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbccc8),
	.w1(32'hbba6dd5d),
	.w2(32'hbb71188c),
	.w3(32'h3b9be8d9),
	.w4(32'h3bc75b5b),
	.w5(32'hbb6027ff),
	.w6(32'hbc3766f2),
	.w7(32'h3b927052),
	.w8(32'hbbe2b6ab),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072de8),
	.w1(32'hbb54a81a),
	.w2(32'hbbd121e0),
	.w3(32'hbb864fcd),
	.w4(32'hbc05de6b),
	.w5(32'h3c83b169),
	.w6(32'hbaaf9a6c),
	.w7(32'h3c426d09),
	.w8(32'h3c21ded8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130f9b),
	.w1(32'h3b30278c),
	.w2(32'h3c778a1d),
	.w3(32'hbb8b7eb3),
	.w4(32'h3c2c267e),
	.w5(32'hbbe7d533),
	.w6(32'hbbf0fbd0),
	.w7(32'hbb81909b),
	.w8(32'hbb9a020d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65e145),
	.w1(32'h3b542d83),
	.w2(32'hbc2e7d13),
	.w3(32'hbb427703),
	.w4(32'hbb80c48d),
	.w5(32'h3bd13e90),
	.w6(32'h3bd0215f),
	.w7(32'h3c3260bf),
	.w8(32'h3be6dbc8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac53cf),
	.w1(32'h3c0d4c64),
	.w2(32'hbc5c3c77),
	.w3(32'hb923d566),
	.w4(32'hbc5bff21),
	.w5(32'hbb89e73b),
	.w6(32'hbbcb5346),
	.w7(32'hbb8c6886),
	.w8(32'h3be6bba4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9f9e5),
	.w1(32'hbb345f9f),
	.w2(32'h3bef67d3),
	.w3(32'h3c09beb6),
	.w4(32'h3a9006f1),
	.w5(32'h3b76d258),
	.w6(32'hbb9516cd),
	.w7(32'hbad31b75),
	.w8(32'h3ac811d5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00225d),
	.w1(32'hbbe3d107),
	.w2(32'hbcda68f5),
	.w3(32'h3a0b400b),
	.w4(32'hbc806125),
	.w5(32'h3d14eea0),
	.w6(32'h3a4fbffa),
	.w7(32'hb8143b1f),
	.w8(32'h3c1ff294),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae13aa4),
	.w1(32'h3b233bd5),
	.w2(32'hba9eb834),
	.w3(32'h3c0a927e),
	.w4(32'h3a0d7029),
	.w5(32'hbb2489f5),
	.w6(32'hbba830a3),
	.w7(32'h3b0339f4),
	.w8(32'h3be2191a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf480dd),
	.w1(32'h3b75863a),
	.w2(32'h3bcf9c87),
	.w3(32'h39d0829c),
	.w4(32'h3c09d863),
	.w5(32'hbbb95dce),
	.w6(32'hbbc11cc5),
	.w7(32'hbbefa02a),
	.w8(32'hbadc2e71),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22f5b),
	.w1(32'h3a2b434c),
	.w2(32'h3bb40619),
	.w3(32'h3b5301a6),
	.w4(32'h39470970),
	.w5(32'h3bdfbb1f),
	.w6(32'h3be268da),
	.w7(32'hbb181de1),
	.w8(32'h3b007bba),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa8771),
	.w1(32'h3a37aa72),
	.w2(32'hbb866097),
	.w3(32'h3baffd7a),
	.w4(32'hbbf407e3),
	.w5(32'h3c7cf7a4),
	.w6(32'h3bdf4717),
	.w7(32'hbba7b2dd),
	.w8(32'h3bbb148b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcab1b8),
	.w1(32'hbb570a68),
	.w2(32'h3a832416),
	.w3(32'h3bb09fe5),
	.w4(32'hbc2cc5df),
	.w5(32'h3a58efc2),
	.w6(32'hbbafa21c),
	.w7(32'hbbd40ba1),
	.w8(32'h3b3d76dd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a409c2),
	.w1(32'h3c10330e),
	.w2(32'hb7c14ee4),
	.w3(32'h3a311cce),
	.w4(32'hbb8cf3e8),
	.w5(32'hbcda11a4),
	.w6(32'h3bc26de8),
	.w7(32'hbc66b690),
	.w8(32'hbbe3cc41),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38d36e),
	.w1(32'hbbd123a9),
	.w2(32'hbc1e12de),
	.w3(32'hbbae0b8f),
	.w4(32'hbb98de8b),
	.w5(32'h3c0e1f6b),
	.w6(32'h3c549fb1),
	.w7(32'h3c11f4ba),
	.w8(32'h3c036577),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6520c8),
	.w1(32'h3b29529e),
	.w2(32'hbbac7406),
	.w3(32'hb97b1dd4),
	.w4(32'hbc24756a),
	.w5(32'h3b7b23e3),
	.w6(32'hbb6a3ae6),
	.w7(32'hbb877f57),
	.w8(32'hbb483a3e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4ff9a),
	.w1(32'hbb30639d),
	.w2(32'h3bd3ade6),
	.w3(32'h3b92f5cd),
	.w4(32'h3b08af78),
	.w5(32'hb99da24d),
	.w6(32'h3bb4fd99),
	.w7(32'h3b2adae2),
	.w8(32'h3b2d1cd1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4658e5),
	.w1(32'h3c180569),
	.w2(32'h3c23e21f),
	.w3(32'hb8f877af),
	.w4(32'h3c50b53d),
	.w5(32'hbc0b6f74),
	.w6(32'h3b501ab1),
	.w7(32'h3a62be09),
	.w8(32'hbc17efa3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb645665),
	.w1(32'h3b35afec),
	.w2(32'hbbec43a4),
	.w3(32'hbb878d27),
	.w4(32'h3b86f4b2),
	.w5(32'hbc40e9cb),
	.w6(32'h3ba33d81),
	.w7(32'h3b8d08a4),
	.w8(32'hbb9560f4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0de345),
	.w1(32'h39eabf46),
	.w2(32'hbb169c07),
	.w3(32'hbbb80afb),
	.w4(32'hbbfd4fb3),
	.w5(32'h3a878e43),
	.w6(32'hbb2ee286),
	.w7(32'h3b260656),
	.w8(32'h3a80fdfe),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8d46a),
	.w1(32'h3b2ed3eb),
	.w2(32'hbb114938),
	.w3(32'hbba8fec0),
	.w4(32'hbb84e7ef),
	.w5(32'h3b6db827),
	.w6(32'hbb86ccdd),
	.w7(32'h3bcb9ba0),
	.w8(32'h3ac6b029),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec06e2),
	.w1(32'h3b16fd93),
	.w2(32'h3b1ca149),
	.w3(32'hba99511a),
	.w4(32'h3bf7f8ac),
	.w5(32'hbb18c4a7),
	.w6(32'hb8888c43),
	.w7(32'hbb7c6fe6),
	.w8(32'hbbadb838),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14cb8f),
	.w1(32'h3b8ee265),
	.w2(32'h3b55efe4),
	.w3(32'h3ace431f),
	.w4(32'h3bbce6fd),
	.w5(32'h39f66620),
	.w6(32'hb9d0552c),
	.w7(32'h3b8f9cbc),
	.w8(32'hbb0ae9c5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a691ccb),
	.w1(32'h3baa841e),
	.w2(32'h3b6ecfe1),
	.w3(32'h3ab189d8),
	.w4(32'h38ed3989),
	.w5(32'hbac07b61),
	.w6(32'h39c13024),
	.w7(32'h3aa36543),
	.w8(32'h3b517fc8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359e61),
	.w1(32'h3a3fe2a9),
	.w2(32'h3b90cb07),
	.w3(32'hbb84b666),
	.w4(32'h3bb0da91),
	.w5(32'h3c073fb3),
	.w6(32'hbc082c7a),
	.w7(32'h3aa3a7d5),
	.w8(32'hbae3025b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b697c1a),
	.w1(32'h3919fe62),
	.w2(32'hbb191e95),
	.w3(32'h3bec387c),
	.w4(32'h3c01c421),
	.w5(32'hbb1ceda2),
	.w6(32'h3b644e3c),
	.w7(32'h39cf4df2),
	.w8(32'h3a88d6b1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6441cc),
	.w1(32'h3bb7a551),
	.w2(32'h3c13faad),
	.w3(32'hba960931),
	.w4(32'h3c2ed356),
	.w5(32'hbc5abf27),
	.w6(32'h39769de8),
	.w7(32'h3b6b7891),
	.w8(32'hbb5c1569),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45db84),
	.w1(32'hbb76f6d8),
	.w2(32'hbca783dc),
	.w3(32'hbbec31fa),
	.w4(32'hbaea8eea),
	.w5(32'h3cae66f3),
	.w6(32'h3b3decf4),
	.w7(32'hba20bf5c),
	.w8(32'h3ba332be),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9558ab),
	.w1(32'h3b82a978),
	.w2(32'h3b96de39),
	.w3(32'h3c247985),
	.w4(32'h3b9ce892),
	.w5(32'hbc084040),
	.w6(32'hbae375eb),
	.w7(32'hbb1adea5),
	.w8(32'hbb90593c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8085c),
	.w1(32'h3b7a6f6e),
	.w2(32'hbb8a423c),
	.w3(32'hbb7d55be),
	.w4(32'h3b57a8b9),
	.w5(32'h3bdbf280),
	.w6(32'h39569e6b),
	.w7(32'h3b680a97),
	.w8(32'h3b9e891c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe11a),
	.w1(32'h3b14a7fd),
	.w2(32'h3beb29bb),
	.w3(32'h3bb1a258),
	.w4(32'h3c0c0312),
	.w5(32'hbcaad1bb),
	.w6(32'h39cedeb0),
	.w7(32'hbc7274bc),
	.w8(32'hbc275bce),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88346b),
	.w1(32'hbbfb1277),
	.w2(32'hbbb7aaa7),
	.w3(32'hbbfa6d57),
	.w4(32'hbc03594f),
	.w5(32'h3b951394),
	.w6(32'h3bb22a79),
	.w7(32'h3b383104),
	.w8(32'h3c1d7ec0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8792b),
	.w1(32'h3b96ca0e),
	.w2(32'h3ab3641c),
	.w3(32'h3b720e4b),
	.w4(32'hbba8290e),
	.w5(32'h3c44385b),
	.w6(32'h3c15adb7),
	.w7(32'hbbaee065),
	.w8(32'h3c59d4ff),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdab7e),
	.w1(32'h3ba0ba19),
	.w2(32'hbc13647d),
	.w3(32'h3c62ff0d),
	.w4(32'hbba7bbf4),
	.w5(32'h3b64e7a1),
	.w6(32'h3c3bf462),
	.w7(32'h3b3bf3dd),
	.w8(32'hba159fab),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b170),
	.w1(32'h3b73c42b),
	.w2(32'hba8a184c),
	.w3(32'hba467c0e),
	.w4(32'h3b966200),
	.w5(32'h3a212af6),
	.w6(32'hbbd2772e),
	.w7(32'hb94cfa9a),
	.w8(32'hbb830176),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b58ea),
	.w1(32'hbb37d467),
	.w2(32'hbac03dab),
	.w3(32'hb9618c2d),
	.w4(32'hbb585363),
	.w5(32'h3ae63be2),
	.w6(32'hbba6fa7e),
	.w7(32'h3a5c7e88),
	.w8(32'h3b95547f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160283),
	.w1(32'hbac9eae2),
	.w2(32'hbbbb9fc2),
	.w3(32'h3c0adacc),
	.w4(32'h39272470),
	.w5(32'h3b73d207),
	.w6(32'h3bf77bc6),
	.w7(32'h3baf3322),
	.w8(32'h3b731514),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07391d),
	.w1(32'hbbb175eb),
	.w2(32'hbc0198f3),
	.w3(32'h3b6881b6),
	.w4(32'hbbd7507d),
	.w5(32'hbc03dd80),
	.w6(32'h3a26e85d),
	.w7(32'hbbd71c7c),
	.w8(32'hbc1c4afa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba23aeb),
	.w1(32'hbc30ea7a),
	.w2(32'hba810417),
	.w3(32'hbbf79e68),
	.w4(32'hbc7dfce1),
	.w5(32'hbbf2f148),
	.w6(32'hbc0271c3),
	.w7(32'hbca5169d),
	.w8(32'hbc0374ad),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeaae1),
	.w1(32'h3af9f0f2),
	.w2(32'h3c004e93),
	.w3(32'hbc820fe6),
	.w4(32'hbbc1fc33),
	.w5(32'hbb4fb55c),
	.w6(32'hbc9809f7),
	.w7(32'hb936d43b),
	.w8(32'h3bb4f5eb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe83f8),
	.w1(32'hb92b4d38),
	.w2(32'hbc0c2e41),
	.w3(32'h396cd059),
	.w4(32'hbae87a69),
	.w5(32'hbbc14cba),
	.w6(32'h3bbd757f),
	.w7(32'hbc100638),
	.w8(32'hbbe784c0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28be9e),
	.w1(32'h3a9c70be),
	.w2(32'hb9ef2790),
	.w3(32'hbbac50f0),
	.w4(32'hb9676dd5),
	.w5(32'h3ad6f01b),
	.w6(32'hbb7c2c38),
	.w7(32'hbb349291),
	.w8(32'hb98a9c37),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fbd34),
	.w1(32'h3b137fb7),
	.w2(32'h3b980f60),
	.w3(32'h3b428f38),
	.w4(32'h3bc8ba4c),
	.w5(32'h3c01be86),
	.w6(32'h3acd8a26),
	.w7(32'h3b2f44db),
	.w8(32'h3b98e51d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23a0db),
	.w1(32'hba8b5546),
	.w2(32'h3ab9bc8e),
	.w3(32'h3c0f7295),
	.w4(32'h3ab30bab),
	.w5(32'h3ba00dad),
	.w6(32'h3b724021),
	.w7(32'hbb64403d),
	.w8(32'h3b7562e0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9cb3f),
	.w1(32'h3a6b255a),
	.w2(32'hb9b9afe1),
	.w3(32'h3bacacaf),
	.w4(32'hbb7195a6),
	.w5(32'h39516f7c),
	.w6(32'h3aca29c0),
	.w7(32'hbab1d61c),
	.w8(32'hbb4d6783),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b569e9e),
	.w1(32'h3b8593b5),
	.w2(32'h3b11e0f3),
	.w3(32'h39448635),
	.w4(32'h3b4d5cd5),
	.w5(32'h3add7909),
	.w6(32'h3a0f6b71),
	.w7(32'h3b8640ef),
	.w8(32'h3b303a88),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2972de),
	.w1(32'hbc0f3fe4),
	.w2(32'hbc096d14),
	.w3(32'h3b151f6a),
	.w4(32'hbc296fab),
	.w5(32'hbc48cb8e),
	.w6(32'h3b9b5cb4),
	.w7(32'hbc0d11e0),
	.w8(32'hbc1892e6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf55bd5),
	.w1(32'h3c34095b),
	.w2(32'h3bb6e03a),
	.w3(32'hbc4beb9a),
	.w4(32'h3c81bb54),
	.w5(32'h3c075668),
	.w6(32'hbc1d0cc3),
	.w7(32'h3c82fafd),
	.w8(32'h3b2a393b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04a1c9),
	.w1(32'hbad29758),
	.w2(32'hb98fe328),
	.w3(32'h3c02d6ac),
	.w4(32'h3aaed79d),
	.w5(32'h3a513107),
	.w6(32'h3a2f84c9),
	.w7(32'h3a6e7f05),
	.w8(32'h3b3efb8d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbc52c),
	.w1(32'hbc4f8a5a),
	.w2(32'h39c24c85),
	.w3(32'hbb269e84),
	.w4(32'hbc6439b6),
	.w5(32'hbabcb86f),
	.w6(32'h3ad7c4b9),
	.w7(32'hbc5223c9),
	.w8(32'h3b04cec2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b65e5),
	.w1(32'h3b8e5e7c),
	.w2(32'hb9a79a76),
	.w3(32'hba00b0dc),
	.w4(32'h3ba3e02a),
	.w5(32'h3b28077f),
	.w6(32'h3b2347ae),
	.w7(32'h3b998f3f),
	.w8(32'h3b7f48bb),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63ed58),
	.w1(32'hbc1ad1ae),
	.w2(32'hbba248bb),
	.w3(32'hbb57aabe),
	.w4(32'hbbef5c81),
	.w5(32'hbb009c31),
	.w6(32'hba7ca6f8),
	.w7(32'hbb4913a2),
	.w8(32'hbc10ec41),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238241),
	.w1(32'hb91ceaea),
	.w2(32'hbbdd2659),
	.w3(32'h3b033690),
	.w4(32'hba3eab57),
	.w5(32'hbbe69152),
	.w6(32'hba5640b3),
	.w7(32'h3b93b28e),
	.w8(32'hbb4187b7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa292ea),
	.w1(32'hbacccbb1),
	.w2(32'hbace5e96),
	.w3(32'h39bcde57),
	.w4(32'h3ab0a5df),
	.w5(32'h3b310997),
	.w6(32'h3bbd304b),
	.w7(32'hba1b5dee),
	.w8(32'h3af16fa8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c98cdc),
	.w1(32'hbc1a6b5e),
	.w2(32'hbbaf5f63),
	.w3(32'h391b85f1),
	.w4(32'hbbe10d30),
	.w5(32'hbab6a3ca),
	.w6(32'h3b76924d),
	.w7(32'hbc21975d),
	.w8(32'hbc051384),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac43705),
	.w1(32'hbabc608a),
	.w2(32'hbb29090e),
	.w3(32'h3b4e1918),
	.w4(32'h3ad31dd5),
	.w5(32'h3b087fae),
	.w6(32'hbb2bb7c6),
	.w7(32'hb9eec1f9),
	.w8(32'h3a4da00e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b033703),
	.w1(32'h3af81840),
	.w2(32'h3ac1e37f),
	.w3(32'hbb517417),
	.w4(32'h3b28c4db),
	.w5(32'h3790ac29),
	.w6(32'hbb6870ba),
	.w7(32'h39ef1d09),
	.w8(32'h3ba994d4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04602),
	.w1(32'h3a6730c5),
	.w2(32'h3b02a348),
	.w3(32'hba11242c),
	.w4(32'h3b31305d),
	.w5(32'h3b5a65ed),
	.w6(32'h3b27b869),
	.w7(32'h3b082642),
	.w8(32'h3b8b6729),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11bf83),
	.w1(32'hbb69849b),
	.w2(32'h3b1d6e9a),
	.w3(32'h3b73cca5),
	.w4(32'h3a39b58b),
	.w5(32'h3c0a3907),
	.w6(32'h3b8bead1),
	.w7(32'hbad4c7fa),
	.w8(32'h3bbc95bc),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d24c1),
	.w1(32'hba265c19),
	.w2(32'hbba03ab8),
	.w3(32'h3bf5eda0),
	.w4(32'hbb712fa7),
	.w5(32'hbc0bbd72),
	.w6(32'h3bc64ba3),
	.w7(32'h3ba60afe),
	.w8(32'hbb0d812a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa716e4),
	.w1(32'h3c378aaf),
	.w2(32'h3a94777d),
	.w3(32'hbc0b9c74),
	.w4(32'h3bafc070),
	.w5(32'hbbcb9949),
	.w6(32'hbba478d3),
	.w7(32'hbb73d01e),
	.w8(32'hbbbd4302),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9dd9e),
	.w1(32'h3a82dbe7),
	.w2(32'h3b1946ee),
	.w3(32'hbb85e43e),
	.w4(32'hbb3084bb),
	.w5(32'h38635cc5),
	.w6(32'hbacec11c),
	.w7(32'hbbdcff7d),
	.w8(32'h3b2edbeb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380321ab),
	.w1(32'hbc26f180),
	.w2(32'hbc4d6c74),
	.w3(32'hbbe192f7),
	.w4(32'hbc0d3a1d),
	.w5(32'hbbac9a96),
	.w6(32'hbbc0833c),
	.w7(32'hbbc5f569),
	.w8(32'hbbfe75e3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb601d33),
	.w1(32'hbb2be40f),
	.w2(32'hbb44f0b3),
	.w3(32'h3b18a537),
	.w4(32'h3a290a68),
	.w5(32'hbab9ae58),
	.w6(32'h3a09ab21),
	.w7(32'h3ab11ebf),
	.w8(32'hbb4d2e3f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeec013),
	.w1(32'h39b3cd3e),
	.w2(32'h3a8a969d),
	.w3(32'hbc157dcd),
	.w4(32'hba86bffb),
	.w5(32'h3a140f2f),
	.w6(32'hbc10e653),
	.w7(32'hbaaea70f),
	.w8(32'h3a804680),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b29719),
	.w1(32'hbb9d7bf6),
	.w2(32'h3a84a51d),
	.w3(32'h391dd0ea),
	.w4(32'hbbae8512),
	.w5(32'h3bc62b06),
	.w6(32'hbb3491d1),
	.w7(32'hbc0aa14d),
	.w8(32'h3ba9985a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157c2a),
	.w1(32'hbbd9e512),
	.w2(32'hbbb09b14),
	.w3(32'h3bc6f42a),
	.w4(32'hbc2480bb),
	.w5(32'hbb52c300),
	.w6(32'h3bd05c98),
	.w7(32'hbc0e13a1),
	.w8(32'hbb318b97),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a940a),
	.w1(32'hbb504b75),
	.w2(32'hbc80dd4e),
	.w3(32'h3ba87dba),
	.w4(32'h3ae971ee),
	.w5(32'hbbf1a884),
	.w6(32'h3a620dbb),
	.w7(32'h3c413445),
	.w8(32'hbbb533a5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7b8cf),
	.w1(32'hbc85a6ce),
	.w2(32'h3bc75098),
	.w3(32'h3c187cae),
	.w4(32'hbc8f9f08),
	.w5(32'h3c3d9824),
	.w6(32'h3b533cc3),
	.w7(32'hbc90c49f),
	.w8(32'h3c7adc91),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab494),
	.w1(32'h3c00cf69),
	.w2(32'h3bac3202),
	.w3(32'hbbd23fa8),
	.w4(32'h3c25188a),
	.w5(32'h3bc9b1ce),
	.w6(32'hbc14b8d4),
	.w7(32'h3b70fb62),
	.w8(32'hba8fdffe),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e58b9),
	.w1(32'h3a195406),
	.w2(32'hbbac933c),
	.w3(32'hbb7b6424),
	.w4(32'h3ad41783),
	.w5(32'hbbb2ce6f),
	.w6(32'hbb84c480),
	.w7(32'h3ae97677),
	.w8(32'hbb5e2e4b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedfc1e),
	.w1(32'h3a991286),
	.w2(32'hbb0557d3),
	.w3(32'hbc22f97c),
	.w4(32'h3a7e4022),
	.w5(32'hbb45686a),
	.w6(32'hbbb5350c),
	.w7(32'hbbad68d9),
	.w8(32'hbbf7c940),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43b913),
	.w1(32'hbaeeff2f),
	.w2(32'h3a9107cb),
	.w3(32'hba21f9ec),
	.w4(32'hbb383d80),
	.w5(32'h3a89adb1),
	.w6(32'hbb179b7b),
	.w7(32'hb9e4ad2d),
	.w8(32'hbaca34ce),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1ade1),
	.w1(32'h3a870446),
	.w2(32'hbb3f8756),
	.w3(32'hbb8efbaf),
	.w4(32'hbb3489b3),
	.w5(32'hbbf86b6e),
	.w6(32'hbb59acbf),
	.w7(32'hbb4eed95),
	.w8(32'hbbfcf768),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa4a1),
	.w1(32'h3b0bb236),
	.w2(32'hba96d0ad),
	.w3(32'hbbbe9475),
	.w4(32'h3b856521),
	.w5(32'hbb7f3165),
	.w6(32'hbbe386bf),
	.w7(32'h3c0d1a8a),
	.w8(32'hbb2d795c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a2e34),
	.w1(32'h381914a7),
	.w2(32'h3b4d74bf),
	.w3(32'h3c0e4af8),
	.w4(32'hbb4712eb),
	.w5(32'h3b61749c),
	.w6(32'h3bfc2ca3),
	.w7(32'hbba24f82),
	.w8(32'h3b3d4ad1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c62722),
	.w1(32'h3c035d0c),
	.w2(32'h3a839ea5),
	.w3(32'hb7f1a809),
	.w4(32'h3bb909b9),
	.w5(32'h3b0fe3c3),
	.w6(32'hba0c3c6a),
	.w7(32'h3bc33446),
	.w8(32'h3b006804),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5e958),
	.w1(32'hbc04b5eb),
	.w2(32'hbb867219),
	.w3(32'hbbc96bfa),
	.w4(32'hbc10dc27),
	.w5(32'hbb559ac0),
	.w6(32'hbbb1c2ed),
	.w7(32'hba925ee8),
	.w8(32'h3a02fe54),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada79fa),
	.w1(32'hbb2b2cf1),
	.w2(32'h3b7ed19b),
	.w3(32'h3ae1626b),
	.w4(32'hba9feca7),
	.w5(32'h3c1055c8),
	.w6(32'h39bf1313),
	.w7(32'hbbf210a3),
	.w8(32'h3c06be3f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f3894),
	.w1(32'hbb39b4b6),
	.w2(32'h3b14eede),
	.w3(32'hbc85cbfd),
	.w4(32'hb88cf8e1),
	.w5(32'h3c4a7822),
	.w6(32'hbc64adca),
	.w7(32'hbb50e2b4),
	.w8(32'h3bd6006f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70b01c),
	.w1(32'h3a2d4193),
	.w2(32'hb9af91c5),
	.w3(32'h3b6da96f),
	.w4(32'hbb862f6b),
	.w5(32'hbafa9552),
	.w6(32'hbaaa9524),
	.w7(32'hba74d92d),
	.w8(32'h3aaa0fbf),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c523),
	.w1(32'h3b080ab6),
	.w2(32'hbb692876),
	.w3(32'h3a011357),
	.w4(32'h3bc07c94),
	.w5(32'hbb65c811),
	.w6(32'h3ade35ab),
	.w7(32'h3b31baca),
	.w8(32'h3aec4cfc),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25f60d),
	.w1(32'hbbe57a39),
	.w2(32'hbbe2341e),
	.w3(32'hbb4130de),
	.w4(32'hbbf97d1e),
	.w5(32'hbb51a3f4),
	.w6(32'h3a505a3d),
	.w7(32'hbbda7251),
	.w8(32'hb9962c20),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34b524),
	.w1(32'hb9b51f52),
	.w2(32'h3b30b8fe),
	.w3(32'hbb923e88),
	.w4(32'h3a95a525),
	.w5(32'h39999d2a),
	.w6(32'hbb25c32e),
	.w7(32'h3b9a697f),
	.w8(32'h3b6fdcaf),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf89c),
	.w1(32'hba452397),
	.w2(32'h3c06b943),
	.w3(32'h3bbca034),
	.w4(32'h3c656b13),
	.w5(32'h3d294d06),
	.w6(32'h3bb31feb),
	.w7(32'h3c3815e4),
	.w8(32'h3cbd4d8d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1a65c),
	.w1(32'h3b99ce62),
	.w2(32'h3b18e693),
	.w3(32'h3cc5f841),
	.w4(32'h3b969b6c),
	.w5(32'h3bac5ea1),
	.w6(32'h3c6a236f),
	.w7(32'h3b5546db),
	.w8(32'h3b20c8fd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c7215),
	.w1(32'h3b515e18),
	.w2(32'h39c2ab03),
	.w3(32'h3bf816ad),
	.w4(32'h3b2407ad),
	.w5(32'h3a1f6ba8),
	.w6(32'h3bcc5d32),
	.w7(32'hb7bf14f2),
	.w8(32'h3b6852ac),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3ed99),
	.w1(32'h3ba00b39),
	.w2(32'hbbee4035),
	.w3(32'h38ca025e),
	.w4(32'h3b5dd6e0),
	.w5(32'hbc205403),
	.w6(32'hb9e69e46),
	.w7(32'h3ba2eb64),
	.w8(32'hbb717d0a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7fefb),
	.w1(32'h3bb46efd),
	.w2(32'h3a65bca5),
	.w3(32'hbb2d1d63),
	.w4(32'hbb7c8197),
	.w5(32'hbbeaf2a4),
	.w6(32'h3bf6a049),
	.w7(32'hb8807ec6),
	.w8(32'h3add7415),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d583),
	.w1(32'h3baa1733),
	.w2(32'h3a6ce1c9),
	.w3(32'hbac4e4d7),
	.w4(32'hb933d2d4),
	.w5(32'hbb503e8c),
	.w6(32'h3b6f7d17),
	.w7(32'h3b943bc0),
	.w8(32'h3a100106),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5be6),
	.w1(32'h3b9d21cf),
	.w2(32'h3c1bf9be),
	.w3(32'h3b7635bb),
	.w4(32'h3a2a646a),
	.w5(32'h3c4e0173),
	.w6(32'h3b943ab7),
	.w7(32'hbac279a4),
	.w8(32'h3c13dc2e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd2551),
	.w1(32'hbb2a8e5a),
	.w2(32'h3c09563b),
	.w3(32'h3bc83dbc),
	.w4(32'hbb9abc42),
	.w5(32'h3c1d50df),
	.w6(32'h3b508b65),
	.w7(32'hbbd9660a),
	.w8(32'h3b84a570),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b80b),
	.w1(32'hbb806d2e),
	.w2(32'hbbaa6cec),
	.w3(32'h3b172244),
	.w4(32'hbb037c83),
	.w5(32'hbc0eecf0),
	.w6(32'h3a1d3fd6),
	.w7(32'hbb4f339c),
	.w8(32'hbc2928fd),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule