module layer_8_featuremap_38(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910a3f),
	.w1(32'hbbae569e),
	.w2(32'h38b6c1d2),
	.w3(32'hbbf690c4),
	.w4(32'h3839c6da),
	.w5(32'hbc481194),
	.w6(32'hbc01aa62),
	.w7(32'hbb8f336b),
	.w8(32'hbb15bf61),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6b8f9),
	.w1(32'h3a2264c3),
	.w2(32'h3b8b6396),
	.w3(32'hbb932c94),
	.w4(32'h3c1d9cd9),
	.w5(32'h3b820096),
	.w6(32'hbaac7705),
	.w7(32'h3ba3f93a),
	.w8(32'h3b334e47),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15481a),
	.w1(32'h3afd6e90),
	.w2(32'h3b9713e9),
	.w3(32'hbc17809f),
	.w4(32'h3c016581),
	.w5(32'h3b261552),
	.w6(32'hbbf44210),
	.w7(32'h3c0be4de),
	.w8(32'h3bd1aff8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbfecbd),
	.w1(32'h3a33a86c),
	.w2(32'h3c4c2373),
	.w3(32'hbb863bd5),
	.w4(32'hbb6c3a28),
	.w5(32'hbc2fe8fe),
	.w6(32'hbc9fa1c1),
	.w7(32'hbc1153b8),
	.w8(32'hbc5df7c8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8186de),
	.w1(32'hbc5c18f6),
	.w2(32'hbbfc977b),
	.w3(32'hbc042472),
	.w4(32'h3ac6f207),
	.w5(32'hbb111baa),
	.w6(32'hbc261335),
	.w7(32'h3bc521ad),
	.w8(32'h3ba11c1a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5dc69),
	.w1(32'hbc72217e),
	.w2(32'hba2002be),
	.w3(32'hbc95c00b),
	.w4(32'h3cd701d1),
	.w5(32'h3a3073b0),
	.w6(32'hbcaaabdb),
	.w7(32'h3cb25718),
	.w8(32'h3b6da748),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b698f2f),
	.w1(32'hbbe1653f),
	.w2(32'h3aaf64c2),
	.w3(32'hb62f89ea),
	.w4(32'hba0a3c97),
	.w5(32'hbb1e2e73),
	.w6(32'hba727354),
	.w7(32'hbb000862),
	.w8(32'h3ab1b628),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca19d24),
	.w1(32'hbbfba9ce),
	.w2(32'h3c031e9c),
	.w3(32'hbcce20ce),
	.w4(32'hbb32662c),
	.w5(32'hbb1a289a),
	.w6(32'hbc9b56aa),
	.w7(32'h3a88eed5),
	.w8(32'hbb3f760f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c1d45),
	.w1(32'hbc2e2637),
	.w2(32'hbbbc3f0e),
	.w3(32'hbbf839b6),
	.w4(32'hba66bf08),
	.w5(32'hbbdcdb2f),
	.w6(32'hbba98ae2),
	.w7(32'hba1a8a7b),
	.w8(32'hbc1c447b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adccb9d),
	.w1(32'h3c100a77),
	.w2(32'hb9fc8a14),
	.w3(32'hbc393dd0),
	.w4(32'h399091e1),
	.w5(32'h3c35d47d),
	.w6(32'hbd4a053e),
	.w7(32'hbb7ec19d),
	.w8(32'hbc298736),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb453e90),
	.w1(32'h3a8eac64),
	.w2(32'h3b2f2d70),
	.w3(32'hbc4e7ad5),
	.w4(32'hba2ddf2e),
	.w5(32'hbbf215f9),
	.w6(32'hbc0e87f6),
	.w7(32'hbc1b93bf),
	.w8(32'h39971736),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f3668),
	.w1(32'hbc97fb9b),
	.w2(32'hbc25db27),
	.w3(32'hbcb03f34),
	.w4(32'hbc35d062),
	.w5(32'hbca0f40e),
	.w6(32'hbca4e895),
	.w7(32'hbbda0600),
	.w8(32'hbc8f0414),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc520c4c),
	.w1(32'h3aa1a04f),
	.w2(32'h3b23c446),
	.w3(32'hbc8dc9a2),
	.w4(32'h3b96fd8d),
	.w5(32'h3b002c8f),
	.w6(32'hbc67d180),
	.w7(32'h3c06efa2),
	.w8(32'h3bef56d5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cab39),
	.w1(32'hbc907b5e),
	.w2(32'h3c0e4e85),
	.w3(32'h3c4ab534),
	.w4(32'h3c24fb3b),
	.w5(32'hbbb7c079),
	.w6(32'h3bfcb5a7),
	.w7(32'h3c9a76f6),
	.w8(32'h3ba134a6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba11ad5),
	.w1(32'hbc608882),
	.w2(32'h3bb82c43),
	.w3(32'h3c22a634),
	.w4(32'h3b2b2e1f),
	.w5(32'h3a515604),
	.w6(32'h3b2daf34),
	.w7(32'h3c8c48eb),
	.w8(32'hbb7a4643),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ee88),
	.w1(32'h3aec2fb3),
	.w2(32'hbb5b7600),
	.w3(32'h3b363b71),
	.w4(32'h3c32fef8),
	.w5(32'h3ae47e20),
	.w6(32'hb7c9e33d),
	.w7(32'hbb3b9d86),
	.w8(32'hbabcb136),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66759e),
	.w1(32'hbce5ca2b),
	.w2(32'hb9420b32),
	.w3(32'h3c7e7e09),
	.w4(32'h3ca74852),
	.w5(32'h3d073aff),
	.w6(32'h3c6d0d9f),
	.w7(32'h3bc8b87c),
	.w8(32'hbb22b890),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0b219),
	.w1(32'hbc87b5d7),
	.w2(32'hbc34cf2a),
	.w3(32'hbcbb95a7),
	.w4(32'hbbaa4787),
	.w5(32'hbc7043e3),
	.w6(32'hbccfc11f),
	.w7(32'hbbcfd57a),
	.w8(32'hbc7dff9c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5b1d95),
	.w1(32'h38b70e83),
	.w2(32'h3b6faa67),
	.w3(32'hbd6a0ff9),
	.w4(32'hbbf3cf17),
	.w5(32'hbc46f377),
	.w6(32'hbd5a363e),
	.w7(32'hbc5c863b),
	.w8(32'hbb39c4a9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd157bb0),
	.w1(32'hbd1b2018),
	.w2(32'hbd3c6060),
	.w3(32'hbd3066de),
	.w4(32'hbccbb60c),
	.w5(32'hbc342c9d),
	.w6(32'hbd03eaf0),
	.w7(32'hbc34534b),
	.w8(32'hbcac7b2f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf3ff1),
	.w1(32'hbb61020f),
	.w2(32'hbbd25150),
	.w3(32'hbc6b95e8),
	.w4(32'hbb6cc06b),
	.w5(32'h3b8da010),
	.w6(32'hbc485315),
	.w7(32'h3c1efdd7),
	.w8(32'h3c06b82a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ab29),
	.w1(32'h3a92d8f0),
	.w2(32'h3c1b3bf4),
	.w3(32'h3b14d78a),
	.w4(32'h3cb5be12),
	.w5(32'h3c8f3983),
	.w6(32'hbbd66ede),
	.w7(32'h3c98f4f0),
	.w8(32'hb9e0a0a2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb378733),
	.w1(32'h3c8fb46f),
	.w2(32'h3cb1d58d),
	.w3(32'hbc1d1d5a),
	.w4(32'hbc7502e2),
	.w5(32'h3bda54bb),
	.w6(32'hbc07cf47),
	.w7(32'hbb08ec3f),
	.w8(32'h3c2cc975),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28c3c0),
	.w1(32'hbc6f9692),
	.w2(32'hbb5aa1dc),
	.w3(32'hbbb6299e),
	.w4(32'h3c3f1f5e),
	.w5(32'h3b2ac027),
	.w6(32'h38812811),
	.w7(32'hbaf48833),
	.w8(32'hbc7633af),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ca0b),
	.w1(32'hbc681f58),
	.w2(32'hbc208a6d),
	.w3(32'hbbc838d6),
	.w4(32'h3b2220e0),
	.w5(32'h3c042624),
	.w6(32'hbc062602),
	.w7(32'h3ad1b1b2),
	.w8(32'hbc0a2cb6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb31003),
	.w1(32'h3c104b90),
	.w2(32'hbb9a7d0e),
	.w3(32'hbc9de833),
	.w4(32'hbc545b6d),
	.w5(32'hbb9b703a),
	.w6(32'hbc8b2850),
	.w7(32'hbb9ebdcb),
	.w8(32'hbba33493),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8462a),
	.w1(32'h3c2238d8),
	.w2(32'hbbce17f8),
	.w3(32'hbc020ddf),
	.w4(32'hbc26e448),
	.w5(32'hba86f361),
	.w6(32'hbb4557e1),
	.w7(32'hbbfe97a7),
	.w8(32'hbacbb843),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd543527),
	.w1(32'h3d9a0e97),
	.w2(32'h3dc2937d),
	.w3(32'hbd8a5734),
	.w4(32'h3d29d3c4),
	.w5(32'h3d35dee2),
	.w6(32'hbd9948bf),
	.w7(32'h3b0ba153),
	.w8(32'h3c656d24),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb7f1e),
	.w1(32'hbbcfe107),
	.w2(32'hbce309c7),
	.w3(32'hbc9e8450),
	.w4(32'h3c24b61f),
	.w5(32'hbcb54f02),
	.w6(32'hbbcd9318),
	.w7(32'hbc2ee9dd),
	.w8(32'h39c64787),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd06f1),
	.w1(32'hbb974228),
	.w2(32'hb932e544),
	.w3(32'hbbc9d31d),
	.w4(32'h3aee1bb9),
	.w5(32'hbab4026b),
	.w6(32'hbb5a4fef),
	.w7(32'h3b8fc312),
	.w8(32'h3c01b087),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2adec5),
	.w1(32'hbb90c550),
	.w2(32'h3c2d18e9),
	.w3(32'hbca4ab01),
	.w4(32'hbceaa0a1),
	.w5(32'h3b478601),
	.w6(32'h3c203cfd),
	.w7(32'h3c73017f),
	.w8(32'hbc200c06),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc94ebe),
	.w1(32'h3b13e12f),
	.w2(32'hbc7cfeec),
	.w3(32'hbc1df87d),
	.w4(32'h3c0eded9),
	.w5(32'h3c53be49),
	.w6(32'hbc87feb9),
	.w7(32'h3c775e0d),
	.w8(32'hbb5f1f56),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb53fed),
	.w1(32'hbbee43e7),
	.w2(32'h3cd561d8),
	.w3(32'hbc021eb5),
	.w4(32'hba907893),
	.w5(32'h3c0f0b09),
	.w6(32'hbc4ac423),
	.w7(32'hbbc00b78),
	.w8(32'h3cc4dd4d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5989b7),
	.w1(32'hbcbfee57),
	.w2(32'hbc77d9c9),
	.w3(32'h3b5a6035),
	.w4(32'h3ca1199a),
	.w5(32'h3c807b46),
	.w6(32'h3c9f4b88),
	.w7(32'h3ba4551e),
	.w8(32'h3b4e4b91),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc856394),
	.w1(32'hbca53ef3),
	.w2(32'hbc41913f),
	.w3(32'hbc5255a8),
	.w4(32'h3c418b52),
	.w5(32'hbc821bf2),
	.w6(32'hbc3c5d19),
	.w7(32'h3c9f9e1d),
	.w8(32'hbca70ea5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83dd46),
	.w1(32'hbc341003),
	.w2(32'h3b2ac8b4),
	.w3(32'hbc9cce4c),
	.w4(32'hbb994777),
	.w5(32'hbc1f51b7),
	.w6(32'hbc8f003b),
	.w7(32'hbc36a3a3),
	.w8(32'hbbdd7c42),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b5cbb),
	.w1(32'hbbd672bf),
	.w2(32'h398e80d6),
	.w3(32'hbb0bb008),
	.w4(32'h3b9f3575),
	.w5(32'hbb570119),
	.w6(32'h3a94dd72),
	.w7(32'hbbde68de),
	.w8(32'hbb08408b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac92d2),
	.w1(32'hbb7a799b),
	.w2(32'h3ba577aa),
	.w3(32'hba9e8c6a),
	.w4(32'h3b881691),
	.w5(32'h3abd01bd),
	.w6(32'h3b437131),
	.w7(32'h3c2a007d),
	.w8(32'h3cba4a4d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c973b),
	.w1(32'hbce06fd6),
	.w2(32'h3c3c6a72),
	.w3(32'h3ce0e546),
	.w4(32'h3bb8538b),
	.w5(32'h3c11f8a8),
	.w6(32'h3bb59734),
	.w7(32'h3d1869b6),
	.w8(32'hb8bbbe1e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e73f4),
	.w1(32'h3893b54d),
	.w2(32'hb9a2b368),
	.w3(32'h3b7ff5a1),
	.w4(32'hbb1561fd),
	.w5(32'h3bb5c100),
	.w6(32'hbb8ba749),
	.w7(32'h3ba85fd7),
	.w8(32'hbb83f4cc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdb496a4),
	.w1(32'hbc710c77),
	.w2(32'hbd4b0907),
	.w3(32'hbdbec463),
	.w4(32'hbd0cbfaa),
	.w5(32'hbd766be2),
	.w6(32'hbdcdddcc),
	.w7(32'hbca6fbc2),
	.w8(32'hbd2bd414),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37890a),
	.w1(32'h3baeb553),
	.w2(32'h3bfbf151),
	.w3(32'hbc649085),
	.w4(32'h3aaf19bb),
	.w5(32'h3bbbc06a),
	.w6(32'hbc4db538),
	.w7(32'h3a8e2d5b),
	.w8(32'hbb8e02da),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034324),
	.w1(32'hbae3d1ab),
	.w2(32'hba2d9ef0),
	.w3(32'hbbb42e65),
	.w4(32'h3b2d099c),
	.w5(32'hbb89fc3a),
	.w6(32'hbc2027e4),
	.w7(32'hbb19c600),
	.w8(32'h3b311ef2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca08217),
	.w1(32'hbc2265c5),
	.w2(32'hbc2de0e5),
	.w3(32'hbca5534f),
	.w4(32'hbbd11e2c),
	.w5(32'hbc08dc62),
	.w6(32'hbcb6615c),
	.w7(32'hbbd8dac4),
	.w8(32'hbc0938b6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51f9b1),
	.w1(32'h3b373905),
	.w2(32'h3be4026e),
	.w3(32'hbc323d9b),
	.w4(32'h3c1e1801),
	.w5(32'h3bf6a022),
	.w6(32'hbc65ac1d),
	.w7(32'h3b863df9),
	.w8(32'hba9df714),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d084a),
	.w1(32'h3c1f5a99),
	.w2(32'h3c218356),
	.w3(32'hbb976d3a),
	.w4(32'h3bf1e9ff),
	.w5(32'h3c1684d1),
	.w6(32'hbc0e6da6),
	.w7(32'h3b733086),
	.w8(32'h3b51797a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b781006),
	.w1(32'h3c22644a),
	.w2(32'h39d9b695),
	.w3(32'h3c2d822c),
	.w4(32'hb9796273),
	.w5(32'hbabfde8a),
	.w6(32'hba5e5acf),
	.w7(32'h3bcf6f96),
	.w8(32'hbac23301),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996f497),
	.w1(32'h3b88f51c),
	.w2(32'h3bbe186d),
	.w3(32'hba15b04d),
	.w4(32'h3b6402b1),
	.w5(32'h3accf193),
	.w6(32'hbb273cbc),
	.w7(32'h3b351348),
	.w8(32'h3b82774b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8faa7e),
	.w1(32'h3a206e1f),
	.w2(32'h3ab82e07),
	.w3(32'hbc26cfd4),
	.w4(32'h3bfd9fb9),
	.w5(32'h3bb96216),
	.w6(32'hbc60c974),
	.w7(32'h3b560966),
	.w8(32'hbaa24b79),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ee05),
	.w1(32'hbaaeedb5),
	.w2(32'hbc281f88),
	.w3(32'hbc2986b1),
	.w4(32'hbb04e5a3),
	.w5(32'hbc3d10fc),
	.w6(32'hbc85d705),
	.w7(32'hbbc1bc2f),
	.w8(32'hbc23cd9c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a3f8),
	.w1(32'h3c2bf4c6),
	.w2(32'h3c60ab3b),
	.w3(32'hbbcfab9c),
	.w4(32'h3c8c8503),
	.w5(32'h3c93cb9b),
	.w6(32'h3b9248cc),
	.w7(32'h3cc8029d),
	.w8(32'h3cc006b2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8d20ec),
	.w1(32'hbb8b3c88),
	.w2(32'h3bd00f56),
	.w3(32'hbd7a1892),
	.w4(32'h39a1bebe),
	.w5(32'hbc32c1c9),
	.w6(32'hbd7e409c),
	.w7(32'hbad892f0),
	.w8(32'hbc60d71d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1af5a),
	.w1(32'h3b5c53c4),
	.w2(32'hbb977605),
	.w3(32'hbca5f6f5),
	.w4(32'h3bb25e9d),
	.w5(32'hbb141bd5),
	.w6(32'hbc38bf78),
	.w7(32'hb9967b8a),
	.w8(32'hbb943d51),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca329e5),
	.w1(32'hbc234fa5),
	.w2(32'hbc3455ef),
	.w3(32'hbc9a7eb1),
	.w4(32'hbc2f1fb6),
	.w5(32'hbc4b1432),
	.w6(32'hbcdc39b0),
	.w7(32'hbc7fe44c),
	.w8(32'hbca5e25f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873582),
	.w1(32'hbaab4da9),
	.w2(32'hb9a609b1),
	.w3(32'h3b93010c),
	.w4(32'hbbb27f35),
	.w5(32'hbb05123a),
	.w6(32'hbb65e582),
	.w7(32'h3b1a3909),
	.w8(32'h3b2429c8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b9001),
	.w1(32'hbc40e764),
	.w2(32'hbc83c8fe),
	.w3(32'hbc490cfa),
	.w4(32'hbb712b1d),
	.w5(32'hbbd9fd2f),
	.w6(32'hbbbf5a9a),
	.w7(32'h3b4dd342),
	.w8(32'hbc47941b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf452b),
	.w1(32'hbc1d2062),
	.w2(32'hbc0324ae),
	.w3(32'hbc8f460b),
	.w4(32'hba54fdc3),
	.w5(32'hbbffecda),
	.w6(32'hbc8693e9),
	.w7(32'hb90b1a9e),
	.w8(32'hbc95b815),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1806e6),
	.w1(32'hbb7e5f84),
	.w2(32'h3c0db79f),
	.w3(32'hbd1aa2d4),
	.w4(32'hbc00afc3),
	.w5(32'hbb91a236),
	.w6(32'hbd3a06a8),
	.w7(32'hbc18432f),
	.w8(32'hbb9f5559),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ba31),
	.w1(32'h3b8ce7f7),
	.w2(32'h3c4b730c),
	.w3(32'h3b04e790),
	.w4(32'h3bf80bc0),
	.w5(32'h3c2e7ab4),
	.w6(32'h3b49a42a),
	.w7(32'h3be06dfb),
	.w8(32'h3b92a131),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b9c6b),
	.w1(32'hba911734),
	.w2(32'h39c90840),
	.w3(32'hbb9a5881),
	.w4(32'h3af79d59),
	.w5(32'hbc1a3bbf),
	.w6(32'hbbe43d71),
	.w7(32'hb963dcf2),
	.w8(32'hbb5cb875),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfca33b),
	.w1(32'hbc0b1996),
	.w2(32'h3c5fde10),
	.w3(32'h3ab67f82),
	.w4(32'h3c013578),
	.w5(32'hbb52ddc6),
	.w6(32'hbbaa3295),
	.w7(32'hb9a4f66b),
	.w8(32'hbaf811eb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19ec17),
	.w1(32'hb96786a2),
	.w2(32'hbbd65207),
	.w3(32'hba26de12),
	.w4(32'h3aba1206),
	.w5(32'hba2c5c1c),
	.w6(32'h3b123015),
	.w7(32'hbb0eb0e4),
	.w8(32'h3ab2fb5b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd45b056),
	.w1(32'hbbc8ebbe),
	.w2(32'hbc620fee),
	.w3(32'hbd351277),
	.w4(32'h3b28756a),
	.w5(32'hbbf54b25),
	.w6(32'hbd2acf30),
	.w7(32'h3ba8a131),
	.w8(32'hbc4dd04d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2559),
	.w1(32'h3bff137e),
	.w2(32'hbb579caf),
	.w3(32'hbc4df85c),
	.w4(32'h3aa8cfff),
	.w5(32'hbab9351c),
	.w6(32'hbc863187),
	.w7(32'hbbc27b58),
	.w8(32'hbb535782),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab30d8e),
	.w1(32'hb9cf1368),
	.w2(32'h3ad201d5),
	.w3(32'h3ad5c7e9),
	.w4(32'h3a19a01a),
	.w5(32'h3b37480e),
	.w6(32'h3b2a2a80),
	.w7(32'h3adacf23),
	.w8(32'h3a2fa4ce),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3988df),
	.w1(32'h3b442bc8),
	.w2(32'h3c02dc37),
	.w3(32'hbc5b6b07),
	.w4(32'h389aa5e4),
	.w5(32'h3b8b5d01),
	.w6(32'hbc4b02f1),
	.w7(32'h393e2aa4),
	.w8(32'h3b02b135),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5f0b4),
	.w1(32'hbadf1cc7),
	.w2(32'hbb3c167a),
	.w3(32'hbc7b7492),
	.w4(32'h3bec6127),
	.w5(32'h3b59fc7c),
	.w6(32'hbc83b6b8),
	.w7(32'h3c06979f),
	.w8(32'h3b6f3149),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc906353),
	.w1(32'h3bcd0615),
	.w2(32'hbb0a00fb),
	.w3(32'hbc83ffa1),
	.w4(32'h3bfad9bb),
	.w5(32'h3b6c28ff),
	.w6(32'hbc934112),
	.w7(32'h3bbb59b9),
	.w8(32'hba01244c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefd060),
	.w1(32'hbaaba15b),
	.w2(32'hbb073ce2),
	.w3(32'hbb198976),
	.w4(32'hb98387a0),
	.w5(32'h3989f688),
	.w6(32'hba835c09),
	.w7(32'hba741c78),
	.w8(32'h3a99c647),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b2a9a),
	.w1(32'hbb270d02),
	.w2(32'h39a9c71b),
	.w3(32'hbc5eaebb),
	.w4(32'h3c0ebf4b),
	.w5(32'h3b348e24),
	.w6(32'hbc42f2d2),
	.w7(32'h3c375993),
	.w8(32'h3bd2174f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b2cb0),
	.w1(32'hba87859c),
	.w2(32'hba9d7349),
	.w3(32'hbae36ee6),
	.w4(32'hb9efa617),
	.w5(32'h39f79bef),
	.w6(32'hb9b329e4),
	.w7(32'hbaafe5ed),
	.w8(32'hba08dba6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc18d86),
	.w1(32'hbb2076ea),
	.w2(32'hbc1554b8),
	.w3(32'hbc937d6f),
	.w4(32'h3b883eba),
	.w5(32'hba9f6c5c),
	.w6(32'hbcb0575d),
	.w7(32'h3a4db0f3),
	.w8(32'hbc10a13b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefcf0e),
	.w1(32'hbb20018b),
	.w2(32'hbad3cc0a),
	.w3(32'hbb40d48d),
	.w4(32'hbb249f94),
	.w5(32'hb9e28c1e),
	.w6(32'hbaab44df),
	.w7(32'hbb3df23c),
	.w8(32'hbb461670),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9356d),
	.w1(32'h3c397dd8),
	.w2(32'hbbd611fc),
	.w3(32'hbc18c357),
	.w4(32'hbb61f782),
	.w5(32'hbc1821e0),
	.w6(32'hbc94ea31),
	.w7(32'hbbf8c78d),
	.w8(32'hbcb443f3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090166),
	.w1(32'hbae621bf),
	.w2(32'hbac1bd74),
	.w3(32'hbb07d835),
	.w4(32'hbad1e16b),
	.w5(32'hb9c79660),
	.w6(32'hbb019107),
	.w7(32'hba93fe5f),
	.w8(32'hb9396292),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca01c6d),
	.w1(32'hbb975bbd),
	.w2(32'hbbf931da),
	.w3(32'hbc7823df),
	.w4(32'h38953acf),
	.w5(32'hbbba4e03),
	.w6(32'hbc473ff2),
	.w7(32'h3b3d8fc8),
	.w8(32'hbb4ea2fd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90252),
	.w1(32'hbadf2457),
	.w2(32'hbaffcffa),
	.w3(32'hbae93882),
	.w4(32'hba03cb5a),
	.w5(32'hb99b1f1e),
	.w6(32'hba8bbbc7),
	.w7(32'hbad95877),
	.w8(32'h3ab484e5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca359ca),
	.w1(32'hb9af8240),
	.w2(32'hbbc5b5a7),
	.w3(32'hbc958944),
	.w4(32'h3ad96bb8),
	.w5(32'hbb75cccc),
	.w6(32'hbcbde420),
	.w7(32'h3b9a2885),
	.w8(32'hbb26fb4f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8d41),
	.w1(32'hbb022ae0),
	.w2(32'h3bd9b4b3),
	.w3(32'hbc5b92eb),
	.w4(32'h3a94f1cb),
	.w5(32'h3c44c9b1),
	.w6(32'hbc28e47b),
	.w7(32'hbbe86baa),
	.w8(32'hbc231ab6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ab888),
	.w1(32'hbb014bb3),
	.w2(32'hbb23c0d3),
	.w3(32'hbb61359c),
	.w4(32'hbb309692),
	.w5(32'hba88ef0f),
	.w6(32'hbb8c0936),
	.w7(32'hbb132d09),
	.w8(32'hbb9e0cfb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87779c),
	.w1(32'h3b82bfc6),
	.w2(32'h3bba6ff4),
	.w3(32'hbba20287),
	.w4(32'hba923ea2),
	.w5(32'hbbe6b235),
	.w6(32'hbb3fe823),
	.w7(32'hb9dd2cf0),
	.w8(32'hb9b5a65f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0f646),
	.w1(32'hbbd3ff01),
	.w2(32'hbc50e18c),
	.w3(32'hbc29c99c),
	.w4(32'h3c202f9d),
	.w5(32'hba8eb481),
	.w6(32'hbc5265ed),
	.w7(32'h3aaaa68d),
	.w8(32'h39024683),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a4be1),
	.w1(32'hbc0f7a2b),
	.w2(32'hbc46ae0f),
	.w3(32'hbd09b6ac),
	.w4(32'hbc06b50a),
	.w5(32'hbc49531a),
	.w6(32'hbd1bdd42),
	.w7(32'hbb5ba644),
	.w8(32'hbc3b185c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcf6d8d),
	.w1(32'hbc1ea2d5),
	.w2(32'hbd1edbce),
	.w3(32'hbdbc0ece),
	.w4(32'hbbcafb69),
	.w5(32'hbd58c9ba),
	.w6(32'hbdc06537),
	.w7(32'h3a93486e),
	.w8(32'hbd37b3e3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd741fdf),
	.w1(32'hbc9d13e0),
	.w2(32'hbc8292c9),
	.w3(32'hbd70da72),
	.w4(32'hbc607492),
	.w5(32'hbcde663f),
	.w6(32'hbd81f194),
	.w7(32'hbc033881),
	.w8(32'hbc99edf2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eba6c),
	.w1(32'hbc9d3fc4),
	.w2(32'hbcc12332),
	.w3(32'h3b9bd8d8),
	.w4(32'hba93d8e5),
	.w5(32'hbc8b3b9a),
	.w6(32'hbae4c14e),
	.w7(32'hbb4769f2),
	.w8(32'hbbbc8940),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ecde7),
	.w1(32'h3aa81ae0),
	.w2(32'h3b6ddf41),
	.w3(32'h3c0b47f0),
	.w4(32'h3bbf2c74),
	.w5(32'h3ba81a77),
	.w6(32'h3bbb5d9a),
	.w7(32'h3acedadf),
	.w8(32'h3a8e6899),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed1e9b),
	.w1(32'h3a9b40fc),
	.w2(32'h3a2f07a5),
	.w3(32'h39c9e48a),
	.w4(32'hb89b19d3),
	.w5(32'h3a21cb5c),
	.w6(32'h39a0bd89),
	.w7(32'h37bbd6dc),
	.w8(32'hbb99d6d1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040cd7),
	.w1(32'h3afe63d7),
	.w2(32'h3b06cda0),
	.w3(32'h39a95d70),
	.w4(32'h3ac7fd3d),
	.w5(32'hb998960e),
	.w6(32'h398d62f6),
	.w7(32'hba99c68b),
	.w8(32'h3b2bccb9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cddcd),
	.w1(32'hba2c2907),
	.w2(32'h3b244c95),
	.w3(32'h3c0881b2),
	.w4(32'h3b80dcc1),
	.w5(32'h3b360b73),
	.w6(32'h3bad4c30),
	.w7(32'h3a7e1b24),
	.w8(32'hba2addbc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90d164),
	.w1(32'hbbccb8db),
	.w2(32'hbc1b7e5b),
	.w3(32'hbc1ea917),
	.w4(32'h3b0a0cd6),
	.w5(32'hbb999e0c),
	.w6(32'hbc0b68ef),
	.w7(32'hb9843599),
	.w8(32'hbc08211f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba34a9),
	.w1(32'hbbcf8c3b),
	.w2(32'hbb8cefb6),
	.w3(32'hbb3f8201),
	.w4(32'hba9d5105),
	.w5(32'hbaf67787),
	.w6(32'hbb88f1e4),
	.w7(32'hbbb12aae),
	.w8(32'hbb91140b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd02bf10),
	.w1(32'h3aaba1cd),
	.w2(32'hbbbce78c),
	.w3(32'hbcdc8248),
	.w4(32'h3afb891c),
	.w5(32'hbc42c2b2),
	.w6(32'hbcfd5b0f),
	.w7(32'hbb7f81e2),
	.w8(32'hbb861f8f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b04b9),
	.w1(32'h3b29efff),
	.w2(32'hbb07510b),
	.w3(32'hbc435b33),
	.w4(32'h3bfe6648),
	.w5(32'h3aa3295d),
	.w6(32'hbc81fe40),
	.w7(32'h3bdc5123),
	.w8(32'hbae1d33d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadc883),
	.w1(32'hb708a392),
	.w2(32'hbbec1e47),
	.w3(32'hbb30bf5a),
	.w4(32'h3b780845),
	.w5(32'hbbcfbd89),
	.w6(32'hba0f9f3e),
	.w7(32'h3b8e8b6a),
	.w8(32'hbc50db9d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2441a),
	.w1(32'hb9b23bac),
	.w2(32'h3b36d8cd),
	.w3(32'hbcb5225d),
	.w4(32'h39c8f9f4),
	.w5(32'hba241796),
	.w6(32'hbcaf97b3),
	.w7(32'hbc249b80),
	.w8(32'hbaf17013),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd25b25e),
	.w1(32'hbc331f15),
	.w2(32'hbc546ada),
	.w3(32'hbcc4813e),
	.w4(32'h3a4fd9b9),
	.w5(32'hbbc6b538),
	.w6(32'hbcdfde00),
	.w7(32'h3b8896d4),
	.w8(32'hbb8387d2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beacf2e),
	.w1(32'hba560959),
	.w2(32'hbb7a3422),
	.w3(32'hba3c25aa),
	.w4(32'hbbd95310),
	.w5(32'hbba27b91),
	.w6(32'h3c2139e3),
	.w7(32'h3b613db1),
	.w8(32'h3adb0821),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36a9a8),
	.w1(32'hba0bbd4e),
	.w2(32'hbaa5e2c5),
	.w3(32'h3b2d1950),
	.w4(32'h39e10e40),
	.w5(32'h3b337253),
	.w6(32'h3b708dfa),
	.w7(32'h3ab94336),
	.w8(32'h39ad5fdd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20b1ff),
	.w1(32'hb97dd25d),
	.w2(32'hba2b9785),
	.w3(32'hb93a8e2e),
	.w4(32'hba0b23fd),
	.w5(32'h39abea3f),
	.w6(32'hb97c9a94),
	.w7(32'hbaaef601),
	.w8(32'hbb0fbb0b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca390),
	.w1(32'hb8e80fab),
	.w2(32'h3afcce95),
	.w3(32'hbaad4655),
	.w4(32'hb8bc9537),
	.w5(32'hbad3d756),
	.w6(32'hba2667b0),
	.w7(32'hbaa65e3a),
	.w8(32'h3a08a823),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7a46),
	.w1(32'hbac44029),
	.w2(32'hbb9773db),
	.w3(32'hbbad0f69),
	.w4(32'h3a559a14),
	.w5(32'hba95d2b7),
	.w6(32'hbb92950e),
	.w7(32'hb90efcde),
	.w8(32'hbad60f57),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73e9ae7),
	.w1(32'h3a4ecb1c),
	.w2(32'hba9f188d),
	.w3(32'hbae0bf7b),
	.w4(32'h3b0e82bb),
	.w5(32'h3aabac53),
	.w6(32'h38612f17),
	.w7(32'h39f85b38),
	.w8(32'hbb8fe323),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0100b3),
	.w1(32'hbc2da833),
	.w2(32'hbc1da45c),
	.w3(32'hbcce5531),
	.w4(32'h3b5c97e1),
	.w5(32'hbbf22c81),
	.w6(32'hbcd441a3),
	.w7(32'hbbcac535),
	.w8(32'h3adb6433),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4a55),
	.w1(32'hba04ee86),
	.w2(32'hbbeb7454),
	.w3(32'hbbd55364),
	.w4(32'h3ba2a823),
	.w5(32'hbb1eb871),
	.w6(32'hbbf09a1d),
	.w7(32'h39e1779f),
	.w8(32'hbbbd8199),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cd578),
	.w1(32'hbb862e5f),
	.w2(32'h3adcb00f),
	.w3(32'hbc6181bb),
	.w4(32'h3b09474a),
	.w5(32'h3aeca12b),
	.w6(32'hbc8b7ae2),
	.w7(32'hba655a18),
	.w8(32'hbb8eb25d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6b355),
	.w1(32'hbb881328),
	.w2(32'hbb083666),
	.w3(32'h3a392e96),
	.w4(32'hbb2c9356),
	.w5(32'hbb1ad76c),
	.w6(32'hbb6acc47),
	.w7(32'hbb9ca699),
	.w8(32'hbb9cd414),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcace439),
	.w1(32'hbb18e7b8),
	.w2(32'hbc22daed),
	.w3(32'hbc89e0ea),
	.w4(32'h3b868e50),
	.w5(32'hbb584ed5),
	.w6(32'hbc8f5973),
	.w7(32'h3a0db97c),
	.w8(32'hbbbb5a79),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093cde),
	.w1(32'hba6c45de),
	.w2(32'hbc0d3790),
	.w3(32'hbbf94c2d),
	.w4(32'h3ad4d98e),
	.w5(32'hbbd092b6),
	.w6(32'hbbf25bea),
	.w7(32'hbb41b471),
	.w8(32'hbc1b8e2c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5cfdc),
	.w1(32'hbb2d8795),
	.w2(32'hbafcbbce),
	.w3(32'hbb578833),
	.w4(32'h39db406b),
	.w5(32'h3a1c2421),
	.w6(32'h39951c37),
	.w7(32'h3ba692bc),
	.w8(32'h3c0d593c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0aeaa8),
	.w1(32'h3a7c462b),
	.w2(32'hbb42da4a),
	.w3(32'hbcff147b),
	.w4(32'h3baf8131),
	.w5(32'h3a9e0c1d),
	.w6(32'hbcee6774),
	.w7(32'h3bb9585e),
	.w8(32'hbb953dc8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d4aaa),
	.w1(32'hbb791e95),
	.w2(32'hbc3c29ee),
	.w3(32'hbd23576e),
	.w4(32'h3b044290),
	.w5(32'hbbdf2e9f),
	.w6(32'hbd318bda),
	.w7(32'h3943c807),
	.w8(32'hbc085cc2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b3624),
	.w1(32'h3a802a16),
	.w2(32'hbc64bfca),
	.w3(32'hbc2bf59b),
	.w4(32'h3c0ef08b),
	.w5(32'hbb8b15a9),
	.w6(32'hbc632ee4),
	.w7(32'h3b2b2a5f),
	.w8(32'hbc1cdcbd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9298b0),
	.w1(32'hb9359e24),
	.w2(32'hb9703e29),
	.w3(32'h3b6f9cc1),
	.w4(32'hba94c0c3),
	.w5(32'hbab4b5c1),
	.w6(32'h3b623ff8),
	.w7(32'hba942024),
	.w8(32'hbabe3d22),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76fe84),
	.w1(32'hbac601f7),
	.w2(32'hba179d3c),
	.w3(32'h3b22f598),
	.w4(32'hbb23e4db),
	.w5(32'hbb1bc830),
	.w6(32'h3a804911),
	.w7(32'hbb34ab93),
	.w8(32'hbb2eaba1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39a2d4),
	.w1(32'hbb4306ea),
	.w2(32'hbb5c4e47),
	.w3(32'hbb30a9fb),
	.w4(32'hba854bd0),
	.w5(32'hbac1838f),
	.w6(32'hbadba0ca),
	.w7(32'hb9ee7a19),
	.w8(32'hb992c57d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf0e23),
	.w1(32'hba6f7fe6),
	.w2(32'hbbd1a77b),
	.w3(32'hbc887040),
	.w4(32'h3b71102b),
	.w5(32'hbaf719ed),
	.w6(32'hbc9eaea9),
	.w7(32'h3b4b0611),
	.w8(32'hbb6aad9f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbee1e7),
	.w1(32'hbac50c9b),
	.w2(32'hbbc29226),
	.w3(32'hbcc5584a),
	.w4(32'hbb04b588),
	.w5(32'hbc059ef7),
	.w6(32'hbcbb76ed),
	.w7(32'hb9fd498c),
	.w8(32'hbb8075ad),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06a333),
	.w1(32'hbb25dda2),
	.w2(32'hba86a284),
	.w3(32'h3a450097),
	.w4(32'hbad9749a),
	.w5(32'hba95dca1),
	.w6(32'hb9b8b311),
	.w7(32'h3954878b),
	.w8(32'hba2a90a3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29a66),
	.w1(32'hba0dbaea),
	.w2(32'h3ab48dba),
	.w3(32'hba69829b),
	.w4(32'hba43dc39),
	.w5(32'h381b95a4),
	.w6(32'hba518b6e),
	.w7(32'hb9f5d3b4),
	.w8(32'h399721bb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e1698),
	.w1(32'hbc3992c3),
	.w2(32'hbbe57da6),
	.w3(32'hbc0098ed),
	.w4(32'hbad91e64),
	.w5(32'hbc2ddb96),
	.w6(32'hbbe57d49),
	.w7(32'h3977cbe8),
	.w8(32'hbbf494a9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6540b0),
	.w1(32'hbc01c1fb),
	.w2(32'hbc3fec0d),
	.w3(32'hbc67095e),
	.w4(32'hbc39b45b),
	.w5(32'hbc4d2f33),
	.w6(32'hbca337a8),
	.w7(32'hbc3cf3e8),
	.w8(32'hbb6cd735),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b370),
	.w1(32'hb9d5d708),
	.w2(32'hbb25c34b),
	.w3(32'hbab10233),
	.w4(32'hbaaa8c6b),
	.w5(32'hbb28ff6a),
	.w6(32'hbb02a8b3),
	.w7(32'hbada7784),
	.w8(32'hbadd4411),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d8515),
	.w1(32'h3b095aa5),
	.w2(32'hbb04b6a4),
	.w3(32'hbc03acbc),
	.w4(32'h3b3dc19a),
	.w5(32'hbafd3434),
	.w6(32'hbbed3cff),
	.w7(32'h3b41e8c7),
	.w8(32'hbb4b2522),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa50c2c),
	.w1(32'h3a96050e),
	.w2(32'h3b250fb5),
	.w3(32'h3b2a7d1e),
	.w4(32'h3bacea82),
	.w5(32'h3b60a201),
	.w6(32'h3b987c0b),
	.w7(32'h3bc3d4c8),
	.w8(32'h3ba58af4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00b62c),
	.w1(32'h3b3e9c3d),
	.w2(32'hbb3d34ff),
	.w3(32'hbb4da848),
	.w4(32'h3b96da42),
	.w5(32'h39c0c032),
	.w6(32'hbaf22829),
	.w7(32'h3bc9f741),
	.w8(32'h3b61bc28),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06b59c),
	.w1(32'h3b8ac6a8),
	.w2(32'h3b0f847c),
	.w3(32'hbc295ed8),
	.w4(32'h3b751168),
	.w5(32'h3a0ceff1),
	.w6(32'hbc25acd9),
	.w7(32'h3b018763),
	.w8(32'h3a886135),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a993cec),
	.w1(32'h3c43c3e5),
	.w2(32'h3c711223),
	.w3(32'h3ab83559),
	.w4(32'h3c10094d),
	.w5(32'h3c650bd5),
	.w6(32'hba08a494),
	.w7(32'h3ba41ac1),
	.w8(32'h3c2a0511),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule