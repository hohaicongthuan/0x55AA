module layer_10_featuremap_51(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e3931),
	.w1(32'h3a8cbbfc),
	.w2(32'h39aa0396),
	.w3(32'hbc0c6abf),
	.w4(32'hbc1c7f16),
	.w5(32'hbc202370),
	.w6(32'hb9a8cd8a),
	.w7(32'h3b3d6f39),
	.w8(32'hbc0723a3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97f562),
	.w1(32'hbaae512a),
	.w2(32'h3c1788dc),
	.w3(32'hba463801),
	.w4(32'h3b1c1b09),
	.w5(32'h39e70ef1),
	.w6(32'hbb67d19d),
	.w7(32'hbb9ff677),
	.w8(32'hbb0a221f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c035c48),
	.w1(32'hba18350e),
	.w2(32'h399a780d),
	.w3(32'h3bed8613),
	.w4(32'h3b34e29b),
	.w5(32'h3a20fc60),
	.w6(32'h3b97b745),
	.w7(32'h3b38c734),
	.w8(32'h3af1f92b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833889),
	.w1(32'hbc0abef6),
	.w2(32'hbc0a3c9a),
	.w3(32'h3b615d02),
	.w4(32'h3c214b15),
	.w5(32'hbc647ab0),
	.w6(32'hbb0e4cf8),
	.w7(32'h3b5a6a29),
	.w8(32'h3bc6eb85),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc965245),
	.w1(32'hbc13a405),
	.w2(32'h3b49bc91),
	.w3(32'hbc800aca),
	.w4(32'hbc5119c3),
	.w5(32'h3be6ba94),
	.w6(32'hbb4344b9),
	.w7(32'hbbd1592b),
	.w8(32'h3c37ad70),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b523d01),
	.w1(32'h3bc10c08),
	.w2(32'h3ae3f1d1),
	.w3(32'h3a5294c1),
	.w4(32'h3b818f05),
	.w5(32'h3ac16524),
	.w6(32'h3af8f332),
	.w7(32'h3b8c3259),
	.w8(32'h3b405194),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6072ca),
	.w1(32'h3b44d17e),
	.w2(32'h3c50d0ff),
	.w3(32'h3b34bd31),
	.w4(32'hbb5c056e),
	.w5(32'h3bc23856),
	.w6(32'h3aa66907),
	.w7(32'hbba3ed6e),
	.w8(32'h3a06567b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5dbfb),
	.w1(32'hbbfc9ec1),
	.w2(32'hbc83c3c9),
	.w3(32'hbb75120a),
	.w4(32'hbb62e831),
	.w5(32'hbc59fbd6),
	.w6(32'hbc122e1b),
	.w7(32'hbc03942a),
	.w8(32'hbc186a9a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe38959),
	.w1(32'hbb8a8eaf),
	.w2(32'h3acc0977),
	.w3(32'hbc20c33d),
	.w4(32'hbba03eb8),
	.w5(32'hbacff15b),
	.w6(32'hbba51ff8),
	.w7(32'h3b76835a),
	.w8(32'hbb15d1c6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8eff),
	.w1(32'h3b650020),
	.w2(32'hbb70dda9),
	.w3(32'hbbeea395),
	.w4(32'h3b16fd61),
	.w5(32'hbbbaab93),
	.w6(32'hbc43982f),
	.w7(32'hba75b2b3),
	.w8(32'hbc1b9e3f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb906fe9),
	.w1(32'hbabaee63),
	.w2(32'hbb55d663),
	.w3(32'hbaf59840),
	.w4(32'hbadf93ef),
	.w5(32'h3a86a8d6),
	.w6(32'hbb164371),
	.w7(32'h3a062944),
	.w8(32'h3b9ec7a0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba533c18),
	.w1(32'h3b1c78a1),
	.w2(32'hba11dfa7),
	.w3(32'h3c36971a),
	.w4(32'h3b96ffc0),
	.w5(32'h3b9d1bea),
	.w6(32'h3bbc7810),
	.w7(32'h3b004c12),
	.w8(32'h38ac9f7c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42e877),
	.w1(32'hbbca4d17),
	.w2(32'h3c08fdf6),
	.w3(32'hbbb5867c),
	.w4(32'hbb3226ee),
	.w5(32'hba7420f1),
	.w6(32'h3907cf0e),
	.w7(32'h39a2f412),
	.w8(32'hbbcf326d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02e23),
	.w1(32'h3b780daf),
	.w2(32'hbc1893b3),
	.w3(32'h3beafbd9),
	.w4(32'h3934cc1c),
	.w5(32'hbc13ae53),
	.w6(32'h3aba9636),
	.w7(32'hbbcff394),
	.w8(32'hbbdc0c89),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5134f0),
	.w1(32'hbc325189),
	.w2(32'h3bf78f85),
	.w3(32'hbb3252b1),
	.w4(32'hbaeb2190),
	.w5(32'h3c4452a9),
	.w6(32'hbbc79f95),
	.w7(32'hbb98faac),
	.w8(32'h3a548bbb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be98f44),
	.w1(32'h3c194c63),
	.w2(32'h3ad273dd),
	.w3(32'h3c5345ac),
	.w4(32'h3c973985),
	.w5(32'h3ad1b200),
	.w6(32'hbba09874),
	.w7(32'h3a2c7404),
	.w8(32'hbaf66669),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392489e7),
	.w1(32'h3aeb4868),
	.w2(32'hbb45e39b),
	.w3(32'h3a2d518c),
	.w4(32'h3a8ff6b8),
	.w5(32'h3abeb9d6),
	.w6(32'h3a841b2b),
	.w7(32'h3b53e9aa),
	.w8(32'h3b1880b9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc833701),
	.w1(32'hbbbe4af2),
	.w2(32'hba81d7c5),
	.w3(32'hbc9a39bb),
	.w4(32'hbc652f4c),
	.w5(32'h3a9db2f5),
	.w6(32'hbc414e8a),
	.w7(32'hbc97c8b4),
	.w8(32'hbab8a917),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadce472),
	.w1(32'h3b9941d6),
	.w2(32'hba8b1ec1),
	.w3(32'hbbc7e0fb),
	.w4(32'hb9f26973),
	.w5(32'hbbdfe6d2),
	.w6(32'h3982386f),
	.w7(32'h3a43caf7),
	.w8(32'hbc316582),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb798abe),
	.w1(32'hbb805de7),
	.w2(32'hbb076cc5),
	.w3(32'hbbb2565d),
	.w4(32'hbc1acff8),
	.w5(32'hba72e4bc),
	.w6(32'hbc9c7bb6),
	.w7(32'hbc5928c8),
	.w8(32'h3b0b275b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c8c8d),
	.w1(32'hba6732bd),
	.w2(32'h3c011a3e),
	.w3(32'hbb38682d),
	.w4(32'hbb818f45),
	.w5(32'hbb49a1bb),
	.w6(32'hb99176cc),
	.w7(32'h39789fa5),
	.w8(32'h3aef3d22),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a346c20),
	.w1(32'h3b168049),
	.w2(32'hbbda03a7),
	.w3(32'hbaead9f4),
	.w4(32'h3b60217d),
	.w5(32'hbb822f09),
	.w6(32'h3b2969b6),
	.w7(32'h3ba3e15a),
	.w8(32'hbad0927b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9eda10),
	.w1(32'hbbf5cd56),
	.w2(32'hbbf6b0e6),
	.w3(32'hbca47d25),
	.w4(32'hbc13aa44),
	.w5(32'hb9af0143),
	.w6(32'hbc9e99c8),
	.w7(32'hbc761546),
	.w8(32'hbc1d977f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1345bc),
	.w1(32'hbb29ee15),
	.w2(32'h3b8b1d54),
	.w3(32'hbb981067),
	.w4(32'h3aede081),
	.w5(32'h39fd5579),
	.w6(32'hbb694287),
	.w7(32'h3b6e1239),
	.w8(32'hbb3e3664),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c078de4),
	.w1(32'h3c325d4e),
	.w2(32'hbb4f5977),
	.w3(32'h3bc4c643),
	.w4(32'h3c5f214b),
	.w5(32'h3be0addc),
	.w6(32'h3bab1bfc),
	.w7(32'h3b8656c1),
	.w8(32'hb9f67b9a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9c841),
	.w1(32'hbb0d729b),
	.w2(32'hb915203b),
	.w3(32'h3c1a0441),
	.w4(32'h3b7c84ea),
	.w5(32'h3a9f615e),
	.w6(32'h3bc86b93),
	.w7(32'h3c066851),
	.w8(32'hbaa7624d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf5082),
	.w1(32'h3bd72b96),
	.w2(32'hbb4b8bd4),
	.w3(32'hbc1273f2),
	.w4(32'hba900cc1),
	.w5(32'hbab8c8ea),
	.w6(32'hbab1921e),
	.w7(32'h3b647b04),
	.w8(32'hbb498eca),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08b0de),
	.w1(32'h3b096881),
	.w2(32'h3bb75582),
	.w3(32'h3a44f44d),
	.w4(32'h3bc481cd),
	.w5(32'h3c2b83cf),
	.w6(32'h3b3973e7),
	.w7(32'h3b1e0b26),
	.w8(32'h3c072e85),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906e6ed),
	.w1(32'hbb2ff341),
	.w2(32'h38f40889),
	.w3(32'h3c27674c),
	.w4(32'h3bf62aba),
	.w5(32'h3988fccc),
	.w6(32'h3bd72b25),
	.w7(32'h3b82864d),
	.w8(32'h3b4575e0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52ba4),
	.w1(32'h3c7252ac),
	.w2(32'hbd6b1d0c),
	.w3(32'h3c6ce487),
	.w4(32'h3c2e2331),
	.w5(32'hbdc11a8f),
	.w6(32'h3a697628),
	.w7(32'h3ae1b5de),
	.w8(32'hbd878dc2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc950080),
	.w1(32'h3d173989),
	.w2(32'h3bc92eb7),
	.w3(32'hbc03e487),
	.w4(32'h3dc82b3b),
	.w5(32'hb9c5c693),
	.w6(32'hbc3feae2),
	.w7(32'h3d6f65a1),
	.w8(32'h3c34bd76),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59356),
	.w1(32'h3be4c6b4),
	.w2(32'h3b6996d4),
	.w3(32'h3b81f33c),
	.w4(32'h3c3ea459),
	.w5(32'h3ba64867),
	.w6(32'h3c1bfa28),
	.w7(32'h3c08b2cb),
	.w8(32'h3c0d4da3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ffe3e),
	.w1(32'h3ba1b82e),
	.w2(32'hbd803c02),
	.w3(32'h3bb39848),
	.w4(32'h3c46b025),
	.w5(32'hbdc8d324),
	.w6(32'h3b39d954),
	.w7(32'h3b92ecac),
	.w8(32'hbd8a50c2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6555d),
	.w1(32'h3d11f58a),
	.w2(32'hbadc2106),
	.w3(32'h397e300a),
	.w4(32'h3de39ecb),
	.w5(32'hbc26896d),
	.w6(32'hbc1260f3),
	.w7(32'h3d6ed86e),
	.w8(32'hbb92de77),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51034e),
	.w1(32'hb9e329b4),
	.w2(32'h3ce477d5),
	.w3(32'hbb9feac3),
	.w4(32'hbb159774),
	.w5(32'h3d3bd10c),
	.w6(32'h3bc7fbc4),
	.w7(32'h3b475103),
	.w8(32'h3cfd4f75),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeb731),
	.w1(32'hbca7bc2b),
	.w2(32'h3c38a9a4),
	.w3(32'hbad2b42d),
	.w4(32'hbd64fcaf),
	.w5(32'h3b82a59f),
	.w6(32'hb9116960),
	.w7(32'hbd262c0f),
	.w8(32'h3a15f4d6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f684),
	.w1(32'hbc077ede),
	.w2(32'hbd16c027),
	.w3(32'h3b155a96),
	.w4(32'hbbbf514b),
	.w5(32'hbd6a4910),
	.w6(32'hbc11664c),
	.w7(32'hbc0a33c0),
	.w8(32'hbd27d2d8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4a3c0),
	.w1(32'h3ce39fba),
	.w2(32'hb9b6da41),
	.w3(32'h3b1fab3d),
	.w4(32'h3dc31fca),
	.w5(32'h3c3a9281),
	.w6(32'hbc936b5c),
	.w7(32'h3d28ef46),
	.w8(32'h3c13d7ff),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3dd8b),
	.w1(32'h3c8ef759),
	.w2(32'h3b9ecb7a),
	.w3(32'h3d05ae7e),
	.w4(32'h3c6f50de),
	.w5(32'h3b48a4f6),
	.w6(32'h3c9e00d0),
	.w7(32'h3c1f8b7b),
	.w8(32'hbbd7c734),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3274e3),
	.w1(32'h3bbeef5b),
	.w2(32'h3a8e2556),
	.w3(32'hbc80bd7e),
	.w4(32'h3bd89a84),
	.w5(32'hbb9b4dce),
	.w6(32'hbc438af7),
	.w7(32'hbbd7699b),
	.w8(32'hbc430ff8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b7393),
	.w1(32'h3c418051),
	.w2(32'h3b3eea2e),
	.w3(32'h3b0e5ba2),
	.w4(32'h3c558a51),
	.w5(32'h3c01bf82),
	.w6(32'hba1c79fb),
	.w7(32'h3c01139c),
	.w8(32'h3b74b58e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ee465),
	.w1(32'h3bc2aaf8),
	.w2(32'h3a5a5c12),
	.w3(32'h3c37e4d0),
	.w4(32'h3ba809a2),
	.w5(32'hbb63b353),
	.w6(32'h3b89b223),
	.w7(32'h3bcef7bf),
	.w8(32'h3bcc3e1b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0a8ba),
	.w1(32'h3c61746a),
	.w2(32'h3d683edc),
	.w3(32'h3bdd7663),
	.w4(32'h3ba1d2b8),
	.w5(32'h3db3cb44),
	.w6(32'h3c1c9fab),
	.w7(32'h3ad3e8b8),
	.w8(32'h3d6aba69),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc8978),
	.w1(32'hbd3c7584),
	.w2(32'h3aaa4dc1),
	.w3(32'hbcb91921),
	.w4(32'hbdd75e4e),
	.w5(32'hbc5cfd91),
	.w6(32'hbc17ef19),
	.w7(32'hbd7b1b49),
	.w8(32'hbaf9890f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc184933),
	.w1(32'hbb29729a),
	.w2(32'hbb91a6d6),
	.w3(32'hbc0d06f4),
	.w4(32'h3c2b8771),
	.w5(32'hbc52a33c),
	.w6(32'hba2437db),
	.w7(32'h3bb77703),
	.w8(32'hbc2da04c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3caf4),
	.w1(32'hbb5b2341),
	.w2(32'h3aa51587),
	.w3(32'hbbd14ab5),
	.w4(32'h3c073300),
	.w5(32'hbb4df167),
	.w6(32'hbbfa0159),
	.w7(32'hbaaeee44),
	.w8(32'hbb0598ba),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473f62),
	.w1(32'h3aa4317f),
	.w2(32'hbc12f73a),
	.w3(32'hbc377248),
	.w4(32'hbb4c0a30),
	.w5(32'hbc49e672),
	.w6(32'hbb573bbd),
	.w7(32'h3abe6a77),
	.w8(32'hbbd2a54c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c8002),
	.w1(32'h3acdae4c),
	.w2(32'h3d63d25a),
	.w3(32'hbced6976),
	.w4(32'hbb606346),
	.w5(32'h3dc514e1),
	.w6(32'hbca047dc),
	.w7(32'hb95106f1),
	.w8(32'h3d650331),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baacb17),
	.w1(32'hbd667608),
	.w2(32'h3c24cb2a),
	.w3(32'hbbf13ba8),
	.w4(32'hbdfbee7a),
	.w5(32'h3b8430d0),
	.w6(32'hbb40bdcb),
	.w7(32'hbda20d68),
	.w8(32'h3b436318),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70a016),
	.w1(32'h3c1c1ba9),
	.w2(32'h3b50c815),
	.w3(32'h3c7adc57),
	.w4(32'hbae714aa),
	.w5(32'h3bdb3b39),
	.w6(32'hbb29590b),
	.w7(32'hbb139b85),
	.w8(32'h3c1da211),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ab592),
	.w1(32'hbbd7f2c6),
	.w2(32'hbc1329a6),
	.w3(32'h3b64e652),
	.w4(32'h3badcb8a),
	.w5(32'hbaf47c86),
	.w6(32'h3c21807b),
	.w7(32'h3c01817e),
	.w8(32'h3b6070c2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1e884),
	.w1(32'hbca449de),
	.w2(32'h3bc6ae2b),
	.w3(32'hbcdf4fb7),
	.w4(32'hbc5564c4),
	.w5(32'h3c6f0c81),
	.w6(32'hbc261fd9),
	.w7(32'hba4e6e98),
	.w8(32'h3c3f6105),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b855ed4),
	.w1(32'h3b0eb3fc),
	.w2(32'hbb6d05c4),
	.w3(32'h3c4bad0f),
	.w4(32'h3bfc9439),
	.w5(32'hbb006ec2),
	.w6(32'h3c54066f),
	.w7(32'h3acd90dd),
	.w8(32'hbb121b9c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133041),
	.w1(32'hbb5dc01b),
	.w2(32'h3be85ec6),
	.w3(32'hbc36e5ef),
	.w4(32'hba124a98),
	.w5(32'h3b5ffdd4),
	.w6(32'hbc51a84e),
	.w7(32'hba086f17),
	.w8(32'hbc3f05fc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c03be),
	.w1(32'h3c09670f),
	.w2(32'h3c10b98f),
	.w3(32'h3a902c7e),
	.w4(32'hbb2167eb),
	.w5(32'hba9aa581),
	.w6(32'hbc0728c2),
	.w7(32'hbc3588ef),
	.w8(32'hbb112368),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b419391),
	.w1(32'h3b427964),
	.w2(32'h3a443077),
	.w3(32'h3a2ffe7a),
	.w4(32'h3b37dc5d),
	.w5(32'hbb98c390),
	.w6(32'hba8e668e),
	.w7(32'hb9ceb2fb),
	.w8(32'h3b2c7cc6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa4a2c),
	.w1(32'h3b1a4f6f),
	.w2(32'h3bb0360e),
	.w3(32'h395242bb),
	.w4(32'h3aafa3fc),
	.w5(32'h3bb17396),
	.w6(32'hba9aefeb),
	.w7(32'hbb379e7b),
	.w8(32'h3b480f42),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c2cf),
	.w1(32'hbb7fea53),
	.w2(32'hbacdf9b1),
	.w3(32'hbb846805),
	.w4(32'hbbb85d7c),
	.w5(32'hbaeabde8),
	.w6(32'hbb8f0dee),
	.w7(32'hbbdee728),
	.w8(32'hbc061749),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68a54),
	.w1(32'h3c7cd0ec),
	.w2(32'h3c4cb2e2),
	.w3(32'hbbc4478e),
	.w4(32'h3c8e57f8),
	.w5(32'h3be8db6a),
	.w6(32'hbc5772af),
	.w7(32'h3b0e2165),
	.w8(32'h3a6c4f15),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2442ae),
	.w1(32'h3c2f14e3),
	.w2(32'h3c881202),
	.w3(32'h3b3c2c66),
	.w4(32'h3c1559da),
	.w5(32'h3ca7e47e),
	.w6(32'hbb1ca5f5),
	.w7(32'h3b01c90c),
	.w8(32'h3c39b97c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbe424),
	.w1(32'hbb298146),
	.w2(32'hbc4823cf),
	.w3(32'h3a92055f),
	.w4(32'hbc0283b5),
	.w5(32'hbc59630b),
	.w6(32'hbbce4140),
	.w7(32'hbc72e342),
	.w8(32'hbbbf909c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc392e2e),
	.w1(32'h39e13655),
	.w2(32'hbb98d9fd),
	.w3(32'hbcae30bf),
	.w4(32'hbbaca460),
	.w5(32'hbb83e1e4),
	.w6(32'hbbe95b8a),
	.w7(32'h3affe29f),
	.w8(32'hb99490d7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc331db9),
	.w1(32'hbbb5629b),
	.w2(32'h39cf205c),
	.w3(32'h3baf34d2),
	.w4(32'hbb43849e),
	.w5(32'h3aee3e64),
	.w6(32'h3bc0e94d),
	.w7(32'h3bbc0232),
	.w8(32'h3a51e3cb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8552),
	.w1(32'h3c57685c),
	.w2(32'h3a8bbd21),
	.w3(32'h3a5e9f42),
	.w4(32'h3c322271),
	.w5(32'h3b884311),
	.w6(32'h3bcb2cb1),
	.w7(32'h3c7a8526),
	.w8(32'hbb986879),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd6a9),
	.w1(32'hbbe91023),
	.w2(32'h3b142c07),
	.w3(32'h3b346d52),
	.w4(32'hbab59162),
	.w5(32'h3be2fd41),
	.w6(32'hbc02c8dd),
	.w7(32'h3b91b514),
	.w8(32'h3bddbb91),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f769e),
	.w1(32'h3ac46212),
	.w2(32'h3a92208e),
	.w3(32'h3c084cb2),
	.w4(32'h3bd25fb4),
	.w5(32'h3b210962),
	.w6(32'h3c025b3f),
	.w7(32'h3c1f9a5e),
	.w8(32'h3ba49c93),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2836),
	.w1(32'h3ac8ed6c),
	.w2(32'h3bcf8582),
	.w3(32'h3aab26e7),
	.w4(32'h3cb45b9b),
	.w5(32'h3bd21651),
	.w6(32'hbad63b8c),
	.w7(32'h3b0397ad),
	.w8(32'hbb422920),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a969879),
	.w1(32'h3c139f77),
	.w2(32'h38ade723),
	.w3(32'h3bc7be68),
	.w4(32'hba7e550c),
	.w5(32'h3ae39f5e),
	.w6(32'hbb855b62),
	.w7(32'hbb068838),
	.w8(32'h3bbc5192),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9ae5e),
	.w1(32'h3b171e07),
	.w2(32'hbb0485fe),
	.w3(32'hbb82ccec),
	.w4(32'h3ba3e0f9),
	.w5(32'hbaf6b4b8),
	.w6(32'hbb8d6c62),
	.w7(32'hbb8a3754),
	.w8(32'hbb4127b5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb608ec),
	.w1(32'h3c59cc18),
	.w2(32'hbadc4ad3),
	.w3(32'h3c28a514),
	.w4(32'h3c927f9e),
	.w5(32'hbb91a64e),
	.w6(32'h3c32a45b),
	.w7(32'h3c45883d),
	.w8(32'hbb8747f4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc100222),
	.w1(32'h3c29aecb),
	.w2(32'hbb3272de),
	.w3(32'hbc3a3dd3),
	.w4(32'h3c381e30),
	.w5(32'h3ac82088),
	.w6(32'hbb9aba37),
	.w7(32'h3c344548),
	.w8(32'hb9f65b27),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c58df4),
	.w1(32'h3bbd3101),
	.w2(32'h3b0de3b4),
	.w3(32'hbb4dfe76),
	.w4(32'h3c332410),
	.w5(32'h3b206894),
	.w6(32'hbb52cf6b),
	.w7(32'h3ba47c3d),
	.w8(32'hbc1e43dd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab21fdc),
	.w1(32'h3aaecac1),
	.w2(32'hba827410),
	.w3(32'hb9b454eb),
	.w4(32'h3b99b5bb),
	.w5(32'hbb455fbd),
	.w6(32'h3a55d6cd),
	.w7(32'h3c02a72f),
	.w8(32'hb9ea5b9f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab30e),
	.w1(32'hbbe1dde2),
	.w2(32'h3d22fd88),
	.w3(32'hbcb47bcc),
	.w4(32'hbb99e885),
	.w5(32'h3d8a9cef),
	.w6(32'hbc4a1b74),
	.w7(32'h3a139577),
	.w8(32'h3d319005),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19aac4),
	.w1(32'hbcedafb2),
	.w2(32'h395e1d56),
	.w3(32'hbab584a2),
	.w4(32'hbd9cac83),
	.w5(32'hbbecb624),
	.w6(32'h3b3f274f),
	.w7(32'hbd43581f),
	.w8(32'hbbcc3a0f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b50c),
	.w1(32'h3ab780af),
	.w2(32'hbb965383),
	.w3(32'h3b18b14a),
	.w4(32'h3be9618f),
	.w5(32'hbbfe0086),
	.w6(32'hbc248c17),
	.w7(32'h3b5d3a5c),
	.w8(32'hbc19185d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fa31a),
	.w1(32'hbc7b98b9),
	.w2(32'hbc34be47),
	.w3(32'hbca8a031),
	.w4(32'hbcab5a1a),
	.w5(32'hbc60f812),
	.w6(32'hbcbaf5b0),
	.w7(32'hbc0dd160),
	.w8(32'hbba26814),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc541c9c),
	.w1(32'h3aa58ddd),
	.w2(32'hbbc30a26),
	.w3(32'hbbf95be1),
	.w4(32'h3b0621f2),
	.w5(32'hbb03051e),
	.w6(32'h3b9d6ae0),
	.w7(32'h3c49fc53),
	.w8(32'hbb75ced5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c1551),
	.w1(32'h3ba67a9b),
	.w2(32'hbbe30fa6),
	.w3(32'hbbb3b0bd),
	.w4(32'hbb050f6e),
	.w5(32'hbbdce05e),
	.w6(32'hbbf2f67f),
	.w7(32'hbb91196b),
	.w8(32'hbba12767),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af74775),
	.w1(32'hb9c0118e),
	.w2(32'h3c7a2272),
	.w3(32'hbae14ca6),
	.w4(32'h3b0291d9),
	.w5(32'h3c4ce9aa),
	.w6(32'h3bb62be6),
	.w7(32'hba67da90),
	.w8(32'h3b9913bf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf14121),
	.w1(32'hba4e3eb8),
	.w2(32'hbcf6d441),
	.w3(32'hbc5a085d),
	.w4(32'hb9ef0074),
	.w5(32'hbd329039),
	.w6(32'hbb5e2611),
	.w7(32'h3c16e3f4),
	.w8(32'hbceab718),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b8f6b),
	.w1(32'h3c9be395),
	.w2(32'hbc5bc38b),
	.w3(32'hbbf9cea2),
	.w4(32'h3d7aa1f5),
	.w5(32'hbb9f5587),
	.w6(32'hbc2127e7),
	.w7(32'h3d01ce23),
	.w8(32'hbc63a959),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09a079),
	.w1(32'hba867854),
	.w2(32'hbc360505),
	.w3(32'h3c151a1a),
	.w4(32'h3a00f1d5),
	.w5(32'hbc23fdf9),
	.w6(32'hbbf9d587),
	.w7(32'h3b2a4eb3),
	.w8(32'hbb970677),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49bd40),
	.w1(32'hbb1ca1b3),
	.w2(32'h3bac6089),
	.w3(32'hbc95939d),
	.w4(32'hbc1d08b0),
	.w5(32'h3c23bdfc),
	.w6(32'hbc3e4998),
	.w7(32'h39430671),
	.w8(32'hb8bfca22),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5b7b),
	.w1(32'h3a2dcbc3),
	.w2(32'hbc25c415),
	.w3(32'h3c06975f),
	.w4(32'h3ba6c808),
	.w5(32'hbc0ca193),
	.w6(32'h3bfb2685),
	.w7(32'h3c28760f),
	.w8(32'h3b96b4cd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97db3f),
	.w1(32'h3b128bd5),
	.w2(32'hbaaa3820),
	.w3(32'h3bce621f),
	.w4(32'h3bea96cb),
	.w5(32'h3b0a9a68),
	.w6(32'h3c160086),
	.w7(32'h3bf794e4),
	.w8(32'hba1a0988),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9831d0),
	.w1(32'hbb6c0f2d),
	.w2(32'hbb71c254),
	.w3(32'hbc504e5a),
	.w4(32'h3b90357b),
	.w5(32'hbb1f9682),
	.w6(32'hbc610e45),
	.w7(32'hb95697a4),
	.w8(32'hbb853100),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5a7f7),
	.w1(32'h3b7d0eaa),
	.w2(32'h3ba24703),
	.w3(32'h39d5ca1b),
	.w4(32'hba49a296),
	.w5(32'h3aecd3e3),
	.w6(32'h3a580d40),
	.w7(32'hbb07bdee),
	.w8(32'h3bf513ba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd0f9),
	.w1(32'hbc494436),
	.w2(32'h3c4d6978),
	.w3(32'hbbacd6a2),
	.w4(32'hba04a9f4),
	.w5(32'h3bc06780),
	.w6(32'h3bf12380),
	.w7(32'h3bda7e3e),
	.w8(32'h3c0331ae),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ea690),
	.w1(32'hbc37c4ba),
	.w2(32'h3adf2d4c),
	.w3(32'hbc07211c),
	.w4(32'hbb9758ee),
	.w5(32'h3c6b9c77),
	.w6(32'hbc7ecd31),
	.w7(32'hbc37ab33),
	.w8(32'hb9aa6d90),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb5035),
	.w1(32'h3a1f115f),
	.w2(32'h3c9446e0),
	.w3(32'h3c6d2390),
	.w4(32'h3b39affd),
	.w5(32'h3d2f63d4),
	.w6(32'h3b091d50),
	.w7(32'h3acc5300),
	.w8(32'h3cc7e323),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a296f1),
	.w1(32'hb88acc04),
	.w2(32'h3b6c09bb),
	.w3(32'h3c841c11),
	.w4(32'h3bfbc4c7),
	.w5(32'hbb0afccf),
	.w6(32'h3b8b36ce),
	.w7(32'hbb9a0b3c),
	.w8(32'hbb9cb503),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7db9e),
	.w1(32'h3c0a9b57),
	.w2(32'h3c488e7e),
	.w3(32'hba098e2d),
	.w4(32'h3bcc8921),
	.w5(32'h3c95b91c),
	.w6(32'h3b683668),
	.w7(32'h3b33e149),
	.w8(32'h3bdb824c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc37ba8),
	.w1(32'hbc6c17f4),
	.w2(32'hbbe612a5),
	.w3(32'hbc477734),
	.w4(32'hbccef6fa),
	.w5(32'hb9cead9c),
	.w6(32'hbb909bf1),
	.w7(32'hbc91aa71),
	.w8(32'hbbf175c6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064d78),
	.w1(32'h3a2a27b0),
	.w2(32'h3af376e3),
	.w3(32'h3c0e0bbb),
	.w4(32'h3c2e92cb),
	.w5(32'h3b77f497),
	.w6(32'h3a4a5384),
	.w7(32'h3b2c0e33),
	.w8(32'hbad29baf),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b726834),
	.w1(32'hbc0c86ac),
	.w2(32'h3c0cd4ee),
	.w3(32'h3c694b08),
	.w4(32'h3bb3aa20),
	.w5(32'hbb62e7f7),
	.w6(32'h3accc6ab),
	.w7(32'hbc520f99),
	.w8(32'hb98959fd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7df2a5),
	.w1(32'h3bbe1bfd),
	.w2(32'h3a90302f),
	.w3(32'h3aa94d02),
	.w4(32'hbbd10666),
	.w5(32'h3c5367b5),
	.w6(32'hbc030065),
	.w7(32'hbb435551),
	.w8(32'h3c17b210),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c8684),
	.w1(32'h3b158f63),
	.w2(32'hbba7b887),
	.w3(32'hbbfb07ee),
	.w4(32'h3b270bff),
	.w5(32'hbc2ed8c2),
	.w6(32'hba9864fa),
	.w7(32'hbadb5286),
	.w8(32'h3b7b824e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ed992),
	.w1(32'hbbe1b1b0),
	.w2(32'h3c970928),
	.w3(32'hbc7f4735),
	.w4(32'h3ba5fcc9),
	.w5(32'h3cca97c6),
	.w6(32'h39fee518),
	.w7(32'h3b9e6d84),
	.w8(32'h3c409ce7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20595c),
	.w1(32'hbc1c4f7a),
	.w2(32'hbc2a0cbd),
	.w3(32'hbc5a5100),
	.w4(32'hbc25ad4f),
	.w5(32'hbba6b256),
	.w6(32'hbcbe6722),
	.w7(32'hbc869f87),
	.w8(32'hbb30091f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891fa2),
	.w1(32'h3bfe5b7d),
	.w2(32'hbc026d55),
	.w3(32'h3c08fca9),
	.w4(32'h3c0c2aca),
	.w5(32'hbc123a5c),
	.w6(32'hbbce7f7b),
	.w7(32'h3b2abe3e),
	.w8(32'hbb7c5f2e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b434ae0),
	.w1(32'h3b91c77a),
	.w2(32'hbbd6073d),
	.w3(32'hb875132d),
	.w4(32'h3c0bf1f7),
	.w5(32'hbba52e71),
	.w6(32'h3b805b3d),
	.w7(32'h3c0b0d4b),
	.w8(32'h38e320ce),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc794fae),
	.w1(32'h3b55930d),
	.w2(32'h3b08d851),
	.w3(32'hbc2bf5c6),
	.w4(32'h3b7cb9c5),
	.w5(32'h3a7fbf64),
	.w6(32'hbca4d44b),
	.w7(32'hbbea0498),
	.w8(32'hbbe42936),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a243),
	.w1(32'h3b1624f2),
	.w2(32'hbc279d38),
	.w3(32'hbc791046),
	.w4(32'hbaa1680d),
	.w5(32'hbbbb28e9),
	.w6(32'h3acb4c56),
	.w7(32'h3c1ab554),
	.w8(32'hbb76e676),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7ebf8),
	.w1(32'hbcff03b1),
	.w2(32'hbd20ab3d),
	.w3(32'hbd073055),
	.w4(32'hbc99df87),
	.w5(32'hbc785e45),
	.w6(32'hbcc5074b),
	.w7(32'hbc48779e),
	.w8(32'hbc6342ce),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf547),
	.w1(32'hbbd3144d),
	.w2(32'hbc196731),
	.w3(32'hbbdc49a7),
	.w4(32'h3bccd632),
	.w5(32'hbc7ec88d),
	.w6(32'h3c1ec71e),
	.w7(32'h3bec691b),
	.w8(32'hbc290e7e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17232),
	.w1(32'h3ad46002),
	.w2(32'hbaef0da8),
	.w3(32'hbc4df095),
	.w4(32'h3c17d0e2),
	.w5(32'h3bd007eb),
	.w6(32'h38bcf2ca),
	.w7(32'h3c4257cb),
	.w8(32'h3c5fc17c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0c58),
	.w1(32'h3bc911dd),
	.w2(32'hbb8da89d),
	.w3(32'h3aa108ad),
	.w4(32'h3c1500b0),
	.w5(32'hb9ac971b),
	.w6(32'h3a1b2ee5),
	.w7(32'hba8c340b),
	.w8(32'h3af57638),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9b9cb),
	.w1(32'h3c10db4f),
	.w2(32'h3c108fb1),
	.w3(32'hbbebee7a),
	.w4(32'hbb898f19),
	.w5(32'h3bd8660c),
	.w6(32'hbba76684),
	.w7(32'h3b398be7),
	.w8(32'h3b28ad88),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e4038),
	.w1(32'h3c92acdf),
	.w2(32'hbc08d24f),
	.w3(32'h3c39cce3),
	.w4(32'h3c112bf6),
	.w5(32'h3bb286b4),
	.w6(32'h3bf456a6),
	.w7(32'h3b9ced10),
	.w8(32'h3c46a0c5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba62ed6),
	.w1(32'hbb4df9d5),
	.w2(32'hbbf1e65f),
	.w3(32'hbb8daeeb),
	.w4(32'hbb8dac18),
	.w5(32'hbc077d68),
	.w6(32'hbb37754e),
	.w7(32'h3adda0bd),
	.w8(32'h3b19b0d0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ea37),
	.w1(32'h3b70bf10),
	.w2(32'h3b46e925),
	.w3(32'hbc13de5d),
	.w4(32'h3a4bfbab),
	.w5(32'hbb6b2702),
	.w6(32'hba9def7c),
	.w7(32'h3b73e0e2),
	.w8(32'hbc0013e5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58b96c),
	.w1(32'hbb27f33d),
	.w2(32'hbb75df30),
	.w3(32'hbcaf0630),
	.w4(32'hbc39e3eb),
	.w5(32'hbbe10982),
	.w6(32'hbc5d270a),
	.w7(32'hba677dc6),
	.w8(32'h3c2cc54f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38ddc1),
	.w1(32'h3bf1cd4d),
	.w2(32'hbb375a4f),
	.w3(32'hbc3962ad),
	.w4(32'h3976e203),
	.w5(32'h3b0c9561),
	.w6(32'hbc2a7ff2),
	.w7(32'hbb1e03e7),
	.w8(32'h3c0cc758),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf989f8),
	.w1(32'hba297f65),
	.w2(32'h3b06ffc2),
	.w3(32'h3b9143f6),
	.w4(32'hb8548673),
	.w5(32'h3b5fb295),
	.w6(32'h3c2df893),
	.w7(32'h3c3292a8),
	.w8(32'h3b9c72aa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e64b4),
	.w1(32'h3b5fab9c),
	.w2(32'hbb8b0112),
	.w3(32'hbb13d92f),
	.w4(32'h3b971015),
	.w5(32'h3bf26008),
	.w6(32'hba5a8dd8),
	.w7(32'hbb2f3edf),
	.w8(32'h3c2a41af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc601e80),
	.w1(32'hbc0efdcd),
	.w2(32'h3b32231a),
	.w3(32'hbb278417),
	.w4(32'h3a3f8ff2),
	.w5(32'h3b983bf1),
	.w6(32'h3b165860),
	.w7(32'h3b7bfe61),
	.w8(32'hbaefeaef),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38220d),
	.w1(32'h3b9402ad),
	.w2(32'h3b7828f1),
	.w3(32'h3b19de4c),
	.w4(32'h3b82c88f),
	.w5(32'h3b64b33d),
	.w6(32'hbbc71a5a),
	.w7(32'hbbda9174),
	.w8(32'h3c449040),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb146a5b),
	.w1(32'h3a8f3e79),
	.w2(32'h3b08da71),
	.w3(32'h3ab98d52),
	.w4(32'h3c1d25ac),
	.w5(32'h3ab9fe79),
	.w6(32'h3b96c9d5),
	.w7(32'h3b94fd93),
	.w8(32'hbb0a0200),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b354401),
	.w1(32'hba2f394d),
	.w2(32'hbb8a1d21),
	.w3(32'hbacb8cc1),
	.w4(32'h3ba5c11a),
	.w5(32'hbbe0f2f0),
	.w6(32'h3b0af76c),
	.w7(32'h3bab5131),
	.w8(32'h39998e4b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb858da4),
	.w1(32'hbb8b231b),
	.w2(32'hbc16376d),
	.w3(32'hbb62d7ed),
	.w4(32'h38e0fc38),
	.w5(32'hbc9779f2),
	.w6(32'h3b1b3566),
	.w7(32'h3ac84aee),
	.w8(32'hbc2f5c05),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2f8d0),
	.w1(32'h3c26012c),
	.w2(32'hbcc21a49),
	.w3(32'hbb3d8a89),
	.w4(32'h3c879174),
	.w5(32'hbd2639a5),
	.w6(32'hbb942158),
	.w7(32'h3c1e281b),
	.w8(32'hbce4e4e2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c1e0a),
	.w1(32'h3cd64149),
	.w2(32'hbc0d3338),
	.w3(32'h3bdbbf83),
	.w4(32'h3d66a033),
	.w5(32'hbc825890),
	.w6(32'hb9444848),
	.w7(32'h3cf565a7),
	.w8(32'hbcbad5c0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc775eaf),
	.w1(32'hbb184a7d),
	.w2(32'h3ab05621),
	.w3(32'hbd046c5d),
	.w4(32'h3ae57011),
	.w5(32'h3b3ec37f),
	.w6(32'hbc2e0042),
	.w7(32'h3c27abbc),
	.w8(32'h3b99543b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6fd4),
	.w1(32'h3bed7b2c),
	.w2(32'hbc382551),
	.w3(32'h3c02cf64),
	.w4(32'h3c1d8b7d),
	.w5(32'hbc9691aa),
	.w6(32'h3bafbf84),
	.w7(32'h3bb6a2ab),
	.w8(32'hbb4d566c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc899c78),
	.w1(32'hbc1fb0c3),
	.w2(32'hbafe98c7),
	.w3(32'hbcabeff8),
	.w4(32'hbc006dff),
	.w5(32'hbafb5476),
	.w6(32'hbc55f9da),
	.w7(32'h39f16bbf),
	.w8(32'hba19083e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4df38),
	.w1(32'hbae822d5),
	.w2(32'h3ba0ab1b),
	.w3(32'hbc5df9aa),
	.w4(32'hbb5ea9e0),
	.w5(32'h3bd40ac7),
	.w6(32'hbc0f84df),
	.w7(32'hba45b1a4),
	.w8(32'hbb7007f7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacced32),
	.w1(32'hbb593562),
	.w2(32'hb9333862),
	.w3(32'h3b13167f),
	.w4(32'hbbb27fb0),
	.w5(32'hbc2bc38a),
	.w6(32'hbb9b5626),
	.w7(32'h3a013ea1),
	.w8(32'h3c87b3fe),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1ae60),
	.w1(32'h3b42901e),
	.w2(32'hbb86064c),
	.w3(32'hbb814926),
	.w4(32'h3c2bfddb),
	.w5(32'hbbcd7a6d),
	.w6(32'h3b8ad8f1),
	.w7(32'h3c2c8a55),
	.w8(32'hbaa47bcb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35c0f),
	.w1(32'h3b713856),
	.w2(32'hba31ac5d),
	.w3(32'hbb6b5635),
	.w4(32'hbb5f3fbf),
	.w5(32'h3b99a077),
	.w6(32'hbbf02880),
	.w7(32'hbc1597f3),
	.w8(32'hba0c8638),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba771ec4),
	.w1(32'hb7d0d040),
	.w2(32'hbbf05086),
	.w3(32'hba49e3bb),
	.w4(32'h3aa4396f),
	.w5(32'hb83ddaa9),
	.w6(32'h39220249),
	.w7(32'hba13e277),
	.w8(32'h399da427),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ad4cf),
	.w1(32'h3a9f33e4),
	.w2(32'hbbd1f46e),
	.w3(32'hbba0049f),
	.w4(32'h3b84a245),
	.w5(32'h3b990268),
	.w6(32'hba5a6b00),
	.w7(32'hb7fec551),
	.w8(32'h3b611f12),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d9034),
	.w1(32'hbb9d6ef7),
	.w2(32'hbc360a15),
	.w3(32'hb9148cb2),
	.w4(32'h3b5a7272),
	.w5(32'hbc992d68),
	.w6(32'h3bf205dc),
	.w7(32'hba387c57),
	.w8(32'hbcb881dc),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84cb1d),
	.w1(32'hbb18c4cb),
	.w2(32'h3d07d31a),
	.w3(32'hbcb5847d),
	.w4(32'hb98f4f6c),
	.w5(32'h3d8774e9),
	.w6(32'hbcc0d4a4),
	.w7(32'hbc1d2fda),
	.w8(32'h3d18f170),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37e92b),
	.w1(32'hbd2405cc),
	.w2(32'hbb7499fd),
	.w3(32'hbcb3877c),
	.w4(32'hbdab19c3),
	.w5(32'h3b050a21),
	.w6(32'hbc7b8a60),
	.w7(32'hbd652fb8),
	.w8(32'hbb24654a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1398e4),
	.w1(32'h3b1728e0),
	.w2(32'hbb2d63e1),
	.w3(32'h3bad3f07),
	.w4(32'h3c16b674),
	.w5(32'h3b19b09d),
	.w6(32'h3bde4c1f),
	.w7(32'h3b76a953),
	.w8(32'hbb854c74),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde0942),
	.w1(32'h3b3951c1),
	.w2(32'h3afdd1be),
	.w3(32'hbbe22679),
	.w4(32'h3c043d38),
	.w5(32'h3bdf9d6b),
	.w6(32'hbbbbbad6),
	.w7(32'h3aa452b3),
	.w8(32'hba8c138f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9473),
	.w1(32'hbbf2c7c3),
	.w2(32'hbd14633a),
	.w3(32'h3b36bf8f),
	.w4(32'hbadad7af),
	.w5(32'hbd41da5c),
	.w6(32'hbbf5d154),
	.w7(32'hbc67c4a7),
	.w8(32'hbd141122),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe62f2b),
	.w1(32'h3cdaf1a2),
	.w2(32'h3a22972e),
	.w3(32'h3a8ebeec),
	.w4(32'h3d80f2d6),
	.w5(32'hbbd633ab),
	.w6(32'hbb94303b),
	.w7(32'h3d17c468),
	.w8(32'hbb4d43ea),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ade8),
	.w1(32'hbb807322),
	.w2(32'h3c6453a5),
	.w3(32'hbb385bfe),
	.w4(32'h3bff7f6e),
	.w5(32'h3cbff52a),
	.w6(32'h3b7457fb),
	.w7(32'hb9c8133a),
	.w8(32'h3c2b96af),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3df7a3),
	.w1(32'hbc6ac26c),
	.w2(32'hba885721),
	.w3(32'hbbc0c91e),
	.w4(32'hbcf41a46),
	.w5(32'hbb592d14),
	.w6(32'hbbeeb68b),
	.w7(32'hbcb9e373),
	.w8(32'hbb68898a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f82c3),
	.w1(32'hbabdbcc2),
	.w2(32'h3bcf7da5),
	.w3(32'hbc2a41e5),
	.w4(32'hbbad48bf),
	.w5(32'hbc2792ec),
	.w6(32'hbc1c21dc),
	.w7(32'hbba457c8),
	.w8(32'hbaf00903),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17f05d),
	.w1(32'hbb8f088e),
	.w2(32'h3b5877e1),
	.w3(32'hbc9c663e),
	.w4(32'hbb884213),
	.w5(32'h3b8d10f9),
	.w6(32'hbc247946),
	.w7(32'h3aac1101),
	.w8(32'hba2f8596),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e09f),
	.w1(32'h3baea2d9),
	.w2(32'hbcb5b7e1),
	.w3(32'hbab1184d),
	.w4(32'hba8baef8),
	.w5(32'hbcfbd801),
	.w6(32'hbbea66dd),
	.w7(32'hbc2fb0d0),
	.w8(32'hbcb88ec1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e400),
	.w1(32'h3c71ff8a),
	.w2(32'h3c21a6a7),
	.w3(32'hba53df75),
	.w4(32'h3d1adf8c),
	.w5(32'h3c0469de),
	.w6(32'hbad717c4),
	.w7(32'h3cb8d62f),
	.w8(32'h3bbca390),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9a3ad),
	.w1(32'h3b8afec8),
	.w2(32'hbb2caee5),
	.w3(32'h3aaf8966),
	.w4(32'h3ab8fc55),
	.w5(32'hbbbf7096),
	.w6(32'hbb5e4de0),
	.w7(32'hb95cde30),
	.w8(32'hbbdef091),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc504028),
	.w1(32'hbb7a7fb0),
	.w2(32'hbbe90d7c),
	.w3(32'hbc5326a0),
	.w4(32'hbbfef2b4),
	.w5(32'h3b56b534),
	.w6(32'hbc82ee06),
	.w7(32'hbc70be06),
	.w8(32'hbc09e0a4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080ebe),
	.w1(32'h3bbba747),
	.w2(32'h3b1929ef),
	.w3(32'hbbe4d5c0),
	.w4(32'h3b369e25),
	.w5(32'h39cc3f92),
	.w6(32'hba982b57),
	.w7(32'hbb00536a),
	.w8(32'hbb9a73ff),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c05c9),
	.w1(32'h3b25d643),
	.w2(32'h3bae4bea),
	.w3(32'hbc067702),
	.w4(32'hbb0af07b),
	.w5(32'h3c10f64e),
	.w6(32'hbbb50e6d),
	.w7(32'h3ae578ad),
	.w8(32'h3b25e1aa),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4d92),
	.w1(32'hbb02a012),
	.w2(32'hbb89b106),
	.w3(32'hbb658358),
	.w4(32'hbb09ef17),
	.w5(32'h3b731d1d),
	.w6(32'hbaa4ca35),
	.w7(32'h3b563b3c),
	.w8(32'h3bda944f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83a9cb),
	.w1(32'hbb9d7bac),
	.w2(32'hbcdb70c8),
	.w3(32'hba9bace0),
	.w4(32'hbaf63d32),
	.w5(32'hbd569b30),
	.w6(32'h3c6072ec),
	.w7(32'h3b325083),
	.w8(32'hbd0f4d83),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cdeae),
	.w1(32'h3c658467),
	.w2(32'hbbc68fd2),
	.w3(32'hbc293a78),
	.w4(32'h3d48ca21),
	.w5(32'hba7f6a52),
	.w6(32'hbcc120e2),
	.w7(32'h3c90e95f),
	.w8(32'hbac0d5b4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38a461),
	.w1(32'h3aa2d149),
	.w2(32'hbb3c2715),
	.w3(32'hbc318382),
	.w4(32'h3c568da7),
	.w5(32'h3c63038c),
	.w6(32'hbc1e5124),
	.w7(32'hbbcde0d0),
	.w8(32'h3c06a6f1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e244d),
	.w1(32'h3c4d82b5),
	.w2(32'hbbb83c0d),
	.w3(32'h3c71673c),
	.w4(32'h3c1c1bf5),
	.w5(32'hbb9ef975),
	.w6(32'h3c05b545),
	.w7(32'h3ba30f60),
	.w8(32'h38f8710d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cf7aa),
	.w1(32'h39431816),
	.w2(32'h3a1b2756),
	.w3(32'h3b18b431),
	.w4(32'h3bc1fa25),
	.w5(32'h3c038c13),
	.w6(32'hbaf38000),
	.w7(32'h3c4edc76),
	.w8(32'h3ba6d4b4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb855ae0),
	.w1(32'hba95abf5),
	.w2(32'hbbb2f3f9),
	.w3(32'h3ad17198),
	.w4(32'h3b995b19),
	.w5(32'hba7e938e),
	.w6(32'hba707f6d),
	.w7(32'h3b0a4df3),
	.w8(32'h3bf3e00d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9c8e3),
	.w1(32'hbbdbdb09),
	.w2(32'hbae21e62),
	.w3(32'h3c1c520d),
	.w4(32'h3c0592d5),
	.w5(32'hbba8e819),
	.w6(32'h3c534d91),
	.w7(32'h3bbd54f0),
	.w8(32'hbc32f302),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd8da1),
	.w1(32'h3c2af056),
	.w2(32'hbbc0f37a),
	.w3(32'hbbc95808),
	.w4(32'hba0f8e23),
	.w5(32'hbb6e1294),
	.w6(32'hbba54b7a),
	.w7(32'hbb5a295a),
	.w8(32'hbbb4f191),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbad92),
	.w1(32'hbba43e9d),
	.w2(32'hba2f2836),
	.w3(32'hbb8563c1),
	.w4(32'hbb102ab3),
	.w5(32'h3b9f1828),
	.w6(32'hbbeb4775),
	.w7(32'hbb588f4f),
	.w8(32'h3a216a0a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4516be),
	.w1(32'h3abe0107),
	.w2(32'hbc35e087),
	.w3(32'h3bab62bf),
	.w4(32'h3c262131),
	.w5(32'hbc31f65a),
	.w6(32'h3a603e48),
	.w7(32'h3c0ab1da),
	.w8(32'hbb9fbd02),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91088a),
	.w1(32'hbc010a9c),
	.w2(32'hbaaf18bd),
	.w3(32'hbcd39ba3),
	.w4(32'hbc6997b9),
	.w5(32'h3c2f18ce),
	.w6(32'hbb72a80d),
	.w7(32'hbad0f4a7),
	.w8(32'h3ba62977),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad4d0f),
	.w1(32'hbb26ce7e),
	.w2(32'hbb7591d2),
	.w3(32'h3c9763a8),
	.w4(32'h3c28f529),
	.w5(32'hbbe8193a),
	.w6(32'h3c5e278b),
	.w7(32'h3bcaeae4),
	.w8(32'hbc48a3f2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86132b),
	.w1(32'hbb65f8c0),
	.w2(32'h3bbf4ef1),
	.w3(32'hbc716739),
	.w4(32'h39a9b012),
	.w5(32'h3c26a320),
	.w6(32'hbc16e93e),
	.w7(32'hbba5f61b),
	.w8(32'h3c5f46dd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e5372),
	.w1(32'h3c0f7978),
	.w2(32'h3c3e2728),
	.w3(32'h3c4b6029),
	.w4(32'h3c60c615),
	.w5(32'h3c50db02),
	.w6(32'h3c892d48),
	.w7(32'h3c6587fb),
	.w8(32'h3ab1ca0d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7662f4),
	.w1(32'h3c460c6a),
	.w2(32'hbc28a7a8),
	.w3(32'h3c4ac547),
	.w4(32'h3b89eb94),
	.w5(32'hbbdbc163),
	.w6(32'h3b59c8f1),
	.w7(32'hba83d01a),
	.w8(32'hbc39aab9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63dec1),
	.w1(32'hbc7055dd),
	.w2(32'hbb873acb),
	.w3(32'hbc29cc7d),
	.w4(32'hbbf55964),
	.w5(32'hbc7e2358),
	.w6(32'hbbd7f977),
	.w7(32'hbc12178d),
	.w8(32'hbbde0b5c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf636a3),
	.w1(32'hbbe592dc),
	.w2(32'hbbe573ac),
	.w3(32'hbc4bd456),
	.w4(32'hbb1dcc5c),
	.w5(32'hbb72a8f3),
	.w6(32'hbba6ff05),
	.w7(32'hbafc35ac),
	.w8(32'hbb9ffb2b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd36b1),
	.w1(32'hbca6b051),
	.w2(32'hbc015248),
	.w3(32'hbcdd05ea),
	.w4(32'hbc95c602),
	.w5(32'hbbe1d48a),
	.w6(32'hbc6f3f7e),
	.w7(32'hbc3792b8),
	.w8(32'hbb1a6786),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9155de),
	.w1(32'hbb2e1144),
	.w2(32'hbc740f27),
	.w3(32'hbb8db28b),
	.w4(32'hbc0d8643),
	.w5(32'hbca8bf3e),
	.w6(32'hbc5ea7ad),
	.w7(32'hbc0e6c4e),
	.w8(32'hbcb5530b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210a50),
	.w1(32'hbbd124bd),
	.w2(32'h3bca6871),
	.w3(32'hbc26198e),
	.w4(32'hbbcc5893),
	.w5(32'h3c2d5137),
	.w6(32'hbbc94a49),
	.w7(32'hbb480897),
	.w8(32'h3bb27fef),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f6f6d),
	.w1(32'h3c3a33a7),
	.w2(32'hbb6ee3fe),
	.w3(32'h3c88eb08),
	.w4(32'h3c86cb7a),
	.w5(32'hbaa86c41),
	.w6(32'h3c6c399d),
	.w7(32'h3c157106),
	.w8(32'h3a085192),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44c305),
	.w1(32'hbaa60452),
	.w2(32'h3b42430c),
	.w3(32'hbae1549e),
	.w4(32'h3b191b74),
	.w5(32'hbc1e6e31),
	.w6(32'hba7b192e),
	.w7(32'hba801790),
	.w8(32'hbc0c8678),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91a8f7),
	.w1(32'h3a8ca057),
	.w2(32'hbb57b417),
	.w3(32'hbc86b3fb),
	.w4(32'hbb9d6128),
	.w5(32'hbc63e128),
	.w6(32'hbc9c661f),
	.w7(32'hbc16f1c2),
	.w8(32'hbc86a281),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c0efa),
	.w1(32'hbb3b3663),
	.w2(32'hbb9de228),
	.w3(32'hbc336f28),
	.w4(32'hbaffcacb),
	.w5(32'hbb0a39dc),
	.w6(32'hbc0bdaa8),
	.w7(32'hbbb049ae),
	.w8(32'h3be52e30),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbda1c),
	.w1(32'h3b935f17),
	.w2(32'hbc5dbc1f),
	.w3(32'hbb0cd81a),
	.w4(32'h3b40c263),
	.w5(32'hbc88478f),
	.w6(32'h3ae461d2),
	.w7(32'hba3f7b31),
	.w8(32'hbc8b321b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23d1df),
	.w1(32'hb928e962),
	.w2(32'hbb91bc69),
	.w3(32'hbb96a962),
	.w4(32'hbc1822f2),
	.w5(32'hbbd5c59d),
	.w6(32'hbb78c63c),
	.w7(32'hbc07221c),
	.w8(32'h3a596da9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d0bef),
	.w1(32'hbb3aa4ac),
	.w2(32'hbaa186e5),
	.w3(32'hbc71fffa),
	.w4(32'hbb5ffee1),
	.w5(32'h3c3f37d5),
	.w6(32'hbc00ebe7),
	.w7(32'hba81a828),
	.w8(32'h3bc3ea83),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0144b),
	.w1(32'h3ac50e6e),
	.w2(32'h3c1514f3),
	.w3(32'h3cac9201),
	.w4(32'h3c3a2e7b),
	.w5(32'h3c16f47d),
	.w6(32'h3c4f8daa),
	.w7(32'h3c465aa0),
	.w8(32'h3b6a980f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c982c84),
	.w1(32'h3c30478d),
	.w2(32'h3ab7837d),
	.w3(32'h3c8505f9),
	.w4(32'h3c8df02e),
	.w5(32'h39d5317c),
	.w6(32'h3c724986),
	.w7(32'h3c802911),
	.w8(32'hbbac099c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a767300),
	.w1(32'h3ac551ef),
	.w2(32'h3c780690),
	.w3(32'hbc30ce74),
	.w4(32'hbb91499c),
	.w5(32'h3bf2725c),
	.w6(32'hbc09e550),
	.w7(32'hbc076cdf),
	.w8(32'h3b40209f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea6f45),
	.w1(32'h3c13f4aa),
	.w2(32'hbbc40a6d),
	.w3(32'h3c4a1e0a),
	.w4(32'h3c4185d3),
	.w5(32'h3b209f6d),
	.w6(32'hbafe7aa3),
	.w7(32'h3a9be332),
	.w8(32'hbb1ab737),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12d348),
	.w1(32'h3b591647),
	.w2(32'hbaf08c4d),
	.w3(32'h3bded32b),
	.w4(32'h3b35762a),
	.w5(32'h3a55c76d),
	.w6(32'hbb84f8c9),
	.w7(32'hbb362129),
	.w8(32'hbc1320b8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7dfeb0),
	.w1(32'hba3e008e),
	.w2(32'hbc892d7e),
	.w3(32'hbb0cd729),
	.w4(32'h39cb7875),
	.w5(32'hbca745d2),
	.w6(32'hbbaef5c7),
	.w7(32'h3ba1b751),
	.w8(32'hbc8700b0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbad981),
	.w1(32'hbc6035c8),
	.w2(32'hbc0021a5),
	.w3(32'hbcd7402a),
	.w4(32'hbca4cc46),
	.w5(32'h3baf1bc1),
	.w6(32'hbcc75084),
	.w7(32'hbc62a382),
	.w8(32'hbb827ac6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2b72e),
	.w1(32'hbc415ad1),
	.w2(32'hbc349d94),
	.w3(32'h3b8394f3),
	.w4(32'hbc482844),
	.w5(32'hbc1acf4a),
	.w6(32'h3bb33bcd),
	.w7(32'hbc38ef58),
	.w8(32'hbc3c66fa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9df65c),
	.w1(32'hbc6499fa),
	.w2(32'h3b833987),
	.w3(32'hbc916cf4),
	.w4(32'hbc24898d),
	.w5(32'h3c0c997a),
	.w6(32'hbc877fef),
	.w7(32'hbbbcde42),
	.w8(32'h3cd5258c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72bb3c),
	.w1(32'h3c512ef4),
	.w2(32'hbc0d8a50),
	.w3(32'h3bb85e5f),
	.w4(32'h3c7c1529),
	.w5(32'hbba2da65),
	.w6(32'h3cfa66ef),
	.w7(32'h3d19818b),
	.w8(32'hbbbbb58e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf4014),
	.w1(32'hbbd37460),
	.w2(32'hbc0d4a42),
	.w3(32'hbc3e4f5f),
	.w4(32'hbbae5ccc),
	.w5(32'hbc38ae3e),
	.w6(32'hbb8dd2d6),
	.w7(32'h3b7a215e),
	.w8(32'hbbc914fa),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab63d82),
	.w1(32'h3b0bff3a),
	.w2(32'hbbc361b3),
	.w3(32'hb8f792ee),
	.w4(32'h3ca288c1),
	.w5(32'hbb31e937),
	.w6(32'hbb580f3b),
	.w7(32'h3b8f2e65),
	.w8(32'hbc0b499f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a159f17),
	.w1(32'h3b262301),
	.w2(32'hbab036bf),
	.w3(32'h39bed1ab),
	.w4(32'h3ba8d3f6),
	.w5(32'h3c248049),
	.w6(32'hbaf830f0),
	.w7(32'h3a793ce9),
	.w8(32'h3baea4af),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f8df4),
	.w1(32'h3bf33278),
	.w2(32'hbca68526),
	.w3(32'h3c9dcb0f),
	.w4(32'h3c23aeb3),
	.w5(32'hbc21a79f),
	.w6(32'h3c6527ac),
	.w7(32'h3bcdcbc9),
	.w8(32'hbc546966),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2d8d9),
	.w1(32'hbc2feb6e),
	.w2(32'h3bd8113b),
	.w3(32'hbc59606d),
	.w4(32'hbbc22949),
	.w5(32'h3c5d0c0c),
	.w6(32'hbcaac6aa),
	.w7(32'hbc80e90a),
	.w8(32'h3c2b2e43),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9232a),
	.w1(32'h3bdbe2d7),
	.w2(32'hbbea0b37),
	.w3(32'h3c9435f8),
	.w4(32'h3c1f4aa5),
	.w5(32'hbc357e80),
	.w6(32'h3c24fe32),
	.w7(32'h3c303bca),
	.w8(32'hbc5b5ada),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3653c5),
	.w1(32'hbc0804c0),
	.w2(32'hbafe56ce),
	.w3(32'hbc47684a),
	.w4(32'hbc537f6e),
	.w5(32'h3b107bd1),
	.w6(32'hbc73b902),
	.w7(32'hbc449a0e),
	.w8(32'hba403acd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc214370),
	.w1(32'hbc26dac0),
	.w2(32'h3c24c47d),
	.w3(32'hbba7248a),
	.w4(32'hbb92a45e),
	.w5(32'h3c8a1944),
	.w6(32'hbc02aa24),
	.w7(32'hbc642786),
	.w8(32'h3c17508a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c985563),
	.w1(32'h3c2e1404),
	.w2(32'hbaa4bda1),
	.w3(32'h3d083573),
	.w4(32'h3ca271f9),
	.w5(32'h3c1ee858),
	.w6(32'h3c8e5b4d),
	.w7(32'h3c5fa6ce),
	.w8(32'h3b01bf91),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cb924),
	.w1(32'h3a5a6fd1),
	.w2(32'hbc895f42),
	.w3(32'h3cc272ae),
	.w4(32'h3c6e99cd),
	.w5(32'hbcb2b1af),
	.w6(32'h3c444a79),
	.w7(32'h3bd45769),
	.w8(32'hbca0596a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf07d8e),
	.w1(32'hbc77ccac),
	.w2(32'hbb8ab0e9),
	.w3(32'hbd0a6038),
	.w4(32'hbca1874e),
	.w5(32'hbb75694a),
	.w6(32'hbd05cfa3),
	.w7(32'hbcb5277b),
	.w8(32'hbbf6fdb0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93335c),
	.w1(32'hbc72beaf),
	.w2(32'h3b703960),
	.w3(32'hbb5dee02),
	.w4(32'hbc86d2b0),
	.w5(32'h3bb5907b),
	.w6(32'hbc245184),
	.w7(32'hbc79079a),
	.w8(32'h3b9f5c98),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7df96),
	.w1(32'h3a632bf1),
	.w2(32'hba030eb4),
	.w3(32'h3b9b36fe),
	.w4(32'h3ac8a0f2),
	.w5(32'h3c5db539),
	.w6(32'h3be5c651),
	.w7(32'h3b83932d),
	.w8(32'h3c67a7e1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e93d8),
	.w1(32'hba98cecb),
	.w2(32'hbc272664),
	.w3(32'h3ca1bb11),
	.w4(32'h3bec422a),
	.w5(32'hbc593e7b),
	.w6(32'h3c838687),
	.w7(32'h3af5b4cb),
	.w8(32'hbc4c16b7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd518d1),
	.w1(32'h3b33a96f),
	.w2(32'hb8d806fe),
	.w3(32'hbc797a41),
	.w4(32'hbaaf47db),
	.w5(32'hba87d077),
	.w6(32'hbc064913),
	.w7(32'h3bafd4d6),
	.w8(32'h3b5fc67c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb851f8c),
	.w1(32'h3b9775eb),
	.w2(32'h3b9ef5b2),
	.w3(32'hbc0ce574),
	.w4(32'h3b9b1bb9),
	.w5(32'h3cb73479),
	.w6(32'hbb3ad884),
	.w7(32'h3baa1959),
	.w8(32'h3c473b9b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c848a50),
	.w1(32'h3bb15746),
	.w2(32'h3a981a58),
	.w3(32'h3d45418f),
	.w4(32'h3d0b1978),
	.w5(32'h3c12cebb),
	.w6(32'h3cf5ce7f),
	.w7(32'h3c9ff8ea),
	.w8(32'h3a1d03f3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75e16d),
	.w1(32'h3c0591cf),
	.w2(32'h3c0cd902),
	.w3(32'h3cd5dd5c),
	.w4(32'h3cb87370),
	.w5(32'h3c5fd079),
	.w6(32'h3c14d357),
	.w7(32'h3c654c95),
	.w8(32'hbadb543f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae9169),
	.w1(32'h3c407620),
	.w2(32'h3bd21ce6),
	.w3(32'h3cb3c40c),
	.w4(32'h3cae4475),
	.w5(32'h3bac9387),
	.w6(32'h3c2c7e61),
	.w7(32'h3c696e06),
	.w8(32'hba9aca84),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819b9b),
	.w1(32'h3b7f5cc3),
	.w2(32'h39292419),
	.w3(32'h3c3c917c),
	.w4(32'h3b8e1771),
	.w5(32'h3b0d21cb),
	.w6(32'h3b5c8a2b),
	.w7(32'h3ba3de8f),
	.w8(32'hb91d0ef9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfdf81),
	.w1(32'h39deb87d),
	.w2(32'hbc000b91),
	.w3(32'hbbd0dee6),
	.w4(32'h3aa592ae),
	.w5(32'hbbc0f941),
	.w6(32'hbb9f2968),
	.w7(32'h3a95327d),
	.w8(32'hbb8be138),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b7eb0),
	.w1(32'hbbcb866a),
	.w2(32'hbbe1f65b),
	.w3(32'hbb937e39),
	.w4(32'hbbb770ec),
	.w5(32'h3b538589),
	.w6(32'hba4a5e72),
	.w7(32'hbb471c75),
	.w8(32'hbbab2369),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7519),
	.w1(32'hbbb077df),
	.w2(32'h3c0a1854),
	.w3(32'h3bb189d6),
	.w4(32'h3ba11eb3),
	.w5(32'h3c416c50),
	.w6(32'h3adcc182),
	.w7(32'hb98af4cb),
	.w8(32'h3be6a915),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3763a3),
	.w1(32'h3bbc0e84),
	.w2(32'h3ba52d77),
	.w3(32'h3a275482),
	.w4(32'hb95fe4fd),
	.w5(32'hba02b0b8),
	.w6(32'h3b0fcfd2),
	.w7(32'h3af97f96),
	.w8(32'hbb890551),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c347747),
	.w1(32'h3b8829b0),
	.w2(32'h3c054802),
	.w3(32'h3c4f6cd6),
	.w4(32'h3b9f8ae3),
	.w5(32'h3c821b1c),
	.w6(32'h3bcfcf65),
	.w7(32'h3bfb2aae),
	.w8(32'h3c159dd3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21fb40),
	.w1(32'h3b7bdbfa),
	.w2(32'hbc045fc0),
	.w3(32'h3c71a698),
	.w4(32'h3b625554),
	.w5(32'hbc41de0b),
	.w6(32'h3bddd244),
	.w7(32'hbabc2a99),
	.w8(32'hbc8fe752),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac8b9b),
	.w1(32'hbc09f7b5),
	.w2(32'hbc074e2a),
	.w3(32'hbc4468c1),
	.w4(32'hbc9bbf9b),
	.w5(32'hbc2453c9),
	.w6(32'hbc63619c),
	.w7(32'hbc73fb82),
	.w8(32'hbc1e9fb0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08ba4d),
	.w1(32'hbb0afad4),
	.w2(32'h3b302c0a),
	.w3(32'h3960f17c),
	.w4(32'h3b4f865e),
	.w5(32'h3be43924),
	.w6(32'hbb5e1da5),
	.w7(32'hbc05a329),
	.w8(32'hbb953b9c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5314f0),
	.w1(32'hbaf9b846),
	.w2(32'h3bd7408d),
	.w3(32'hbba6f6e2),
	.w4(32'hbb9e44d7),
	.w5(32'h3c1806fa),
	.w6(32'hbb6b8b46),
	.w7(32'hbb16a08c),
	.w8(32'h3b6414ce),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57eaa2),
	.w1(32'h3bcb9cb6),
	.w2(32'hbc7f6f64),
	.w3(32'h3c768a3a),
	.w4(32'h3c4b7355),
	.w5(32'hbc4db99e),
	.w6(32'h3c1db11a),
	.w7(32'h3bd7ba0d),
	.w8(32'hbc49a346),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ba637),
	.w1(32'hbc49272f),
	.w2(32'h3b7e60e7),
	.w3(32'hbc178fe4),
	.w4(32'hbc505c47),
	.w5(32'h3b2a8527),
	.w6(32'hbc50775d),
	.w7(32'hbba6b4e4),
	.w8(32'hbbcbb6f5),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6506b),
	.w1(32'hbac36897),
	.w2(32'h3b2506dc),
	.w3(32'hbc08b50e),
	.w4(32'hbb86364d),
	.w5(32'hbb781d36),
	.w6(32'hbc915f29),
	.w7(32'hbc6bfcf9),
	.w8(32'hbaa44748),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc003327),
	.w1(32'hba4c6f91),
	.w2(32'hbba1125e),
	.w3(32'hbcc167a1),
	.w4(32'hbc068115),
	.w5(32'hb93199a6),
	.w6(32'hbc6ae779),
	.w7(32'h3953dfd1),
	.w8(32'hbb86407c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb319ee),
	.w1(32'hb9b7610f),
	.w2(32'hbb3c6c6d),
	.w3(32'hbaba1b34),
	.w4(32'h3b6de33b),
	.w5(32'hbb76dc82),
	.w6(32'hbb58e86f),
	.w7(32'hbab1a180),
	.w8(32'hbb942226),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1479f8),
	.w1(32'hbb0a6096),
	.w2(32'hb9e88d52),
	.w3(32'hbc226d26),
	.w4(32'hbb0b5e48),
	.w5(32'h3c28a89b),
	.w6(32'hbc0f40d9),
	.w7(32'hbb6fb60b),
	.w8(32'h3b25d1c6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b0cff),
	.w1(32'h3b6062d3),
	.w2(32'h3b1f2ab5),
	.w3(32'h3cd15371),
	.w4(32'h3c21bd41),
	.w5(32'hbc0f006a),
	.w6(32'h3c5863ab),
	.w7(32'h3c185dab),
	.w8(32'hbb8f8c86),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb756),
	.w1(32'h3a8baed2),
	.w2(32'hbb93148e),
	.w3(32'hbb868024),
	.w4(32'hbc79991d),
	.w5(32'h3bd1b6fe),
	.w6(32'hbc129074),
	.w7(32'hbb80c655),
	.w8(32'h3b17659b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39f5bf),
	.w1(32'hbbd6b345),
	.w2(32'h3b9b5c30),
	.w3(32'h3c9c6256),
	.w4(32'h3b9f9f14),
	.w5(32'h3c3a833b),
	.w6(32'h3b4b0f72),
	.w7(32'h39581c50),
	.w8(32'h3c189bc3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab2aba),
	.w1(32'h3bf78004),
	.w2(32'hbb26c95c),
	.w3(32'h3cbf24ce),
	.w4(32'h3cabd211),
	.w5(32'hbbcc1d58),
	.w6(32'h3c83bc66),
	.w7(32'h3c7e28ec),
	.w8(32'hbb494b45),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd7014),
	.w1(32'h3c45bce6),
	.w2(32'h3b00ccb3),
	.w3(32'hb917f10f),
	.w4(32'h3b30b330),
	.w5(32'h3c0c581a),
	.w6(32'hbaddc5e5),
	.w7(32'h3c123d49),
	.w8(32'h3c1d30ff),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c23e),
	.w1(32'hbbf10918),
	.w2(32'hbbee7fbc),
	.w3(32'hbb93c24e),
	.w4(32'hbc0a6884),
	.w5(32'hbb6dcf75),
	.w6(32'hbbb2d0e5),
	.w7(32'hbbd0db9b),
	.w8(32'hbb87acd4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1c10),
	.w1(32'h3b93d1b3),
	.w2(32'hbb642c0e),
	.w3(32'h3b95c006),
	.w4(32'h3bf62d67),
	.w5(32'h3be6360d),
	.w6(32'h3baa8e56),
	.w7(32'h3c174e34),
	.w8(32'hb9e73db0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ddecd),
	.w1(32'hbb346442),
	.w2(32'hbbc0dbe6),
	.w3(32'h3c560381),
	.w4(32'h3c186ec6),
	.w5(32'hbbf6a614),
	.w6(32'h3bc8f70b),
	.w7(32'h3b2309b6),
	.w8(32'hba88da7b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5875af),
	.w1(32'hbbe063ca),
	.w2(32'hbade0dbc),
	.w3(32'hbc8fe29c),
	.w4(32'hbc689548),
	.w5(32'hbabd544f),
	.w6(32'hbc6e0a52),
	.w7(32'hbc1ffbd6),
	.w8(32'hbc1f1a66),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e07503),
	.w1(32'hbab5ad40),
	.w2(32'h3c0bb728),
	.w3(32'hbba67aae),
	.w4(32'hbc199aae),
	.w5(32'h3c14e94c),
	.w6(32'hbc82b584),
	.w7(32'hbc8f7346),
	.w8(32'h3b666e8f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2fbbd),
	.w1(32'h3b88de77),
	.w2(32'hbacd077d),
	.w3(32'h3b1bd5af),
	.w4(32'hbbee27d0),
	.w5(32'h3b3d85e5),
	.w6(32'h3afff412),
	.w7(32'hbbca6deb),
	.w8(32'h3bda7c0d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53c69),
	.w1(32'hbbc8e3b2),
	.w2(32'hbbaf15d5),
	.w3(32'hbb8826e2),
	.w4(32'hbc0e5245),
	.w5(32'hbb840ac7),
	.w6(32'hbb09daf9),
	.w7(32'hbb8ca741),
	.w8(32'hbb8fdffa),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24df7e),
	.w1(32'hbadaf674),
	.w2(32'h39eae91d),
	.w3(32'h39aef913),
	.w4(32'hbac93211),
	.w5(32'h3a9cf755),
	.w6(32'h39d865bb),
	.w7(32'hbabefd94),
	.w8(32'h3bb62eb6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71ef39),
	.w1(32'hbc6a84f0),
	.w2(32'hbac57d5e),
	.w3(32'hbbf576a3),
	.w4(32'hbc773685),
	.w5(32'h3c2b0e25),
	.w6(32'hbb5aa21f),
	.w7(32'hbab85efc),
	.w8(32'h3c612ac9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4313f),
	.w1(32'h3c0736d0),
	.w2(32'hbb58d0b9),
	.w3(32'h3c087b62),
	.w4(32'h3b27d188),
	.w5(32'h3b61d8eb),
	.w6(32'h3c4cf181),
	.w7(32'h3b83d5af),
	.w8(32'hbb4c09ad),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3a4da),
	.w1(32'hbafb49cf),
	.w2(32'h3babe1e0),
	.w3(32'h3b5c1e59),
	.w4(32'h3c4b367d),
	.w5(32'h3c1c97bf),
	.w6(32'h3afb01fb),
	.w7(32'h3b570cb8),
	.w8(32'h3b90551d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42d762),
	.w1(32'h3c79eafd),
	.w2(32'h3993685a),
	.w3(32'h3c9a2a13),
	.w4(32'h3c855f06),
	.w5(32'hbaf7b722),
	.w6(32'h3c2a31fc),
	.w7(32'h3c39a4cc),
	.w8(32'h3ba0d4cf),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67875e),
	.w1(32'hbb9742ad),
	.w2(32'hbc440702),
	.w3(32'hbc7b34fa),
	.w4(32'hbba93d18),
	.w5(32'hbc22a622),
	.w6(32'hbc31522a),
	.w7(32'hbc54a633),
	.w8(32'hbbffce15),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592462),
	.w1(32'hbc230c39),
	.w2(32'h3a95c913),
	.w3(32'hbbe24453),
	.w4(32'hbc1cba03),
	.w5(32'h3bb53200),
	.w6(32'hbbd0df70),
	.w7(32'hbc1e3a84),
	.w8(32'h3aa98943),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f6169),
	.w1(32'hba4cd805),
	.w2(32'hbc315f4e),
	.w3(32'h3adb6c4a),
	.w4(32'h3c7ab92c),
	.w5(32'hbc03fd01),
	.w6(32'h3bd52ab1),
	.w7(32'h3c46f99b),
	.w8(32'hbca19a25),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6f75),
	.w1(32'hbb597ad3),
	.w2(32'h3a936aed),
	.w3(32'hbc848cbc),
	.w4(32'hbb21c46b),
	.w5(32'h390f3020),
	.w6(32'hbc0a6de7),
	.w7(32'h3af80f5d),
	.w8(32'h39751cd1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab79ec),
	.w1(32'h38a00b44),
	.w2(32'h3a3e790f),
	.w3(32'hbb154a2e),
	.w4(32'h3911693e),
	.w5(32'h3b575bc7),
	.w6(32'hbb04e176),
	.w7(32'h39f34e5e),
	.w8(32'hbbb1ae70),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43fa49),
	.w1(32'hbb7426a3),
	.w2(32'hbbd1b46e),
	.w3(32'hbad900e2),
	.w4(32'hbc216c5d),
	.w5(32'hbb92333a),
	.w6(32'hbc314349),
	.w7(32'hbc47209b),
	.w8(32'h3b9cc19a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfac50f),
	.w1(32'hbb58bf8d),
	.w2(32'hbba16ef2),
	.w3(32'hb8a89cdc),
	.w4(32'hbaa303e3),
	.w5(32'hbaa58029),
	.w6(32'h3bdc07f4),
	.w7(32'h3bf81688),
	.w8(32'hbbbbf808),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb080),
	.w1(32'hbbb715bc),
	.w2(32'hbbbbffdd),
	.w3(32'hbbda1f26),
	.w4(32'hbab1368b),
	.w5(32'h3c03d657),
	.w6(32'hbc234dc0),
	.w7(32'hbb1e0e4b),
	.w8(32'h3b5ab6c9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2a2b7),
	.w1(32'hbb8e83b2),
	.w2(32'h3bb602e0),
	.w3(32'h3c814187),
	.w4(32'h3c224e6a),
	.w5(32'h3c26066f),
	.w6(32'h3c64be69),
	.w7(32'h3b97b541),
	.w8(32'h3b67b24d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55a4d1),
	.w1(32'h3bbb92b8),
	.w2(32'hbb19e721),
	.w3(32'h3cf19e18),
	.w4(32'h3c90f78b),
	.w5(32'hbbc4bb3f),
	.w6(32'h3c9acf85),
	.w7(32'h3c0751b2),
	.w8(32'hbb22033f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafc4f1),
	.w1(32'hbb026454),
	.w2(32'h3a95ea6a),
	.w3(32'hbc04fc1b),
	.w4(32'hbb995e97),
	.w5(32'h3b9177dd),
	.w6(32'hbba9928a),
	.w7(32'hba8df3cd),
	.w8(32'h3b723cbb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01d783),
	.w1(32'h3bc41050),
	.w2(32'hbb57eb23),
	.w3(32'h3c718b1b),
	.w4(32'h3c1e9354),
	.w5(32'hbc846310),
	.w6(32'h3c0f0fbf),
	.w7(32'h3bf12e48),
	.w8(32'hbc28b9e4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b4cfb),
	.w1(32'hbb9e1fd4),
	.w2(32'hbc2ced8d),
	.w3(32'hbb2016ed),
	.w4(32'hba17a247),
	.w5(32'hbc3bf1fa),
	.w6(32'h3aa561fb),
	.w7(32'hbbaeaf68),
	.w8(32'hbb63fd04),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24eff1),
	.w1(32'hbc0afb7a),
	.w2(32'h3bb6e5b1),
	.w3(32'hbc174c03),
	.w4(32'hbc14f0e0),
	.w5(32'h3b6590a4),
	.w6(32'hbb5755f9),
	.w7(32'hbbc042b0),
	.w8(32'h3b87a6df),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8438a1),
	.w1(32'h3c3d4f98),
	.w2(32'h3b45be87),
	.w3(32'hbbda9ff3),
	.w4(32'h3c5dc61b),
	.w5(32'h3bae1e14),
	.w6(32'hbb8d91c3),
	.w7(32'hbbbcb725),
	.w8(32'h3be52e8c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6ea9),
	.w1(32'h3c0aa7fb),
	.w2(32'h3bb22272),
	.w3(32'h3cc20e1b),
	.w4(32'h3bcd9fda),
	.w5(32'h3c59ef4d),
	.w6(32'h3c895380),
	.w7(32'h3a98fc96),
	.w8(32'h3c1cce5a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf7bbd),
	.w1(32'h3b9dc2a2),
	.w2(32'hbc53a0cf),
	.w3(32'h3cc07c71),
	.w4(32'h3c43f87c),
	.w5(32'hba8efabb),
	.w6(32'h3c6036cb),
	.w7(32'h3c02ee8b),
	.w8(32'hbb320e63),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule