module layer_10_featuremap_345(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4192b5),
	.w1(32'h3b84f3a1),
	.w2(32'h38034def),
	.w3(32'h3af9e572),
	.w4(32'hbad804c5),
	.w5(32'hbb65413e),
	.w6(32'h3b5095e0),
	.w7(32'h3a98feff),
	.w8(32'hbb39269c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c3b0),
	.w1(32'hbc3095e6),
	.w2(32'hbc57673e),
	.w3(32'hbbc5db01),
	.w4(32'hbb41cc31),
	.w5(32'hbb8a9431),
	.w6(32'h3b4c03ab),
	.w7(32'hba591298),
	.w8(32'hb95c28a3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d94cb),
	.w1(32'hba86147b),
	.w2(32'hbb20ac61),
	.w3(32'hb9f3cf7d),
	.w4(32'hba5d2d75),
	.w5(32'hb9837cd9),
	.w6(32'hbb6961d4),
	.w7(32'hbb4276d5),
	.w8(32'h37cda9a7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f9a580),
	.w1(32'h3ac493e3),
	.w2(32'h3a88e960),
	.w3(32'h39c101a6),
	.w4(32'h3ae31911),
	.w5(32'h39fb316a),
	.w6(32'h3aa92efb),
	.w7(32'h3b561ed0),
	.w8(32'hba9c7ba8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcbb77),
	.w1(32'h3b9c58d6),
	.w2(32'h3c3af74c),
	.w3(32'hbae4a79b),
	.w4(32'h3962dee2),
	.w5(32'h3b050ca2),
	.w6(32'hbac66ae7),
	.w7(32'h3b3359b9),
	.w8(32'h3afb38b2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3954e),
	.w1(32'h3b42bea3),
	.w2(32'h3a8b05a1),
	.w3(32'hb941d4df),
	.w4(32'hba1b8931),
	.w5(32'h3ac4721c),
	.w6(32'h3ac57d0c),
	.w7(32'h3b1117d0),
	.w8(32'hba7d0a91),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394baf),
	.w1(32'h3b0719b2),
	.w2(32'h3bdd400c),
	.w3(32'h3ab9e216),
	.w4(32'hba604d99),
	.w5(32'h3bb515fb),
	.w6(32'hbc1f7fea),
	.w7(32'h3afe5ea8),
	.w8(32'h3c0adae9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b51fc),
	.w1(32'h3c56db81),
	.w2(32'h3cc30bd7),
	.w3(32'hbc0a0c57),
	.w4(32'h3b356961),
	.w5(32'h3c659d79),
	.w6(32'hbc4a6de7),
	.w7(32'h3b361ade),
	.w8(32'h3b839cf6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fc25e),
	.w1(32'h3b8e4ba7),
	.w2(32'h3ba3ca6d),
	.w3(32'h3b9fa4d1),
	.w4(32'h3bc68029),
	.w5(32'h3ab529f6),
	.w6(32'h3ad35a7f),
	.w7(32'h3b8690a7),
	.w8(32'h3b3c777a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d496),
	.w1(32'h3c70054b),
	.w2(32'h3c357d12),
	.w3(32'h3b11805a),
	.w4(32'h3ba2f4d1),
	.w5(32'h3bf7c376),
	.w6(32'hbba03e01),
	.w7(32'hba05c51c),
	.w8(32'hb94bf4e6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31a3ec),
	.w1(32'h3b1dd29e),
	.w2(32'h3a41a008),
	.w3(32'hba5bd29a),
	.w4(32'hba3c8385),
	.w5(32'h3b32c74c),
	.w6(32'hbb171cae),
	.w7(32'h3ac500c9),
	.w8(32'hb9837ad1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d4dc4),
	.w1(32'h3c0a5af4),
	.w2(32'h3c4446f4),
	.w3(32'h3b5cf78f),
	.w4(32'hb88c980d),
	.w5(32'h3a23d367),
	.w6(32'hbc09021d),
	.w7(32'hbba242b1),
	.w8(32'hbb2a3caf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52d3a0),
	.w1(32'h3c8de25f),
	.w2(32'h3c538d04),
	.w3(32'h3b6f3378),
	.w4(32'h3c0458b2),
	.w5(32'h3bbdba9d),
	.w6(32'hbba4ef64),
	.w7(32'hbb2f58c3),
	.w8(32'hbb2a3277),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad8fbe),
	.w1(32'h3b1ba710),
	.w2(32'h3baa1dc4),
	.w3(32'hba903372),
	.w4(32'h3b676e78),
	.w5(32'h3c2c4610),
	.w6(32'hbb680820),
	.w7(32'h3b3c04cf),
	.w8(32'h3bf84de3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3d5ca),
	.w1(32'hbb73aa24),
	.w2(32'hbad52d90),
	.w3(32'h3b59a0eb),
	.w4(32'h3b19faa6),
	.w5(32'hbbb028ad),
	.w6(32'h3b5f63d3),
	.w7(32'h3ba475e8),
	.w8(32'hbb8ed70b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03e8a2),
	.w1(32'h3bb4b168),
	.w2(32'h3ba94eb6),
	.w3(32'hbb9ed623),
	.w4(32'h38e3a7f7),
	.w5(32'h3bda0a3c),
	.w6(32'hbbc9ec49),
	.w7(32'hbbd4fc4e),
	.w8(32'hb9b551bf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944036),
	.w1(32'h3beb0993),
	.w2(32'h3b172011),
	.w3(32'h3a9e1a6c),
	.w4(32'h3ac59f11),
	.w5(32'hb962e57a),
	.w6(32'h3a9d081c),
	.w7(32'h3b048f5f),
	.w8(32'hba2994e4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31660b),
	.w1(32'h3c914942),
	.w2(32'h3c5fa697),
	.w3(32'hbbe30e57),
	.w4(32'h3c18ea6f),
	.w5(32'h3b950aac),
	.w6(32'hbc3819c2),
	.w7(32'hbb5592ba),
	.w8(32'hbb274fea),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d7ea),
	.w1(32'h3bfe8e9d),
	.w2(32'h3be4ddbc),
	.w3(32'hb986320c),
	.w4(32'h3bb282a8),
	.w5(32'h3b249814),
	.w6(32'hbbc3fc1a),
	.w7(32'hbb27810c),
	.w8(32'hbb0ae3c4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad3cf5),
	.w1(32'hb9365db7),
	.w2(32'hbaf86cc2),
	.w3(32'hbb8e1ae5),
	.w4(32'hbbd60170),
	.w5(32'hbb6a6548),
	.w6(32'hbade7c8b),
	.w7(32'hbb66186d),
	.w8(32'hbb6e4b7f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7ffa6),
	.w1(32'hba64ead7),
	.w2(32'hba95f0b4),
	.w3(32'hba5d4579),
	.w4(32'hb96ddef1),
	.w5(32'h3b1fbf7e),
	.w6(32'hba52ebc2),
	.w7(32'hbaed4304),
	.w8(32'h3a4fde44),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75f035),
	.w1(32'hbb16d9bc),
	.w2(32'hbadefefa),
	.w3(32'h3b787e92),
	.w4(32'h3b643074),
	.w5(32'hbb82c501),
	.w6(32'h3b9cc7fd),
	.w7(32'h3bae1377),
	.w8(32'hbb0023b0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c729a24),
	.w1(32'h3b6bf7c0),
	.w2(32'h3c87b9b5),
	.w3(32'hbc015397),
	.w4(32'h3a0a995d),
	.w5(32'h3bbd090e),
	.w6(32'hbcbad856),
	.w7(32'hbc92deb1),
	.w8(32'hbb96bdcc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe6d8b),
	.w1(32'hbaf690e6),
	.w2(32'h394ffbaa),
	.w3(32'hbbf8d6b3),
	.w4(32'hbbcda20b),
	.w5(32'hbbcc67d7),
	.w6(32'hbc51093f),
	.w7(32'hbbfe0c7f),
	.w8(32'hbbd2b909),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc287a1d),
	.w1(32'hbcd03eec),
	.w2(32'hbcdaa993),
	.w3(32'hbb991ae2),
	.w4(32'hbc65429c),
	.w5(32'hbc273f2d),
	.w6(32'h3bda39ec),
	.w7(32'h3b69ab75),
	.w8(32'h39c500d4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a395680),
	.w1(32'hb9121b99),
	.w2(32'h3ae08e1b),
	.w3(32'h3a983e4f),
	.w4(32'h3b0a333c),
	.w5(32'h3af2143d),
	.w6(32'hba1a8986),
	.w7(32'h3b601531),
	.w8(32'h3a4361c4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af27264),
	.w1(32'hb8e55035),
	.w2(32'h3b1418c2),
	.w3(32'h382488d5),
	.w4(32'h392084ab),
	.w5(32'hb9d80dc1),
	.w6(32'hbad0155c),
	.w7(32'h3a1eee53),
	.w8(32'h3b557cd2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca85329),
	.w1(32'h3c1fbadd),
	.w2(32'hbbe9dd02),
	.w3(32'h3c60572d),
	.w4(32'h3d08d191),
	.w5(32'h3ba3c7d2),
	.w6(32'h3c3a13dc),
	.w7(32'h3cbd274f),
	.w8(32'h3bddd274),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ca4b9),
	.w1(32'hbb1a0b97),
	.w2(32'hbb4cd985),
	.w3(32'hbb7e564e),
	.w4(32'hbc03541e),
	.w5(32'hbb84683c),
	.w6(32'hba22a12a),
	.w7(32'hbb7948c0),
	.w8(32'hbb5781aa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d43cb3),
	.w1(32'hbbe44a4c),
	.w2(32'hbc530c12),
	.w3(32'h3b537f42),
	.w4(32'h3c3e625a),
	.w5(32'h39902d8a),
	.w6(32'h3c0103a8),
	.w7(32'h3c763945),
	.w8(32'h3c509f07),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba666862),
	.w1(32'hbb8fbc14),
	.w2(32'h3a845d74),
	.w3(32'hbb7ec6dd),
	.w4(32'hbb198206),
	.w5(32'hba160689),
	.w6(32'hb9cb4026),
	.w7(32'hb9cdba31),
	.w8(32'hbb4e3d93),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2d2d),
	.w1(32'hbb0ca9d7),
	.w2(32'hbb3ff6ef),
	.w3(32'h3b25c800),
	.w4(32'h3ba9071f),
	.w5(32'h37f85c86),
	.w6(32'hbb80bc01),
	.w7(32'hbb2e79f0),
	.w8(32'h3b175bd6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121b1a),
	.w1(32'h3a8858f3),
	.w2(32'h3b96eca6),
	.w3(32'hbbbfa8cb),
	.w4(32'hbad13ef8),
	.w5(32'hb9ce70d3),
	.w6(32'hbc053f8d),
	.w7(32'hbb9510f9),
	.w8(32'hbbcc9a02),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2dcdc),
	.w1(32'hbbec69d5),
	.w2(32'hbbc925bd),
	.w3(32'hbb322d69),
	.w4(32'hbb8c872d),
	.w5(32'hba0d3fad),
	.w6(32'h3a829d59),
	.w7(32'hb96cf1a8),
	.w8(32'h3b2e74ad),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ee918),
	.w1(32'h3ab0d820),
	.w2(32'h3a770c7c),
	.w3(32'h3ad4ac21),
	.w4(32'h3a51d9b1),
	.w5(32'hbb821a19),
	.w6(32'h3b04cf31),
	.w7(32'h3b09336e),
	.w8(32'hba883ce8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0664),
	.w1(32'hb8cfd461),
	.w2(32'hba00e9c3),
	.w3(32'hbb1786ce),
	.w4(32'hbb295ec1),
	.w5(32'h3b7b16c9),
	.w6(32'hbba4f607),
	.w7(32'hbb366900),
	.w8(32'h3a9fc3f5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ea279),
	.w1(32'hbc369ab8),
	.w2(32'h3c4aa7d9),
	.w3(32'hbc4c0084),
	.w4(32'hbcbb1eb4),
	.w5(32'hba854ff5),
	.w6(32'hbca30f46),
	.w7(32'hbcac838c),
	.w8(32'hb9bca10c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba18cd0),
	.w1(32'hbc6f7311),
	.w2(32'hbce9b207),
	.w3(32'h3c165b23),
	.w4(32'h3b2c5f6c),
	.w5(32'hbc3b6d7a),
	.w6(32'h3ce91285),
	.w7(32'h3c89a3a8),
	.w8(32'hbb3eaf3a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5841e),
	.w1(32'h3adf7b33),
	.w2(32'hbcac9ead),
	.w3(32'h3c272768),
	.w4(32'h3c9a910c),
	.w5(32'hbb24583b),
	.w6(32'h3c6507ef),
	.w7(32'h3c9f83b1),
	.w8(32'h3bd6ae57),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca813),
	.w1(32'hba6fa7aa),
	.w2(32'hbb878593),
	.w3(32'hba1668bd),
	.w4(32'hbb9e533c),
	.w5(32'hb82aef30),
	.w6(32'h3b6bd1b6),
	.w7(32'hbad9e758),
	.w8(32'h3839cb12),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97abe1),
	.w1(32'h3a4d629d),
	.w2(32'hba28b2f0),
	.w3(32'h3b002166),
	.w4(32'h3a0b8a36),
	.w5(32'h3b3b1d83),
	.w6(32'h3adcb600),
	.w7(32'hbaad52ec),
	.w8(32'hba06c970),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba322f5f),
	.w1(32'hba06239f),
	.w2(32'h3afd091c),
	.w3(32'h3ac67ba2),
	.w4(32'h3a878d5f),
	.w5(32'h3aa92e60),
	.w6(32'hbacc66c9),
	.w7(32'h3ade8bc1),
	.w8(32'h3ac641c4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8147),
	.w1(32'hbb7737cb),
	.w2(32'hbb0ee1f9),
	.w3(32'h3af4a5e8),
	.w4(32'h378ff2d1),
	.w5(32'hbbbda0f8),
	.w6(32'h3b4e8d9b),
	.w7(32'h3aae61c8),
	.w8(32'hbb62cd8e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce5ae8b),
	.w1(32'h3c8fa4f3),
	.w2(32'h3c172b09),
	.w3(32'hbb2d8195),
	.w4(32'h3b9ed20b),
	.w5(32'h3c566e79),
	.w6(32'hbc22b8f8),
	.w7(32'hbc02b377),
	.w8(32'h3b11af5f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b2eb),
	.w1(32'hbaf34fbf),
	.w2(32'hba3b4843),
	.w3(32'h3baf4592),
	.w4(32'h3b2b68e8),
	.w5(32'hbbb2437c),
	.w6(32'h3aa8d3ff),
	.w7(32'h3a7f16b1),
	.w8(32'hbbddf8a5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46e34),
	.w1(32'hbb9130c3),
	.w2(32'hb7c2d1e8),
	.w3(32'hbbb0fb49),
	.w4(32'hbc096f15),
	.w5(32'hbb237850),
	.w6(32'hbbe541f7),
	.w7(32'hbbc61193),
	.w8(32'hbc3ea641),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b888354),
	.w1(32'h3acf51aa),
	.w2(32'hbb2c89ad),
	.w3(32'hbae565fc),
	.w4(32'hbac9f217),
	.w5(32'h3b879ed5),
	.w6(32'hbbb88728),
	.w7(32'hbbb7fe7c),
	.w8(32'h399a6d65),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd1a5),
	.w1(32'h3cec7c6e),
	.w2(32'h3cd66940),
	.w3(32'h3be3385f),
	.w4(32'h3cab2c84),
	.w5(32'h3c7e4e95),
	.w6(32'hbc5a2a7d),
	.w7(32'h3723e0f0),
	.w8(32'h3b264f2c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a07f6),
	.w1(32'hbac4488c),
	.w2(32'hbae0a9e1),
	.w3(32'h3a9ba4cd),
	.w4(32'h3a1f9f1c),
	.w5(32'h3b860701),
	.w6(32'h3a9a1618),
	.w7(32'hb8f7dfc5),
	.w8(32'h3ad654e0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84caba),
	.w1(32'h3b8468b4),
	.w2(32'h3bd97977),
	.w3(32'h3bc2e19e),
	.w4(32'h3be184fb),
	.w5(32'h3b8b1dac),
	.w6(32'h3b192e3b),
	.w7(32'h3ba9dccf),
	.w8(32'h3bd32e91),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b82ce),
	.w1(32'hbb8ebb59),
	.w2(32'hbb3f6fd1),
	.w3(32'hbc085318),
	.w4(32'hbbc8e060),
	.w5(32'hbaf42a4c),
	.w6(32'hbbeb24e0),
	.w7(32'hbba340e6),
	.w8(32'hbb330df1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54e6d6),
	.w1(32'h3b187ea1),
	.w2(32'hbad6fdc9),
	.w3(32'hbaa8414c),
	.w4(32'hbb0e8c31),
	.w5(32'hbac9b690),
	.w6(32'hbb686be5),
	.w7(32'hba156854),
	.w8(32'hba888057),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5f4e7),
	.w1(32'hb999c80d),
	.w2(32'h3a0d52e8),
	.w3(32'hbae7806e),
	.w4(32'hba1aa0ee),
	.w5(32'hba94e14f),
	.w6(32'hbb6e909e),
	.w7(32'h39f7668b),
	.w8(32'hbb1e56fa),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c931522),
	.w1(32'h3ce6dd79),
	.w2(32'h3ccef32b),
	.w3(32'h3b5d218f),
	.w4(32'h3bde8104),
	.w5(32'h3c01e354),
	.w6(32'hbc19a168),
	.w7(32'hbbc4e07e),
	.w8(32'hbbbefefe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af934ba),
	.w1(32'h3a2fe1ca),
	.w2(32'hb6a13c57),
	.w3(32'hba450e17),
	.w4(32'hbb0d00ae),
	.w5(32'hbb37d788),
	.w6(32'h39f6dae7),
	.w7(32'hbb358028),
	.w8(32'hba9ec350),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad231a9),
	.w1(32'hbb7abbf5),
	.w2(32'hbb6aaaaf),
	.w3(32'hbb7b7aab),
	.w4(32'hbba1452e),
	.w5(32'hba76ea6c),
	.w6(32'hbb579c20),
	.w7(32'hbb80678c),
	.w8(32'h3a2c3f98),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9061b73),
	.w1(32'hbaa01867),
	.w2(32'hbb225d96),
	.w3(32'h3a01cfd1),
	.w4(32'hba1b7d08),
	.w5(32'hbaee7964),
	.w6(32'hba98cdaa),
	.w7(32'hbb1b51c9),
	.w8(32'hba492653),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900fa79),
	.w1(32'h3b9dd2d1),
	.w2(32'hb98bd915),
	.w3(32'hba8a5eb8),
	.w4(32'hbab16e83),
	.w5(32'h3bd9e753),
	.w6(32'h3b3a3ae8),
	.w7(32'h3a16d514),
	.w8(32'h3b69a968),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a1437),
	.w1(32'h3a092dbe),
	.w2(32'h3bb46a59),
	.w3(32'h3bce42fb),
	.w4(32'h3bef15b2),
	.w5(32'h3b961886),
	.w6(32'h3ac886ca),
	.w7(32'h3bd758da),
	.w8(32'hb9f66eef),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860727),
	.w1(32'hbb5df520),
	.w2(32'h3a80837b),
	.w3(32'h3be5b779),
	.w4(32'h3b149e6d),
	.w5(32'hba5a9aa8),
	.w6(32'hb9899128),
	.w7(32'h3b845c4f),
	.w8(32'h39e539f0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84f8e1),
	.w1(32'h3b8f6dca),
	.w2(32'h3b72d38f),
	.w3(32'hbb5050fd),
	.w4(32'hba46fdaa),
	.w5(32'hbad5be7e),
	.w6(32'hbb7fb322),
	.w7(32'hbb4a41bd),
	.w8(32'hbba79f93),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca61a67),
	.w1(32'h3bce829c),
	.w2(32'hbbe57179),
	.w3(32'h39838cd7),
	.w4(32'h3b9c0127),
	.w5(32'hbbde3d2e),
	.w6(32'h3beb970d),
	.w7(32'h3be9b29e),
	.w8(32'hbb1a3b2d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdbe47),
	.w1(32'h3a0c0079),
	.w2(32'h3aa8d05e),
	.w3(32'hbab33156),
	.w4(32'hbb0ce26f),
	.w5(32'hb9c5df16),
	.w6(32'hbac05fd7),
	.w7(32'h39bb8e53),
	.w8(32'h3a63ed13),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5e062),
	.w1(32'hba032070),
	.w2(32'hba6fff7e),
	.w3(32'hba13ff33),
	.w4(32'hba2ee2ec),
	.w5(32'h3abfe661),
	.w6(32'hba3d418d),
	.w7(32'hbac1c2a2),
	.w8(32'h3b3bf177),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29bf7b),
	.w1(32'hba4e4b4c),
	.w2(32'hba92f322),
	.w3(32'hbb22a601),
	.w4(32'hbb5f9804),
	.w5(32'h3ab0daca),
	.w6(32'hba900941),
	.w7(32'hbb291cda),
	.w8(32'hba8797f4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23b0e3),
	.w1(32'hbb1c56fd),
	.w2(32'hbb8131c3),
	.w3(32'h3afeb1d3),
	.w4(32'h3a0a5406),
	.w5(32'hbb64f2fb),
	.w6(32'hba1f65e7),
	.w7(32'hb9e7c895),
	.w8(32'hbb8da974),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6f8c),
	.w1(32'h3ce34896),
	.w2(32'h3c798671),
	.w3(32'hbb8c32aa),
	.w4(32'h3b986c11),
	.w5(32'h3ba5267c),
	.w6(32'hbc1005f9),
	.w7(32'h3b226baf),
	.w8(32'h3bc3193e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1399cc),
	.w1(32'h3b831173),
	.w2(32'h3c8c669f),
	.w3(32'hbaeaee26),
	.w4(32'h3c243cd9),
	.w5(32'h3bedb7c2),
	.w6(32'hbb876ee8),
	.w7(32'h3b01a522),
	.w8(32'hbb69748b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8adda9),
	.w1(32'h3b3b7461),
	.w2(32'h3a0462a1),
	.w3(32'hbc1d93ea),
	.w4(32'hbb7e1987),
	.w5(32'hbc0223c8),
	.w6(32'hbc25dae0),
	.w7(32'hbb879637),
	.w8(32'hbb717e32),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e88ca),
	.w1(32'hbca71565),
	.w2(32'hbcd6e531),
	.w3(32'hbb01c6f9),
	.w4(32'hbb9a6cb1),
	.w5(32'hbbe6661c),
	.w6(32'h3c2f116c),
	.w7(32'h3bef64fd),
	.w8(32'h39a03ba5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45e2e9),
	.w1(32'hb7f4e986),
	.w2(32'h3b15e369),
	.w3(32'h3a82aaac),
	.w4(32'h3b30e9f6),
	.w5(32'hbb79dba3),
	.w6(32'h3aa65b51),
	.w7(32'h3b570e32),
	.w8(32'hbaa2cda0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5aaf7b),
	.w1(32'h3b8984ea),
	.w2(32'h39a7f2db),
	.w3(32'hbaa275f8),
	.w4(32'h3988e49e),
	.w5(32'hb9a36bc7),
	.w6(32'h38c0767d),
	.w7(32'hbb1b7471),
	.w8(32'h3afd96a3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9dd4),
	.w1(32'h398fab9e),
	.w2(32'hbb16f3d7),
	.w3(32'h3b6c71ad),
	.w4(32'h3b350a76),
	.w5(32'hbaf8b38e),
	.w6(32'hba62e962),
	.w7(32'hbb2618a7),
	.w8(32'hbac605b6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac635da),
	.w1(32'h3b46cdea),
	.w2(32'h3b40a1eb),
	.w3(32'h3875cdf8),
	.w4(32'h3b214198),
	.w5(32'h3b524c83),
	.w6(32'h3b2e37a8),
	.w7(32'h3aa71b63),
	.w8(32'hbad1040c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba635f),
	.w1(32'h3c089888),
	.w2(32'h3b3ba403),
	.w3(32'h3a232222),
	.w4(32'hbb031128),
	.w5(32'h39dbae1f),
	.w6(32'h3b6f5eca),
	.w7(32'h3a7d9938),
	.w8(32'h39a051ed),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2e92a),
	.w1(32'h3c3db486),
	.w2(32'h3bdcaedc),
	.w3(32'h3b560df6),
	.w4(32'h3b8351cf),
	.w5(32'h3ba71db8),
	.w6(32'hbbb52de6),
	.w7(32'hbb700f0d),
	.w8(32'hbb62329c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a34ba),
	.w1(32'h3c17b3ac),
	.w2(32'h3c3914f6),
	.w3(32'hbc4c5b5a),
	.w4(32'hbb2f9b38),
	.w5(32'h3c10c4f3),
	.w6(32'hbc91e740),
	.w7(32'hbab1b0b0),
	.w8(32'h3a9540c6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b742ac6),
	.w1(32'hbbb00895),
	.w2(32'hbba3e2ec),
	.w3(32'h3b276184),
	.w4(32'hb922dd18),
	.w5(32'hbb69a5bf),
	.w6(32'h39957460),
	.w7(32'h39c1a19a),
	.w8(32'hbb299f0d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beae255),
	.w1(32'h3c111b55),
	.w2(32'h3be68ced),
	.w3(32'hbbd4dbf0),
	.w4(32'h3ab0e2f7),
	.w5(32'h399a54e8),
	.w6(32'hbbc21546),
	.w7(32'hba741bc3),
	.w8(32'hb9e3b229),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe12e7),
	.w1(32'h3c437dca),
	.w2(32'h3bbefaef),
	.w3(32'hbab77566),
	.w4(32'h3a9aed55),
	.w5(32'h3ba5d75d),
	.w6(32'hbb45eea7),
	.w7(32'hb90e46e8),
	.w8(32'h3be36ed7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be07904),
	.w1(32'h3b2c9161),
	.w2(32'h3b3a9d56),
	.w3(32'h3ba2a37a),
	.w4(32'h3be489db),
	.w5(32'h39003cf7),
	.w6(32'h3b1546b4),
	.w7(32'h3b886732),
	.w8(32'h3b11f2b8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e2fb),
	.w1(32'h3bbd4554),
	.w2(32'h3bc4aaa1),
	.w3(32'h3a1137fa),
	.w4(32'h3b98b3b9),
	.w5(32'h3bc7c171),
	.w6(32'hbba76a82),
	.w7(32'hbac5de40),
	.w8(32'h3b268768),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c58e0),
	.w1(32'hb9ba1ed8),
	.w2(32'hba043dd3),
	.w3(32'hbb1a2bd0),
	.w4(32'hbaec7bcb),
	.w5(32'h3bdb7d74),
	.w6(32'hbaecbce1),
	.w7(32'hbadc297c),
	.w8(32'h3ba7f54e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30d82),
	.w1(32'h3c2fd379),
	.w2(32'h3bc453f2),
	.w3(32'h3bef52ff),
	.w4(32'h3c057c2a),
	.w5(32'hbabb88b1),
	.w6(32'h3c21fa54),
	.w7(32'h3c02bc36),
	.w8(32'hba9ba06d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45d0b4),
	.w1(32'h39ae0f7e),
	.w2(32'hbacea667),
	.w3(32'hbad4c5e9),
	.w4(32'hb98b71f3),
	.w5(32'hbb42f5f5),
	.w6(32'hb92f0d18),
	.w7(32'hba7827e0),
	.w8(32'hbac27278),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257a30),
	.w1(32'hbbb36c09),
	.w2(32'hbb8dbf36),
	.w3(32'hbb31f534),
	.w4(32'hbb3d250f),
	.w5(32'hb954b154),
	.w6(32'hbb84d819),
	.w7(32'h3aca5b70),
	.w8(32'h3ac43b38),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b185838),
	.w1(32'hbbd1b16f),
	.w2(32'hbb9e2457),
	.w3(32'hbab7111a),
	.w4(32'hbb27fea9),
	.w5(32'hbb6fbdaf),
	.w6(32'h3b7a5374),
	.w7(32'h3a2879f5),
	.w8(32'hbb5da9f9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0667b5),
	.w1(32'hbb859e34),
	.w2(32'hbba585b3),
	.w3(32'hbb1b9087),
	.w4(32'hbb6e42b3),
	.w5(32'h3b10c8a7),
	.w6(32'hba8f4c29),
	.w7(32'hbb2c38d7),
	.w8(32'hba9e65f9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3db0d9),
	.w1(32'hbbe81912),
	.w2(32'hba7cd2c0),
	.w3(32'hb9ffb3e1),
	.w4(32'hbb56ff3e),
	.w5(32'hbb4da513),
	.w6(32'hbba2d7ce),
	.w7(32'hbae8a0ad),
	.w8(32'hbbbca51a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee30e1),
	.w1(32'h3c87887b),
	.w2(32'h3c0e494c),
	.w3(32'hbbcf48c6),
	.w4(32'h3a3e1415),
	.w5(32'h3be50bc6),
	.w6(32'hbc5c03c8),
	.w7(32'hbace6e5b),
	.w8(32'h3af63c04),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38d00e),
	.w1(32'hb99466a6),
	.w2(32'hbbc1f267),
	.w3(32'h3c03cbd6),
	.w4(32'h3be48aed),
	.w5(32'hbb00226c),
	.w6(32'h3ba632be),
	.w7(32'h3ac83b32),
	.w8(32'hbb12ae4d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc54bbb),
	.w1(32'h3c5f306f),
	.w2(32'h3c8a3a7f),
	.w3(32'hbc37732e),
	.w4(32'hbbe56426),
	.w5(32'h3b8bfa33),
	.w6(32'hbc64fe36),
	.w7(32'hbbdd77ed),
	.w8(32'hbb72e8b4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9e2dd),
	.w1(32'hba9a70de),
	.w2(32'hbb106a25),
	.w3(32'hba9c8786),
	.w4(32'h3a5aee31),
	.w5(32'hb97ea37b),
	.w6(32'hbad10708),
	.w7(32'hb848a6f2),
	.w8(32'hbb2e536e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c153d5f),
	.w1(32'h3c2be016),
	.w2(32'h3bc87a88),
	.w3(32'hbc390b67),
	.w4(32'h3b0411fc),
	.w5(32'hba432be2),
	.w6(32'hbc5d5990),
	.w7(32'hbb890100),
	.w8(32'h3a8f203d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad47de5),
	.w1(32'hbaed2821),
	.w2(32'hbb1d2a05),
	.w3(32'hbbb0eb37),
	.w4(32'hbb9b38e2),
	.w5(32'h3bd42b41),
	.w6(32'hbb4c537d),
	.w7(32'hbc00fdc5),
	.w8(32'hbb46dc8d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4d1d),
	.w1(32'hbc09c1b4),
	.w2(32'hbc6622a8),
	.w3(32'h3c20145f),
	.w4(32'h3c2b7243),
	.w5(32'hbb88e55d),
	.w6(32'h3badcdab),
	.w7(32'h3bf6d87b),
	.w8(32'h3991eeb3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba4d56),
	.w1(32'hbac3ce13),
	.w2(32'h3a416311),
	.w3(32'hbb93865f),
	.w4(32'hbb270085),
	.w5(32'h3a319a63),
	.w6(32'hbb4a89ae),
	.w7(32'hbb1ac2b2),
	.w8(32'h3b891619),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc9bcf),
	.w1(32'h3bafe10f),
	.w2(32'h3c05a54b),
	.w3(32'hbbf7d961),
	.w4(32'h3b0f9acf),
	.w5(32'h3c254d28),
	.w6(32'hbc6019b6),
	.w7(32'hbbb634fe),
	.w8(32'h3b82f69e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99201d),
	.w1(32'h3cad9f1b),
	.w2(32'h3c627a32),
	.w3(32'h3c06462a),
	.w4(32'h3a4d9d90),
	.w5(32'hbb28a83e),
	.w6(32'hbad8cf3d),
	.w7(32'hbb1e803d),
	.w8(32'hbbae96be),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a066),
	.w1(32'hbc71be87),
	.w2(32'h38af3177),
	.w3(32'hbb506ead),
	.w4(32'hbc56faf2),
	.w5(32'h3b3d5b5a),
	.w6(32'hbc618b08),
	.w7(32'hbc4a7f85),
	.w8(32'hba165f90),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d8bf1),
	.w1(32'hbc8fd689),
	.w2(32'hbc38d5b1),
	.w3(32'h3c36e20c),
	.w4(32'hbbf9c48a),
	.w5(32'hbbb737e7),
	.w6(32'h3ce3e12c),
	.w7(32'h3c6a066a),
	.w8(32'hbbf3d05a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63bc14),
	.w1(32'hbc6c0ca7),
	.w2(32'hbc2c8890),
	.w3(32'h3b3d2ebe),
	.w4(32'hbb8bd57f),
	.w5(32'hbae22942),
	.w6(32'h3baf430f),
	.w7(32'hbc3b13f1),
	.w8(32'hbb1517c7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1495c0),
	.w1(32'h3c92c63a),
	.w2(32'h3c4c100e),
	.w3(32'h3a3ec21c),
	.w4(32'hbb03994a),
	.w5(32'h3c08c248),
	.w6(32'hbc7a706d),
	.w7(32'hbbc5800e),
	.w8(32'h3b45f70f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b360823),
	.w1(32'h3a8c85c2),
	.w2(32'h3b97b490),
	.w3(32'h3b609d27),
	.w4(32'hbaa535d6),
	.w5(32'h3b19befe),
	.w6(32'h3a531d80),
	.w7(32'hbb01b423),
	.w8(32'h3b473fed),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcacabd),
	.w1(32'h3ba6c0f5),
	.w2(32'h3b7de878),
	.w3(32'h3a93ebe0),
	.w4(32'hbbe85669),
	.w5(32'h3a2b241a),
	.w6(32'hbc39d2eb),
	.w7(32'hbc8bf042),
	.w8(32'hbc8b863b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e4724),
	.w1(32'h3c1ff74e),
	.w2(32'h3c41a012),
	.w3(32'hbb8bc229),
	.w4(32'hba3b724c),
	.w5(32'h3b8093b9),
	.w6(32'hbaf9d0af),
	.w7(32'hbb19faa1),
	.w8(32'hbba8a6af),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92bc05),
	.w1(32'hbb2c75d8),
	.w2(32'hbb2bb4ed),
	.w3(32'h3b777b7e),
	.w4(32'h3b60e443),
	.w5(32'h3b60b14b),
	.w6(32'h3b1e4e5b),
	.w7(32'h3b6a5bb6),
	.w8(32'h3b0c606e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85924a),
	.w1(32'hbc106140),
	.w2(32'hb75cbb30),
	.w3(32'h39888f54),
	.w4(32'hbaa214d1),
	.w5(32'h3b31fd1e),
	.w6(32'h3c937e11),
	.w7(32'h3c6aafd4),
	.w8(32'h3b22ed39),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aec98),
	.w1(32'h3bf6eefe),
	.w2(32'h3bd18c4b),
	.w3(32'hbb39e910),
	.w4(32'h3b4afa5a),
	.w5(32'h3cb27e80),
	.w6(32'hbb2525d3),
	.w7(32'hbb2481bc),
	.w8(32'h3b9c631a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96323c),
	.w1(32'h3bd63147),
	.w2(32'hbac65643),
	.w3(32'h3bddb0fd),
	.w4(32'h3b100ee8),
	.w5(32'hbc280a91),
	.w6(32'h3c142d6f),
	.w7(32'h3be65b5a),
	.w8(32'hbbeef932),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9e536),
	.w1(32'h3c15ac63),
	.w2(32'h3a4028b5),
	.w3(32'hb88dfbe2),
	.w4(32'h3c514570),
	.w5(32'h3b6a760f),
	.w6(32'h3acd0333),
	.w7(32'h3be10f46),
	.w8(32'h3a60ef1c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7be0f5),
	.w1(32'hbaef6eee),
	.w2(32'hbb8e04de),
	.w3(32'h3b94118e),
	.w4(32'hbab89e17),
	.w5(32'h3c023ba1),
	.w6(32'h3c0be2e3),
	.w7(32'h3b1510df),
	.w8(32'h3bd177ec),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c362b),
	.w1(32'hbc3ddffc),
	.w2(32'hbc115240),
	.w3(32'h3a406010),
	.w4(32'hbc088b88),
	.w5(32'hba9b5076),
	.w6(32'hbc1914e7),
	.w7(32'hbc073035),
	.w8(32'hbc3dd18d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2051c),
	.w1(32'h3ba52552),
	.w2(32'h3c00f73c),
	.w3(32'h3c123a6e),
	.w4(32'h3bd19c38),
	.w5(32'h3bf0ffa2),
	.w6(32'hbbc411e7),
	.w7(32'h3aad04a0),
	.w8(32'h3bc3dd59),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9535de),
	.w1(32'hbb1d9f21),
	.w2(32'h3b0c6700),
	.w3(32'hbac0db74),
	.w4(32'hbaa52163),
	.w5(32'hbac5371a),
	.w6(32'hbbf58362),
	.w7(32'hbb984288),
	.w8(32'hbb91b226),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545f67),
	.w1(32'hbb8250b0),
	.w2(32'h3989ed4e),
	.w3(32'h3b8deff6),
	.w4(32'h3b12a988),
	.w5(32'hba85ec5f),
	.w6(32'h3b1f37de),
	.w7(32'hba7b7592),
	.w8(32'h39e87b6d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e2b14),
	.w1(32'h3b153240),
	.w2(32'h3c3e00d4),
	.w3(32'h37b09f7e),
	.w4(32'h3b908b48),
	.w5(32'hbb9262d5),
	.w6(32'hbb662299),
	.w7(32'h3c12d9a8),
	.w8(32'hbbdaf52c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39feff),
	.w1(32'hbb66ec07),
	.w2(32'hbab589c2),
	.w3(32'hbbc8536a),
	.w4(32'hbba9711a),
	.w5(32'h3b7343bb),
	.w6(32'hbc06f6b1),
	.w7(32'hbbb7e7d3),
	.w8(32'hbb16ba37),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fce069),
	.w1(32'hbb6f01ac),
	.w2(32'hbbac21cd),
	.w3(32'hba4740be),
	.w4(32'hbbb1c10b),
	.w5(32'h3b4dabcd),
	.w6(32'hbb758f43),
	.w7(32'hbc000109),
	.w8(32'h3bbe9846),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab289a0),
	.w1(32'hb9a35753),
	.w2(32'h39da1f5f),
	.w3(32'h39fd8693),
	.w4(32'hbb90d074),
	.w5(32'hb9cc8164),
	.w6(32'h3b943103),
	.w7(32'hbb56c162),
	.w8(32'hbbb53c8a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffefa7),
	.w1(32'h3b04adb2),
	.w2(32'h38ee62de),
	.w3(32'h3a99dcca),
	.w4(32'hbb35c1b3),
	.w5(32'hbb2f748c),
	.w6(32'h3b320f93),
	.w7(32'hba92d340),
	.w8(32'hbaf2cc07),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b811173),
	.w1(32'h3b687dae),
	.w2(32'h3addc50e),
	.w3(32'hbb47b682),
	.w4(32'hbb6aa0e6),
	.w5(32'h3b9a4c37),
	.w6(32'hbc81046e),
	.w7(32'hbc104b54),
	.w8(32'h3a48bd66),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99276b),
	.w1(32'hbcbabb85),
	.w2(32'hbcdec313),
	.w3(32'hb909ed6f),
	.w4(32'hbb85c01a),
	.w5(32'hbcac1669),
	.w6(32'h3d0bc0aa),
	.w7(32'h3c95243f),
	.w8(32'hb99bf6a1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea49ab),
	.w1(32'hbb107b9b),
	.w2(32'h398de0bb),
	.w3(32'hbc86396a),
	.w4(32'hbc2b9d28),
	.w5(32'h3a8911c7),
	.w6(32'h3aaaadfe),
	.w7(32'hbc0483e9),
	.w8(32'hba9bded8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3e5d5),
	.w1(32'h3c7f99dc),
	.w2(32'h3aa3a411),
	.w3(32'h3c0a6acf),
	.w4(32'hbaeddb46),
	.w5(32'hbaac8783),
	.w6(32'h3ba6b4ea),
	.w7(32'h3a6883bb),
	.w8(32'hbb0f06eb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90dbb0d),
	.w1(32'h3ae1af60),
	.w2(32'hbb3eec79),
	.w3(32'h3905e518),
	.w4(32'hba9d8054),
	.w5(32'hbbdce6d8),
	.w6(32'hba99b4ae),
	.w7(32'hbb45132e),
	.w8(32'h3be0db9e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814151),
	.w1(32'hbbcc03d1),
	.w2(32'hbb920b90),
	.w3(32'hbc2fb2fe),
	.w4(32'hbb9ac65b),
	.w5(32'hbaccbd75),
	.w6(32'h3c9adf1e),
	.w7(32'h3b87981f),
	.w8(32'h3afa147d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e922e),
	.w1(32'hbba44623),
	.w2(32'h3b8ca543),
	.w3(32'hbb62ee5f),
	.w4(32'hbb6bc47f),
	.w5(32'h3cd5b795),
	.w6(32'hbc04c35c),
	.w7(32'h3abb285a),
	.w8(32'h3c18ad27),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c885926),
	.w1(32'h3ba01dfc),
	.w2(32'h3c338b72),
	.w3(32'h3be84674),
	.w4(32'h3caf65cc),
	.w5(32'hba5efacd),
	.w6(32'hbb375bbc),
	.w7(32'h3aba0394),
	.w8(32'hbc0af16e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05e8dd),
	.w1(32'hbb956992),
	.w2(32'hbb9043b2),
	.w3(32'hba14ca14),
	.w4(32'hbaeb0310),
	.w5(32'h3b4538e0),
	.w6(32'hb9ede284),
	.w7(32'hbbac74f2),
	.w8(32'hba328534),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c59d6),
	.w1(32'h3b3f54ed),
	.w2(32'hbb664182),
	.w3(32'hb8fd644a),
	.w4(32'hbc03d439),
	.w5(32'hbb386643),
	.w6(32'h3b7ba455),
	.w7(32'h3b249977),
	.w8(32'hbb926834),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7107da),
	.w1(32'hbb8a037c),
	.w2(32'hbb01e0bf),
	.w3(32'hbb5c9f05),
	.w4(32'hba5d5648),
	.w5(32'h385394e5),
	.w6(32'hbaf7471f),
	.w7(32'hb9f08a15),
	.w8(32'hbc5153f5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f2e6),
	.w1(32'h3a8377a4),
	.w2(32'h3b6fb40a),
	.w3(32'hbadbd451),
	.w4(32'hbbb1c51a),
	.w5(32'h3b0ed46c),
	.w6(32'hbb19c932),
	.w7(32'hbc32b124),
	.w8(32'hbb38ac8c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dc672),
	.w1(32'hba125fad),
	.w2(32'h3b295d19),
	.w3(32'h3b0cd647),
	.w4(32'h3b63a96d),
	.w5(32'hbbe809bf),
	.w6(32'hb941ec34),
	.w7(32'h3bacb542),
	.w8(32'hb90c5482),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006833),
	.w1(32'h3c577670),
	.w2(32'h3c9725a9),
	.w3(32'hbbb23d98),
	.w4(32'h3b9fe190),
	.w5(32'h3c6d8030),
	.w6(32'hbaa7a463),
	.w7(32'h3b68b7a2),
	.w8(32'h3a7bf695),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70aa75),
	.w1(32'hbc633453),
	.w2(32'hbc014ea0),
	.w3(32'h3c88ba98),
	.w4(32'h3c6ecd40),
	.w5(32'hbaba98da),
	.w6(32'h3b894255),
	.w7(32'hb9c1b30b),
	.w8(32'hba8b6501),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c74c),
	.w1(32'h3b31e09d),
	.w2(32'h3c10974f),
	.w3(32'h3816f2f0),
	.w4(32'h3b0b4c75),
	.w5(32'h3b8943a1),
	.w6(32'hbc7f3cdc),
	.w7(32'h3a59d905),
	.w8(32'h3b11eaa0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77849c),
	.w1(32'h3c4978c1),
	.w2(32'h3c8b75a6),
	.w3(32'hbbb878cb),
	.w4(32'hbb29a2da),
	.w5(32'h3b87e670),
	.w6(32'hbc2e0a61),
	.w7(32'hbbba8de9),
	.w8(32'hbb080b91),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d7fe7),
	.w1(32'hbc90a856),
	.w2(32'hbc158782),
	.w3(32'hbc1cb217),
	.w4(32'hbc51051a),
	.w5(32'hbb102f49),
	.w6(32'hbabc494d),
	.w7(32'h38267c6a),
	.w8(32'hbbb450c6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0427a2),
	.w1(32'h3b7ec755),
	.w2(32'h3b952d8e),
	.w3(32'h3b61b257),
	.w4(32'hbb58c0b3),
	.w5(32'h3be6806a),
	.w6(32'hbb8cdb25),
	.w7(32'h3babb348),
	.w8(32'h3bb1dd59),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec0c25),
	.w1(32'hbb1474ff),
	.w2(32'hba808bc8),
	.w3(32'hbb0a2777),
	.w4(32'h3b02afa4),
	.w5(32'h3a80a356),
	.w6(32'h3a5f07c3),
	.w7(32'hbb8ffdba),
	.w8(32'hb89467ff),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabeea2),
	.w1(32'hbb01d6ae),
	.w2(32'hbc3c38f3),
	.w3(32'h3b8c1bb5),
	.w4(32'h3c62f6eb),
	.w5(32'hbc466552),
	.w6(32'hbb831fac),
	.w7(32'h3bf2fe42),
	.w8(32'hbbf979cb),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbc847),
	.w1(32'hbba8f499),
	.w2(32'hbbb11c8a),
	.w3(32'hbc0a34c6),
	.w4(32'hbbe7a57f),
	.w5(32'hb918d867),
	.w6(32'hbae03677),
	.w7(32'hbba7d17a),
	.w8(32'hbc27da24),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28db86),
	.w1(32'hbb8bcd31),
	.w2(32'hb7721127),
	.w3(32'hbc53e923),
	.w4(32'h39498199),
	.w5(32'hbb129168),
	.w6(32'hbbf0d943),
	.w7(32'hbc31b66b),
	.w8(32'hbb60c6a7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41b931),
	.w1(32'hbbc0995a),
	.w2(32'hbb4eee2c),
	.w3(32'h3925f952),
	.w4(32'h3b658a8b),
	.w5(32'hbb07a349),
	.w6(32'h3c80e236),
	.w7(32'h3bf19fc4),
	.w8(32'hbb443357),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a73b2c),
	.w1(32'h3b4d5909),
	.w2(32'hba20999e),
	.w3(32'hbb070795),
	.w4(32'hbaad1462),
	.w5(32'hbac65d8f),
	.w6(32'hbae4fe77),
	.w7(32'hbad6a524),
	.w8(32'hbbf645a9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf822),
	.w1(32'hbc144f04),
	.w2(32'hbc13e685),
	.w3(32'h3b0f7249),
	.w4(32'hbb2c7849),
	.w5(32'hbbe63518),
	.w6(32'h3ae7d64f),
	.w7(32'hbadcf487),
	.w8(32'hbb9dd430),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006b18),
	.w1(32'h3c532200),
	.w2(32'h3b8d1f6a),
	.w3(32'hb99cc24d),
	.w4(32'h3be7e88c),
	.w5(32'h3c0e1e0f),
	.w6(32'hbc093d37),
	.w7(32'hbb645917),
	.w8(32'hbc3c5303),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f311d),
	.w1(32'hbb9a5931),
	.w2(32'hbb8bdd31),
	.w3(32'hbc8a9fe9),
	.w4(32'hbb103860),
	.w5(32'h3a1e9622),
	.w6(32'hbc8c3bd7),
	.w7(32'hbc744392),
	.w8(32'h3b679158),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987a97),
	.w1(32'h3c8214f8),
	.w2(32'h3c493b13),
	.w3(32'h3b0185d9),
	.w4(32'h3c02844c),
	.w5(32'h3c1ce3a1),
	.w6(32'hbb28f712),
	.w7(32'hbb4b9160),
	.w8(32'hbadbe477),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1750fc),
	.w1(32'h3ad2f321),
	.w2(32'hbb40b75a),
	.w3(32'h3ae223ff),
	.w4(32'hbb6ec49b),
	.w5(32'hbba6d6bf),
	.w6(32'hbbdafda9),
	.w7(32'hbb562bb2),
	.w8(32'hbb8651a7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8685bf),
	.w1(32'hbbc94eff),
	.w2(32'h3c59b474),
	.w3(32'hbc6409e8),
	.w4(32'h3b5e33f7),
	.w5(32'h3b59370a),
	.w6(32'hbc8ef4da),
	.w7(32'hbc2ba7d2),
	.w8(32'hbba85d75),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c145380),
	.w1(32'h3c408dc8),
	.w2(32'hbb2825b8),
	.w3(32'h3bd0ee51),
	.w4(32'h3ca7df27),
	.w5(32'hbbcb6e2d),
	.w6(32'h3c63a406),
	.w7(32'h3c531b31),
	.w8(32'h3bc0ef3b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1134f7),
	.w1(32'hbc150f7d),
	.w2(32'hbc0b37af),
	.w3(32'hbc68eeb3),
	.w4(32'hbc152c90),
	.w5(32'hbb47be2e),
	.w6(32'h3c751e77),
	.w7(32'h3c033605),
	.w8(32'h39e2d71e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6d338),
	.w1(32'hbba55b40),
	.w2(32'hbb30f374),
	.w3(32'hbbc5813f),
	.w4(32'hbb41f61a),
	.w5(32'h3c33fbcb),
	.w6(32'hbae8109b),
	.w7(32'hbb00fd63),
	.w8(32'h3b6b074d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78249a),
	.w1(32'h3c3726b1),
	.w2(32'h3be46090),
	.w3(32'h3bc2ac71),
	.w4(32'h3b0ceb93),
	.w5(32'hbc3ce000),
	.w6(32'h3b61582c),
	.w7(32'h3b62fb15),
	.w8(32'hbbf3b7a2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c9ef),
	.w1(32'h38c82c7e),
	.w2(32'hbb94672a),
	.w3(32'hbbe5bba1),
	.w4(32'hbb2eacb4),
	.w5(32'hbb539e95),
	.w6(32'hbb54844e),
	.w7(32'h3a1ba284),
	.w8(32'hbb5811a5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a60ec),
	.w1(32'hbc64418c),
	.w2(32'hbc0d0a1a),
	.w3(32'hbb8aca91),
	.w4(32'h3b4fe681),
	.w5(32'hbb9a38f6),
	.w6(32'hbb5e5794),
	.w7(32'hbb64060d),
	.w8(32'hbab5f41c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6c7af),
	.w1(32'h3c794cbd),
	.w2(32'h3c3b3bde),
	.w3(32'h3b7876e8),
	.w4(32'h3bc1c4e3),
	.w5(32'h3bb95e0d),
	.w6(32'hbb840b8f),
	.w7(32'hba1731f6),
	.w8(32'h3a90ede6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47080d),
	.w1(32'h3ae59a00),
	.w2(32'h3b814438),
	.w3(32'h3c968cf6),
	.w4(32'h3bab7e89),
	.w5(32'hbb2af3f0),
	.w6(32'h3a820c99),
	.w7(32'h3bf0fa82),
	.w8(32'hbbb28e45),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe01af),
	.w1(32'h3c1e2647),
	.w2(32'h3b94fe56),
	.w3(32'hb9a3cead),
	.w4(32'h3b3d20df),
	.w5(32'h3a345108),
	.w6(32'hbbabd117),
	.w7(32'hbb8041a5),
	.w8(32'hbc314e8b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f66fb),
	.w1(32'h3ae8080a),
	.w2(32'h3a86a13e),
	.w3(32'hbb01b7c1),
	.w4(32'h39b01a05),
	.w5(32'hbb010d84),
	.w6(32'hbb295011),
	.w7(32'hbb86d031),
	.w8(32'hba952100),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4156ec),
	.w1(32'h3a9e7561),
	.w2(32'hbc01e7f2),
	.w3(32'h3ad4b138),
	.w4(32'hbb83c86f),
	.w5(32'hbb3309f1),
	.w6(32'hbb06ae64),
	.w7(32'hbbecd744),
	.w8(32'hbc1f50b8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12f6ba),
	.w1(32'hbab475aa),
	.w2(32'hb98c9fa2),
	.w3(32'h3ad21f0f),
	.w4(32'h3acb4302),
	.w5(32'h3b116e50),
	.w6(32'h3bee843a),
	.w7(32'h3aec5a1b),
	.w8(32'hbbd5c449),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc495730),
	.w1(32'h3babc41d),
	.w2(32'hbb504678),
	.w3(32'hbba8ee24),
	.w4(32'h3b119266),
	.w5(32'h3bebd54f),
	.w6(32'h3a955a6d),
	.w7(32'h3bbda7fb),
	.w8(32'h3bf81bd8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c153235),
	.w1(32'hba795605),
	.w2(32'h3bf74e9f),
	.w3(32'hbc1cfb75),
	.w4(32'hbb93ffd4),
	.w5(32'hbc1a9d37),
	.w6(32'hbc9cf1b0),
	.w7(32'hbb4064a5),
	.w8(32'h3b192af5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51b33b),
	.w1(32'hbb40922a),
	.w2(32'hbb62fba3),
	.w3(32'hbbc8c1f5),
	.w4(32'hbbc204be),
	.w5(32'h3b36a31f),
	.w6(32'h3cd0f4b7),
	.w7(32'h3be4c3a7),
	.w8(32'h3bafc63e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07fb06),
	.w1(32'hbbc5f452),
	.w2(32'hbb6da7e9),
	.w3(32'hbb95733a),
	.w4(32'h3b0aac84),
	.w5(32'h3b35caa0),
	.w6(32'hbaf86e02),
	.w7(32'hbc169c93),
	.w8(32'h3ba266b5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4473a),
	.w1(32'h3c31eb11),
	.w2(32'h3c2d8812),
	.w3(32'h3aba15fb),
	.w4(32'h3a1c5207),
	.w5(32'hbbb16268),
	.w6(32'hbc47c6a0),
	.w7(32'hbbc0cbee),
	.w8(32'hbab41bb0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28751a),
	.w1(32'hbc14f397),
	.w2(32'hbc256caa),
	.w3(32'hbc8a5fb3),
	.w4(32'hbc4b6dba),
	.w5(32'h3c204862),
	.w6(32'h3c630fb1),
	.w7(32'h3a4dac55),
	.w8(32'h3c2b1187),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1110ea),
	.w1(32'h3b0a5a29),
	.w2(32'h3ba65e60),
	.w3(32'h3bbca355),
	.w4(32'h3bc0b288),
	.w5(32'hbb03618c),
	.w6(32'hba31bece),
	.w7(32'h3c81b8ab),
	.w8(32'hba31341d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca3897),
	.w1(32'h3c0833ea),
	.w2(32'h3ac52911),
	.w3(32'h3b2a3458),
	.w4(32'h3b8c8fe4),
	.w5(32'h3b9ab5cd),
	.w6(32'h3bd101c0),
	.w7(32'h3ba53a5f),
	.w8(32'h3c15a194),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd6edf),
	.w1(32'h3cace8fa),
	.w2(32'h3bef1b4d),
	.w3(32'hba9efa51),
	.w4(32'h3b46357c),
	.w5(32'h3b964309),
	.w6(32'h3bd5d77c),
	.w7(32'hbb37ff84),
	.w8(32'h3c1b2c75),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c070906),
	.w1(32'h3b3fd16a),
	.w2(32'h3be03292),
	.w3(32'h3a08d530),
	.w4(32'hb9b41146),
	.w5(32'hbbc8af95),
	.w6(32'h3cf28aba),
	.w7(32'h3c656d3b),
	.w8(32'hbb96c094),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd51728),
	.w1(32'h3b467ad5),
	.w2(32'h3b992842),
	.w3(32'hbc3cd554),
	.w4(32'hbbddc9d7),
	.w5(32'h3b816d31),
	.w6(32'hbc1ca206),
	.w7(32'hbc381c75),
	.w8(32'hbaea6b0e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35ca49),
	.w1(32'h3bc16b98),
	.w2(32'h3beb6e16),
	.w3(32'h3b42aca0),
	.w4(32'h3b8fd78d),
	.w5(32'hbc1fa83b),
	.w6(32'hbbcd5e60),
	.w7(32'h3b3df6bd),
	.w8(32'hb9c5c10e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e574e5),
	.w1(32'hbbc84b40),
	.w2(32'hbbd9510d),
	.w3(32'hbc32655f),
	.w4(32'hbbd357db),
	.w5(32'h3a703c45),
	.w6(32'hbc077e3f),
	.w7(32'hbb842949),
	.w8(32'h3b9c9bc9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e3582),
	.w1(32'h3a5e3164),
	.w2(32'h3b8e792d),
	.w3(32'hbb36cbd8),
	.w4(32'h3aa945cc),
	.w5(32'h3b9ac52e),
	.w6(32'h3b2d041f),
	.w7(32'hbba859ef),
	.w8(32'h394fee3f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a5a03),
	.w1(32'h3bf54f09),
	.w2(32'hba701e6f),
	.w3(32'h3c68afd2),
	.w4(32'h39952afb),
	.w5(32'hbb5ed640),
	.w6(32'h3b42bf24),
	.w7(32'hbacab542),
	.w8(32'hbbbf71d1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded0b2),
	.w1(32'hbb390b42),
	.w2(32'hbb74502c),
	.w3(32'hba6841c1),
	.w4(32'hbb9f746c),
	.w5(32'hb9b2c0cf),
	.w6(32'hbb0915be),
	.w7(32'hb933f0df),
	.w8(32'hbb2032ea),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76092a),
	.w1(32'h3b0b7165),
	.w2(32'h3b4300f3),
	.w3(32'hbb0e3359),
	.w4(32'h3b3471ee),
	.w5(32'h3b529ed4),
	.w6(32'h3acd56b4),
	.w7(32'h3aeb04a7),
	.w8(32'hbb490ee3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82785e),
	.w1(32'hbb7d1110),
	.w2(32'hbba74f6f),
	.w3(32'h386d3cfe),
	.w4(32'hba8e7d16),
	.w5(32'hbb89dcf9),
	.w6(32'h38d39308),
	.w7(32'hbad4d772),
	.w8(32'h3a0e4cd4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1224d),
	.w1(32'h3bd69299),
	.w2(32'h3bc62bcb),
	.w3(32'hbb79dbb1),
	.w4(32'hbaa8c997),
	.w5(32'hbb3d9a2a),
	.w6(32'h3b7c0b3c),
	.w7(32'h3ade8e13),
	.w8(32'hb74bfa23),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b8f56),
	.w1(32'h3aeedb39),
	.w2(32'h3b256f67),
	.w3(32'hbc0c672f),
	.w4(32'hbb5fa0f5),
	.w5(32'h3bb83b46),
	.w6(32'hb9f63232),
	.w7(32'hbab41c25),
	.w8(32'h3b48d8af),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c344c10),
	.w1(32'h3c823590),
	.w2(32'h3c94ea81),
	.w3(32'h39fa2dab),
	.w4(32'hbabdfc2c),
	.w5(32'h3b68c854),
	.w6(32'hbc099d8d),
	.w7(32'hb9b61e9a),
	.w8(32'h3c7a3ed9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7486f8),
	.w1(32'hba8c2b78),
	.w2(32'h3c047ebe),
	.w3(32'h39c9fb4b),
	.w4(32'h3ae88ff9),
	.w5(32'hbb386daa),
	.w6(32'h3a328e0b),
	.w7(32'hbb080500),
	.w8(32'hbbc0dd76),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7f287),
	.w1(32'hba4d275a),
	.w2(32'h3ad5d315),
	.w3(32'hbb8f058b),
	.w4(32'hbadc68b1),
	.w5(32'hbbb3a7a5),
	.w6(32'hbab46c43),
	.w7(32'h3a6c07fc),
	.w8(32'hbb57fd08),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68461d),
	.w1(32'h3d1d167e),
	.w2(32'h3c86b1e8),
	.w3(32'hba5548ee),
	.w4(32'hbb0d07fa),
	.w5(32'hbbaf8873),
	.w6(32'hbb132d93),
	.w7(32'hba956148),
	.w8(32'hbb5a1cb6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a18b7),
	.w1(32'h3c6862e4),
	.w2(32'hbb17ea76),
	.w3(32'hbbcefa59),
	.w4(32'h3c2c071e),
	.w5(32'h3958ebc8),
	.w6(32'h3ca695d4),
	.w7(32'h3c435619),
	.w8(32'h3be83088),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33cd64),
	.w1(32'h3998277e),
	.w2(32'h3bb4e138),
	.w3(32'hbc73ccc0),
	.w4(32'h3a6b0d19),
	.w5(32'h3ba8ea22),
	.w6(32'h3ccff0ff),
	.w7(32'h3c087e71),
	.w8(32'hbb60b850),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7dcc5),
	.w1(32'hbb2edbc2),
	.w2(32'hbb126f32),
	.w3(32'h3a62211c),
	.w4(32'hbabfdc33),
	.w5(32'hba0a1c62),
	.w6(32'h3a2fbeae),
	.w7(32'hbb94ba49),
	.w8(32'hba8fdb79),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b1124),
	.w1(32'h3b14813f),
	.w2(32'hb9e8dd0c),
	.w3(32'hba4a2173),
	.w4(32'hbb09ac8c),
	.w5(32'hbbbe2927),
	.w6(32'hbb18bca7),
	.w7(32'hbb2bd15f),
	.w8(32'hbab07bdc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c06c),
	.w1(32'h3be40430),
	.w2(32'h3bfbbc46),
	.w3(32'hbb5ca5a3),
	.w4(32'h3a89def7),
	.w5(32'hbb6c5d55),
	.w6(32'hba01e3cc),
	.w7(32'h3b87db43),
	.w8(32'hbbb228ac),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99fdc3),
	.w1(32'h3ad3851a),
	.w2(32'h3b67cfef),
	.w3(32'hbbd43a5a),
	.w4(32'hbbdf43ec),
	.w5(32'h3c04331e),
	.w6(32'hbb7b1347),
	.w7(32'hbbf14f46),
	.w8(32'h3bb0eb31),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62ef11),
	.w1(32'hbb842787),
	.w2(32'hbbb89df6),
	.w3(32'h3b557182),
	.w4(32'h3c48a075),
	.w5(32'hbb88c745),
	.w6(32'h3b26b71a),
	.w7(32'h3b8d8ce6),
	.w8(32'h3b3929b3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18fa96),
	.w1(32'hbc3c7b70),
	.w2(32'hbca336cc),
	.w3(32'h3b878707),
	.w4(32'hbc0da4a3),
	.w5(32'hbbff5195),
	.w6(32'hb8a5e2ba),
	.w7(32'h3c06b629),
	.w8(32'hbbb2def3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b651c),
	.w1(32'hba03e442),
	.w2(32'h393ac721),
	.w3(32'h3ae0fb81),
	.w4(32'hbb94a06f),
	.w5(32'hbaf92aa6),
	.w6(32'hbb3cc351),
	.w7(32'hba1d6136),
	.w8(32'h3a9578b4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69d0ef),
	.w1(32'h3b804018),
	.w2(32'h3c3c535c),
	.w3(32'hbb97a5d0),
	.w4(32'h39467cc2),
	.w5(32'h3c0e6453),
	.w6(32'hbc13e970),
	.w7(32'hbb5b134f),
	.w8(32'h3afd75f5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a4d11),
	.w1(32'hba15277e),
	.w2(32'h3b53e318),
	.w3(32'h3b67ff54),
	.w4(32'h3b1730ee),
	.w5(32'h3b8375d8),
	.w6(32'h3b766d5c),
	.w7(32'h3b292041),
	.w8(32'hbc041e49),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba690df),
	.w1(32'hbc71177e),
	.w2(32'hbb9dce4c),
	.w3(32'hb9c4bd2c),
	.w4(32'h3c1e3e57),
	.w5(32'hbbc62025),
	.w6(32'h3ba4130d),
	.w7(32'hbbe111ab),
	.w8(32'h3adf54d3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a7807),
	.w1(32'hbab978b8),
	.w2(32'h3a7ab22b),
	.w3(32'hbc07d337),
	.w4(32'hba5c4d1c),
	.w5(32'h3bebd8d5),
	.w6(32'h3cfae29f),
	.w7(32'h3c5050f5),
	.w8(32'hbb58ef19),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a717625),
	.w1(32'h3b30f0c9),
	.w2(32'h3b4c50b5),
	.w3(32'hbb41d3ea),
	.w4(32'h3a487755),
	.w5(32'h3bf6230f),
	.w6(32'hbae1cb65),
	.w7(32'hbb449e5d),
	.w8(32'h3c24214a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0295f),
	.w1(32'hbadbe15f),
	.w2(32'hbb59b11b),
	.w3(32'hbbc4a403),
	.w4(32'hb91093ce),
	.w5(32'h3af8a513),
	.w6(32'hbc0b6d22),
	.w7(32'h3b8eeec2),
	.w8(32'h3a26a1fa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18f98c),
	.w1(32'hbb211c3a),
	.w2(32'hbb9a77fe),
	.w3(32'hba46cc9e),
	.w4(32'h3b1422ce),
	.w5(32'hbb2d8fab),
	.w6(32'h3b820a15),
	.w7(32'h3c3fc867),
	.w8(32'hba5c9d1e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88b160),
	.w1(32'hbb04e580),
	.w2(32'hbbb86616),
	.w3(32'h3aed9173),
	.w4(32'hba7f8c9f),
	.w5(32'hbb488693),
	.w6(32'h3a633bb1),
	.w7(32'hbad3a01b),
	.w8(32'hbbe35881),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5227c6),
	.w1(32'hbb91882e),
	.w2(32'hbb311a73),
	.w3(32'hbb968279),
	.w4(32'hbbec8d53),
	.w5(32'hbaff4864),
	.w6(32'h3a217afd),
	.w7(32'hbbd6b800),
	.w8(32'hbbd42a52),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb206),
	.w1(32'hbc6009f8),
	.w2(32'hbc00edac),
	.w3(32'h3b0fa521),
	.w4(32'hb9a31c42),
	.w5(32'h3b028e07),
	.w6(32'hba9ea18a),
	.w7(32'hbb0389cc),
	.w8(32'hbb07396f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27bb41),
	.w1(32'h3b9dbbaa),
	.w2(32'h3b84e86b),
	.w3(32'h3b50faa4),
	.w4(32'h3bc2de50),
	.w5(32'h3be099d2),
	.w6(32'h3c372e6e),
	.w7(32'h3badfb38),
	.w8(32'hbc03965e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4f455),
	.w1(32'h3b8c0d95),
	.w2(32'h3c581555),
	.w3(32'h3bd9bcf2),
	.w4(32'h3c721a9b),
	.w5(32'hba78a2ea),
	.w6(32'hbd0efbba),
	.w7(32'hbc15a24d),
	.w8(32'h3910ca64),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eaea7),
	.w1(32'h39d4d4e9),
	.w2(32'hb988edbf),
	.w3(32'hbb756899),
	.w4(32'hba4735f0),
	.w5(32'h38542ad2),
	.w6(32'h3b7f770d),
	.w7(32'h3b10dd26),
	.w8(32'h3b958707),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd781),
	.w1(32'hbc0c387c),
	.w2(32'hbba27950),
	.w3(32'h3be030ea),
	.w4(32'h3b8f1ed3),
	.w5(32'hbc0f703b),
	.w6(32'h3b31d053),
	.w7(32'hbab6a66a),
	.w8(32'hbbf643bc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96f488),
	.w1(32'hbb6d386f),
	.w2(32'h3adbb306),
	.w3(32'hbbb0a99c),
	.w4(32'hbb30a5f2),
	.w5(32'h3bc42dd5),
	.w6(32'hbc0b4b6f),
	.w7(32'hbaba56e0),
	.w8(32'hbb7d047b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3a21e),
	.w1(32'h3b5dac1e),
	.w2(32'h3c057e63),
	.w3(32'hbb3809c3),
	.w4(32'h3a3bbf89),
	.w5(32'hbb02c446),
	.w6(32'hbc180746),
	.w7(32'hbb4763e8),
	.w8(32'h3b814b23),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a8ff),
	.w1(32'hbb4e8614),
	.w2(32'hbbc305ba),
	.w3(32'hbb5e45fa),
	.w4(32'hbc3c2b83),
	.w5(32'hbbf88f6d),
	.w6(32'h3c879e50),
	.w7(32'h3c4489df),
	.w8(32'hbb90a15c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9caa449),
	.w1(32'h3b35d9e8),
	.w2(32'h3974788e),
	.w3(32'hbb963065),
	.w4(32'hbbf7e7b0),
	.w5(32'h3af9ef54),
	.w6(32'h3b01b8ce),
	.w7(32'hbbc0a594),
	.w8(32'hbb8cf2e5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b849c),
	.w1(32'hbb3c2183),
	.w2(32'hbb4733e4),
	.w3(32'h3aaf49f5),
	.w4(32'h3ba25dab),
	.w5(32'hb98eee9c),
	.w6(32'hbb76277d),
	.w7(32'hbb11e8ca),
	.w8(32'h3acdb6c6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1afea0),
	.w1(32'h3b3b89dd),
	.w2(32'h3baa1062),
	.w3(32'h3a8c68be),
	.w4(32'h3bc82451),
	.w5(32'h3bbce34e),
	.w6(32'h3b23abaf),
	.w7(32'h3b922330),
	.w8(32'hbbd5da8f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f4381),
	.w1(32'hbc79b2d8),
	.w2(32'h3c92866d),
	.w3(32'h3bb94cca),
	.w4(32'hb98c3c2e),
	.w5(32'h3c0fbcde),
	.w6(32'hbc6c9a99),
	.w7(32'h3bd4e56e),
	.w8(32'hbbc4e8df),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c525776),
	.w1(32'h3b22e8b2),
	.w2(32'h3a9d39f1),
	.w3(32'hbc392c1a),
	.w4(32'h3b5d3367),
	.w5(32'hbaaa78b4),
	.w6(32'hbcdd2cd4),
	.w7(32'hbc0ba4d4),
	.w8(32'hbb7dccf1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5861),
	.w1(32'h3b763bcc),
	.w2(32'h3c09ca6e),
	.w3(32'hbc09ad56),
	.w4(32'hbad7bce8),
	.w5(32'h3c078141),
	.w6(32'hbc8be057),
	.w7(32'hbc415817),
	.w8(32'hbc06687a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c600),
	.w1(32'hbc096be1),
	.w2(32'hbc1d608e),
	.w3(32'h3c0b8038),
	.w4(32'h3b68cfdf),
	.w5(32'hbb9f3aef),
	.w6(32'h3c0bd34d),
	.w7(32'hb98295e5),
	.w8(32'hbb44675f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5a4cb),
	.w1(32'hbb99550a),
	.w2(32'hbcae40c2),
	.w3(32'h3c119001),
	.w4(32'h3b1194b9),
	.w5(32'h3bb98e5d),
	.w6(32'h3c00efcb),
	.w7(32'h385698dc),
	.w8(32'h3b4fc8d9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f9cb5),
	.w1(32'hbb7e5156),
	.w2(32'h3b2c78db),
	.w3(32'hbbb5dad5),
	.w4(32'h3bd784c3),
	.w5(32'h39607c66),
	.w6(32'hbc47bcd3),
	.w7(32'hbadc1c89),
	.w8(32'h3b6ee833),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c235825),
	.w1(32'h3bdc6878),
	.w2(32'hbb0dac6c),
	.w3(32'hb9cab082),
	.w4(32'hbbcf1855),
	.w5(32'hbbc2c480),
	.w6(32'hbb581170),
	.w7(32'h3c7bbbf8),
	.w8(32'hbbb421fa),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4580f),
	.w1(32'h3bdbdfdd),
	.w2(32'h3b1891c5),
	.w3(32'h3b84b2df),
	.w4(32'h39d0cd22),
	.w5(32'h3b047abd),
	.w6(32'h3ae9a724),
	.w7(32'hbb79ecaf),
	.w8(32'hbb5ef294),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a91ab),
	.w1(32'h3b18067d),
	.w2(32'h3c02ab5f),
	.w3(32'h3bf17547),
	.w4(32'h3c1fdf80),
	.w5(32'hba5c74ca),
	.w6(32'hbbc61210),
	.w7(32'h3b7cdcd3),
	.w8(32'hba8ce19f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b893137),
	.w1(32'h3bb6689f),
	.w2(32'h3b5e596a),
	.w3(32'hba4c8faf),
	.w4(32'h3af00915),
	.w5(32'h3c2b4d4b),
	.w6(32'hbb90a37a),
	.w7(32'hbaefc8dc),
	.w8(32'h3b394f80),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03d063),
	.w1(32'hba410a93),
	.w2(32'hb89ad6c7),
	.w3(32'hbb90cf48),
	.w4(32'hbb60c2f3),
	.w5(32'hba8c89d7),
	.w6(32'hbc352467),
	.w7(32'hbbc08696),
	.w8(32'h39afe12e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f64d8),
	.w1(32'hba599c5f),
	.w2(32'h3b51a1e3),
	.w3(32'hbb690330),
	.w4(32'h3ae3919a),
	.w5(32'hbc40ba1c),
	.w6(32'hbbad2bdd),
	.w7(32'h3ba0dda6),
	.w8(32'hbc4fe47d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1a30),
	.w1(32'hbc0a7a19),
	.w2(32'hbc30e924),
	.w3(32'hbbe7c411),
	.w4(32'hbc37a36d),
	.w5(32'h3a8fb874),
	.w6(32'hbbe8d9ff),
	.w7(32'hbc840985),
	.w8(32'hbb39e9dc),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c3f1c),
	.w1(32'h3bda9cf0),
	.w2(32'h3b85dbdf),
	.w3(32'hbc920c49),
	.w4(32'h3bd456f7),
	.w5(32'h3b1bc8bf),
	.w6(32'hbcb3dd8b),
	.w7(32'hbb5008fb),
	.w8(32'hbb73e7cb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a696834),
	.w1(32'h3b123f32),
	.w2(32'h3a33fb19),
	.w3(32'hb899b0e8),
	.w4(32'h39d0a96e),
	.w5(32'h3c106a8a),
	.w6(32'hbbe4a5d8),
	.w7(32'hbb83f5f0),
	.w8(32'h3aa2771e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a436),
	.w1(32'hb99aedb7),
	.w2(32'hbaedc484),
	.w3(32'h3ac95107),
	.w4(32'hba924271),
	.w5(32'hbb070921),
	.w6(32'h3b60a8c0),
	.w7(32'h3b8fd070),
	.w8(32'hbbc4b7b2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b5706),
	.w1(32'h3c0baf99),
	.w2(32'h3c14df0d),
	.w3(32'hbb69405e),
	.w4(32'h3bc75b8f),
	.w5(32'h3ba923ea),
	.w6(32'hbc0bf6ca),
	.w7(32'hb95a841e),
	.w8(32'h3b739f62),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba342017),
	.w1(32'hbbf780f4),
	.w2(32'hbc052b5c),
	.w3(32'hbc0cb338),
	.w4(32'hbb9011e2),
	.w5(32'h3b61131e),
	.w6(32'hbb9c402f),
	.w7(32'hba895a93),
	.w8(32'h3ba9adf7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4cf64),
	.w1(32'hbc05d5c7),
	.w2(32'h39210149),
	.w3(32'hbbf48faf),
	.w4(32'hba148b71),
	.w5(32'hbb0220f5),
	.w6(32'hbbbe4ffb),
	.w7(32'hb912acec),
	.w8(32'hba1112bc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb916ec),
	.w1(32'h3b2692d0),
	.w2(32'hbb55be8b),
	.w3(32'hbb44fbb5),
	.w4(32'hba38d698),
	.w5(32'h3a113a1a),
	.w6(32'hbbdb32df),
	.w7(32'hbb947d69),
	.w8(32'hbb187720),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a113cc),
	.w1(32'h3a8acec8),
	.w2(32'hba493f50),
	.w3(32'h3abdb222),
	.w4(32'h3a4a0b0f),
	.w5(32'h395e01d8),
	.w6(32'hbae6f60b),
	.w7(32'hb8c05764),
	.w8(32'hba4341c5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2a36d),
	.w1(32'hbb22aba3),
	.w2(32'hbc016976),
	.w3(32'h3a9307af),
	.w4(32'hbb710b3e),
	.w5(32'hbb1500ba),
	.w6(32'h3b0577a2),
	.w7(32'hbae044fb),
	.w8(32'h3bbacaa0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3ee9a),
	.w1(32'h3c4907d7),
	.w2(32'h3c64c62c),
	.w3(32'h3c1a59ce),
	.w4(32'h3ca04ee1),
	.w5(32'h3c064077),
	.w6(32'hbc89c0d0),
	.w7(32'h3bd11733),
	.w8(32'h3b382a4e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09b923),
	.w1(32'h3c2fcc99),
	.w2(32'h3c027146),
	.w3(32'hbba59fd4),
	.w4(32'h3aa67a68),
	.w5(32'h3b9fe6b5),
	.w6(32'hbc56ec05),
	.w7(32'hbbb9ed59),
	.w8(32'h3c857f54),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d14236c),
	.w1(32'h3cb8e9bb),
	.w2(32'h3c920f54),
	.w3(32'hba9f7080),
	.w4(32'h3c4d5e1e),
	.w5(32'hb8a92204),
	.w6(32'h3b60b123),
	.w7(32'h3c9e9398),
	.w8(32'hbadd6dc2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59559c),
	.w1(32'h3b150471),
	.w2(32'hbb139097),
	.w3(32'hbb037ac4),
	.w4(32'hbaabedcc),
	.w5(32'hbaea9763),
	.w6(32'hb9e289f4),
	.w7(32'hbaa8c463),
	.w8(32'hbb50f2e1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00d0b),
	.w1(32'hbb01688d),
	.w2(32'hbb2f24f1),
	.w3(32'h3b81a760),
	.w4(32'h3b76397c),
	.w5(32'h3a65b5e6),
	.w6(32'hbc0ca17d),
	.w7(32'hbbc21b22),
	.w8(32'h3a87cb3b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba909283),
	.w1(32'hba26e962),
	.w2(32'h395917af),
	.w3(32'hba2024b9),
	.w4(32'h3b0e9d80),
	.w5(32'h3b634e32),
	.w6(32'h3ac2c81f),
	.w7(32'h3b0874c2),
	.w8(32'hbab85c8f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39950cad),
	.w1(32'h3a7f07eb),
	.w2(32'h3ba47943),
	.w3(32'h3c126199),
	.w4(32'hba093236),
	.w5(32'h3aa8cae4),
	.w6(32'h3c152dce),
	.w7(32'h3ba0aeb5),
	.w8(32'h3b073e91),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3df2),
	.w1(32'h3c0a9944),
	.w2(32'h3c1b0a6c),
	.w3(32'hbbb5567d),
	.w4(32'hbab4a336),
	.w5(32'h3b289fe6),
	.w6(32'hbb928603),
	.w7(32'hba68b865),
	.w8(32'hbb990789),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc267c9),
	.w1(32'h3b5d8159),
	.w2(32'hbb4e9fca),
	.w3(32'h394a9a81),
	.w4(32'h3b9cadc8),
	.w5(32'hbb068863),
	.w6(32'hbbcaada0),
	.w7(32'hbbb022be),
	.w8(32'hbb16e00c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39b4a7),
	.w1(32'hbc03c9bc),
	.w2(32'h3a0d7517),
	.w3(32'hbb9c14ef),
	.w4(32'h3c368e27),
	.w5(32'h3aad71eb),
	.w6(32'hbc22a961),
	.w7(32'h3b07eb6b),
	.w8(32'hba6bbe5c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b887ce6),
	.w1(32'h3a908f5b),
	.w2(32'h3bf9f050),
	.w3(32'h3beea617),
	.w4(32'hb9ffbfa5),
	.w5(32'hb80e86d4),
	.w6(32'h3c049db2),
	.w7(32'h3bd1e46f),
	.w8(32'hbb864907),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a439),
	.w1(32'hbaa53320),
	.w2(32'hba88c1f0),
	.w3(32'h3a9756e6),
	.w4(32'h3ae1e7ab),
	.w5(32'hba647a0d),
	.w6(32'h3b9508cd),
	.w7(32'hbb23632d),
	.w8(32'h3b028fec),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5afae),
	.w1(32'h3bd147e8),
	.w2(32'h3b6c0896),
	.w3(32'hbb81cc38),
	.w4(32'hbb04f123),
	.w5(32'hbab33e88),
	.w6(32'h3c356044),
	.w7(32'h3aa21cea),
	.w8(32'hbb3a11b9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926c5d),
	.w1(32'h3b565614),
	.w2(32'hbac534d0),
	.w3(32'hbb081b57),
	.w4(32'hbb9ea6c6),
	.w5(32'hba2ada7c),
	.w6(32'hbb71f6f8),
	.w7(32'hbba72ffe),
	.w8(32'h3c8520a8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d161276),
	.w1(32'h3cb3d276),
	.w2(32'h3bb7b456),
	.w3(32'h3c92176a),
	.w4(32'h3cde013b),
	.w5(32'h39613878),
	.w6(32'h3b23b61b),
	.w7(32'h3cc92c3c),
	.w8(32'hbb8906ef),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a298cfb),
	.w1(32'hbb221c44),
	.w2(32'hbb790b29),
	.w3(32'hb98d625f),
	.w4(32'h395d3364),
	.w5(32'h3a80eb4e),
	.w6(32'hbb0e410e),
	.w7(32'h3a0bb5b2),
	.w8(32'h3c8aecb0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951789),
	.w1(32'h3bd2eb1f),
	.w2(32'hbb2db3a7),
	.w3(32'hbb714d5c),
	.w4(32'hbc432dc2),
	.w5(32'hbbcabdc3),
	.w6(32'hbb40c525),
	.w7(32'hbc3e8fe5),
	.w8(32'hbc7ce7c6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule