module layer_8_featuremap_30(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ab8a),
	.w1(32'hb88df0e2),
	.w2(32'hb9fac4d1),
	.w3(32'hba24fc23),
	.w4(32'hb9b5d9df),
	.w5(32'hba54a953),
	.w6(32'h396113d2),
	.w7(32'hb9a3cc76),
	.w8(32'hb988d789),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2f95f),
	.w1(32'h37e4dc59),
	.w2(32'hb9e9d59e),
	.w3(32'hb92fbdf8),
	.w4(32'hb8fa37ae),
	.w5(32'hba098954),
	.w6(32'h38969b2c),
	.w7(32'hb9b5eabf),
	.w8(32'hba0020c0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba468bc2),
	.w1(32'hb98390da),
	.w2(32'hb9b4df7d),
	.w3(32'hba06f7e5),
	.w4(32'hb99a8d57),
	.w5(32'hba00ec93),
	.w6(32'hb8a87bf5),
	.w7(32'hb92463e2),
	.w8(32'h3aa2697b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37bdcd),
	.w1(32'hba76b60a),
	.w2(32'hba925cca),
	.w3(32'hbaeb1703),
	.w4(32'hbb702c55),
	.w5(32'hbb1d0d46),
	.w6(32'hb9d7a05c),
	.w7(32'hba8cd21a),
	.w8(32'hba1664d6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b2df1),
	.w1(32'hb900cf17),
	.w2(32'hb919170b),
	.w3(32'hb9e697d2),
	.w4(32'hb985bd45),
	.w5(32'hb8bdcad5),
	.w6(32'h3944ca1d),
	.w7(32'h38ddbcc5),
	.w8(32'h388a9542),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a19d15),
	.w1(32'h39aed4f2),
	.w2(32'hbb00cb48),
	.w3(32'h3a51a424),
	.w4(32'hb73ebe49),
	.w5(32'hbb0553da),
	.w6(32'h3a17b342),
	.w7(32'hbab4ae76),
	.w8(32'hba625889),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d41e6),
	.w1(32'hba095185),
	.w2(32'hba3ac4e6),
	.w3(32'hba4458e9),
	.w4(32'hba1eb422),
	.w5(32'hba558b00),
	.w6(32'h384b875c),
	.w7(32'hba1a4560),
	.w8(32'hba56aef7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bb556),
	.w1(32'hb9bbe336),
	.w2(32'hb98e2ef0),
	.w3(32'hba1f728a),
	.w4(32'hba1a6bd1),
	.w5(32'hb9225469),
	.w6(32'h39559057),
	.w7(32'hb8825e68),
	.w8(32'hba9a119d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fd739),
	.w1(32'hba168d5d),
	.w2(32'hba9e6fa4),
	.w3(32'hba6f787e),
	.w4(32'hba604200),
	.w5(32'hbaafc63a),
	.w6(32'hb954d827),
	.w7(32'hba72fa74),
	.w8(32'h39f84b30),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7238b3),
	.w1(32'hbae8b7f5),
	.w2(32'hbabf3d31),
	.w3(32'hba842653),
	.w4(32'hbbc3c1ce),
	.w5(32'hbaf9c9df),
	.w6(32'h3a96cad1),
	.w7(32'hbac480b9),
	.w8(32'hba5bf104),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c76d1),
	.w1(32'hb9b9e108),
	.w2(32'hba06057e),
	.w3(32'hbab7da66),
	.w4(32'hba76d62a),
	.w5(32'hb9e639a2),
	.w6(32'h395617b3),
	.w7(32'hb930f6f7),
	.w8(32'hba74cf31),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f2316),
	.w1(32'hb98bf84e),
	.w2(32'hb986d7f7),
	.w3(32'hba2c65a1),
	.w4(32'hb9b771a6),
	.w5(32'hba15deb0),
	.w6(32'hb86d62f7),
	.w7(32'hb98f4a1b),
	.w8(32'hba6faf8a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73e28a),
	.w1(32'hba168fed),
	.w2(32'hba6e6ed3),
	.w3(32'hba6bccc8),
	.w4(32'hba290079),
	.w5(32'hba295286),
	.w6(32'hb90a1ddf),
	.w7(32'hba27393a),
	.w8(32'hb801cf31),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b342e),
	.w1(32'h39afd6d8),
	.w2(32'hbb14356b),
	.w3(32'h3a8e765d),
	.w4(32'h3984e9de),
	.w5(32'hbb0bc1e6),
	.w6(32'h3a235951),
	.w7(32'hbadd2a05),
	.w8(32'hb9827ed3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9050719),
	.w1(32'h3965a01e),
	.w2(32'hba2f9a63),
	.w3(32'h38cacc80),
	.w4(32'hb92ef977),
	.w5(32'hba8af53e),
	.w6(32'h3a3c828e),
	.w7(32'hb8d58007),
	.w8(32'h39b7c471),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c093d6),
	.w1(32'hb941f831),
	.w2(32'h392b19cb),
	.w3(32'h393e1432),
	.w4(32'h38ec5036),
	.w5(32'hb9106bd0),
	.w6(32'hb985db82),
	.w7(32'hb9fb3aaa),
	.w8(32'h39659295),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32e6d5),
	.w1(32'hbb86cd88),
	.w2(32'hbba08750),
	.w3(32'h3b869585),
	.w4(32'hb9cc5bd1),
	.w5(32'hbbaaf257),
	.w6(32'hbb17e74e),
	.w7(32'hbb27f191),
	.w8(32'hba90ab9d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e88c5),
	.w1(32'hb6f7d4da),
	.w2(32'hb9b8dd4b),
	.w3(32'hba73ce04),
	.w4(32'h39364275),
	.w5(32'hb98ac109),
	.w6(32'h39d693bb),
	.w7(32'h3968526d),
	.w8(32'hba892fcb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba388888),
	.w1(32'h3a50e6cc),
	.w2(32'h3a1032b4),
	.w3(32'hb9d3ed37),
	.w4(32'h39a32a73),
	.w5(32'h3a738a4f),
	.w6(32'h3a0834ac),
	.w7(32'h39890539),
	.w8(32'hbafbe8fd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35c57b),
	.w1(32'hb9b6da0d),
	.w2(32'hba93f7d7),
	.w3(32'h3aed7e09),
	.w4(32'h3b6e67be),
	.w5(32'h3ab659fe),
	.w6(32'hbbaecdf6),
	.w7(32'hbb924f8e),
	.w8(32'hbad032c4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba956f9d),
	.w1(32'hb8532322),
	.w2(32'h39e60258),
	.w3(32'hba9e9060),
	.w4(32'hb94d55f5),
	.w5(32'h39f95f1c),
	.w6(32'hb933a454),
	.w7(32'h39472437),
	.w8(32'hb9e3c021),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ab607),
	.w1(32'h38125572),
	.w2(32'h393c7f27),
	.w3(32'h387a519a),
	.w4(32'hb91517cb),
	.w5(32'hb80f4335),
	.w6(32'h3a78149d),
	.w7(32'h3a3ffbb6),
	.w8(32'hba915d81),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba222e8c),
	.w1(32'hba56d772),
	.w2(32'h3a36e407),
	.w3(32'h3a7cc944),
	.w4(32'h3b0708c6),
	.w5(32'h3b243715),
	.w6(32'hba76d7d1),
	.w7(32'hb9ed40b4),
	.w8(32'hbacad345),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e2812),
	.w1(32'h3903eb0a),
	.w2(32'hba05b349),
	.w3(32'hba867323),
	.w4(32'h398a0aee),
	.w5(32'hb9c6fe9f),
	.w6(32'h3a07b859),
	.w7(32'hb958151b),
	.w8(32'h3a5dc602),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78c1a7),
	.w1(32'h3a9c002d),
	.w2(32'hb9e73c5b),
	.w3(32'h3accb44d),
	.w4(32'h397449d3),
	.w5(32'h3a1b5cfd),
	.w6(32'h3a0545d9),
	.w7(32'hba417c7a),
	.w8(32'hba40a515),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa07c9),
	.w1(32'hba113c84),
	.w2(32'h3a4c41e8),
	.w3(32'h3a75d84e),
	.w4(32'h3b06c4de),
	.w5(32'h3b25392a),
	.w6(32'hba68aa1b),
	.w7(32'hb99523a3),
	.w8(32'hba4135b5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e777f7),
	.w1(32'hb9ff0213),
	.w2(32'h3a3b3f09),
	.w3(32'h3a37e6d3),
	.w4(32'h3ae0c282),
	.w5(32'h3b0d3b57),
	.w6(32'hba526adc),
	.w7(32'hb987a7c6),
	.w8(32'hbaca2b33),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab879ae),
	.w1(32'h390dd36c),
	.w2(32'h3aa249e7),
	.w3(32'hbae12b13),
	.w4(32'h394d19cb),
	.w5(32'h3a6de446),
	.w6(32'h38b4b517),
	.w7(32'h3a1c659e),
	.w8(32'hb9e8e901),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae57360),
	.w1(32'hbb15b2f2),
	.w2(32'hb949ebca),
	.w3(32'hba6f6f5c),
	.w4(32'hbb73eb30),
	.w5(32'h3a9676ef),
	.w6(32'hbb902a6f),
	.w7(32'hbb8678f5),
	.w8(32'hb9c066f0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd4728),
	.w1(32'hb941eeb5),
	.w2(32'hb98e777c),
	.w3(32'hb9ae9c1e),
	.w4(32'hb999f59e),
	.w5(32'hb9db2666),
	.w6(32'h38810751),
	.w7(32'hb912137d),
	.w8(32'hbafa02a7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bb0ca),
	.w1(32'hba8e2cd9),
	.w2(32'hbaf90fd5),
	.w3(32'hba786f81),
	.w4(32'hba9456e5),
	.w5(32'hbaec9c75),
	.w6(32'hbb46edb0),
	.w7(32'hba87db00),
	.w8(32'hbb57826e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14bd01),
	.w1(32'hbab5bbda),
	.w2(32'hbac9bbe0),
	.w3(32'hbb116994),
	.w4(32'hbaae108c),
	.w5(32'hb98837d6),
	.w6(32'hba8c99dd),
	.w7(32'hba464ab0),
	.w8(32'hbb091b27),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b73bd),
	.w1(32'hba8ffe6d),
	.w2(32'hba593e7d),
	.w3(32'hba958a9f),
	.w4(32'hba5cab6d),
	.w5(32'hbaca51cf),
	.w6(32'hbb08cfea),
	.w7(32'hba991b8d),
	.w8(32'h3aed61c9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acc780),
	.w1(32'hbb0f04de),
	.w2(32'hbae9dfdd),
	.w3(32'hba5cdb06),
	.w4(32'hba8094f6),
	.w5(32'hbab52f65),
	.w6(32'h3a627d7c),
	.w7(32'h3a33daab),
	.w8(32'h37c0b64e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998804a),
	.w1(32'h39903302),
	.w2(32'hbb055e66),
	.w3(32'h3a73b560),
	.w4(32'h392004d3),
	.w5(32'hbaff6192),
	.w6(32'h3a0adc2c),
	.w7(32'hbac99588),
	.w8(32'hba8f15d8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97c853),
	.w1(32'h395de28d),
	.w2(32'hb9d150b3),
	.w3(32'hba0f8174),
	.w4(32'h3935f452),
	.w5(32'hba1825d1),
	.w6(32'hb835a0fd),
	.w7(32'hb9927c89),
	.w8(32'hba8acabe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a031d),
	.w1(32'h3ad407d4),
	.w2(32'h39c80a1f),
	.w3(32'hb96a2412),
	.w4(32'h3ab97069),
	.w5(32'hb900cb62),
	.w6(32'hba2986fc),
	.w7(32'hba72a627),
	.w8(32'hba33bf53),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba978cf5),
	.w1(32'hb9e6f24c),
	.w2(32'hb9b9c21b),
	.w3(32'hba618a14),
	.w4(32'hb9e7b338),
	.w5(32'hba21661b),
	.w6(32'hb8b6508e),
	.w7(32'hb888b107),
	.w8(32'hba40ead6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888d0f2),
	.w1(32'h3a593764),
	.w2(32'hba22d2a0),
	.w3(32'h39acac5b),
	.w4(32'hb9464b33),
	.w5(32'hbaa932c5),
	.w6(32'h3adeb3c5),
	.w7(32'h3a0ab0c2),
	.w8(32'hb9bc074f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a5f9c),
	.w1(32'h3a442e09),
	.w2(32'h39b295d0),
	.w3(32'hb9d0621d),
	.w4(32'h3a505d6c),
	.w5(32'h39cebc02),
	.w6(32'h39d11f36),
	.w7(32'h3990c6e1),
	.w8(32'hb99db315),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd2ec9),
	.w1(32'hb9354fb2),
	.w2(32'h39d515b9),
	.w3(32'h39d1a992),
	.w4(32'h3a57e676),
	.w5(32'h3a8abf86),
	.w6(32'hb99c8e43),
	.w7(32'hb810a6ad),
	.w8(32'hba0b575a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba125861),
	.w1(32'hba5bf5a4),
	.w2(32'hb93f2ce4),
	.w3(32'hb92f8eea),
	.w4(32'hb8368a7c),
	.w5(32'hb945f836),
	.w6(32'hba41c524),
	.w7(32'h39159b78),
	.w8(32'hba367a0e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31d5e7),
	.w1(32'h39ea0fbd),
	.w2(32'hba496f2b),
	.w3(32'hbabdbb0c),
	.w4(32'hba206753),
	.w5(32'hbb4511a0),
	.w6(32'hb99d20be),
	.w7(32'hba789289),
	.w8(32'hba730856),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44c1a2),
	.w1(32'hba743111),
	.w2(32'hb99e647b),
	.w3(32'hba0162af),
	.w4(32'hba2c7bb9),
	.w5(32'hb9fbd9e0),
	.w6(32'hba888902),
	.w7(32'hb94141ec),
	.w8(32'hbab4f005),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba461120),
	.w1(32'hba9da810),
	.w2(32'hba2610ac),
	.w3(32'hb9932854),
	.w4(32'hba5f1e37),
	.w5(32'hba9375ec),
	.w6(32'hbab955b7),
	.w7(32'hba585d9f),
	.w8(32'hbaf6ceb4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec94ae),
	.w1(32'hbb0cd41f),
	.w2(32'hbb191749),
	.w3(32'hba4f0cbe),
	.w4(32'hbaaeea74),
	.w5(32'hba856c75),
	.w6(32'hbb422185),
	.w7(32'hbb1427f6),
	.w8(32'hbb5dec98),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa06f80),
	.w1(32'h3b81cca6),
	.w2(32'hba6410b1),
	.w3(32'h3a67a98d),
	.w4(32'h3b1088d5),
	.w5(32'h3b2c34fe),
	.w6(32'hba974aa0),
	.w7(32'hbb49ba18),
	.w8(32'hb9ed0523),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874f77e),
	.w1(32'hbac20f1b),
	.w2(32'hba926c9e),
	.w3(32'hbab3d1b4),
	.w4(32'hbb3002ae),
	.w5(32'hbae95a36),
	.w6(32'hb9dc9cf3),
	.w7(32'hb95f54b7),
	.w8(32'h3b0065d1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3df9c),
	.w1(32'h39b872de),
	.w2(32'h3a75be13),
	.w3(32'h3ad2db0d),
	.w4(32'h3a7c5ff3),
	.w5(32'h3ace8011),
	.w6(32'h3a883af7),
	.w7(32'h3a8399c6),
	.w8(32'hbabdd4de),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba756996),
	.w1(32'hbacd493f),
	.w2(32'hba74fd72),
	.w3(32'hb9d9962a),
	.w4(32'hba4f32a7),
	.w5(32'hba816fc8),
	.w6(32'hbaf3d759),
	.w7(32'hba83c979),
	.w8(32'hb9f88873),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12fd8f),
	.w1(32'hba28ab22),
	.w2(32'hb953d5a4),
	.w3(32'hb9b7bbaf),
	.w4(32'hb9e1a013),
	.w5(32'hb9b13038),
	.w6(32'hba144310),
	.w7(32'hb91d3b99),
	.w8(32'hba795d57),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52880c),
	.w1(32'hba89f4ae),
	.w2(32'hba57519f),
	.w3(32'hb9b0cae3),
	.w4(32'hba2374e4),
	.w5(32'hba9a0200),
	.w6(32'hba5e44a2),
	.w7(32'hb9a32698),
	.w8(32'hba954a3b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac764be),
	.w1(32'hba8eb8ac),
	.w2(32'h3a9757ae),
	.w3(32'h3adbdca4),
	.w4(32'hbb1992b5),
	.w5(32'hb879555a),
	.w6(32'hba398b07),
	.w7(32'h3958c92f),
	.w8(32'hb998566b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8165e75),
	.w1(32'hba19a256),
	.w2(32'hb8a9a5aa),
	.w3(32'h3a2a879c),
	.w4(32'h399678d9),
	.w5(32'h39e4c09c),
	.w6(32'hba0f0c4d),
	.w7(32'hb9af6c5e),
	.w8(32'hbaaa1469),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ad41d),
	.w1(32'hbb12fa4c),
	.w2(32'hbb0560fe),
	.w3(32'hbb12974d),
	.w4(32'hbadc8f8b),
	.w5(32'hb976593a),
	.w6(32'hbb74cb0c),
	.w7(32'hbb371251),
	.w8(32'hbb640a23),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fbd51),
	.w1(32'hbb7c8091),
	.w2(32'hbb081c87),
	.w3(32'hbb2f2ee7),
	.w4(32'hba82b341),
	.w5(32'hba44887c),
	.w6(32'hbb5498bd),
	.w7(32'hbb24584a),
	.w8(32'hb82775ad),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87ebf52),
	.w1(32'h3af2748e),
	.w2(32'h3a34cd1d),
	.w3(32'h39933414),
	.w4(32'h3a8bc70a),
	.w5(32'h38fe7625),
	.w6(32'hb9ec08b1),
	.w7(32'hb9fc105a),
	.w8(32'hb9c98c2f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe9749),
	.w1(32'h3afab351),
	.w2(32'hb7a19b30),
	.w3(32'hbb013089),
	.w4(32'h3aa3012e),
	.w5(32'hbb2339fd),
	.w6(32'h3a541a56),
	.w7(32'hbad20a22),
	.w8(32'h3a3ad6ba),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b4fe0),
	.w1(32'hb9c808bb),
	.w2(32'h3958b9e6),
	.w3(32'h3a41c674),
	.w4(32'h385fd08a),
	.w5(32'h37e01333),
	.w6(32'h38fd9e12),
	.w7(32'h39742046),
	.w8(32'hbb85794d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb556ab7),
	.w1(32'hbb851584),
	.w2(32'hbba42931),
	.w3(32'hbb8610d9),
	.w4(32'hbbad7989),
	.w5(32'hbb94c1c3),
	.w6(32'hbbabfe2b),
	.w7(32'hbb9e93fc),
	.w8(32'h3a5ca3a8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4103),
	.w1(32'h3b827f9a),
	.w2(32'h3ac847f0),
	.w3(32'h3a5c7ab2),
	.w4(32'h3b9e97f1),
	.w5(32'h3b56c7e7),
	.w6(32'hbaf05e09),
	.w7(32'hbac0b433),
	.w8(32'hba92e90d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81c7bd),
	.w1(32'hbb08eb3f),
	.w2(32'hbb31c1a6),
	.w3(32'hbb0de247),
	.w4(32'hbb2b061a),
	.w5(32'hbaf1eeaa),
	.w6(32'hbb13602b),
	.w7(32'hbb0eb9f5),
	.w8(32'hbac8063a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc4b1),
	.w1(32'hbadf7163),
	.w2(32'hba050e78),
	.w3(32'hb987fac3),
	.w4(32'hb9cd6a8f),
	.w5(32'hba3a083a),
	.w6(32'hbad1307c),
	.w7(32'hba0b28be),
	.w8(32'h392a9014),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7c00),
	.w1(32'h3bac5e62),
	.w2(32'h3b0a3ebc),
	.w3(32'h38cd6d2a),
	.w4(32'h3b16fabc),
	.w5(32'hbab0fdb7),
	.w6(32'h3b84c9f0),
	.w7(32'h394d4c3e),
	.w8(32'hba623a4c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a5bb3),
	.w1(32'hba84923e),
	.w2(32'h3901bbec),
	.w3(32'hba0235a0),
	.w4(32'hba430938),
	.w5(32'hb92d43bb),
	.w6(32'hba83556c),
	.w7(32'h38abfd06),
	.w8(32'hb9b82a84),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9923990),
	.w1(32'hb9b8232d),
	.w2(32'hb8e9f0f5),
	.w3(32'hb91d2fa9),
	.w4(32'hb91a0054),
	.w5(32'hb991f1a8),
	.w6(32'hb9b5bd76),
	.w7(32'hb86edd71),
	.w8(32'hb9f79077),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c89a0d),
	.w1(32'hb9f07801),
	.w2(32'hb9c09213),
	.w3(32'hb8b671f1),
	.w4(32'hb9b7d2f5),
	.w5(32'hb9f82542),
	.w6(32'hb9c2377d),
	.w7(32'hb946379b),
	.w8(32'h3a511b35),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925b435),
	.w1(32'hba77a64c),
	.w2(32'hbb51458f),
	.w3(32'hb9e5e1b0),
	.w4(32'hba873945),
	.w5(32'hba521c82),
	.w6(32'h3a625287),
	.w7(32'hb62d8a0e),
	.w8(32'hba9b84b2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54ed68),
	.w1(32'hba9ec379),
	.w2(32'hba2bcc37),
	.w3(32'hb9ee6f95),
	.w4(32'hba51a806),
	.w5(32'hba5cf6f0),
	.w6(32'hbab2a25b),
	.w7(32'hba5e1114),
	.w8(32'hba65088b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928faae),
	.w1(32'hba4680e6),
	.w2(32'hba409fb5),
	.w3(32'hb8d272cb),
	.w4(32'hba2f8371),
	.w5(32'hbac9f4ed),
	.w6(32'hba3132a8),
	.w7(32'hba1f469b),
	.w8(32'hba3f1259),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06f9f0),
	.w1(32'hba55d54b),
	.w2(32'hb871deec),
	.w3(32'hb88b7561),
	.w4(32'hb98b679e),
	.w5(32'hb9d30743),
	.w6(32'hba2b3fdb),
	.w7(32'h3906c881),
	.w8(32'hbaba507c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82b78e),
	.w1(32'hbacf60a8),
	.w2(32'hba8e15f1),
	.w3(32'hba1ef71d),
	.w4(32'hba7ff79f),
	.w5(32'hba834074),
	.w6(32'hbae49ecc),
	.w7(32'hba8bab64),
	.w8(32'hba86788d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131523),
	.w1(32'hba82d300),
	.w2(32'hb8f4490b),
	.w3(32'hb85b1d46),
	.w4(32'hba0935be),
	.w5(32'hba17e210),
	.w6(32'hba8a23cc),
	.w7(32'hb902d9cd),
	.w8(32'hbaa96140),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ca913),
	.w1(32'h395076b9),
	.w2(32'hbabc8701),
	.w3(32'hbab38403),
	.w4(32'hba35ecb0),
	.w5(32'hbac10447),
	.w6(32'h3aa46b9d),
	.w7(32'hbb01d247),
	.w8(32'hbad1349b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab88e66),
	.w1(32'hba9afd78),
	.w2(32'hbad3800b),
	.w3(32'hba5b567b),
	.w4(32'hba998c43),
	.w5(32'hbab998c9),
	.w6(32'hbaafcf9b),
	.w7(32'hbabd2a71),
	.w8(32'hb9dc0cea),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fd1b4),
	.w1(32'hba2dfb5c),
	.w2(32'hb9909250),
	.w3(32'hb7b01446),
	.w4(32'hb98c3019),
	.w5(32'hba02d272),
	.w6(32'hba25d3ca),
	.w7(32'hb812f50a),
	.w8(32'hba879892),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56a055),
	.w1(32'hba83be7a),
	.w2(32'hba5e5e5e),
	.w3(32'hba048e6f),
	.w4(32'hba35cf99),
	.w5(32'hba4fd91e),
	.w6(32'hba84cfbd),
	.w7(32'hb9ff01f8),
	.w8(32'hba2ee7fe),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8f536),
	.w1(32'hba778c04),
	.w2(32'hba476622),
	.w3(32'h381c9a09),
	.w4(32'hba45f5b4),
	.w5(32'hbad5812a),
	.w6(32'hba4ac118),
	.w7(32'hba39bbe1),
	.w8(32'hba9834f0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22b564),
	.w1(32'hba8db4d6),
	.w2(32'hba499947),
	.w3(32'hb9c3df6a),
	.w4(32'hba1b37eb),
	.w5(32'hba949207),
	.w6(32'hba44401f),
	.w7(32'hba344d5d),
	.w8(32'hba1570a5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8931e1),
	.w1(32'hbaae7394),
	.w2(32'hba5e2902),
	.w3(32'hba93532c),
	.w4(32'hbad920e0),
	.w5(32'hba2856df),
	.w6(32'hba9dbd13),
	.w7(32'hba2e5852),
	.w8(32'h3ad7cb4b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39144774),
	.w1(32'h37f4f2ba),
	.w2(32'hbb36303e),
	.w3(32'h398db285),
	.w4(32'h39f0ed22),
	.w5(32'hbb3f1e7e),
	.w6(32'h3a15fdd3),
	.w7(32'h3a6c37b7),
	.w8(32'hba225d5e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba484850),
	.w1(32'hba86b25f),
	.w2(32'hba80ee46),
	.w3(32'hb9f97c56),
	.w4(32'hba6f0937),
	.w5(32'hba72dc7c),
	.w6(32'hba6791da),
	.w7(32'hba4b0d4e),
	.w8(32'hbb2f0133),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb059e78),
	.w1(32'hbb3ffead),
	.w2(32'hbb1f0e16),
	.w3(32'hbacf7859),
	.w4(32'hbb2cdb4d),
	.w5(32'hbb0558d5),
	.w6(32'hbb6e3898),
	.w7(32'hbb1b4d66),
	.w8(32'h39fdeeb0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92c7c1),
	.w1(32'h3a968081),
	.w2(32'hbb180e81),
	.w3(32'hbb1c42bb),
	.w4(32'hbb229353),
	.w5(32'hb77afb4f),
	.w6(32'hbb1c390a),
	.w7(32'hbb80cbf6),
	.w8(32'hbac1973b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba755f29),
	.w1(32'hbb04323a),
	.w2(32'hbaeb75cf),
	.w3(32'hb8a1c59c),
	.w4(32'hbabb1b82),
	.w5(32'hbaa87038),
	.w6(32'hbb02903b),
	.w7(32'hbaf16dfc),
	.w8(32'hbac8d130),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d7d76),
	.w1(32'hbaade926),
	.w2(32'hba379683),
	.w3(32'hb9b71572),
	.w4(32'hba319137),
	.w5(32'hba86debb),
	.w6(32'hbabb6b7a),
	.w7(32'hba2e5c5d),
	.w8(32'h3b36db39),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae669c8),
	.w1(32'h39dc0ca5),
	.w2(32'h3aa01732),
	.w3(32'h3b084ea9),
	.w4(32'h3aa51d84),
	.w5(32'h3b09fb9a),
	.w6(32'h3ab0f7d5),
	.w7(32'h3aaeff3d),
	.w8(32'hba3d2397),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c45273),
	.w1(32'hbabe8926),
	.w2(32'hb9bfd759),
	.w3(32'hba0fc679),
	.w4(32'hbaa89d5f),
	.w5(32'hb9d76ea1),
	.w6(32'hbad8126c),
	.w7(32'hb97a3726),
	.w8(32'hbb5b7b84),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ebfcd),
	.w1(32'hbb240fd0),
	.w2(32'hbb93c0f0),
	.w3(32'hbb4e1ff5),
	.w4(32'hbb810270),
	.w5(32'hbb863aa3),
	.w6(32'hbb8eabbe),
	.w7(32'hbb85d67f),
	.w8(32'h3b2b1dac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addffbd),
	.w1(32'h39e36a99),
	.w2(32'h3a98575a),
	.w3(32'h3b01a416),
	.w4(32'h3a9dc710),
	.w5(32'h3aff5e06),
	.w6(32'h3aaa198a),
	.w7(32'h3aa6a57e),
	.w8(32'h3b10c424),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3807a),
	.w1(32'h39db450c),
	.w2(32'h3a880934),
	.w3(32'h3ae43308),
	.w4(32'h3a8c657b),
	.w5(32'h3adfe9cf),
	.w6(32'h3a966379),
	.w7(32'h3a936ee2),
	.w8(32'hba54a132),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45575b),
	.w1(32'hba98ac62),
	.w2(32'hba31a89e),
	.w3(32'hb97bff92),
	.w4(32'hba437c5b),
	.w5(32'hba3aaf6e),
	.w6(32'hbaabf574),
	.w7(32'hba55ba89),
	.w8(32'hb97e17a0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba977dc9),
	.w1(32'hbaab9ce0),
	.w2(32'hb9c13ae5),
	.w3(32'hba69e1d0),
	.w4(32'hbb89e380),
	.w5(32'hbaf35e52),
	.w6(32'hba302078),
	.w7(32'hb9197380),
	.w8(32'hb9a95bc9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a2e7f),
	.w1(32'hb911cb5f),
	.w2(32'hb9886a21),
	.w3(32'h38db0195),
	.w4(32'hb7ff4f6b),
	.w5(32'hb9a13d8f),
	.w6(32'h370e1c00),
	.w7(32'h38450f44),
	.w8(32'h3ad385dc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64e953),
	.w1(32'h3a4907ea),
	.w2(32'hbb10b3ad),
	.w3(32'hbaec9dc4),
	.w4(32'hba9dbb4a),
	.w5(32'hbafe4f46),
	.w6(32'hb9cb9bc6),
	.w7(32'hba139e92),
	.w8(32'hbb8763f7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d9c35),
	.w1(32'hbbb56eb2),
	.w2(32'hbb8ee088),
	.w3(32'hbad438a9),
	.w4(32'hbb6ab3ee),
	.w5(32'hbb6169f4),
	.w6(32'hbba80a0c),
	.w7(32'hbb8dd611),
	.w8(32'h3ae87bed),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae28ea6),
	.w1(32'hb94cdbf3),
	.w2(32'hba8a5195),
	.w3(32'hb9f21fcb),
	.w4(32'h39db1c89),
	.w5(32'h37f73c8f),
	.w6(32'h3aa71440),
	.w7(32'h3aa466b4),
	.w8(32'hba05b539),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5694ec),
	.w1(32'h3b4e46fd),
	.w2(32'h39456ec1),
	.w3(32'h3947bceb),
	.w4(32'hbaaeb468),
	.w5(32'h3a70c985),
	.w6(32'h3b08da74),
	.w7(32'hbabad508),
	.w8(32'hba16c807),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9234af0),
	.w1(32'hba5bdd9d),
	.w2(32'hba25367d),
	.w3(32'hb74146ae),
	.w4(32'hba2f5b21),
	.w5(32'hbab09e68),
	.w6(32'hba3a3a8f),
	.w7(32'hba1dfa3c),
	.w8(32'hbaa84642),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7de6e8),
	.w1(32'hbab9e594),
	.w2(32'hb9776c3e),
	.w3(32'hba3be94e),
	.w4(32'hba993447),
	.w5(32'hb9d9e7e7),
	.w6(32'hbb058562),
	.w7(32'hba35b137),
	.w8(32'hbb35fd68),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5f2e),
	.w1(32'hbb3fc97f),
	.w2(32'hbb887136),
	.w3(32'hbb0d7bb9),
	.w4(32'hbb33a8b2),
	.w5(32'hbb4c52d7),
	.w6(32'hbb8aef3e),
	.w7(32'hbb769bc7),
	.w8(32'hba1270c5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb93d6),
	.w1(32'hba3243e8),
	.w2(32'hba005ca1),
	.w3(32'hb9728bf8),
	.w4(32'hba01223f),
	.w5(32'hba22eeff),
	.w6(32'hba1015bd),
	.w7(32'hb97b3f4e),
	.w8(32'hbb2f2098),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d4db),
	.w1(32'hbb0d8ed3),
	.w2(32'hbab6586d),
	.w3(32'hba7456aa),
	.w4(32'hba6067be),
	.w5(32'hbb110fbb),
	.w6(32'hbada2795),
	.w7(32'hbab390cf),
	.w8(32'hbb23cd01),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f9a9),
	.w1(32'hbb264b7f),
	.w2(32'hbb1fab63),
	.w3(32'hbab9c5e5),
	.w4(32'hbb09b3a4),
	.w5(32'hbb02191c),
	.w6(32'hbb2725f2),
	.w7(32'hbb2657e1),
	.w8(32'h3a83a103),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a318229),
	.w1(32'h3941908b),
	.w2(32'h39e19b33),
	.w3(32'h3a49a7de),
	.w4(32'h39fba12e),
	.w5(32'h3a494b23),
	.w6(32'h3a070ebe),
	.w7(32'h3a03afa9),
	.w8(32'h398e3a11),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a7d8b),
	.w1(32'hba2435c7),
	.w2(32'hb9d7e8ed),
	.w3(32'hb9e308ad),
	.w4(32'hb999e204),
	.w5(32'hba15ee84),
	.w6(32'h39980e3f),
	.w7(32'hb9a1c759),
	.w8(32'h3acdcf40),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f429),
	.w1(32'hba53b5a0),
	.w2(32'hb9c9848a),
	.w3(32'h3ad2d02f),
	.w4(32'hbb69ec24),
	.w5(32'hbb64a57a),
	.w6(32'hbb88da5d),
	.w7(32'hba2acc31),
	.w8(32'h3850b25e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b07ffa),
	.w1(32'hb9e861ff),
	.w2(32'h39000808),
	.w3(32'hba184672),
	.w4(32'hb7462965),
	.w5(32'h394eac26),
	.w6(32'h3992d480),
	.w7(32'hb7e9fdff),
	.w8(32'h391d7e94),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96102af),
	.w1(32'h395f5e8e),
	.w2(32'h39939137),
	.w3(32'hba1efc25),
	.w4(32'h39844f84),
	.w5(32'h39b83c03),
	.w6(32'h3a1cb2db),
	.w7(32'h39983b87),
	.w8(32'hbab99454),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08dd9c),
	.w1(32'hbaf2ce22),
	.w2(32'hbac1c8c6),
	.w3(32'hbabfc43f),
	.w4(32'hba779daa),
	.w5(32'hbaca5ef8),
	.w6(32'hba880b9a),
	.w7(32'hba811078),
	.w8(32'h391675ea),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abba21d),
	.w1(32'hbbb0e53f),
	.w2(32'hbb18cc56),
	.w3(32'hba95a8a5),
	.w4(32'hbbe36a4f),
	.w5(32'hbba629e4),
	.w6(32'h3ae7f0a1),
	.w7(32'h3a4a29f9),
	.w8(32'hba7c781a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a74c3),
	.w1(32'hb7ab0694),
	.w2(32'hbab90995),
	.w3(32'hb924e8bf),
	.w4(32'h39fb1a09),
	.w5(32'hbaa944b2),
	.w6(32'h398aa258),
	.w7(32'hb96a5297),
	.w8(32'h3a12d8af),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3867327f),
	.w1(32'hb9d360d8),
	.w2(32'hba3d3fcd),
	.w3(32'h3a2ceee1),
	.w4(32'h3934614b),
	.w5(32'h38b952f9),
	.w6(32'hb9879712),
	.w7(32'hbaa9f1c7),
	.w8(32'hb881965f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ddb19),
	.w1(32'hba46c746),
	.w2(32'hb8aab8fe),
	.w3(32'hba68e2d2),
	.w4(32'hb92e90a7),
	.w5(32'hb92daeda),
	.w6(32'h39438458),
	.w7(32'h39d090fb),
	.w8(32'h39e09f7c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386ed29d),
	.w1(32'hb9034b90),
	.w2(32'h39867e1f),
	.w3(32'hb87da5af),
	.w4(32'h395fb95e),
	.w5(32'h39e92f8e),
	.w6(32'h39bad17d),
	.w7(32'h39d005ed),
	.w8(32'h3a599ede),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bf35a),
	.w1(32'hb9ea3d4e),
	.w2(32'h39169b68),
	.w3(32'hb957a097),
	.w4(32'h37f98a58),
	.w5(32'h3a0a4a30),
	.w6(32'h3a5dead2),
	.w7(32'h3a007041),
	.w8(32'h39cfac2b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f220e),
	.w1(32'h3a074ce5),
	.w2(32'h3b01dec4),
	.w3(32'h3b222576),
	.w4(32'h3aafa352),
	.w5(32'h3ac03ae2),
	.w6(32'hbaacad76),
	.w7(32'h3b142b40),
	.w8(32'h3af44d8d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256b6e),
	.w1(32'h3942d214),
	.w2(32'h3a1cd6ab),
	.w3(32'h3abb2d04),
	.w4(32'h3a866e23),
	.w5(32'h3aeb8744),
	.w6(32'h3aa01cc0),
	.w7(32'h39bdb9c0),
	.w8(32'hbb25948c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a61c5),
	.w1(32'hbaeb2e4b),
	.w2(32'hb9ace5f6),
	.w3(32'hba82234e),
	.w4(32'hbb479732),
	.w5(32'hbb7c656a),
	.w6(32'hb90029da),
	.w7(32'h3b1555a0),
	.w8(32'hb9e9aa71),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376656),
	.w1(32'hbae527ee),
	.w2(32'hbab8e8cd),
	.w3(32'h3ad29f82),
	.w4(32'h39dfe6b6),
	.w5(32'h394fa4d3),
	.w6(32'hba2d027b),
	.w7(32'hb91f9790),
	.w8(32'hba4a7c34),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f4e54),
	.w1(32'hba954281),
	.w2(32'h3b3664cf),
	.w3(32'h3a907a98),
	.w4(32'h3ae81c26),
	.w5(32'h39eafd47),
	.w6(32'hbabb7ff6),
	.w7(32'h3b179484),
	.w8(32'hbab1785d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a5775),
	.w1(32'h3a5b40f8),
	.w2(32'hba26ab21),
	.w3(32'h399c6f59),
	.w4(32'hbb463ad1),
	.w5(32'hbb2c1394),
	.w6(32'hbb4e83be),
	.w7(32'h393d796c),
	.w8(32'h3a974386),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94b595),
	.w1(32'hb878b6b4),
	.w2(32'h3a53608b),
	.w3(32'h3aa98d67),
	.w4(32'h3a1af849),
	.w5(32'h3a5e487e),
	.w6(32'h3a1d3ee1),
	.w7(32'h3a461b34),
	.w8(32'hb95b8403),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01c08d),
	.w1(32'hba2101c6),
	.w2(32'hbafcca72),
	.w3(32'hbab9c2c8),
	.w4(32'hbb091974),
	.w5(32'hbb00dba8),
	.w6(32'hba72beee),
	.w7(32'hbb15e821),
	.w8(32'h3988ea11),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31d4bd),
	.w1(32'hbab7a32f),
	.w2(32'h3b7c7800),
	.w3(32'h3a1f302a),
	.w4(32'h3a68ed98),
	.w5(32'hbb172dbc),
	.w6(32'hbb328212),
	.w7(32'h3a7dfbca),
	.w8(32'hbaf89a83),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab509b3),
	.w1(32'hbb588662),
	.w2(32'hbb392d87),
	.w3(32'hbb0130cd),
	.w4(32'hbb0c649c),
	.w5(32'hbb4d919b),
	.w6(32'hba440c09),
	.w7(32'hbab6ae88),
	.w8(32'h3b1204b3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16ed63),
	.w1(32'hba3152aa),
	.w2(32'h3a868f94),
	.w3(32'h399d9788),
	.w4(32'h39d1708f),
	.w5(32'h3ac44f77),
	.w6(32'h3a6bdcc6),
	.w7(32'h3aa95cf8),
	.w8(32'hbb44ade4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f8bb),
	.w1(32'hbb298dfd),
	.w2(32'hbb23f3cb),
	.w3(32'h3af4fc0d),
	.w4(32'hb90d9f29),
	.w5(32'h3a4fc119),
	.w6(32'hbaf42744),
	.w7(32'hba13c85a),
	.w8(32'h38fadc7e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule