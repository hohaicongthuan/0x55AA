module layer_8_featuremap_1(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bda24),
	.w1(32'h3b5371ea),
	.w2(32'hbbcc62d7),
	.w3(32'hbc70b83b),
	.w4(32'h3b467b38),
	.w5(32'hbb1bea21),
	.w6(32'hbbcbdca9),
	.w7(32'hba911d28),
	.w8(32'hbbea37d7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea548),
	.w1(32'hbbf847e9),
	.w2(32'hb97be1ee),
	.w3(32'h3c196291),
	.w4(32'hbbcb21ef),
	.w5(32'hbb0ea285),
	.w6(32'h3aa0e4dd),
	.w7(32'hbb28fcb8),
	.w8(32'hbadda6ce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abebea5),
	.w1(32'hbbc660fa),
	.w2(32'h3a60ca59),
	.w3(32'hba6e564d),
	.w4(32'hbc022f1e),
	.w5(32'h3af94de7),
	.w6(32'hbb2378ed),
	.w7(32'hbbf37044),
	.w8(32'hba670970),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc8ff4),
	.w1(32'hb9ba37e6),
	.w2(32'h3b68f364),
	.w3(32'h3bdcc342),
	.w4(32'hbb70ec20),
	.w5(32'h3b0cb21e),
	.w6(32'h3b4064d6),
	.w7(32'hbaefa23f),
	.w8(32'hbb86fa5f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd08bae),
	.w1(32'hbb82449b),
	.w2(32'hbc0b8e83),
	.w3(32'h3c017953),
	.w4(32'hbb9c693b),
	.w5(32'hbb82fa89),
	.w6(32'hba94f0a8),
	.w7(32'hba804a80),
	.w8(32'hbbbfb7ed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840790),
	.w1(32'h3be5e381),
	.w2(32'h3a46d359),
	.w3(32'h3b9446d5),
	.w4(32'hba5b6fdb),
	.w5(32'hbc43b429),
	.w6(32'hbb047eba),
	.w7(32'hbc8b3482),
	.w8(32'hbb9d56d1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf43848),
	.w1(32'hbbc5fc5f),
	.w2(32'hbb034ebf),
	.w3(32'hbc4b921b),
	.w4(32'hbac5a96e),
	.w5(32'h3a5c4441),
	.w6(32'h398f220a),
	.w7(32'hbb75a370),
	.w8(32'h3b0cb1d6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4ac73),
	.w1(32'h3c6e1626),
	.w2(32'hbc213d09),
	.w3(32'h3bd04afb),
	.w4(32'h3c8fb899),
	.w5(32'h3b123696),
	.w6(32'h3be5ddbd),
	.w7(32'hbb85b9d3),
	.w8(32'h3c45b73c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc321f53),
	.w1(32'h3bed8ef8),
	.w2(32'h3c3e7724),
	.w3(32'hbc93736e),
	.w4(32'h3c007e53),
	.w5(32'h3c67f388),
	.w6(32'hbbcda6ac),
	.w7(32'h3c429da4),
	.w8(32'h3c8850d6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c744ac9),
	.w1(32'hbbc95f37),
	.w2(32'hbd24e454),
	.w3(32'h3c9adf5d),
	.w4(32'hbd457cef),
	.w5(32'hbd5f0fd2),
	.w6(32'h3c63f5ea),
	.w7(32'hbc7d03e2),
	.w8(32'hbb5d206c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b3d82),
	.w1(32'hbabeba95),
	.w2(32'hbc05d369),
	.w3(32'hbc5603e4),
	.w4(32'hbbb9b27c),
	.w5(32'hb9878ba0),
	.w6(32'h3c8cb615),
	.w7(32'hbc0a9121),
	.w8(32'hb964576a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93ed2a),
	.w1(32'h3c4874fa),
	.w2(32'hbc8a8298),
	.w3(32'hbbec9e62),
	.w4(32'h3c256ff5),
	.w5(32'hbd019cc7),
	.w6(32'hbbd24a53),
	.w7(32'h3c5a04cd),
	.w8(32'hbca9b1d6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99b12b),
	.w1(32'hbc92be3a),
	.w2(32'h3c0f9c7f),
	.w3(32'hbd052185),
	.w4(32'hbc994a83),
	.w5(32'h3ba3388a),
	.w6(32'hbcb51d9b),
	.w7(32'hbcca64f9),
	.w8(32'hbd2ec0a1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdec9f2),
	.w1(32'hbc010c8f),
	.w2(32'hbb5a2930),
	.w3(32'h3cff9d31),
	.w4(32'hb949645c),
	.w5(32'h3c0254fe),
	.w6(32'hbc1eb4fc),
	.w7(32'hbb80cf7f),
	.w8(32'h3b9cbfb8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027af5),
	.w1(32'h3a819ff4),
	.w2(32'h3ba4d792),
	.w3(32'h3ae4d8d2),
	.w4(32'h3ae46717),
	.w5(32'hba6001f0),
	.w6(32'h3b8b65df),
	.w7(32'h3b005e05),
	.w8(32'h3b11bb8d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01bf5d),
	.w1(32'h3be9c035),
	.w2(32'h3c01803f),
	.w3(32'h39acf214),
	.w4(32'h3c39c9fc),
	.w5(32'h3c7c27f5),
	.w6(32'h3b1fbc1f),
	.w7(32'h3c56393a),
	.w8(32'h3c624f46),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c394a71),
	.w1(32'h3cc934cb),
	.w2(32'h3c81084b),
	.w3(32'h3c93cd94),
	.w4(32'h3ccb72c6),
	.w5(32'hbc260717),
	.w6(32'h3c11cbd8),
	.w7(32'hbc819a36),
	.w8(32'hbd2f79ff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc966f7d),
	.w1(32'h3a24f534),
	.w2(32'h3accb874),
	.w3(32'hbd64eb48),
	.w4(32'h3ad75178),
	.w5(32'h3a9a47fe),
	.w6(32'hbd2f1133),
	.w7(32'h39910134),
	.w8(32'hb9108210),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95183a),
	.w1(32'h3c8df8bc),
	.w2(32'hbb9a1196),
	.w3(32'h3c168cdf),
	.w4(32'h3c9e5f3c),
	.w5(32'hbb5cb4cd),
	.w6(32'h3bd327be),
	.w7(32'h3bb4bffb),
	.w8(32'h3c5cf626),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd60e4),
	.w1(32'hbc92446a),
	.w2(32'hbc14d2e8),
	.w3(32'hbc2bf2b8),
	.w4(32'hbc375895),
	.w5(32'hbb2344d1),
	.w6(32'hbb25299a),
	.w7(32'hbbdae69f),
	.w8(32'hba95833c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12b72e),
	.w1(32'hbbb8dc74),
	.w2(32'h3b4025aa),
	.w3(32'h38828ec7),
	.w4(32'h3aa9472a),
	.w5(32'h3c3bc592),
	.w6(32'hb7faf28d),
	.w7(32'hbbb28b89),
	.w8(32'h3b5f4046),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a8b3),
	.w1(32'hbb214542),
	.w2(32'hbc727c5b),
	.w3(32'h3bc35143),
	.w4(32'hbb4a4d1c),
	.w5(32'h3b5cde95),
	.w6(32'h3bf42991),
	.w7(32'h3cbdba9e),
	.w8(32'h3d1b1ac0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe934ae),
	.w1(32'hbc52c252),
	.w2(32'hbc01a1f8),
	.w3(32'hbb25a8f9),
	.w4(32'h3bfe19d7),
	.w5(32'h3b595e74),
	.w6(32'h3c0dc783),
	.w7(32'h3b0ae66f),
	.w8(32'hbca4ec90),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391d9c),
	.w1(32'hbc9ad8b4),
	.w2(32'hbc0b11b9),
	.w3(32'hbbdc2aeb),
	.w4(32'hbc31ab6c),
	.w5(32'hbb2cdac7),
	.w6(32'hbbccf33b),
	.w7(32'hbbfef39f),
	.w8(32'h3a4b6d36),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d8af),
	.w1(32'h3b93a7ae),
	.w2(32'hbbae38ad),
	.w3(32'hbb768962),
	.w4(32'hb932bc9a),
	.w5(32'hbca1754a),
	.w6(32'hba868281),
	.w7(32'hbca0fd6a),
	.w8(32'hbd118ef0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd28c4e0),
	.w1(32'h3bb410cd),
	.w2(32'h3a8d6bd7),
	.w3(32'hbd2150e3),
	.w4(32'h3c88dda3),
	.w5(32'h3c078e8c),
	.w6(32'hbc1bc0a8),
	.w7(32'h3c90a15c),
	.w8(32'h3c448b14),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd408d),
	.w1(32'hbae658e6),
	.w2(32'h3c8c591b),
	.w3(32'h3c27a92b),
	.w4(32'h3ba7ad07),
	.w5(32'h3cb087a6),
	.w6(32'h3ca4cc31),
	.w7(32'h3b157ad0),
	.w8(32'h3c803f42),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e4d09),
	.w1(32'h3cff5c7b),
	.w2(32'h3d098002),
	.w3(32'h3c714544),
	.w4(32'h3d2d0cc9),
	.w5(32'h3d58a7fc),
	.w6(32'h3ceaafe4),
	.w7(32'h3d5ee87a),
	.w8(32'h3cfebe6c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca69241),
	.w1(32'h3bf15718),
	.w2(32'hbaa3374a),
	.w3(32'h3c8c055e),
	.w4(32'h3bc099c6),
	.w5(32'hbc3ffa44),
	.w6(32'h3c0b2093),
	.w7(32'h3c8c423b),
	.w8(32'h3b956229),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb231ea5),
	.w1(32'h3b9cd6b4),
	.w2(32'h3bdb10a4),
	.w3(32'hbc09d6a3),
	.w4(32'h3c00b3b0),
	.w5(32'h3c1bd7ad),
	.w6(32'h3bfd3557),
	.w7(32'h3b62514a),
	.w8(32'h3a3b14d6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0067a9),
	.w1(32'h3cb1dd3e),
	.w2(32'hbc26501f),
	.w3(32'h3b029fd0),
	.w4(32'h3cd4bf19),
	.w5(32'hbc8a3285),
	.w6(32'hbadcade5),
	.w7(32'h3cc7b268),
	.w8(32'h3b931be1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfabc0),
	.w1(32'hbbc4f36b),
	.w2(32'h3b0e000a),
	.w3(32'hbc91e397),
	.w4(32'hbb3d462f),
	.w5(32'h3bd6f0d9),
	.w6(32'hbbb43112),
	.w7(32'h3a88a973),
	.w8(32'h3c40da04),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54f114),
	.w1(32'h3bda2cf2),
	.w2(32'h3c0bc968),
	.w3(32'h3bc0fa7b),
	.w4(32'h3c37873c),
	.w5(32'h3c5bbfa5),
	.w6(32'h3bba6ac0),
	.w7(32'h3c25b3a9),
	.w8(32'h3c4d68d0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbaf17),
	.w1(32'hbb8f87b9),
	.w2(32'hbc898dbf),
	.w3(32'h3c20447b),
	.w4(32'hbbd5151b),
	.w5(32'hbcf92091),
	.w6(32'h3c0e60b5),
	.w7(32'h3a73b080),
	.w8(32'hbc97c866),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e85b3),
	.w1(32'h3b88d43f),
	.w2(32'hbb3eeba5),
	.w3(32'hbca62022),
	.w4(32'h3a8634f6),
	.w5(32'hbbc84678),
	.w6(32'hbcbad651),
	.w7(32'h3ba06092),
	.w8(32'hba2be8f3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b93c6),
	.w1(32'h3b300f69),
	.w2(32'hbcc903ce),
	.w3(32'h3bec24b7),
	.w4(32'hbba024ba),
	.w5(32'hbd16f7fb),
	.w6(32'h3c061c79),
	.w7(32'hbb7493d7),
	.w8(32'hbcf57b7f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc14f7e),
	.w1(32'hbc9db87c),
	.w2(32'hbc2be3c5),
	.w3(32'hbd26bf50),
	.w4(32'hbce3675a),
	.w5(32'hbcee16b8),
	.w6(32'hbcfc14a6),
	.w7(32'hbc7e263d),
	.w8(32'hbcbdf496),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6283f9),
	.w1(32'hbc6cf9f4),
	.w2(32'hbb37ab3b),
	.w3(32'hbca52e26),
	.w4(32'hbc193bc7),
	.w5(32'hbb4934e8),
	.w6(32'hbcbaef86),
	.w7(32'h3b96e0e8),
	.w8(32'h3b61f5c0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c065fa1),
	.w1(32'hbae7fcfa),
	.w2(32'hbb8c6064),
	.w3(32'h3cb7e79f),
	.w4(32'h3c1d61ae),
	.w5(32'h3b26a2b9),
	.w6(32'h3bd2ebfa),
	.w7(32'h3c62feb6),
	.w8(32'h3c0ee0cb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a2a62),
	.w1(32'h3bd6de38),
	.w2(32'hbcb67131),
	.w3(32'h3cbede2c),
	.w4(32'hb8ea5952),
	.w5(32'hbd05c847),
	.w6(32'h3c9f974b),
	.w7(32'h3a446c38),
	.w8(32'hbcc0e376),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b647a),
	.w1(32'h3b71c165),
	.w2(32'hbb84b522),
	.w3(32'hba8c3932),
	.w4(32'h3ca3f4bc),
	.w5(32'hbafc1fed),
	.w6(32'hbab93e6d),
	.w7(32'hb9efb086),
	.w8(32'hbc02ec84),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ccc3),
	.w1(32'hbbcaceb7),
	.w2(32'hbaf87175),
	.w3(32'hbb3eb384),
	.w4(32'hba1ac82c),
	.w5(32'h3bddaae4),
	.w6(32'h3bc86340),
	.w7(32'hbb1e3672),
	.w8(32'h3b9913fc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc5f3),
	.w1(32'h3c750773),
	.w2(32'h3b83455c),
	.w3(32'hba4df37a),
	.w4(32'h3c19cf6c),
	.w5(32'hbb1281af),
	.w6(32'hba666c9d),
	.w7(32'h3c273068),
	.w8(32'hb98498e4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1738ef),
	.w1(32'h3905b4a7),
	.w2(32'h3be3f681),
	.w3(32'h3b88d21a),
	.w4(32'h3bf256b0),
	.w5(32'hbbb9043e),
	.w6(32'h3bda1afc),
	.w7(32'h3c43a191),
	.w8(32'h3add7fe4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60785f),
	.w1(32'h3c274145),
	.w2(32'h3c9510d8),
	.w3(32'hbc2da359),
	.w4(32'h3c9344dd),
	.w5(32'h3beba541),
	.w6(32'hbc91e849),
	.w7(32'hbc316ea5),
	.w8(32'hbc32f1b6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398c30),
	.w1(32'hbc00d9de),
	.w2(32'hbb10cf5f),
	.w3(32'hba8c05e2),
	.w4(32'hbc587e34),
	.w5(32'hbb626106),
	.w6(32'hbc283711),
	.w7(32'hbc46bb2c),
	.w8(32'h3c048fd0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb765d),
	.w1(32'h3c5db560),
	.w2(32'hbd0117b1),
	.w3(32'hbbdbfc08),
	.w4(32'h3992d72f),
	.w5(32'hbd54b002),
	.w6(32'h3cca14dd),
	.w7(32'hbc827533),
	.w8(32'hbd662cd8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d6fcf),
	.w1(32'h39b79733),
	.w2(32'hbb133b5e),
	.w3(32'hbd39686f),
	.w4(32'h3ca97a75),
	.w5(32'hbc419269),
	.w6(32'hbd438676),
	.w7(32'h3c98455b),
	.w8(32'h3b422e22),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f368b),
	.w1(32'hbb2fb9b4),
	.w2(32'hbb70de9a),
	.w3(32'hbce312f0),
	.w4(32'hbaf763b4),
	.w5(32'hbb6bd9db),
	.w6(32'hbce4fcfa),
	.w7(32'h3bc27006),
	.w8(32'h3b56ab5b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8fb1c),
	.w1(32'h3c55ac2b),
	.w2(32'h3c35e7a4),
	.w3(32'h3bc050b3),
	.w4(32'h3c23b76b),
	.w5(32'h3c955f88),
	.w6(32'h3bec1984),
	.w7(32'h3bb19476),
	.w8(32'h3c3f9f3b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ef1a2),
	.w1(32'hbbcc0c62),
	.w2(32'h3abad566),
	.w3(32'hbc5a0a62),
	.w4(32'hbb9fd42c),
	.w5(32'hba9601ca),
	.w6(32'hbc2412dc),
	.w7(32'hbba151aa),
	.w8(32'h39694afa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc903ce),
	.w1(32'hb9f49174),
	.w2(32'hbc27a284),
	.w3(32'hbacbf490),
	.w4(32'h3bebc03f),
	.w5(32'h3b254b50),
	.w6(32'h3a0f9d74),
	.w7(32'h3ba39ae1),
	.w8(32'hba9970bf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b9216),
	.w1(32'h3c17a5b5),
	.w2(32'h3c5e1d4d),
	.w3(32'h3bb0ff75),
	.w4(32'h3c64e7cf),
	.w5(32'h3b81a632),
	.w6(32'h3b9c9888),
	.w7(32'hbbd73648),
	.w8(32'hbba0c232),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7daf1),
	.w1(32'h3c77f20a),
	.w2(32'h3c5fd5cb),
	.w3(32'hba23c003),
	.w4(32'h3c38053a),
	.w5(32'h3c8623f5),
	.w6(32'hbac6ba7d),
	.w7(32'hbc91390c),
	.w8(32'hbc2873db),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53aa20),
	.w1(32'hbc98c71c),
	.w2(32'hbd23dfd0),
	.w3(32'hbb827c33),
	.w4(32'hbd242398),
	.w5(32'hbd36ffb9),
	.w6(32'hbc498076),
	.w7(32'hbcba72e3),
	.w8(32'hbcff92dd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba987e79),
	.w1(32'h3c0486c1),
	.w2(32'h3b49d81d),
	.w3(32'h3cca6735),
	.w4(32'h3bdad221),
	.w5(32'h3b9b9dd8),
	.w6(32'h3c3c61b8),
	.w7(32'h3ad547a9),
	.w8(32'hbb070ed9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba3d18),
	.w1(32'h3af7a06e),
	.w2(32'hbb4fbaf7),
	.w3(32'hba15030d),
	.w4(32'hbbca0b08),
	.w5(32'hbc72b0d2),
	.w6(32'hbb72b237),
	.w7(32'hbb7880a1),
	.w8(32'hbbf38fcf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846aac),
	.w1(32'h3c8849a0),
	.w2(32'hbbc4d3c5),
	.w3(32'hbba432df),
	.w4(32'h3b6dff87),
	.w5(32'hbb94534b),
	.w6(32'h3b86172b),
	.w7(32'h3b4ae54e),
	.w8(32'h3b2262da),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8a85),
	.w1(32'h3c14f3aa),
	.w2(32'h3c1cd653),
	.w3(32'hbbb4a144),
	.w4(32'h3baec34f),
	.w5(32'h3ba898d9),
	.w6(32'h3c2d8a61),
	.w7(32'h3b9837f8),
	.w8(32'h3b239793),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960287),
	.w1(32'h3c30c374),
	.w2(32'hbd08ce53),
	.w3(32'h39451767),
	.w4(32'hbd1ba36f),
	.w5(32'hbda52b2a),
	.w6(32'h3b189c45),
	.w7(32'hbdab24a0),
	.w8(32'hbdaca2f3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd965edc),
	.w1(32'hbc00492f),
	.w2(32'hbb7a8558),
	.w3(32'hbdaaec71),
	.w4(32'h39afbe3e),
	.w5(32'h3c536623),
	.w6(32'hbc708a85),
	.w7(32'h3c68cbe5),
	.w8(32'h3cace0cc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28192f),
	.w1(32'h3b24e487),
	.w2(32'hbd19c8b7),
	.w3(32'h3c752ca1),
	.w4(32'hbc1c3b9e),
	.w5(32'hbd6d4827),
	.w6(32'h3c5bb462),
	.w7(32'h3c2868da),
	.w8(32'hbd086e76),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a4f8d),
	.w1(32'hbb9f56cb),
	.w2(32'h3af97bd6),
	.w3(32'hbcc57439),
	.w4(32'h3b02876f),
	.w5(32'h3c15b018),
	.w6(32'hbcfccd7d),
	.w7(32'h3acf50dc),
	.w8(32'h3b921c2f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24b79),
	.w1(32'hbc251d8a),
	.w2(32'hb9a844b2),
	.w3(32'h3bbeccb5),
	.w4(32'hbbd25523),
	.w5(32'hbc695552),
	.w6(32'h3a8a4a83),
	.w7(32'hbc91c3d5),
	.w8(32'hbc3cebad),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7040e1),
	.w1(32'h3c1f25fe),
	.w2(32'h3c082c30),
	.w3(32'hbc0f24e9),
	.w4(32'h3c050401),
	.w5(32'h3c06c0b8),
	.w6(32'hbaf9abc2),
	.w7(32'h3c14dadf),
	.w8(32'h3c054825),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b25a6),
	.w1(32'hbbc09e21),
	.w2(32'h3b79a6c5),
	.w3(32'h3b792e31),
	.w4(32'hbc29c05c),
	.w5(32'hbb33e09d),
	.w6(32'h3a7bc3f4),
	.w7(32'hbc004b79),
	.w8(32'hbb154a1c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a183485),
	.w1(32'hbb5520d4),
	.w2(32'h3b5f4cf9),
	.w3(32'hbbbcf256),
	.w4(32'hba6dce94),
	.w5(32'h3bc7ec2e),
	.w6(32'hbb674ee4),
	.w7(32'hba9da55b),
	.w8(32'h3b47ceb6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed8913),
	.w1(32'hbc2564c5),
	.w2(32'hbb9e005d),
	.w3(32'h3b197846),
	.w4(32'hbc27acb5),
	.w5(32'hbbe9fbae),
	.w6(32'h3a8b2de5),
	.w7(32'hbbb46a61),
	.w8(32'hbbadecf8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6558f),
	.w1(32'hb9ad8416),
	.w2(32'h3b1902a4),
	.w3(32'hbb096bee),
	.w4(32'h3b3c848a),
	.w5(32'h3c154ae9),
	.w6(32'hbb20b2c4),
	.w7(32'h3b4a38c7),
	.w8(32'h3bf72dba),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf0d10),
	.w1(32'hba8a1b68),
	.w2(32'hbc1377dd),
	.w3(32'h3c6b44c1),
	.w4(32'h3bdeccf0),
	.w5(32'hbb0d947e),
	.w6(32'h3c28e052),
	.w7(32'h3c3c4dd2),
	.w8(32'hbc11212c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc367ae6),
	.w1(32'h3b40995b),
	.w2(32'h3acdcef6),
	.w3(32'hbbecf283),
	.w4(32'h3b3f89de),
	.w5(32'hbb0e6afe),
	.w6(32'hbc2ac209),
	.w7(32'hbb7333e0),
	.w8(32'hba7b0c8a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3c5e1),
	.w1(32'h3bd6564c),
	.w2(32'h3b5386dc),
	.w3(32'h3b08dd09),
	.w4(32'hbc48327b),
	.w5(32'hbbefa338),
	.w6(32'h3a977f60),
	.w7(32'h3b5314c9),
	.w8(32'h3bbf2ee3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64c7ca),
	.w1(32'hba9d1b0b),
	.w2(32'hba34bd71),
	.w3(32'h3ba9dd15),
	.w4(32'hba0a5b45),
	.w5(32'hbb45fc39),
	.w6(32'hbbd2c939),
	.w7(32'h3a6885c9),
	.w8(32'hbb1d531a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf960a3),
	.w1(32'h3cab669e),
	.w2(32'h3ccf8b54),
	.w3(32'hb9114f83),
	.w4(32'h3c5f0dc1),
	.w5(32'h3c9a8ac2),
	.w6(32'hbb60fad9),
	.w7(32'h3bd656fb),
	.w8(32'h3b077c72),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810eaf),
	.w1(32'hbb23a050),
	.w2(32'hbb68e409),
	.w3(32'h3c770fc1),
	.w4(32'hbbdef7dd),
	.w5(32'hbc08da32),
	.w6(32'hbab41567),
	.w7(32'hbb523965),
	.w8(32'hbbbd292c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5d3aa),
	.w1(32'h3b34d19c),
	.w2(32'h3c174325),
	.w3(32'hbc116cc2),
	.w4(32'h3ad8d0c0),
	.w5(32'h3a693505),
	.w6(32'hbc36344a),
	.w7(32'hbb92b1d8),
	.w8(32'h3c4c6cf1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b8aa5),
	.w1(32'h3cb2f490),
	.w2(32'h3c984b7c),
	.w3(32'hbb64fbc1),
	.w4(32'hbb6d62aa),
	.w5(32'hbcf9a7e0),
	.w6(32'h3bacc23f),
	.w7(32'h3c13f49c),
	.w8(32'h3b24dcc4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56b6bb),
	.w1(32'hba908d1e),
	.w2(32'hbb4ae57c),
	.w3(32'h3a4cb747),
	.w4(32'h3a4f6fe3),
	.w5(32'h3ac1136f),
	.w6(32'hbc193325),
	.w7(32'h3b3e8387),
	.w8(32'h3a9dc865),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a89c4),
	.w1(32'h3bb55514),
	.w2(32'h3bb2b72c),
	.w3(32'hba2b58d7),
	.w4(32'h3c04d33d),
	.w5(32'h3b7e2693),
	.w6(32'hbb997ecb),
	.w7(32'hbab4839d),
	.w8(32'h3aacc409),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f190),
	.w1(32'hbc57ce14),
	.w2(32'hbbb2dc38),
	.w3(32'h3ba03a39),
	.w4(32'hbba9276e),
	.w5(32'hbc8d0476),
	.w6(32'hbad43e70),
	.w7(32'h3c0cb52a),
	.w8(32'h3b990de1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ac04),
	.w1(32'h3b01dd6f),
	.w2(32'h3c929aec),
	.w3(32'hbc8e9c6c),
	.w4(32'hbc7dc67d),
	.w5(32'hbc18f2e4),
	.w6(32'hba706e2e),
	.w7(32'h3bb165c3),
	.w8(32'h3c5c1d8e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b4d7f),
	.w1(32'h3b56f03f),
	.w2(32'h3a01ba4c),
	.w3(32'hbbbeb212),
	.w4(32'h3ba04d3f),
	.w5(32'h3b71cf68),
	.w6(32'h3bc74835),
	.w7(32'h3b9ad04d),
	.w8(32'h3b56ca22),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2a214),
	.w1(32'hbd2ffb70),
	.w2(32'h3d10fa74),
	.w3(32'h3b9fc42a),
	.w4(32'h3ce4dd08),
	.w5(32'hbda2dba0),
	.w6(32'h3b0ba1c7),
	.w7(32'hbb88a754),
	.w8(32'h3c9f379f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c640c77),
	.w1(32'h3a7f2013),
	.w2(32'hb8fcd777),
	.w3(32'hbd83db6d),
	.w4(32'h3bd68e69),
	.w5(32'h3b191cb9),
	.w6(32'h3d2e9a28),
	.w7(32'h3b16eaf0),
	.w8(32'h3ba0219e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b896d07),
	.w1(32'hb9de2458),
	.w2(32'hbb724963),
	.w3(32'h3c12983a),
	.w4(32'h3bdba947),
	.w5(32'h3bf68a52),
	.w6(32'h3b9bb5b6),
	.w7(32'h3b86fc08),
	.w8(32'hbb4e96fa),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d12c),
	.w1(32'hbc8efca6),
	.w2(32'hba764dab),
	.w3(32'hbab5fbb5),
	.w4(32'hbb0de480),
	.w5(32'hbb8b2098),
	.w6(32'hbbaf33e6),
	.w7(32'h3a8d75fb),
	.w8(32'h39d7b19e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dbe90),
	.w1(32'hbd88627b),
	.w2(32'h3c12bf1e),
	.w3(32'hbc691bb2),
	.w4(32'h3da558a8),
	.w5(32'h3cb1d278),
	.w6(32'hbaaa8b37),
	.w7(32'hbcbbfb0c),
	.w8(32'hbce0af92),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa3647),
	.w1(32'h3ab436a4),
	.w2(32'h3b0583f4),
	.w3(32'hbda35f15),
	.w4(32'h39fcbe8d),
	.w5(32'h3b071d71),
	.w6(32'h3d4226e7),
	.w7(32'h3b08507c),
	.w8(32'h3afa339e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f9d74),
	.w1(32'hbc145fe7),
	.w2(32'hbbb4d909),
	.w3(32'h3b552648),
	.w4(32'hbbf6b7b0),
	.w5(32'hbc14b163),
	.w6(32'h3af80280),
	.w7(32'h3bd4b8fa),
	.w8(32'hbbe1e943),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb374197),
	.w1(32'h3ac89119),
	.w2(32'h3b9a1015),
	.w3(32'hbc30c427),
	.w4(32'h3bb816d4),
	.w5(32'h3ad8831a),
	.w6(32'hba0d6934),
	.w7(32'hbb033ee8),
	.w8(32'h3bc8d397),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a96cd),
	.w1(32'hbb010837),
	.w2(32'h3ab89c14),
	.w3(32'hbb62202b),
	.w4(32'hb9ea0ad9),
	.w5(32'h3a849b06),
	.w6(32'h3b381034),
	.w7(32'h3b0c8afe),
	.w8(32'hb826fc2a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7da378),
	.w1(32'h3c83587b),
	.w2(32'h3ceff384),
	.w3(32'hbaae3ee2),
	.w4(32'h3d3287d8),
	.w5(32'hbd352328),
	.w6(32'h3b4ee8b4),
	.w7(32'hbd030e7d),
	.w8(32'h3d188641),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba1591),
	.w1(32'hbbf0f43b),
	.w2(32'hbc11278d),
	.w3(32'h3cda8feb),
	.w4(32'hbb53e9c7),
	.w5(32'h3b6d00cd),
	.w6(32'h3d32bb27),
	.w7(32'hbbc4067e),
	.w8(32'hbc01fc89),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a69e6),
	.w1(32'hbb8a9bcc),
	.w2(32'hbbbd55ad),
	.w3(32'hbaebca1e),
	.w4(32'h3a181be7),
	.w5(32'h3b23e566),
	.w6(32'hbbf795f3),
	.w7(32'hb982b3cc),
	.w8(32'hbb6f525f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a76a),
	.w1(32'hbc364517),
	.w2(32'hbc871e94),
	.w3(32'hbab9f169),
	.w4(32'hbc485e04),
	.w5(32'hbcf033fd),
	.w6(32'hbb4db128),
	.w7(32'hbc0983f8),
	.w8(32'hbc11a1a6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85f6d7),
	.w1(32'h3b7b0c0c),
	.w2(32'hbb931331),
	.w3(32'hbb3a3ae1),
	.w4(32'hbad83567),
	.w5(32'h3c3cbc58),
	.w6(32'hbbebcd66),
	.w7(32'h3b51ee0a),
	.w8(32'hb9c1538e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aff90),
	.w1(32'h3b2b6930),
	.w2(32'h3abefb0d),
	.w3(32'h3c135e83),
	.w4(32'h3b921f3c),
	.w5(32'h3a722abe),
	.w6(32'h3b666d7a),
	.w7(32'h3a91619c),
	.w8(32'h3aba2344),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a852c36),
	.w1(32'hbb3f16e5),
	.w2(32'h380a4f96),
	.w3(32'hba0e3442),
	.w4(32'hb91de0c2),
	.w5(32'hbbb24c9e),
	.w6(32'hbac9999b),
	.w7(32'hbc025160),
	.w8(32'hbb6fb8b2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b1a06),
	.w1(32'h3a27191a),
	.w2(32'hbb309ffe),
	.w3(32'h3be13042),
	.w4(32'h39b7a621),
	.w5(32'hbab198f7),
	.w6(32'hbc82d4d3),
	.w7(32'h390b2a99),
	.w8(32'h3adf796f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83e779),
	.w1(32'h3b589db3),
	.w2(32'hbbd76bd2),
	.w3(32'hbb170a78),
	.w4(32'h3b91b66c),
	.w5(32'h3b2e6b3b),
	.w6(32'hba1511ea),
	.w7(32'h3c0c0bb7),
	.w8(32'h3b8bb0d2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae64365),
	.w1(32'h3cc6051a),
	.w2(32'hbac6db61),
	.w3(32'hbbc69dd1),
	.w4(32'hbbbb6f79),
	.w5(32'hbc4f7e3a),
	.w6(32'hb9bb31aa),
	.w7(32'h3bc6ffcc),
	.w8(32'hbbb8c183),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e4f9),
	.w1(32'h3ca0e987),
	.w2(32'hbc80dd28),
	.w3(32'hbb6f421c),
	.w4(32'hbc406807),
	.w5(32'h3cd7dd95),
	.w6(32'hbb6b1570),
	.w7(32'hbbd09c7d),
	.w8(32'hbb9f2bff),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc969703),
	.w1(32'hbb7f60d1),
	.w2(32'hbbaffcba),
	.w3(32'h3ce60a25),
	.w4(32'hbc73c052),
	.w5(32'h3b8e5ba1),
	.w6(32'hbc87693f),
	.w7(32'h3bbb2647),
	.w8(32'h3c4ed23e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb21a47),
	.w1(32'h3b98ef18),
	.w2(32'hbc30f03f),
	.w3(32'h3c80abc3),
	.w4(32'hbae0189c),
	.w5(32'hbc1a339e),
	.w6(32'hbb73e32a),
	.w7(32'hbbf8857d),
	.w8(32'hbb79203e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1f9b2),
	.w1(32'h3b991970),
	.w2(32'h376a9e42),
	.w3(32'hbc0ebb7d),
	.w4(32'h3c186913),
	.w5(32'h3ba2bf66),
	.w6(32'hbc076aa5),
	.w7(32'hbbc74b07),
	.w8(32'h3addfc6e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab06895),
	.w1(32'h3aba9bf0),
	.w2(32'h3a1969c5),
	.w3(32'h3c641758),
	.w4(32'h3b6854fe),
	.w5(32'h3b87080f),
	.w6(32'h3bc47fa2),
	.w7(32'h3b26fb0b),
	.w8(32'h3b677f24),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b572094),
	.w1(32'h3b8e27b8),
	.w2(32'h3b5c0034),
	.w3(32'h3ab0f2d6),
	.w4(32'h3bcdc52c),
	.w5(32'h3b998ac0),
	.w6(32'h3a6c347d),
	.w7(32'h3bd30dd7),
	.w8(32'h3bc64614),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd46e),
	.w1(32'h3c42c3ed),
	.w2(32'h3b89e87b),
	.w3(32'h39acf847),
	.w4(32'h3c15faaf),
	.w5(32'h3d691464),
	.w6(32'h3b6f22f9),
	.w7(32'h3d2266f9),
	.w8(32'h3c15e432),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3c94a),
	.w1(32'hbaaa5cea),
	.w2(32'hbb87bf7c),
	.w3(32'h3c6771bb),
	.w4(32'hb96f9a38),
	.w5(32'hbb4f6286),
	.w6(32'h3c242add),
	.w7(32'h3c9e813d),
	.w8(32'hbc7d5e5e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce02f0),
	.w1(32'hbca01995),
	.w2(32'hbc9f5b33),
	.w3(32'h3a576de7),
	.w4(32'hbbba685b),
	.w5(32'h3c6a9552),
	.w6(32'hbaf95b75),
	.w7(32'h3a84798f),
	.w8(32'hbc402f54),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e1649),
	.w1(32'hbc51b84c),
	.w2(32'hbcb3cf03),
	.w3(32'h3c196a3c),
	.w4(32'hbb8794e5),
	.w5(32'h3c8e8bc5),
	.w6(32'hbc0a6f00),
	.w7(32'h3c020fe4),
	.w8(32'hbc539192),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2403f2),
	.w1(32'hbc49ef3e),
	.w2(32'h3c72a555),
	.w3(32'h3b9d63d0),
	.w4(32'h3cbe773c),
	.w5(32'hbce7773a),
	.w6(32'hbc1391cc),
	.w7(32'hbc8602bc),
	.w8(32'h3cca3683),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c5449),
	.w1(32'h3b1f62dc),
	.w2(32'h3afc72b8),
	.w3(32'h3c81b026),
	.w4(32'h3a7fe451),
	.w5(32'hbb60eeaa),
	.w6(32'hbc4bafd2),
	.w7(32'hb9a6f3ea),
	.w8(32'h3a2813c2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf29db),
	.w1(32'h3c34c5b3),
	.w2(32'hbb80abb7),
	.w3(32'h3a8a5679),
	.w4(32'h3b6b038c),
	.w5(32'h3963a63a),
	.w6(32'h3ae6ab92),
	.w7(32'hba5db277),
	.w8(32'hbaff1b10),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe0d4a),
	.w1(32'h374e4e26),
	.w2(32'h3b7d256a),
	.w3(32'h3c122cbf),
	.w4(32'h3b39168e),
	.w5(32'hbc36dc84),
	.w6(32'hbad2b204),
	.w7(32'hbbf52a43),
	.w8(32'hb9be9eb1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991dc10),
	.w1(32'h3b2ae7c7),
	.w2(32'h3baae111),
	.w3(32'h3b3fe111),
	.w4(32'h3b3e43f9),
	.w5(32'h3b42dc1a),
	.w6(32'h3abafb29),
	.w7(32'h3b95a36b),
	.w8(32'h3bde7f99),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56e97e),
	.w1(32'hbbec57de),
	.w2(32'hbc11c580),
	.w3(32'h3b18eecc),
	.w4(32'h3b8f20c9),
	.w5(32'h3c1e9f44),
	.w6(32'h3a4f07cf),
	.w7(32'hbc42b1b6),
	.w8(32'hbacd351f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0d16),
	.w1(32'hbd80b38c),
	.w2(32'hbcbdd0da),
	.w3(32'h3c44bef6),
	.w4(32'h3d92c15c),
	.w5(32'h3d030b7e),
	.w6(32'h3bac3846),
	.w7(32'hbb9a112d),
	.w8(32'hbc204f92),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a4372),
	.w1(32'hbc96790e),
	.w2(32'h39a2d0c5),
	.w3(32'hbd190e3e),
	.w4(32'h3c85deb4),
	.w5(32'h3c054a6c),
	.w6(32'h3c8a50f0),
	.w7(32'h3c1d3881),
	.w8(32'hbbad1016),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d331e),
	.w1(32'h3b4bcd1e),
	.w2(32'h3a0727ba),
	.w3(32'hbcc7aca5),
	.w4(32'h3a8c268d),
	.w5(32'h3acc6804),
	.w6(32'h3cd4ad37),
	.w7(32'h3b0dbbc8),
	.w8(32'hb94eb6da),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2720f4),
	.w1(32'hba32416d),
	.w2(32'h3b722794),
	.w3(32'h39e04c7c),
	.w4(32'h3bd20d6c),
	.w5(32'h3a1a1a28),
	.w6(32'hbb9d4975),
	.w7(32'hbbd34510),
	.w8(32'hbbbe263a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab35491),
	.w1(32'hbb48468c),
	.w2(32'hbb31f4df),
	.w3(32'h3ad3136b),
	.w4(32'h3b57efdf),
	.w5(32'h37a80909),
	.w6(32'hbb924014),
	.w7(32'hbc00d988),
	.w8(32'hbbfc3363),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9f08),
	.w1(32'hbb32d06c),
	.w2(32'hba8b8869),
	.w3(32'hb8df327b),
	.w4(32'hbac45077),
	.w5(32'h39c4151a),
	.w6(32'hbbe9aaa5),
	.w7(32'h3abccc8c),
	.w8(32'hba805b80),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9b16a),
	.w1(32'hbba70cc1),
	.w2(32'hbc7f3346),
	.w3(32'hba7b378b),
	.w4(32'hbcbd906f),
	.w5(32'hbc8dc593),
	.w6(32'hbb813ac8),
	.w7(32'h38ca981f),
	.w8(32'hbc1fd99a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392759f7),
	.w1(32'hbc283eba),
	.w2(32'hbb7ac407),
	.w3(32'hba579281),
	.w4(32'hbb7a175f),
	.w5(32'h3bd9041e),
	.w6(32'hbc74e29b),
	.w7(32'h3c4ebc9d),
	.w8(32'h3be16ec5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d7639),
	.w1(32'h3c459cfd),
	.w2(32'hbc4cc73a),
	.w3(32'h398bab4e),
	.w4(32'h3b59086d),
	.w5(32'h3bb5ce1e),
	.w6(32'h3c206583),
	.w7(32'hbc3e8fc6),
	.w8(32'h3c210f82),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f97f4),
	.w1(32'h39f3f0b2),
	.w2(32'h3adf6d72),
	.w3(32'h3c04e04e),
	.w4(32'h3a322706),
	.w5(32'hba712594),
	.w6(32'hbc16af86),
	.w7(32'h3b50fd1d),
	.w8(32'hbb1ee5a0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d75fe),
	.w1(32'h3d6e6622),
	.w2(32'h3c566f71),
	.w3(32'hbb339889),
	.w4(32'hbda4ca7c),
	.w5(32'hbc853b10),
	.w6(32'hbad25498),
	.w7(32'h3cabf6a5),
	.w8(32'h3cd6e807),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule