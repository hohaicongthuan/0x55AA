module layer_8_featuremap_59(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5576),
	.w1(32'hbb19c69a),
	.w2(32'h39b6f828),
	.w3(32'hba982b00),
	.w4(32'hbb5c8fad),
	.w5(32'h39fd3dc6),
	.w6(32'hb9f89fbb),
	.w7(32'h3b48eb74),
	.w8(32'hbb524544),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae147e4),
	.w1(32'hbb1abc01),
	.w2(32'hbb0e1d0f),
	.w3(32'hb7ea819f),
	.w4(32'hbb52339c),
	.w5(32'h39d0347f),
	.w6(32'h3ad24ed8),
	.w7(32'h3a84b5d9),
	.w8(32'hbaf331ec),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157523),
	.w1(32'h3aa9d323),
	.w2(32'h39705476),
	.w3(32'h3acc43f6),
	.w4(32'h395b4003),
	.w5(32'h3abf487a),
	.w6(32'h3aec589c),
	.w7(32'h3b37d614),
	.w8(32'h3a1217aa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d375a),
	.w1(32'h3c9232be),
	.w2(32'hbc740ce4),
	.w3(32'h3c2a550a),
	.w4(32'h3c4b465f),
	.w5(32'h3bd3fe2f),
	.w6(32'h3c0f1f83),
	.w7(32'hbc246e2a),
	.w8(32'hbb1ef996),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06e97a),
	.w1(32'hba9a0a6b),
	.w2(32'hbbb2d6de),
	.w3(32'h3a4a5730),
	.w4(32'hbb6a9259),
	.w5(32'hbbb6447a),
	.w6(32'h3ae0fbe7),
	.w7(32'h3a0b36f1),
	.w8(32'h3cb09da5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3b98f),
	.w1(32'hbc0119bb),
	.w2(32'hbcac4017),
	.w3(32'hb8e51666),
	.w4(32'hbcbdfdfc),
	.w5(32'hbbf768c8),
	.w6(32'h3cc1ba69),
	.w7(32'hbab50795),
	.w8(32'hbbc8738a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21ee93),
	.w1(32'hbb79d987),
	.w2(32'hbb133f44),
	.w3(32'h3b8c6e6b),
	.w4(32'h3a62acfc),
	.w5(32'h3a52139f),
	.w6(32'h39bbd547),
	.w7(32'h3b646de5),
	.w8(32'hbb3cede9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37240e),
	.w1(32'hb93aed7f),
	.w2(32'hbbbf2b41),
	.w3(32'hba10a64f),
	.w4(32'hbb71c19e),
	.w5(32'hbbcc9cbd),
	.w6(32'h3a850020),
	.w7(32'hba3b1d67),
	.w8(32'hbc068adb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6220a),
	.w1(32'hbb0b6928),
	.w2(32'hb98899e8),
	.w3(32'h3ab46a66),
	.w4(32'hbb04aa66),
	.w5(32'h3b0e4060),
	.w6(32'h3a703e49),
	.w7(32'h3bf6f6dd),
	.w8(32'hbbc3bce8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2123c4),
	.w1(32'h3cff98df),
	.w2(32'h3ccd4b8a),
	.w3(32'h3c1be1d1),
	.w4(32'hbc83f2ed),
	.w5(32'hbc751b3f),
	.w6(32'hbc6cf490),
	.w7(32'hbbd2a9ce),
	.w8(32'hbb1a4bbf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17d489),
	.w1(32'h3b89b00d),
	.w2(32'h3b74e5ad),
	.w3(32'h3af8e568),
	.w4(32'h3ad6c8fc),
	.w5(32'h3bbae5eb),
	.w6(32'h3be96b47),
	.w7(32'h3bac2fd1),
	.w8(32'hbb90e25b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97963c),
	.w1(32'hbaee6acc),
	.w2(32'hbb65819f),
	.w3(32'h3ad48c79),
	.w4(32'hbb4005ab),
	.w5(32'h3a38f1c2),
	.w6(32'h3a87c050),
	.w7(32'h3a89580f),
	.w8(32'hbb8d045d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb3684),
	.w1(32'hbb76873a),
	.w2(32'hbabd1604),
	.w3(32'h3b20bdbb),
	.w4(32'h3a8c51ea),
	.w5(32'h3baeab26),
	.w6(32'h3a3fe7e3),
	.w7(32'h3b6b3454),
	.w8(32'h3ccc8a13),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccca329),
	.w1(32'hbc320864),
	.w2(32'hbcc68227),
	.w3(32'h3ae674c5),
	.w4(32'hbcd16e73),
	.w5(32'hbbf848cc),
	.w6(32'h3cd6e193),
	.w7(32'hbae1b45c),
	.w8(32'h3c22c29d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9419ec),
	.w1(32'hbb6ec574),
	.w2(32'hbc7da225),
	.w3(32'h3a50f9ae),
	.w4(32'hbc8c1535),
	.w5(32'hbc4dbc2c),
	.w6(32'h3c91df24),
	.w7(32'hbb9344b5),
	.w8(32'h3ab4f8bb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a00cf8),
	.w1(32'hbb0b70bc),
	.w2(32'h3b16d54b),
	.w3(32'hbb8ed2f6),
	.w4(32'hbbf71873),
	.w5(32'h3b8ff7d5),
	.w6(32'h3b665c33),
	.w7(32'hbad8c3f2),
	.w8(32'hbb288c7e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0c911),
	.w1(32'h3ca5ff41),
	.w2(32'h3c431464),
	.w3(32'hbc3b111b),
	.w4(32'hbab5b83a),
	.w5(32'hbc818f60),
	.w6(32'hbb8bb785),
	.w7(32'h39c5e312),
	.w8(32'hbbc85cb0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f468),
	.w1(32'hbb0092af),
	.w2(32'hbb74dc8b),
	.w3(32'hb6fdc3d1),
	.w4(32'hba76d760),
	.w5(32'h3b87f38a),
	.w6(32'hbb66a237),
	.w7(32'hb900f4be),
	.w8(32'hbc19017d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a314c),
	.w1(32'hbb9d5cde),
	.w2(32'hbb93f69c),
	.w3(32'hbbc3c24d),
	.w4(32'hbc2364bd),
	.w5(32'h3b654d2d),
	.w6(32'hbc2c130c),
	.w7(32'hbb634625),
	.w8(32'hbc10a94e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a03a9),
	.w1(32'h3b21eb66),
	.w2(32'hbd0c3f6b),
	.w3(32'hbcc28a72),
	.w4(32'hbd1cd6d8),
	.w5(32'hbbce2e48),
	.w6(32'hbc414fe1),
	.w7(32'hbc7e9a5a),
	.w8(32'hbaaa621c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185aab),
	.w1(32'h3a9c59d7),
	.w2(32'hbaf4803b),
	.w3(32'h3b2c9840),
	.w4(32'h3bb42a0a),
	.w5(32'hbbc1bc67),
	.w6(32'hbb45c314),
	.w7(32'hb8d006ad),
	.w8(32'h3b07d741),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38dfd),
	.w1(32'hbbbd6c33),
	.w2(32'hbbf08c10),
	.w3(32'h3b9fcb4c),
	.w4(32'hbb9f69c9),
	.w5(32'hbbe6141a),
	.w6(32'h3b546c12),
	.w7(32'h3b61a8f7),
	.w8(32'hbbf787ec),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9be994),
	.w1(32'hbc31b32c),
	.w2(32'h3c31b736),
	.w3(32'h3c64d6ca),
	.w4(32'h3cc30b68),
	.w5(32'h3c6c306b),
	.w6(32'hbcc1b62d),
	.w7(32'h3b98b5b5),
	.w8(32'hbc6dfdea),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e79c),
	.w1(32'hbaf682be),
	.w2(32'h3aca28fe),
	.w3(32'hbc28d40f),
	.w4(32'hbc0291c0),
	.w5(32'h3a96a75e),
	.w6(32'h3a460068),
	.w7(32'h3b4ce052),
	.w8(32'h3c4b7724),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301100),
	.w1(32'hbba2bd4d),
	.w2(32'hbbff3e81),
	.w3(32'hbb2281e9),
	.w4(32'hbafd7a63),
	.w5(32'hbc276a4b),
	.w6(32'h3b2e4b1d),
	.w7(32'h3a696024),
	.w8(32'hbbe5f537),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9349ff),
	.w1(32'hbc2f55ff),
	.w2(32'h3c3301a4),
	.w3(32'h3c5915cd),
	.w4(32'h3cb9e0d4),
	.w5(32'h3c6a054b),
	.w6(32'hbcb4b317),
	.w7(32'h3b976ac7),
	.w8(32'hbbdcf2d3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79f2d7),
	.w1(32'hbc0f4509),
	.w2(32'h3c1e807b),
	.w3(32'h3c3b80e7),
	.w4(32'h3ca04ea3),
	.w5(32'h3c4b04fa),
	.w6(32'hbc956efe),
	.w7(32'h3b9a8b04),
	.w8(32'hbb95d3bc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab225a),
	.w1(32'hbbcea83e),
	.w2(32'hbbf073f2),
	.w3(32'h3c350fba),
	.w4(32'h3b6a165c),
	.w5(32'hbc224970),
	.w6(32'hbbcbcc84),
	.w7(32'hbb2de791),
	.w8(32'h3ca6a819),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be97d70),
	.w1(32'h3bfbf39c),
	.w2(32'h3ca51dd8),
	.w3(32'hbcb27bf9),
	.w4(32'hbd179c1b),
	.w5(32'h3bf58466),
	.w6(32'h3b3fe9e2),
	.w7(32'hbd06e2c8),
	.w8(32'hba6edbb7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c08b6),
	.w1(32'h39fe8c48),
	.w2(32'h388dfbe7),
	.w3(32'h3a8293ea),
	.w4(32'hba85bb6f),
	.w5(32'h3ad8a0d1),
	.w6(32'h3b1c727a),
	.w7(32'h3ad35ffa),
	.w8(32'h3a6c933e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb6c1d),
	.w1(32'h3c347277),
	.w2(32'hbc47a4d3),
	.w3(32'hbd055448),
	.w4(32'hb964adfc),
	.w5(32'h3b36e253),
	.w6(32'h3bb486e6),
	.w7(32'hbc73fac3),
	.w8(32'hbb8a22fb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc566530),
	.w1(32'hbbd6a014),
	.w2(32'h3b967d1c),
	.w3(32'h3baecefb),
	.w4(32'h3bc56c94),
	.w5(32'hbbfb0e0e),
	.w6(32'h3b00e144),
	.w7(32'h3c477ccd),
	.w8(32'h3c26a6d6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c660a44),
	.w1(32'hb9f00147),
	.w2(32'hbcb8968d),
	.w3(32'hbc4ecc02),
	.w4(32'hbb1b06af),
	.w5(32'hbc0169ad),
	.w6(32'h3c649f93),
	.w7(32'hbc818922),
	.w8(32'hbbb67849),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9219c2),
	.w1(32'h3bb23317),
	.w2(32'hbb06a679),
	.w3(32'hbbf8cff1),
	.w4(32'hbbfeb3bd),
	.w5(32'h3c76082c),
	.w6(32'hbaaa5c60),
	.w7(32'hbc86ae66),
	.w8(32'h3cb43ea4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5a5da),
	.w1(32'hbc14f1eb),
	.w2(32'hbcaaecc6),
	.w3(32'h3acee28b),
	.w4(32'hbcb6bb13),
	.w5(32'hbbd2f864),
	.w6(32'h3cbe29fc),
	.w7(32'hba8d2fda),
	.w8(32'hbc3eca04),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd98f20),
	.w1(32'hbb75b56f),
	.w2(32'hbb658826),
	.w3(32'hbba9a223),
	.w4(32'hbbe84df3),
	.w5(32'h3a990bed),
	.w6(32'hbb7c6249),
	.w7(32'h3a3f05e3),
	.w8(32'h38437bb8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc4f95),
	.w1(32'h38de1b10),
	.w2(32'hbb478ca8),
	.w3(32'h3ae375b8),
	.w4(32'hbb01335e),
	.w5(32'hbc18bc1d),
	.w6(32'hbb04e57a),
	.w7(32'h3a1a2533),
	.w8(32'hb952c387),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc25b44),
	.w1(32'h3b31ae4b),
	.w2(32'h3abfcddd),
	.w3(32'h3b632f07),
	.w4(32'h396e013f),
	.w5(32'h3b006bae),
	.w6(32'h3b8cc04d),
	.w7(32'h3b96b50c),
	.w8(32'h3c8cb68f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d14ded4),
	.w1(32'hbbb7a4c6),
	.w2(32'hbd0a956f),
	.w3(32'h3b285063),
	.w4(32'hbd0253bb),
	.w5(32'hbcef5b39),
	.w6(32'h3d20023f),
	.w7(32'hbc33c56a),
	.w8(32'hbb897a80),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba35f3),
	.w1(32'hbafdc5a5),
	.w2(32'hbb4edfe3),
	.w3(32'h3bb13c7a),
	.w4(32'h3ae02097),
	.w5(32'hbbece378),
	.w6(32'hbb1ba605),
	.w7(32'h3ad9b433),
	.w8(32'hbb594af8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eda2e),
	.w1(32'hbb998940),
	.w2(32'h3b7dd01a),
	.w3(32'h3b1b3af5),
	.w4(32'h3be69725),
	.w5(32'h3b849d8a),
	.w6(32'hbc44412c),
	.w7(32'hba6348cc),
	.w8(32'hbbcbc3b1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48cef7),
	.w1(32'hbb81ce58),
	.w2(32'h3a7a453a),
	.w3(32'h39a9185b),
	.w4(32'h3a6340f0),
	.w5(32'hbb45cdcc),
	.w6(32'hbb04e7c0),
	.w7(32'h3b61dc83),
	.w8(32'h3bcd7c8c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb867),
	.w1(32'h3b4cad92),
	.w2(32'h3ae65af4),
	.w3(32'hbc9c7aea),
	.w4(32'hbc3509b8),
	.w5(32'hbaafe27f),
	.w6(32'hbad8945f),
	.w7(32'hbc82422a),
	.w8(32'hbc2b7acf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074c62),
	.w1(32'hbbab45ba),
	.w2(32'h3b362fc4),
	.w3(32'h3a5119d1),
	.w4(32'h3b8edfe5),
	.w5(32'h3b193e0f),
	.w6(32'hbc3e3d6c),
	.w7(32'hbacf11f8),
	.w8(32'hbc193456),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4318),
	.w1(32'hbb853ef3),
	.w2(32'h3b0aa590),
	.w3(32'h3a4a6f35),
	.w4(32'h3b6d2bbf),
	.w5(32'h3b03a86e),
	.w6(32'hbc1ecb43),
	.w7(32'hbb2e7374),
	.w8(32'h3b882f04),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba617b8e),
	.w1(32'hbb5c8a9e),
	.w2(32'hbbb8c7df),
	.w3(32'hba82b844),
	.w4(32'hbbe91ea3),
	.w5(32'hbc27f6b3),
	.w6(32'h3ace17b8),
	.w7(32'h3b051695),
	.w8(32'hbc96b36a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a962),
	.w1(32'hbbde51a3),
	.w2(32'hbca540c7),
	.w3(32'hbc7aa0e0),
	.w4(32'hbc61cd67),
	.w5(32'hbc619946),
	.w6(32'hbc2763ee),
	.w7(32'hbc815507),
	.w8(32'h3a61f62d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab12bdb),
	.w1(32'hbbb1e5de),
	.w2(32'hba24aa7a),
	.w3(32'h3b346f74),
	.w4(32'h3bdedd40),
	.w5(32'hbb231949),
	.w6(32'hbb5de7a2),
	.w7(32'h3a811b63),
	.w8(32'h3d337229),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d031f5f),
	.w1(32'h3b83c145),
	.w2(32'hbca99598),
	.w3(32'h3a85f52a),
	.w4(32'hbcdc4046),
	.w5(32'hbd10054c),
	.w6(32'h3cea69a0),
	.w7(32'h3b99daba),
	.w8(32'hbbe1e68c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11f10),
	.w1(32'hbbdc7b9e),
	.w2(32'h3aef8fbf),
	.w3(32'h3a79b85d),
	.w4(32'h3ad76d0c),
	.w5(32'h3aa22648),
	.w6(32'hbc1314c4),
	.w7(32'h3a01b3f5),
	.w8(32'hbc091a5f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06650),
	.w1(32'hbae3e033),
	.w2(32'h3b094100),
	.w3(32'hba235c60),
	.w4(32'h3b6141ef),
	.w5(32'h3b91a761),
	.w6(32'hbbb326b9),
	.w7(32'hba8253f6),
	.w8(32'hbc8c1921),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc646dab),
	.w1(32'hbb71b137),
	.w2(32'h3b8cb909),
	.w3(32'hbafae9c6),
	.w4(32'h3be56bd0),
	.w5(32'h3b8dab6f),
	.w6(32'hbc47afcf),
	.w7(32'hbba754ba),
	.w8(32'h3a6f6d6e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f1655),
	.w1(32'hb993a708),
	.w2(32'h3bf6bea9),
	.w3(32'hbaaf67ce),
	.w4(32'hbcb4a133),
	.w5(32'hbb9402a0),
	.w6(32'h3c8f48d3),
	.w7(32'h3c53b134),
	.w8(32'h3d241bef),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf77015),
	.w1(32'h3be7ed9d),
	.w2(32'hbc865510),
	.w3(32'h3baf4384),
	.w4(32'hbc8620d4),
	.w5(32'hbcffc3c1),
	.w6(32'h3cd06722),
	.w7(32'h3b3a51e1),
	.w8(32'hbb080403),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba508c03),
	.w1(32'hbc2fc966),
	.w2(32'hbbdf64b2),
	.w3(32'hbc7440ed),
	.w4(32'hbc168d7a),
	.w5(32'hb9c2efe9),
	.w6(32'hbcbe6961),
	.w7(32'hbca26d9e),
	.w8(32'h3c324b3b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f195e),
	.w1(32'h3b2a2676),
	.w2(32'h3c6c8d88),
	.w3(32'h3c38464e),
	.w4(32'h3c476789),
	.w5(32'h3bdd70ff),
	.w6(32'hbb445c8f),
	.w7(32'h3c135215),
	.w8(32'hbae54188),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a7fc),
	.w1(32'hbc0b8b9d),
	.w2(32'hbb03c05c),
	.w3(32'h3c07b329),
	.w4(32'hbc26abe7),
	.w5(32'hbbff593a),
	.w6(32'hbc8392e1),
	.w7(32'h3bd645ff),
	.w8(32'h3c16de26),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2f609),
	.w1(32'hbbd4d161),
	.w2(32'h3bc62507),
	.w3(32'hbb602abe),
	.w4(32'hbba4aa50),
	.w5(32'h3974d66d),
	.w6(32'hbc1621a7),
	.w7(32'h3bb22391),
	.w8(32'hbc3a4091),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7888e),
	.w1(32'hba1ca083),
	.w2(32'h3c823361),
	.w3(32'h3b45d111),
	.w4(32'h3c12f88f),
	.w5(32'h3c9abb1a),
	.w6(32'hbc06e51b),
	.w7(32'h3c069e39),
	.w8(32'h3bfaa502),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e8fe1),
	.w1(32'hbbf0d4f4),
	.w2(32'hbc369880),
	.w3(32'hbc0b8d5d),
	.w4(32'hbcb566cd),
	.w5(32'hbc922b9d),
	.w6(32'h3b185c99),
	.w7(32'hbb722cb3),
	.w8(32'hbc463a14),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc935cdc),
	.w1(32'h3b913293),
	.w2(32'hb99e1b27),
	.w3(32'hbacbd110),
	.w4(32'hbb9ea600),
	.w5(32'hbc4f80fb),
	.w6(32'hbc68cdfd),
	.w7(32'hbbf5d32e),
	.w8(32'h3b121706),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08b93c),
	.w1(32'hbc2701e0),
	.w2(32'hbbd5c705),
	.w3(32'hbb7bc00e),
	.w4(32'hbc08859a),
	.w5(32'hbc6093cd),
	.w6(32'hbb2d02ca),
	.w7(32'h3b31e5a4),
	.w8(32'hbc860aca),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27bb9b),
	.w1(32'hba0b58bf),
	.w2(32'h3c078e05),
	.w3(32'hba593285),
	.w4(32'h3c09409c),
	.w5(32'h3c27d30d),
	.w6(32'hbc21ef36),
	.w7(32'h38b280f6),
	.w8(32'h3c4d1898),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0edb5),
	.w1(32'h3be0945d),
	.w2(32'hbb5429dc),
	.w3(32'h3c390591),
	.w4(32'h3baeebaf),
	.w5(32'hbc4600c8),
	.w6(32'h3bd2fc50),
	.w7(32'h3b92196d),
	.w8(32'hbb5e2291),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0743ff),
	.w1(32'hbba51b46),
	.w2(32'h38333ab8),
	.w3(32'h3b3dbe5c),
	.w4(32'hb9ad69ed),
	.w5(32'hba3cca31),
	.w6(32'hbc0bbea8),
	.w7(32'hb985e9a9),
	.w8(32'hbbc8126d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80b16f),
	.w1(32'hba4e4b60),
	.w2(32'h3b0d0d9e),
	.w3(32'h3a78111b),
	.w4(32'h3b562ae9),
	.w5(32'h3ac863d4),
	.w6(32'hbb98d3de),
	.w7(32'hba29a244),
	.w8(32'hbbb1a4cd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807f00),
	.w1(32'hbaca2011),
	.w2(32'h3aab9eae),
	.w3(32'hb9afa8af),
	.w4(32'h3a83de39),
	.w5(32'h3a2566ee),
	.w6(32'hbb7c53b4),
	.w7(32'hb9fceb40),
	.w8(32'h3c2fc0db),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e5bb7),
	.w1(32'h3b95ca4c),
	.w2(32'hba75c240),
	.w3(32'hbc87d007),
	.w4(32'hbaafc13b),
	.w5(32'hbba33ab6),
	.w6(32'h3b8323f5),
	.w7(32'hbc1029bc),
	.w8(32'hbbd09e01),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb776470),
	.w1(32'hbb880011),
	.w2(32'h3ad463b5),
	.w3(32'h3a37ac1d),
	.w4(32'h3b21c51c),
	.w5(32'h3b345a4f),
	.w6(32'hbbe5483d),
	.w7(32'h38dca845),
	.w8(32'hbd854bc4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd39c07a),
	.w1(32'hbba9f9c9),
	.w2(32'h3d46d07c),
	.w3(32'h3b8f893f),
	.w4(32'h3d34575c),
	.w5(32'h3d90390c),
	.w6(32'hbd33f919),
	.w7(32'h3c265c69),
	.w8(32'hbbcff85d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789045),
	.w1(32'hbb4b25bb),
	.w2(32'h3a89cf11),
	.w3(32'h39e47638),
	.w4(32'h3aa58cd2),
	.w5(32'hbac567b6),
	.w6(32'hbb8093a7),
	.w7(32'h3affee86),
	.w8(32'hbb937a58),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e489),
	.w1(32'hbbc804e0),
	.w2(32'h3a92c452),
	.w3(32'h3abe24f9),
	.w4(32'h3b27f563),
	.w5(32'h3acdc077),
	.w6(32'hbbe9fb36),
	.w7(32'h3a1cfc57),
	.w8(32'hbc093638),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98e9a6),
	.w1(32'hbb885d7c),
	.w2(32'hba14e263),
	.w3(32'h3a1b976e),
	.w4(32'h3a09e198),
	.w5(32'hbb41a92d),
	.w6(32'hbbc3de3e),
	.w7(32'hb88b209a),
	.w8(32'h3c68d5ca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e1974),
	.w1(32'hbc186bb9),
	.w2(32'hbc2f8791),
	.w3(32'hbc169652),
	.w4(32'h3b9ce878),
	.w5(32'hbaabd381),
	.w6(32'h3ca4ae35),
	.w7(32'hbba67765),
	.w8(32'hbb5e7efe),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb416c39),
	.w1(32'hbb9281ab),
	.w2(32'hbb0e2622),
	.w3(32'hba9e8d4e),
	.w4(32'hb8fb4bb5),
	.w5(32'hbb82a8c8),
	.w6(32'hbb95d58d),
	.w7(32'hbb1ae4dc),
	.w8(32'hbbf491f3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d378),
	.w1(32'hbb3a0cd1),
	.w2(32'h3b108f37),
	.w3(32'h39fa6de4),
	.w4(32'h3b474d8a),
	.w5(32'h3ab50140),
	.w6(32'hbbc940d1),
	.w7(32'h38d3f15c),
	.w8(32'hbb9af78b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b0e7e),
	.w1(32'hbb9f6a04),
	.w2(32'hbb11e746),
	.w3(32'hbb02c42d),
	.w4(32'hba1b67a9),
	.w5(32'hbb928aac),
	.w6(32'hbb60e362),
	.w7(32'hb98baa68),
	.w8(32'hbd9545d9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4b5b32),
	.w1(32'hbbad1ae5),
	.w2(32'h3d69fe02),
	.w3(32'h3baed38f),
	.w4(32'h3d4c741b),
	.w5(32'h3da7f557),
	.w6(32'hbd4b9f49),
	.w7(32'h3c4d12d7),
	.w8(32'hbd26592b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceef8a0),
	.w1(32'hbb903304),
	.w2(32'h3ce1791b),
	.w3(32'h3a7e41b4),
	.w4(32'h3cdb243a),
	.w5(32'h3d2bcb64),
	.w6(32'hbce63a46),
	.w7(32'h3b85660a),
	.w8(32'hba58652a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a0797),
	.w1(32'hbb83b62c),
	.w2(32'h3b4bbae1),
	.w3(32'h3bbb0b6a),
	.w4(32'h3b1923f3),
	.w5(32'hbae904c8),
	.w6(32'hbb99e4fd),
	.w7(32'h39b12d3f),
	.w8(32'hbbc48419),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf1b24),
	.w1(32'h3ab203b9),
	.w2(32'hbc0c7ae2),
	.w3(32'hbb8611f7),
	.w4(32'hbb14243f),
	.w5(32'hba774afb),
	.w6(32'hbc19532a),
	.w7(32'hbc77d38e),
	.w8(32'hbb35f973),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88be82),
	.w1(32'hbbb7f4d9),
	.w2(32'hbbdfd266),
	.w3(32'hbb7579bb),
	.w4(32'hbba4a6eb),
	.w5(32'hbbf2309b),
	.w6(32'hbb5355bc),
	.w7(32'hbae2b7ce),
	.w8(32'hbb0c3b6d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb982bf5),
	.w1(32'hbc6c57da),
	.w2(32'hbc0a4074),
	.w3(32'h3aca59f6),
	.w4(32'hbba6da2d),
	.w5(32'hbc58f1f1),
	.w6(32'hbc2df2f6),
	.w7(32'hbb9da60d),
	.w8(32'hbc932592),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4972f9),
	.w1(32'hbc842e10),
	.w2(32'hbc948149),
	.w3(32'hbb14994b),
	.w4(32'hbcf819d2),
	.w5(32'hbced9ebe),
	.w6(32'hbc57b279),
	.w7(32'h3abfd282),
	.w8(32'h3cc5cad3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dc528),
	.w1(32'h3a94712b),
	.w2(32'hbc7f79d4),
	.w3(32'h397472b4),
	.w4(32'hbc7eafa7),
	.w5(32'hbcd89442),
	.w6(32'h3c82ee8f),
	.w7(32'h39e539e9),
	.w8(32'hbc52a2a0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbad65),
	.w1(32'hbb479d74),
	.w2(32'h3bb780fe),
	.w3(32'hba82ccd9),
	.w4(32'h3bae3509),
	.w5(32'h3bc784ab),
	.w6(32'hbc146199),
	.w7(32'hb893eac2),
	.w8(32'h3d6f8857),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2d313c),
	.w1(32'h3baaff70),
	.w2(32'hbcdedea2),
	.w3(32'h3ab9eb22),
	.w4(32'hbd11f5d1),
	.w5(32'hbd3da469),
	.w6(32'h3d1b7c11),
	.w7(32'h3bcb3373),
	.w8(32'hba98e593),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bda22),
	.w1(32'hbbd142c0),
	.w2(32'hbbf102f0),
	.w3(32'h3a6ea0aa),
	.w4(32'hbaa1759e),
	.w5(32'hbbdddb88),
	.w6(32'hbc1f00d8),
	.w7(32'hbba51955),
	.w8(32'h3ac7b9c8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaa42c),
	.w1(32'h3af97fd2),
	.w2(32'hbc6f9b88),
	.w3(32'hbbe5b1cc),
	.w4(32'hbc512ea3),
	.w5(32'hbcc4439b),
	.w6(32'h3be68cb9),
	.w7(32'hbbf34fb5),
	.w8(32'h3d60b9f9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d229e46),
	.w1(32'h3ba58109),
	.w2(32'hbcd10341),
	.w3(32'h3ac2335a),
	.w4(32'hbd080c44),
	.w5(32'hbd315d17),
	.w6(32'h3d122960),
	.w7(32'h3bc17444),
	.w8(32'h3d40a0fd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d097629),
	.w1(32'h3b86be82),
	.w2(32'hbcb2df9f),
	.w3(32'h3a07b03c),
	.w4(32'hbcec8aef),
	.w5(32'hbd183e01),
	.w6(32'h3cf52482),
	.w7(32'h3b961ab8),
	.w8(32'h3cce0ec7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82f874),
	.w1(32'h39d97b31),
	.w2(32'hbc93e33b),
	.w3(32'hbb1f2880),
	.w4(32'hbc8fb048),
	.w5(32'hbcde1b33),
	.w6(32'h3c88e888),
	.w7(32'hba65671e),
	.w8(32'hba40796d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ca47),
	.w1(32'hbcb84dda),
	.w2(32'h3b7de3ab),
	.w3(32'h3c00c1b8),
	.w4(32'hbc36372a),
	.w5(32'hbc93efa0),
	.w6(32'hbb67ebb4),
	.w7(32'h3bf19e3f),
	.w8(32'hbbc048c4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96608f),
	.w1(32'hba8be8e6),
	.w2(32'h3adf406e),
	.w3(32'hba2b05f6),
	.w4(32'h3b2ffaca),
	.w5(32'h3b1a9a8a),
	.w6(32'hbb7c88c9),
	.w7(32'hba97a22a),
	.w8(32'hbc88fcc5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c30ef),
	.w1(32'hbc5e3a7b),
	.w2(32'hbccc91d1),
	.w3(32'hbba09218),
	.w4(32'hbc500e0a),
	.w5(32'hbcc2526b),
	.w6(32'hbbc9d68e),
	.w7(32'hbbf98ad4),
	.w8(32'h3ce8d91e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc9cdc9),
	.w1(32'hbb005d4a),
	.w2(32'hbd014da7),
	.w3(32'hbbb66cf6),
	.w4(32'hbcf6b265),
	.w5(32'hbd46cd33),
	.w6(32'h3cc61ed5),
	.w7(32'hbbbf38c1),
	.w8(32'h3a2a325c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3af6b),
	.w1(32'hbbee2a23),
	.w2(32'hbc0c3471),
	.w3(32'hbc6776e4),
	.w4(32'hbb7dd827),
	.w5(32'hbbf170af),
	.w6(32'h3b75ec97),
	.w7(32'h3b347244),
	.w8(32'h3bb2b4d8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f2028),
	.w1(32'h3bc7edaf),
	.w2(32'hbc12f1a5),
	.w3(32'h3aceb2ba),
	.w4(32'h3b881a5c),
	.w5(32'hbab720f8),
	.w6(32'h3b9c594d),
	.w7(32'hbbbf5860),
	.w8(32'hbd82fc8e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2f196a),
	.w1(32'hbb8acee2),
	.w2(32'h3d4fb7f6),
	.w3(32'h3ba24ea0),
	.w4(32'h3d3465c4),
	.w5(32'h3d94b1d3),
	.w6(32'hbd2fbbc2),
	.w7(32'h3c3d884f),
	.w8(32'hbb5c280e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb020673),
	.w1(32'hbbf45e27),
	.w2(32'hbbdd6ff7),
	.w3(32'h3ad799a1),
	.w4(32'hbb276ca5),
	.w5(32'hbc08fee5),
	.w6(32'hbc401924),
	.w7(32'hbb948dae),
	.w8(32'h3ca35729),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7655b),
	.w1(32'hbbc4b60b),
	.w2(32'hbcaf66b7),
	.w3(32'hbc106591),
	.w4(32'hbcde538b),
	.w5(32'hbd0e92f5),
	.w6(32'h3bb06fa1),
	.w7(32'hbba7c79d),
	.w8(32'hbbfdf53e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00429),
	.w1(32'hbad9554a),
	.w2(32'h3b2ea4f8),
	.w3(32'h39c8eb70),
	.w4(32'h3b6d7aa4),
	.w5(32'h3b870d84),
	.w6(32'hbb9ff982),
	.w7(32'hb9db8fc2),
	.w8(32'hbd846e7b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5187b3),
	.w1(32'hbc2c9c41),
	.w2(32'h3d400433),
	.w3(32'hb9f93fff),
	.w4(32'h3d3de943),
	.w5(32'h3d931afb),
	.w6(32'hbd4a08c5),
	.w7(32'h3bd9997d),
	.w8(32'h3cb047f2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63def4),
	.w1(32'hba353b21),
	.w2(32'hbc953261),
	.w3(32'hbbd92ede),
	.w4(32'hbcaab61f),
	.w5(32'hbcffa238),
	.w6(32'h3c703543),
	.w7(32'hbb819ed3),
	.w8(32'h3cb9de84),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c893436),
	.w1(32'h3b0e2e0d),
	.w2(32'hbc37c334),
	.w3(32'h3a12f77d),
	.w4(32'hbc66cd7b),
	.w5(32'hbc9a46af),
	.w6(32'h3c7905f8),
	.w7(32'h3b079350),
	.w8(32'h3980603b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6689f),
	.w1(32'hba010048),
	.w2(32'hba4a1513),
	.w3(32'h38fc22f7),
	.w4(32'h38dd31c2),
	.w5(32'hba091c7f),
	.w6(32'hb97b48e0),
	.w7(32'h38f1b0f0),
	.w8(32'hba10667e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1712b),
	.w1(32'h3b5e0803),
	.w2(32'hb9d7f706),
	.w3(32'hb9f95d5b),
	.w4(32'h3a86417c),
	.w5(32'h394119a8),
	.w6(32'h3a7fedf4),
	.w7(32'hbaa8db38),
	.w8(32'hb888e230),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb302a8f8),
	.w1(32'h396fe3fa),
	.w2(32'h39953836),
	.w3(32'h3961535e),
	.w4(32'h3a0f2e54),
	.w5(32'h3942b00b),
	.w6(32'h39ff83b9),
	.w7(32'h3a03726d),
	.w8(32'h379d6638),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b1bb2),
	.w1(32'h38b920be),
	.w2(32'h3890f06a),
	.w3(32'h3887771a),
	.w4(32'h39d0f3ac),
	.w5(32'h390d9d57),
	.w6(32'h39c72e3f),
	.w7(32'h39ce9f3f),
	.w8(32'hb8e552ff),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eb1ab),
	.w1(32'hba53fc7d),
	.w2(32'hba28a506),
	.w3(32'hba16045e),
	.w4(32'hba64ba70),
	.w5(32'hba472d96),
	.w6(32'hb94cceb4),
	.w7(32'hba2430bc),
	.w8(32'hbb06228f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39885090),
	.w1(32'h3a7e723d),
	.w2(32'h3a6c8927),
	.w3(32'h39d10934),
	.w4(32'hbabb5728),
	.w5(32'hba53204d),
	.w6(32'hb94b34f9),
	.w7(32'h39218652),
	.w8(32'hb9cb9a59),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9911003),
	.w1(32'hba8c8a18),
	.w2(32'h395568c8),
	.w3(32'hb8fb7b45),
	.w4(32'h37ec45f5),
	.w5(32'h38ac6f73),
	.w6(32'hba37a8ca),
	.w7(32'h38288ebf),
	.w8(32'h3934db17),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11f749),
	.w1(32'h38c6f984),
	.w2(32'hb95325e0),
	.w3(32'h3a9db30c),
	.w4(32'h3a1805f8),
	.w5(32'h3a05af58),
	.w6(32'hb918b91f),
	.w7(32'h370c5c41),
	.w8(32'h39ffcae6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902bcaa),
	.w1(32'hb90e49d1),
	.w2(32'h39c78fce),
	.w3(32'h38b39969),
	.w4(32'h399a32aa),
	.w5(32'h39e2b22e),
	.w6(32'h39a98b65),
	.w7(32'h39ca6bdf),
	.w8(32'h393b77ce),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39314c7e),
	.w1(32'h393340fc),
	.w2(32'h390b4004),
	.w3(32'h39b30233),
	.w4(32'h39c650fe),
	.w5(32'h393b363e),
	.w6(32'h39d35e4d),
	.w7(32'h3944db3a),
	.w8(32'h3988a902),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d291c),
	.w1(32'h39859bec),
	.w2(32'hb9665c96),
	.w3(32'h39e093ca),
	.w4(32'h3a398824),
	.w5(32'h38e5b1a2),
	.w6(32'h39e4c6e6),
	.w7(32'h396c1ccd),
	.w8(32'h3a839de9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b231),
	.w1(32'h398ec8c4),
	.w2(32'hba320f47),
	.w3(32'hb91c053a),
	.w4(32'hb92022c4),
	.w5(32'hba138f0e),
	.w6(32'hb994ed8f),
	.w7(32'hba99533f),
	.w8(32'h3a0b2bb2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7cb38),
	.w1(32'hba425744),
	.w2(32'hba1a29cc),
	.w3(32'h38bea892),
	.w4(32'hba17bec8),
	.w5(32'hb95f700b),
	.w6(32'hba3e8357),
	.w7(32'hba17ba8b),
	.w8(32'hbae51df5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d2161),
	.w1(32'h3b08f4d7),
	.w2(32'h3b4f735c),
	.w3(32'hba48898c),
	.w4(32'h38908b2d),
	.w5(32'h3ae90955),
	.w6(32'h3811765f),
	.w7(32'h3b2016a8),
	.w8(32'hba62c14a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba007399),
	.w1(32'hbad5654c),
	.w2(32'hba9d7769),
	.w3(32'hb9da9c00),
	.w4(32'hb890bc87),
	.w5(32'h391e58a6),
	.w6(32'hba8ee66b),
	.w7(32'hba41d398),
	.w8(32'hb99e4669),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a079b9f),
	.w1(32'hb9a6914c),
	.w2(32'hba3b23f9),
	.w3(32'hba8d74cb),
	.w4(32'hbac255c2),
	.w5(32'hbac78a4d),
	.w6(32'hba4326ee),
	.w7(32'hba3f050a),
	.w8(32'hba83f93c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c03bf),
	.w1(32'h397f4d85),
	.w2(32'h3874f059),
	.w3(32'hba8edc06),
	.w4(32'hb9b1dbfc),
	.w5(32'h3a9291dc),
	.w6(32'hbb181a59),
	.w7(32'hba3ddda7),
	.w8(32'h3a17ca6d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50022f),
	.w1(32'h39315ce6),
	.w2(32'h39d4adcd),
	.w3(32'h3ab2e646),
	.w4(32'h3a421396),
	.w5(32'h3a6d44d6),
	.w6(32'hb6e1d6b9),
	.w7(32'h399f1a84),
	.w8(32'h39c81606),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8795ff6),
	.w1(32'h3aa34aa1),
	.w2(32'hb9b405e9),
	.w3(32'hba123b8f),
	.w4(32'hb9adf235),
	.w5(32'hba9effa0),
	.w6(32'h39c73637),
	.w7(32'hba0a6033),
	.w8(32'h39f14be3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b61c0),
	.w1(32'h3b2a858c),
	.w2(32'h3aa6bd72),
	.w3(32'hb9acbc7c),
	.w4(32'h39bb1619),
	.w5(32'hbab4fa7e),
	.w6(32'hba5189f8),
	.w7(32'h3a2293c0),
	.w8(32'hba5851af),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffad49),
	.w1(32'hba2bf373),
	.w2(32'hb9b84395),
	.w3(32'hb9a7a38a),
	.w4(32'hb99e191b),
	.w5(32'hba4f202c),
	.w6(32'hb8d4af18),
	.w7(32'hb9dd2c14),
	.w8(32'h39fb2dff),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887cee2),
	.w1(32'hb7baae3d),
	.w2(32'hb79c449d),
	.w3(32'h39624130),
	.w4(32'h3985107c),
	.w5(32'h39d34853),
	.w6(32'h39c83c68),
	.w7(32'h3a086a71),
	.w8(32'hbae88bbd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa378a),
	.w1(32'hb9b7f187),
	.w2(32'hbafd05b7),
	.w3(32'hbae38c68),
	.w4(32'hbaaa88e8),
	.w5(32'hba7d3a44),
	.w6(32'hba5cf0d3),
	.w7(32'hbb389e4a),
	.w8(32'h39b25677),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule