module layer_8_featuremap_237(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb48b8b),
	.w1(32'h3c07041d),
	.w2(32'hb99defd2),
	.w3(32'h3b9e32d5),
	.w4(32'h3b5884c9),
	.w5(32'hbbea835d),
	.w6(32'h3bcbd62e),
	.w7(32'h3c5b4e70),
	.w8(32'h3c165c24),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf97e31),
	.w1(32'hbb5a8c8d),
	.w2(32'hbb88b460),
	.w3(32'h3bd4374b),
	.w4(32'hbad064de),
	.w5(32'hbb34e572),
	.w6(32'hbb2c82c3),
	.w7(32'hbb6028d5),
	.w8(32'h384718da),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9918514),
	.w1(32'hba357c94),
	.w2(32'h3c388c6b),
	.w3(32'h3a82ae5e),
	.w4(32'h3b303aaf),
	.w5(32'h3c68f454),
	.w6(32'hbab91d54),
	.w7(32'h3b799baa),
	.w8(32'h3a9e5e9a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61958a),
	.w1(32'h3b35e4cb),
	.w2(32'h3befb6b0),
	.w3(32'h3c29887b),
	.w4(32'h3b660f4e),
	.w5(32'h3c7bbb14),
	.w6(32'h3bf075d3),
	.w7(32'h3c03bbfc),
	.w8(32'h39f3480f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8ab87),
	.w1(32'hbbb54842),
	.w2(32'hbbff31b1),
	.w3(32'h3c381aef),
	.w4(32'hbb20ff5e),
	.w5(32'hbb654722),
	.w6(32'h3b1a0dcc),
	.w7(32'hbb2e0dd8),
	.w8(32'h3a4d0025),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5219),
	.w1(32'h3b45eedc),
	.w2(32'hbb7c5273),
	.w3(32'hbabfb381),
	.w4(32'h3b3d474a),
	.w5(32'h39d08e44),
	.w6(32'h3b326501),
	.w7(32'h3986047e),
	.w8(32'hbb7397cb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc21c4d),
	.w1(32'hbbad838c),
	.w2(32'hbb564af6),
	.w3(32'h3c212ed9),
	.w4(32'hbb680f4c),
	.w5(32'hbb8fb680),
	.w6(32'hbbc0adbf),
	.w7(32'hbbd72d82),
	.w8(32'hbbdbcae3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e30d),
	.w1(32'h3bf08c70),
	.w2(32'h3bf801f8),
	.w3(32'hbbc1ea8c),
	.w4(32'hbb2ea3da),
	.w5(32'h3b16904e),
	.w6(32'h3a933ebc),
	.w7(32'h3bb84fe9),
	.w8(32'h3b906f42),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9198f),
	.w1(32'hbc226839),
	.w2(32'h3b6f05d2),
	.w3(32'h3b92da1a),
	.w4(32'hbbb44e9f),
	.w5(32'h3bef252b),
	.w6(32'hbbdc6979),
	.w7(32'h3b8743c5),
	.w8(32'h3b99113c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ed506),
	.w1(32'hbb1d84c4),
	.w2(32'hb94fb3ef),
	.w3(32'h3badee71),
	.w4(32'hbab9ea05),
	.w5(32'hbaee5779),
	.w6(32'h3ba62d6b),
	.w7(32'h3a1d0fd5),
	.w8(32'h3a82f95e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9b942),
	.w1(32'hbb719d51),
	.w2(32'hbbffeed5),
	.w3(32'h3a43d9bc),
	.w4(32'hbb596fe8),
	.w5(32'hbbeb6c7d),
	.w6(32'hbb9035c4),
	.w7(32'hbb9638c8),
	.w8(32'hbb2fa439),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e7fd),
	.w1(32'h3ba1baa5),
	.w2(32'h3c092f55),
	.w3(32'hba00fe42),
	.w4(32'h3b210cf8),
	.w5(32'h3c2ecd97),
	.w6(32'h3afdc758),
	.w7(32'h3c17e5ef),
	.w8(32'h3c0e0ca1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aeb30),
	.w1(32'hbc4dd67d),
	.w2(32'hbc4d22fe),
	.w3(32'h3c66b025),
	.w4(32'hbc3b8bee),
	.w5(32'hbc8664fc),
	.w6(32'hbbe85027),
	.w7(32'hbbcd1a54),
	.w8(32'hbbcad868),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15610e),
	.w1(32'hbc4bcfbe),
	.w2(32'hbc3e1f46),
	.w3(32'hbc2fb2e0),
	.w4(32'hbbfd7ac1),
	.w5(32'hbada60dd),
	.w6(32'h39d1b6eb),
	.w7(32'h3b80cb23),
	.w8(32'h3b746c6f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21a5f4),
	.w1(32'hbbef0f32),
	.w2(32'h3b336c28),
	.w3(32'hba44f769),
	.w4(32'hbbb03909),
	.w5(32'h3b7397dc),
	.w6(32'hbc7b58ff),
	.w7(32'hbbe20602),
	.w8(32'hbc155332),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98636c),
	.w1(32'hba7798d5),
	.w2(32'h3a9811d1),
	.w3(32'h39b99199),
	.w4(32'hba2a9221),
	.w5(32'h380ad6e1),
	.w6(32'hbb4614eb),
	.w7(32'hbbb0ad1d),
	.w8(32'h39b669fd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad80525),
	.w1(32'hbb444a45),
	.w2(32'hbc159a8c),
	.w3(32'h3c087541),
	.w4(32'hbae8341d),
	.w5(32'hbbb5a106),
	.w6(32'hbbb80ca3),
	.w7(32'hbc11acf5),
	.w8(32'hbbdedcd8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2cdbe),
	.w1(32'h3b59fde2),
	.w2(32'h3b36c3ac),
	.w3(32'hbbb478c1),
	.w4(32'h3be439ac),
	.w5(32'h3a9a186d),
	.w6(32'h3948dacb),
	.w7(32'hbc0503e7),
	.w8(32'h3b2d038b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b4b23),
	.w1(32'h3b791106),
	.w2(32'h3b88121a),
	.w3(32'hbafa4a5e),
	.w4(32'h3a651560),
	.w5(32'hbbb79e8d),
	.w6(32'hbbd6b486),
	.w7(32'hbc861ff4),
	.w8(32'hbb8a50af),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7a859),
	.w1(32'hbae66409),
	.w2(32'h3b7cf123),
	.w3(32'hbb34609d),
	.w4(32'hbb2c8a00),
	.w5(32'h3b1b7e25),
	.w6(32'hbc117a65),
	.w7(32'hbb31e501),
	.w8(32'hbb35f257),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b748d0f),
	.w1(32'hbb00c0ca),
	.w2(32'hbb056b1e),
	.w3(32'h39393eb2),
	.w4(32'h3ba687e9),
	.w5(32'h3c805306),
	.w6(32'h3b125341),
	.w7(32'h3b463bce),
	.w8(32'h3b7bfc80),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d2c5d),
	.w1(32'hbcc19ea5),
	.w2(32'hbd37f6a4),
	.w3(32'h3be8fbd6),
	.w4(32'hbc870764),
	.w5(32'hbd1af93e),
	.w6(32'hbc75d872),
	.w7(32'hbd0685e5),
	.w8(32'hbca35eeb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd144450),
	.w1(32'h3c551af7),
	.w2(32'h3b2f3127),
	.w3(32'hbcab1d79),
	.w4(32'h3bcc7370),
	.w5(32'hba34766b),
	.w6(32'h3c0f35d8),
	.w7(32'h3b65397f),
	.w8(32'h3b7884b8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b826fe5),
	.w1(32'hbd3580c8),
	.w2(32'hbd85a466),
	.w3(32'hbb8461ae),
	.w4(32'hbd2cb283),
	.w5(32'hbd656dfb),
	.w6(32'hbcd387bd),
	.w7(32'hbd3ce6ee),
	.w8(32'hbd05a560),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd55d768),
	.w1(32'h3b0a65f0),
	.w2(32'h3bc8822b),
	.w3(32'hbd0f3002),
	.w4(32'hb860b440),
	.w5(32'hbb18c2c0),
	.w6(32'h3b4b66a5),
	.w7(32'h3b9d886e),
	.w8(32'h3ac87179),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a405b),
	.w1(32'h385bc71c),
	.w2(32'hbbf41862),
	.w3(32'hbbf447ed),
	.w4(32'h3c44a34c),
	.w5(32'hba45dd48),
	.w6(32'h3b8b50bb),
	.w7(32'h3be415bc),
	.w8(32'h3b8075c2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc580ead),
	.w1(32'h3c3271eb),
	.w2(32'h3c846954),
	.w3(32'h3c05cf71),
	.w4(32'h3b734f11),
	.w5(32'h3bfe1fad),
	.w6(32'h3bbc08fc),
	.w7(32'h3c2b31f4),
	.w8(32'h3a9641d9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dccb4),
	.w1(32'h3b32e526),
	.w2(32'h3b62b9ad),
	.w3(32'h3b60489c),
	.w4(32'hbb0efff0),
	.w5(32'h3b0faf23),
	.w6(32'h3b0f2ed6),
	.w7(32'h3bc0f4bb),
	.w8(32'h3ba768e7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d8209),
	.w1(32'h3b864e02),
	.w2(32'h3be4ca60),
	.w3(32'hb91835f3),
	.w4(32'h3b33b5d7),
	.w5(32'h3bf164b2),
	.w6(32'hbbb83eb3),
	.w7(32'hb9912f89),
	.w8(32'hbbf15de8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2af1b3),
	.w1(32'h39babad5),
	.w2(32'h3aab430f),
	.w3(32'hbbbc9ad3),
	.w4(32'h3be668ea),
	.w5(32'h3c5951ce),
	.w6(32'h3b7a978c),
	.w7(32'h3ad5e478),
	.w8(32'hbb33e56b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24394a),
	.w1(32'hbb33ecc1),
	.w2(32'h38f8c48b),
	.w3(32'h3c716c59),
	.w4(32'hbb31f8b2),
	.w5(32'h39907587),
	.w6(32'hbbfd9ec9),
	.w7(32'hbb466f69),
	.w8(32'hb8f96ad4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ada9e),
	.w1(32'hbbdc20d4),
	.w2(32'h3aa5a0cb),
	.w3(32'h3aa474d6),
	.w4(32'hbbb099c3),
	.w5(32'h39808f02),
	.w6(32'hbc62ab47),
	.w7(32'hbb36327d),
	.w8(32'hbb43f17b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb18c3),
	.w1(32'hbb176976),
	.w2(32'hbb8139cd),
	.w3(32'h3ba923f3),
	.w4(32'h3b5d75dc),
	.w5(32'hbb1ab400),
	.w6(32'hb90ea766),
	.w7(32'hbba5eb5b),
	.w8(32'h3bbe5902),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1e5b1),
	.w1(32'hbc92ac59),
	.w2(32'hbd01acaf),
	.w3(32'hb7a5ef67),
	.w4(32'hbaec6e94),
	.w5(32'hbcb0007a),
	.w6(32'hbc1e50e1),
	.w7(32'hbca65a52),
	.w8(32'hbbf9bb89),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca4471),
	.w1(32'h3bfd5771),
	.w2(32'h3bfdbfda),
	.w3(32'hbc848769),
	.w4(32'h3c0af3de),
	.w5(32'h3c2ec4fc),
	.w6(32'h3c2b4364),
	.w7(32'h3c119198),
	.w8(32'h3b858039),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be97dd0),
	.w1(32'h3b74220f),
	.w2(32'h3c89bb81),
	.w3(32'h3bbe411d),
	.w4(32'h3ba07e47),
	.w5(32'h3c62ba26),
	.w6(32'h3b0624eb),
	.w7(32'hbb18a7e9),
	.w8(32'hbb6427d0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f2ac3),
	.w1(32'h3b8a7c89),
	.w2(32'h3bc94156),
	.w3(32'h3c4c577a),
	.w4(32'h3b1f0cab),
	.w5(32'h3bc7d32f),
	.w6(32'h3baa8f24),
	.w7(32'h3ba86b34),
	.w8(32'h392375e8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6987f),
	.w1(32'hbc2a9a1f),
	.w2(32'h3b85390c),
	.w3(32'h3b4ecc6e),
	.w4(32'hbbd6cacf),
	.w5(32'h3bd4a8c7),
	.w6(32'hbc3ff525),
	.w7(32'hbb1bcd76),
	.w8(32'hbbad83b2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c755),
	.w1(32'h3c523b71),
	.w2(32'h3c80c40f),
	.w3(32'h3b0e986f),
	.w4(32'h3c44bfdd),
	.w5(32'h3c834fc9),
	.w6(32'h3bb5dbe3),
	.w7(32'h3c4b9815),
	.w8(32'h3c36f8b7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4456b8),
	.w1(32'hbc973a6d),
	.w2(32'hbcfae1e9),
	.w3(32'h3c077e5b),
	.w4(32'hbc609331),
	.w5(32'hbc9f7b48),
	.w6(32'hbbbd2fce),
	.w7(32'hbc46d2aa),
	.w8(32'hbc5321e5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7a8a9),
	.w1(32'h3bd47e58),
	.w2(32'h3ccc378c),
	.w3(32'hbc59e2f7),
	.w4(32'h3c02104a),
	.w5(32'h3ce4a3a5),
	.w6(32'h3aba4c2a),
	.w7(32'h3ca640b1),
	.w8(32'h3c20a935),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c892262),
	.w1(32'hbba4dc26),
	.w2(32'h3ba65253),
	.w3(32'h3ca05141),
	.w4(32'hbb55f2d0),
	.w5(32'h3aac409a),
	.w6(32'hbc46b6cc),
	.w7(32'hbba27501),
	.w8(32'hb9cd82b5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcab77),
	.w1(32'hba968246),
	.w2(32'h3b122e42),
	.w3(32'h3ac31dda),
	.w4(32'hbb77eb57),
	.w5(32'hbb4c23c8),
	.w6(32'hbadf634c),
	.w7(32'hba33175c),
	.w8(32'hbaf97b41),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560c3a),
	.w1(32'h3bd0a732),
	.w2(32'h3cbad0c2),
	.w3(32'hbbb87742),
	.w4(32'h39bcc3ed),
	.w5(32'h3c137778),
	.w6(32'hbbeaa301),
	.w7(32'h3b44b7e4),
	.w8(32'h3c1be2ab),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca50d41),
	.w1(32'hbc9f9e2d),
	.w2(32'hbcefd44d),
	.w3(32'h3c5a4629),
	.w4(32'hbc822226),
	.w5(32'hbc9f6a65),
	.w6(32'hbc190281),
	.w7(32'hbca3d74d),
	.w8(32'hbc840117),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccdaa98),
	.w1(32'hba484c37),
	.w2(32'hbab746e6),
	.w3(32'hbc8d6c70),
	.w4(32'h3a56d15e),
	.w5(32'hbacfb39b),
	.w6(32'hbb835780),
	.w7(32'hbb402efe),
	.w8(32'hbac7aa97),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a0dced),
	.w1(32'hbc2cfbbb),
	.w2(32'hbc404d86),
	.w3(32'hbab5093b),
	.w4(32'hbc211525),
	.w5(32'hbc2e2079),
	.w6(32'hbc7d364e),
	.w7(32'hbc50e02f),
	.w8(32'hbc366dcb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaedeb),
	.w1(32'hbceb48db),
	.w2(32'hbd21c36a),
	.w3(32'hbc3454f7),
	.w4(32'hbcca8cb4),
	.w5(32'hbcfc4ee8),
	.w6(32'hbc0ae9f1),
	.w7(32'hbcb6646d),
	.w8(32'hbc58c26f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb0bb6),
	.w1(32'hbc1ecc8d),
	.w2(32'hbc502d50),
	.w3(32'hbc9e3b5d),
	.w4(32'hbc0ebae9),
	.w5(32'hbbf3743d),
	.w6(32'h3ab3c9fe),
	.w7(32'hbbcc53db),
	.w8(32'h3ae455f4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c263c),
	.w1(32'hbb952a3b),
	.w2(32'hbb280c21),
	.w3(32'hbb55b165),
	.w4(32'hbaa45e2d),
	.w5(32'hbc00aafe),
	.w6(32'hbc3b3d5f),
	.w7(32'h3ab6faa9),
	.w8(32'hba0b63a6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9947ff),
	.w1(32'h3b72cc0b),
	.w2(32'h3b0c5d2c),
	.w3(32'h3aa1f52d),
	.w4(32'h395e73ac),
	.w5(32'h3b396931),
	.w6(32'h3a2a220a),
	.w7(32'h3c0d3db9),
	.w8(32'hbad46857),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0667f0),
	.w1(32'h3b9c562e),
	.w2(32'h3c3b85e6),
	.w3(32'hbaf8f9f0),
	.w4(32'h39b23e63),
	.w5(32'h3bb8b89a),
	.w6(32'h3a34e457),
	.w7(32'h3b29b19f),
	.w8(32'hbab7073a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f862),
	.w1(32'hb89c4990),
	.w2(32'h3aa5c090),
	.w3(32'hbb43023b),
	.w4(32'h3b37aca7),
	.w5(32'h3bbe5543),
	.w6(32'h3b0040da),
	.w7(32'h3b8f7877),
	.w8(32'h3b0bdaad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10a633),
	.w1(32'h3b26d700),
	.w2(32'h3c0b72a6),
	.w3(32'h3bdd1a4c),
	.w4(32'hbb701dc0),
	.w5(32'h3b780613),
	.w6(32'h3af27977),
	.w7(32'hbb872e2a),
	.w8(32'h3bf8c3a3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd70bf9),
	.w1(32'h3c2323f5),
	.w2(32'h3ba33af7),
	.w3(32'h3b33d462),
	.w4(32'h3be793b6),
	.w5(32'h3bb3f1fb),
	.w6(32'h3b7646e6),
	.w7(32'h3b9bd12b),
	.w8(32'h3acc2513),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd48810),
	.w1(32'hbc0addaf),
	.w2(32'hbba3fe17),
	.w3(32'h3bd9c7ac),
	.w4(32'hbab6f5b0),
	.w5(32'hbc361753),
	.w6(32'hbc5824d4),
	.w7(32'hbc4c02d4),
	.w8(32'hbbd227a4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc455b7),
	.w1(32'h3babab3d),
	.w2(32'h3a8f9a99),
	.w3(32'hbc04b2f6),
	.w4(32'h3a39f66b),
	.w5(32'hba1de91d),
	.w6(32'hbbabe33e),
	.w7(32'hbb130725),
	.w8(32'h3abe168b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c325572),
	.w1(32'h3c02d4a6),
	.w2(32'h3ad40d41),
	.w3(32'h3b5537e0),
	.w4(32'h3be104f6),
	.w5(32'h3b42bba3),
	.w6(32'h3bbf35d8),
	.w7(32'hb9893c3e),
	.w8(32'hbab73bf8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2980c4),
	.w1(32'hba6cd4b4),
	.w2(32'hbb2ad07d),
	.w3(32'hbafc9abf),
	.w4(32'hbb2c7b42),
	.w5(32'hbaae5970),
	.w6(32'hbb280f6e),
	.w7(32'hbb1cc4b2),
	.w8(32'hbb7b140f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb534c69),
	.w1(32'hbd0fe1dd),
	.w2(32'hbd4efd1e),
	.w3(32'hbb3edf16),
	.w4(32'hbcaf4bc7),
	.w5(32'hbd0976d6),
	.w6(32'hbcb16cf3),
	.w7(32'hbcf04940),
	.w8(32'hbc95c136),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c2110),
	.w1(32'hbc629a28),
	.w2(32'hbafe72fb),
	.w3(32'hbcc63789),
	.w4(32'hbc73427b),
	.w5(32'hbb354fe1),
	.w6(32'hbc5ea951),
	.w7(32'h38fba093),
	.w8(32'hbbf5a4f2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187511),
	.w1(32'hbbc6d126),
	.w2(32'h3ba9733f),
	.w3(32'hbc1750f4),
	.w4(32'hbb35aafe),
	.w5(32'hbabc6c16),
	.w6(32'hbbb01e07),
	.w7(32'h3b13ef11),
	.w8(32'hbaa405c2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd947f4),
	.w1(32'hbb8ff80d),
	.w2(32'h3bde80b2),
	.w3(32'h3a87c727),
	.w4(32'hbab43455),
	.w5(32'h3c0d7195),
	.w6(32'hbb05dca4),
	.w7(32'h3bf9171d),
	.w8(32'h3b8199b2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc901cc),
	.w1(32'h3b13427f),
	.w2(32'h3bb93204),
	.w3(32'h3c310ccf),
	.w4(32'hbb2613b8),
	.w5(32'h3a9d4226),
	.w6(32'h3a99e19d),
	.w7(32'h3bbcbe95),
	.w8(32'hb9e8805a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13332d),
	.w1(32'h3ac2c2f1),
	.w2(32'h3b9e0ad1),
	.w3(32'hb8a98e1c),
	.w4(32'hbb22eb70),
	.w5(32'h3b44336e),
	.w6(32'hbba7322d),
	.w7(32'hb9583ac5),
	.w8(32'hbabff2cf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80bbbd),
	.w1(32'hbc8abe89),
	.w2(32'hbcd3aa2a),
	.w3(32'h3b1d2591),
	.w4(32'hbc6c7ec2),
	.w5(32'hbcc768fa),
	.w6(32'hbab3799d),
	.w7(32'hbc90c8b2),
	.w8(32'hbc7d06d2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc38162),
	.w1(32'h3c54f6ce),
	.w2(32'h3b84b45c),
	.w3(32'hbc6665fd),
	.w4(32'h3c855e6b),
	.w5(32'h3c5f152e),
	.w6(32'h3c67269f),
	.w7(32'hb9c8e12d),
	.w8(32'h3bd448ba),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e4e98),
	.w1(32'h3bdc673d),
	.w2(32'h3bafadd5),
	.w3(32'h3c808bd6),
	.w4(32'h3b5e3e31),
	.w5(32'h3c179197),
	.w6(32'h3b9101df),
	.w7(32'h3bc37944),
	.w8(32'h3c329421),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba57060),
	.w1(32'hbd55c4ed),
	.w2(32'hbd9dd7ff),
	.w3(32'h3af6c20d),
	.w4(32'hbcfc6534),
	.w5(32'hbd7ce3c8),
	.w6(32'hbd2aec08),
	.w7(32'hbd5f03cd),
	.w8(32'hbd098379),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd78d5f3),
	.w1(32'hbb95452c),
	.w2(32'hbba564fa),
	.w3(32'hbd389d62),
	.w4(32'h3b7eb781),
	.w5(32'hbb24f65b),
	.w6(32'hbb2c2dff),
	.w7(32'hbb97ed3e),
	.w8(32'h3b70a337),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04a3fe),
	.w1(32'h3bac6d69),
	.w2(32'h3bb6d1f4),
	.w3(32'hbb0915ce),
	.w4(32'h3ada6e0f),
	.w5(32'h3b7475d4),
	.w6(32'hba24cd1c),
	.w7(32'h3a82a76b),
	.w8(32'hba9f66b4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb089a9b),
	.w1(32'h3bf792e7),
	.w2(32'h3ca419dd),
	.w3(32'hb9cc6ebd),
	.w4(32'h3a4aa86f),
	.w5(32'h3c6d0d3c),
	.w6(32'h3be41077),
	.w7(32'h3c5469c0),
	.w8(32'h3c654a6c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9dcb3c),
	.w1(32'h3c8238ae),
	.w2(32'h3cd24162),
	.w3(32'h3c138a6d),
	.w4(32'h3baddcc7),
	.w5(32'h3c999dc6),
	.w6(32'h3bb8c2d4),
	.w7(32'h3c5dc8d8),
	.w8(32'h3beb6e42),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafa4f5),
	.w1(32'h3b77051c),
	.w2(32'h3c7b207c),
	.w3(32'h3c54e622),
	.w4(32'h3b4cf9a1),
	.w5(32'h3bdd56a8),
	.w6(32'h3ab3423c),
	.w7(32'h3b0ee5dd),
	.w8(32'h3b823902),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba72a41),
	.w1(32'h3be63b9c),
	.w2(32'h3b9a03f1),
	.w3(32'hb987c130),
	.w4(32'h3c3b6cc9),
	.w5(32'h3a573832),
	.w6(32'h3b3f8b8a),
	.w7(32'h3a35f6d0),
	.w8(32'h3bd7bb8a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb1427),
	.w1(32'h3c241802),
	.w2(32'h3c0be2c1),
	.w3(32'hbbc2eadd),
	.w4(32'h3be49fe6),
	.w5(32'h3a15725a),
	.w6(32'hbba2f5b2),
	.w7(32'h38e9e8fc),
	.w8(32'h3aac8111),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c124873),
	.w1(32'h3b5106ca),
	.w2(32'h3a3f041a),
	.w3(32'h3b3c2870),
	.w4(32'h3b0362ca),
	.w5(32'hbab57f5a),
	.w6(32'hba81a22b),
	.w7(32'hbb9798a1),
	.w8(32'h3b19f756),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac3fcc),
	.w1(32'hb985401f),
	.w2(32'h3b931fae),
	.w3(32'h3b2539af),
	.w4(32'h38ede108),
	.w5(32'hbb398481),
	.w6(32'hbbaf9afb),
	.w7(32'hbb154dda),
	.w8(32'hbb461fa4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2839bd),
	.w1(32'h3bc97133),
	.w2(32'h3a927b12),
	.w3(32'hbab33311),
	.w4(32'h3b65fd7a),
	.w5(32'h3a8c02bd),
	.w6(32'h3b7ef173),
	.w7(32'h3a2e148f),
	.w8(32'h391d1491),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d05ff),
	.w1(32'hbc0652a1),
	.w2(32'hbbd05b3f),
	.w3(32'h3b0aa752),
	.w4(32'hbba45502),
	.w5(32'h3b5acf3d),
	.w6(32'h3a470e4a),
	.w7(32'hbb683998),
	.w8(32'hbaac6379),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc033f08),
	.w1(32'hbb37d2ca),
	.w2(32'h3bb1cc97),
	.w3(32'hbbce8c1b),
	.w4(32'h3a1d8266),
	.w5(32'h3c27dc9d),
	.w6(32'h3adff87f),
	.w7(32'h3c795c32),
	.w8(32'h3c202668),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0840),
	.w1(32'hbd52b92b),
	.w2(32'hbd957249),
	.w3(32'hba5ccb76),
	.w4(32'hbcf911d1),
	.w5(32'hbd6944b6),
	.w6(32'hbd24540c),
	.w7(32'hbd4d52b0),
	.w8(32'hbcf2477c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd51fe62),
	.w1(32'h3c04080d),
	.w2(32'h3ba9957a),
	.w3(32'hbd20b568),
	.w4(32'hbb86fe92),
	.w5(32'hbb15b5af),
	.w6(32'hbbfdece2),
	.w7(32'hbbb443f7),
	.w8(32'h39352986),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c851e93),
	.w1(32'h3af36d63),
	.w2(32'h3a62656a),
	.w3(32'hbb673fda),
	.w4(32'hbb393e70),
	.w5(32'h3a8d96fc),
	.w6(32'h3b17c28e),
	.w7(32'hbbcb7b28),
	.w8(32'hbb991c58),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1be163),
	.w1(32'hbb3658b0),
	.w2(32'hbb915b97),
	.w3(32'hba87f2d1),
	.w4(32'hb94158a0),
	.w5(32'hba11d9de),
	.w6(32'h3beab658),
	.w7(32'hb97293dc),
	.w8(32'h3b9556bc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb33cd),
	.w1(32'h3be0040b),
	.w2(32'h3b65b400),
	.w3(32'h3bde9f22),
	.w4(32'h391f07fc),
	.w5(32'hba9a082c),
	.w6(32'h3be7777f),
	.w7(32'h3be3adda),
	.w8(32'h3bbcfdaa),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f90f9),
	.w1(32'h3b52ce5a),
	.w2(32'h3b9a0bcc),
	.w3(32'h3b4a3d01),
	.w4(32'h3b22d1b5),
	.w5(32'h3ba7b155),
	.w6(32'h3af3176c),
	.w7(32'h3b3bf4ae),
	.w8(32'h3b7c599c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42b81b),
	.w1(32'hbbf66453),
	.w2(32'h3a918271),
	.w3(32'h3b3ac71b),
	.w4(32'hbc122c2d),
	.w5(32'hbaa94197),
	.w6(32'hbc0003e0),
	.w7(32'hba0c36a6),
	.w8(32'hbb27bcb5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfb724),
	.w1(32'hbb87b835),
	.w2(32'hbb98ec01),
	.w3(32'h3990ac5d),
	.w4(32'hbb164b84),
	.w5(32'hba817989),
	.w6(32'h3b0bf316),
	.w7(32'h3b045479),
	.w8(32'h3b0b0b6d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb829a),
	.w1(32'h3aad970d),
	.w2(32'h3c1a089c),
	.w3(32'hbb7b29af),
	.w4(32'h3b464f6a),
	.w5(32'h3bb8ff92),
	.w6(32'h3bcf2b31),
	.w7(32'h3c49f9c9),
	.w8(32'h3bfb08a2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1870cb),
	.w1(32'h3c7c8c47),
	.w2(32'h3cce39f6),
	.w3(32'h3b593346),
	.w4(32'h3c200fb1),
	.w5(32'h3cb1aced),
	.w6(32'hbb812261),
	.w7(32'h3c788c4e),
	.w8(32'h3c5aaf0a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb101a8),
	.w1(32'hbc70938b),
	.w2(32'hbcdebd5a),
	.w3(32'h3c3cbe1c),
	.w4(32'hbc31157b),
	.w5(32'hbcb04a11),
	.w6(32'hbc5e6657),
	.w7(32'hbc5a5e36),
	.w8(32'hbc3c03f1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd07342),
	.w1(32'h3ae996c6),
	.w2(32'hba95feea),
	.w3(32'hbcb5c5c9),
	.w4(32'h3b99e3e2),
	.w5(32'h3a0e2ef2),
	.w6(32'h3b86ff98),
	.w7(32'h3a9177a3),
	.w8(32'h3b48eb0d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d25d8c),
	.w1(32'hb9f6c412),
	.w2(32'hbb86060e),
	.w3(32'h3b3ae688),
	.w4(32'hbadf3971),
	.w5(32'hbba5074b),
	.w6(32'hbb39edaf),
	.w7(32'hbba76749),
	.w8(32'hbadba4fd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebc719),
	.w1(32'h3c00d78e),
	.w2(32'h3bd0de14),
	.w3(32'hba883c2c),
	.w4(32'h3bb2bbae),
	.w5(32'hbb07826f),
	.w6(32'h3afd3b57),
	.w7(32'hbb70066b),
	.w8(32'hba63db17),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b792d0d),
	.w1(32'h3b02e870),
	.w2(32'h3bb01979),
	.w3(32'hbbc29bac),
	.w4(32'h3b503ca3),
	.w5(32'h3b8f95e1),
	.w6(32'h3a431326),
	.w7(32'h3b676da4),
	.w8(32'h3ac53154),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e373d8),
	.w1(32'h3bcdc392),
	.w2(32'h3c0c71b2),
	.w3(32'hbb7d1201),
	.w4(32'h3bca20dc),
	.w5(32'h3ba5fb34),
	.w6(32'hbabfddff),
	.w7(32'h3acb525f),
	.w8(32'h3b9dfc88),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2caac6),
	.w1(32'h3cd38b8a),
	.w2(32'h3cefa750),
	.w3(32'h3c1ca033),
	.w4(32'h3c617359),
	.w5(32'h3ca26b12),
	.w6(32'h3b5372e7),
	.w7(32'h3c1fdea7),
	.w8(32'h3c92fc18),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d080d14),
	.w1(32'h3c98e110),
	.w2(32'h3cbd3c4b),
	.w3(32'h3ca839f5),
	.w4(32'h3bce4786),
	.w5(32'h3c5b1f61),
	.w6(32'h39c6af9d),
	.w7(32'h3c035f55),
	.w8(32'h3bd63bc0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa7745),
	.w1(32'h3942ea75),
	.w2(32'h3bc51690),
	.w3(32'h3c45d081),
	.w4(32'hbc03eda4),
	.w5(32'h3b284faf),
	.w6(32'hbb89d3ec),
	.w7(32'h3b3e101f),
	.w8(32'h3b8a6bfc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ba18),
	.w1(32'h3b00ae27),
	.w2(32'hbba28703),
	.w3(32'hbbceac5e),
	.w4(32'h3c11a008),
	.w5(32'h3bfc743e),
	.w6(32'hb8ba6a4d),
	.w7(32'hbb349a77),
	.w8(32'h3ae2a83f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f92e),
	.w1(32'hbc7b9bd5),
	.w2(32'hbccf042e),
	.w3(32'hbb99b3c4),
	.w4(32'hbc0e298b),
	.w5(32'hbc72f373),
	.w6(32'hbbb155ba),
	.w7(32'hbc9378c5),
	.w8(32'hbc10ab8c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3971cd),
	.w1(32'hbcb0a812),
	.w2(32'hbcd33142),
	.w3(32'hbc142250),
	.w4(32'hbc1a06dc),
	.w5(32'hbc8671f7),
	.w6(32'hbc690cae),
	.w7(32'hbc86f375),
	.w8(32'hbc6dc898),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab6ba9),
	.w1(32'hbb53943f),
	.w2(32'h3b478014),
	.w3(32'hbc82036a),
	.w4(32'hb9f7e09b),
	.w5(32'h3af8dcee),
	.w6(32'hbabb2769),
	.w7(32'h3b8cc049),
	.w8(32'h3bd7044a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae26afb),
	.w1(32'h3c4711e1),
	.w2(32'h3c5ad814),
	.w3(32'h3a30e10c),
	.w4(32'h3b316f0a),
	.w5(32'h3bd208b0),
	.w6(32'hbb1abbf7),
	.w7(32'h3ba50a3a),
	.w8(32'hbba5675f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4adf1),
	.w1(32'hbb426d34),
	.w2(32'h3bbcf89a),
	.w3(32'hbb538e96),
	.w4(32'h3aafb079),
	.w5(32'h3bf7f5f6),
	.w6(32'hbbf821aa),
	.w7(32'h39ce918a),
	.w8(32'hbba810b0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8a1f8),
	.w1(32'hba1649ce),
	.w2(32'hbadc9bf3),
	.w3(32'h3b591330),
	.w4(32'h3a468376),
	.w5(32'hbab639f7),
	.w6(32'hbb43898b),
	.w7(32'hbb55df77),
	.w8(32'hb7ec9fb6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0023a),
	.w1(32'h3b1bc171),
	.w2(32'h3c0b7e5c),
	.w3(32'hbc2e98c9),
	.w4(32'hbb5e0b33),
	.w5(32'h3b38c52d),
	.w6(32'h3b6a1ce2),
	.w7(32'h3bf7a7a5),
	.w8(32'h3afcab0b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cc874),
	.w1(32'h3bc8b4c3),
	.w2(32'h3c09ca38),
	.w3(32'h3bae7b60),
	.w4(32'h3b039f1b),
	.w5(32'h3bc4ea63),
	.w6(32'h3bff4c6e),
	.w7(32'h3c29c2d0),
	.w8(32'h3b22b71c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dc324),
	.w1(32'hbb9040c8),
	.w2(32'hbbb86694),
	.w3(32'h3bbce833),
	.w4(32'hbb57cbef),
	.w5(32'hbb611dcc),
	.w6(32'hbb2b5596),
	.w7(32'hbb669ecb),
	.w8(32'hbaee9f49),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d36b5),
	.w1(32'hbc15d375),
	.w2(32'hbc203f10),
	.w3(32'hba40045d),
	.w4(32'hbc4770f9),
	.w5(32'hbb9de200),
	.w6(32'hbbe3232d),
	.w7(32'hbbf2e14f),
	.w8(32'h3b59bfd2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc497c8),
	.w1(32'h39b384ee),
	.w2(32'h3a81ea7d),
	.w3(32'hbac23b3a),
	.w4(32'hbb873705),
	.w5(32'hbb624966),
	.w6(32'hbb5a7418),
	.w7(32'h3a1e5553),
	.w8(32'hb9c16890),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a638afd),
	.w1(32'hbc558cc5),
	.w2(32'hbd09d5ce),
	.w3(32'hbb23e360),
	.w4(32'hbc575e61),
	.w5(32'hbcd7b22e),
	.w6(32'hbb2ee965),
	.w7(32'hbcb3873f),
	.w8(32'h3b669089),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e73da),
	.w1(32'h3c04933d),
	.w2(32'h3c909d3e),
	.w3(32'hba8a6043),
	.w4(32'h3b7b80fc),
	.w5(32'h3bbe7ac2),
	.w6(32'h3aade0a4),
	.w7(32'h3b350f28),
	.w8(32'h3bd49a69),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f8edf),
	.w1(32'h3aa36009),
	.w2(32'hba3a0c7d),
	.w3(32'h3bce95da),
	.w4(32'h3adce20c),
	.w5(32'h3b122ee0),
	.w6(32'h3a537a24),
	.w7(32'h3b091a27),
	.w8(32'hbbca33da),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a6f7),
	.w1(32'hbadfd2d8),
	.w2(32'h38cf26ea),
	.w3(32'hbb2b79fc),
	.w4(32'hbb0eef5c),
	.w5(32'h3831ecce),
	.w6(32'hbb63a0f4),
	.w7(32'hba1d189b),
	.w8(32'hbb63f9e0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a9102),
	.w1(32'h3ab2be49),
	.w2(32'h3be03554),
	.w3(32'hb96b6e0f),
	.w4(32'h3b94b801),
	.w5(32'h3c1a6c22),
	.w6(32'hbb393de7),
	.w7(32'h3b138fb9),
	.w8(32'h3b7efd1d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb01e7),
	.w1(32'h3b0b0b88),
	.w2(32'hbc1e2056),
	.w3(32'h3c151ceb),
	.w4(32'h3bc37826),
	.w5(32'hbbb2bca2),
	.w6(32'h3bc0114f),
	.w7(32'hbc2f7bc6),
	.w8(32'h3b81ba45),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b045147),
	.w1(32'h3b82e729),
	.w2(32'hbb06dcfa),
	.w3(32'h3bb6cbd2),
	.w4(32'h3c3c8989),
	.w5(32'h3bd84393),
	.w6(32'h3b680d4f),
	.w7(32'h3bcd550a),
	.w8(32'h3c17123a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2123ae),
	.w1(32'h3a301516),
	.w2(32'h3b89aa97),
	.w3(32'h3c30131b),
	.w4(32'h3b877227),
	.w5(32'h3ad30754),
	.w6(32'hba181667),
	.w7(32'h3a329415),
	.w8(32'h3acfb1fc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10e453),
	.w1(32'hbd600885),
	.w2(32'hbd98ce1c),
	.w3(32'hbba4b87e),
	.w4(32'hbcf809c6),
	.w5(32'hbd5df81f),
	.w6(32'hbd152011),
	.w7(32'hbd464e41),
	.w8(32'hbceeceb9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd82e9e8),
	.w1(32'hbac9a602),
	.w2(32'h3b9583b8),
	.w3(32'hbd34ec05),
	.w4(32'hbc14285c),
	.w5(32'h365c470b),
	.w6(32'hbc3c3d1f),
	.w7(32'hbb284537),
	.w8(32'hb874c80b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0749),
	.w1(32'h3a41d9b7),
	.w2(32'hb9497b58),
	.w3(32'hbaa3c876),
	.w4(32'h38379450),
	.w5(32'h3a67e5a3),
	.w6(32'h3b352cce),
	.w7(32'h3b42f5e5),
	.w8(32'hba99af3e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f3ac4),
	.w1(32'hbca6da25),
	.w2(32'hbce20e3f),
	.w3(32'hbb2f93f8),
	.w4(32'hbc99e2ef),
	.w5(32'hbcb1d76b),
	.w6(32'hbc5728d6),
	.w7(32'hbcd5993d),
	.w8(32'hbc27ae3e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e64f8),
	.w1(32'h3c6ecf73),
	.w2(32'h3c1489a6),
	.w3(32'hbb133345),
	.w4(32'h3c296ec9),
	.w5(32'h3bf9d7f1),
	.w6(32'h3c723f34),
	.w7(32'h3c040db7),
	.w8(32'h3bf66d7d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30eaf9),
	.w1(32'hbd13d1d2),
	.w2(32'hbd2c248c),
	.w3(32'h3bd60be9),
	.w4(32'hbcb162a2),
	.w5(32'hbd052ed4),
	.w6(32'hbc9ca8a2),
	.w7(32'hbcdfbf82),
	.w8(32'hbca5f72f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01c7fa),
	.w1(32'hbab1fccd),
	.w2(32'hbb29d019),
	.w3(32'hbcb5d868),
	.w4(32'h3ac8f60f),
	.w5(32'hbb4a6cae),
	.w6(32'h39a1402d),
	.w7(32'hbbacdf5a),
	.w8(32'h3a8fa2e7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba236cd1),
	.w1(32'hbb2f0226),
	.w2(32'hbd1411c5),
	.w3(32'h3afb8f47),
	.w4(32'hbbe4180c),
	.w5(32'hbca779a3),
	.w6(32'h3c8d5629),
	.w7(32'hbac53db3),
	.w8(32'hbbcd6060),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule