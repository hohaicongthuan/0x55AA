module layer_10_featuremap_245(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab00a11),
	.w1(32'hbc2c82f0),
	.w2(32'h3aad64cc),
	.w3(32'hbc259aaf),
	.w4(32'h3aa1bed2),
	.w5(32'hbb2e13b1),
	.w6(32'hbc588ba2),
	.w7(32'hba5f0610),
	.w8(32'hb99570e5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4dfa3),
	.w1(32'h3b77c24f),
	.w2(32'h3c0eab25),
	.w3(32'h39fa7b89),
	.w4(32'h3ba896c7),
	.w5(32'h3bcdc08a),
	.w6(32'h3b4bd6ab),
	.w7(32'h3b4260e3),
	.w8(32'h3c1912b1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d49fc),
	.w1(32'hbbcc2c44),
	.w2(32'hbc0fa12a),
	.w3(32'hbbbbe6c2),
	.w4(32'hbb8679a0),
	.w5(32'hba61fe18),
	.w6(32'h39b8034b),
	.w7(32'hbbaa44e0),
	.w8(32'hba38172b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1eb43),
	.w1(32'hbb8be9ce),
	.w2(32'hbbf9a49f),
	.w3(32'hbba20f0f),
	.w4(32'hbbf8b9e7),
	.w5(32'hbc36becd),
	.w6(32'hba606c20),
	.w7(32'hbbeb922b),
	.w8(32'hbcb0ef6e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc638485),
	.w1(32'h3c3fa7d5),
	.w2(32'hb9600a8e),
	.w3(32'h3cada654),
	.w4(32'h3a914b40),
	.w5(32'h3b070efb),
	.w6(32'h3c85c76f),
	.w7(32'hbb62634f),
	.w8(32'h39bf7216),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62ddf2),
	.w1(32'hbb605f56),
	.w2(32'hba7ce64f),
	.w3(32'hba5ca984),
	.w4(32'h36eb5732),
	.w5(32'hbb2e136a),
	.w6(32'hba32eb7f),
	.w7(32'hbb12f7b0),
	.w8(32'hbb744401),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb709955),
	.w1(32'hbc31aca6),
	.w2(32'hbcdbb07c),
	.w3(32'hbb6d6c6e),
	.w4(32'hbc6d63b0),
	.w5(32'hbcc5c8c8),
	.w6(32'hbb227ea3),
	.w7(32'hbc9da002),
	.w8(32'hbcb08003),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a659),
	.w1(32'h3b235a58),
	.w2(32'h3bce6145),
	.w3(32'hba3fdcd7),
	.w4(32'h3b2e92d2),
	.w5(32'h3ca7c838),
	.w6(32'hbb04d82b),
	.w7(32'hbb1bcfbd),
	.w8(32'h3c1b7b27),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9b436),
	.w1(32'h399bdd83),
	.w2(32'h38dc7e38),
	.w3(32'h3b77d7ec),
	.w4(32'h3b0935e3),
	.w5(32'h3b138e68),
	.w6(32'hba8c003a),
	.w7(32'hba2aa786),
	.w8(32'h3ad4434e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ac54a),
	.w1(32'hbb995324),
	.w2(32'hbb778b1b),
	.w3(32'h3ba5d5b0),
	.w4(32'hba64afaf),
	.w5(32'h3b1414cd),
	.w6(32'h3b8135be),
	.w7(32'hbc3baefb),
	.w8(32'hbbe11712),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c67d2),
	.w1(32'hbb05c086),
	.w2(32'h3aa23fdb),
	.w3(32'h39d2db06),
	.w4(32'h3ac0af0a),
	.w5(32'hb7106eac),
	.w6(32'h3b9c02d6),
	.w7(32'h3b331f61),
	.w8(32'h3b06b424),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c388c2e),
	.w1(32'hbb715f8c),
	.w2(32'hbc82ffcc),
	.w3(32'hb98761bb),
	.w4(32'hbc37d0de),
	.w5(32'hbce0c514),
	.w6(32'h3a84c8a2),
	.w7(32'hbc7ca49b),
	.w8(32'hbcb73f92),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0df258),
	.w1(32'h39f1fc61),
	.w2(32'hbc19f723),
	.w3(32'h3ba85e0c),
	.w4(32'hbc3321e4),
	.w5(32'hbc202287),
	.w6(32'h3a48ac45),
	.w7(32'hbc63b258),
	.w8(32'hbc642a14),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2783fc),
	.w1(32'h3cbd0518),
	.w2(32'hbaa9f4f2),
	.w3(32'h3d121a29),
	.w4(32'hbc07078b),
	.w5(32'h3bca5b9d),
	.w6(32'h3d158182),
	.w7(32'hbc27c120),
	.w8(32'h3bc9132a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeffac),
	.w1(32'h3b7f7381),
	.w2(32'h3c0cfc42),
	.w3(32'h3c03feb8),
	.w4(32'h3b25d8d5),
	.w5(32'h3b922177),
	.w6(32'h3b945a85),
	.w7(32'h3af44ca1),
	.w8(32'h3b38f8b0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0243),
	.w1(32'hb94dd451),
	.w2(32'h3c03de24),
	.w3(32'h3c0fd9e7),
	.w4(32'h3c1b198a),
	.w5(32'h3cb27644),
	.w6(32'h3c097389),
	.w7(32'hbb596f79),
	.w8(32'h3c8207ab),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b662e2e),
	.w1(32'h39aa99c4),
	.w2(32'h3a9fea1e),
	.w3(32'h3b2722bb),
	.w4(32'h3be179f0),
	.w5(32'hbba399d4),
	.w6(32'hbac519bd),
	.w7(32'h3a0d53d1),
	.w8(32'hbb8c0050),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90aad1),
	.w1(32'h3a2d398c),
	.w2(32'hbbcf7cb7),
	.w3(32'h3bd37c08),
	.w4(32'hbaf6bcdf),
	.w5(32'hba6f9c09),
	.w6(32'h3bcce400),
	.w7(32'hbc5a0273),
	.w8(32'hbb66c3cd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888e5b),
	.w1(32'hbb55ae0e),
	.w2(32'hbb6547cc),
	.w3(32'h3b3e0da6),
	.w4(32'hbbeb51ad),
	.w5(32'hbc956afc),
	.w6(32'h3b556d7e),
	.w7(32'hbb89e1d0),
	.w8(32'hbcb6fb88),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc815227),
	.w1(32'hbba8c851),
	.w2(32'hbc82f32c),
	.w3(32'hbb6e9b57),
	.w4(32'hbc9dcd9b),
	.w5(32'hbb53fe51),
	.w6(32'h3a6e7c21),
	.w7(32'hbc852cb2),
	.w8(32'hbb893c21),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92eb5b),
	.w1(32'hbaefa0e2),
	.w2(32'h3b070a7f),
	.w3(32'hbb423ad3),
	.w4(32'h3b78fccb),
	.w5(32'h3b959334),
	.w6(32'h3a5fcad6),
	.w7(32'h3b9727cd),
	.w8(32'h3b4976b1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e31735),
	.w1(32'h3a7c442d),
	.w2(32'h3b6f9ea4),
	.w3(32'hb9a7b0f6),
	.w4(32'h3afabacf),
	.w5(32'h3b55fdcf),
	.w6(32'hbbacfa18),
	.w7(32'hba94cd15),
	.w8(32'hb7dd3d30),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf80ec),
	.w1(32'hbc486b6b),
	.w2(32'hbc7a173a),
	.w3(32'h3c297013),
	.w4(32'hbc4d8bdf),
	.w5(32'hbb84b685),
	.w6(32'h3b9418bd),
	.w7(32'hbce58126),
	.w8(32'hbbd76cff),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d07d2),
	.w1(32'hbad941ed),
	.w2(32'hbb2132e9),
	.w3(32'h3c3d5d7f),
	.w4(32'hbbbbdc6f),
	.w5(32'h3bd1401d),
	.w6(32'h3c9351a4),
	.w7(32'hbc66f27a),
	.w8(32'hba87c5b7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b188f),
	.w1(32'hbbbc85d9),
	.w2(32'h3b989267),
	.w3(32'hbbe123d5),
	.w4(32'hbc35c8e8),
	.w5(32'h3c0ce296),
	.w6(32'hba1857aa),
	.w7(32'hbc3fc2c7),
	.w8(32'h3c01d75f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4f23d),
	.w1(32'hb99c60c4),
	.w2(32'hba01918a),
	.w3(32'hb9062858),
	.w4(32'hb9131dc0),
	.w5(32'h3bcd62d3),
	.w6(32'h3ad62d08),
	.w7(32'hbb88b672),
	.w8(32'h3b5fe962),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21c8f0),
	.w1(32'h3b0827fe),
	.w2(32'hbaca2e86),
	.w3(32'h3b9252aa),
	.w4(32'hbb234e98),
	.w5(32'h3a973b0d),
	.w6(32'h3ad8dabf),
	.w7(32'hbabf0e64),
	.w8(32'hbb79cf5d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005f2f),
	.w1(32'hbc9916fb),
	.w2(32'hbc579ea4),
	.w3(32'hbc04fa70),
	.w4(32'hbbd6de55),
	.w5(32'h3b887fd6),
	.w6(32'hbc25c8fa),
	.w7(32'hbc821a90),
	.w8(32'h3c2e2d17),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1e761),
	.w1(32'h3cb52ed0),
	.w2(32'h3d0a6b5a),
	.w3(32'h3c9611bd),
	.w4(32'h3cb90ae0),
	.w5(32'hbb429095),
	.w6(32'h3d1e5ca6),
	.w7(32'h3d200ed2),
	.w8(32'hbba3db79),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225a9b),
	.w1(32'hbbbb0e64),
	.w2(32'h399bbe9b),
	.w3(32'hbc060ca8),
	.w4(32'hbc514dc1),
	.w5(32'hbc1d4a26),
	.w6(32'h3b58f08d),
	.w7(32'hbc2f89e9),
	.w8(32'hbc060006),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88db7e),
	.w1(32'hbb143cb2),
	.w2(32'hbbacab5f),
	.w3(32'h3ad3ec3e),
	.w4(32'h3ad77e52),
	.w5(32'h3a8b39db),
	.w6(32'h37cd9da3),
	.w7(32'hbb670e21),
	.w8(32'h3a2f12ab),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06781c),
	.w1(32'hba65144a),
	.w2(32'h3beaf3ef),
	.w3(32'hbae20fb1),
	.w4(32'h3bcbf79e),
	.w5(32'hbb6164ac),
	.w6(32'h3ad98aa9),
	.w7(32'h3bc4824e),
	.w8(32'hba40f85a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a489),
	.w1(32'hbc1ed38b),
	.w2(32'hbb6cbd41),
	.w3(32'hba31629c),
	.w4(32'hbb6435c1),
	.w5(32'hbb4188aa),
	.w6(32'h3ab9a414),
	.w7(32'hbc19f814),
	.w8(32'hbb852274),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadee810),
	.w1(32'h3b4c737c),
	.w2(32'hbb261c87),
	.w3(32'h3b0678ae),
	.w4(32'h39d59a71),
	.w5(32'h3af0f2b9),
	.w6(32'h3c07192f),
	.w7(32'hbb800d72),
	.w8(32'hbbd01f04),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf92bd7),
	.w1(32'hbc8168e6),
	.w2(32'hbc3a80e9),
	.w3(32'hbc6761c4),
	.w4(32'hbc88f05d),
	.w5(32'hbb46900b),
	.w6(32'hbba0a6f0),
	.w7(32'hbc643ea0),
	.w8(32'hbb3d4ed5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3070a5),
	.w1(32'hbb7d8c94),
	.w2(32'hbc1dc778),
	.w3(32'h3b7f92de),
	.w4(32'h3997e174),
	.w5(32'hbb233fd0),
	.w6(32'hbaf71428),
	.w7(32'hbbaa5450),
	.w8(32'hbbaf65a9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c745150),
	.w1(32'h3c958337),
	.w2(32'h3b934cd0),
	.w3(32'h3c9d128b),
	.w4(32'h3c7fe739),
	.w5(32'h3c5c0415),
	.w6(32'h3cbdca77),
	.w7(32'h3c3f8bbd),
	.w8(32'hbc9d083e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dcb01),
	.w1(32'hbbf48a51),
	.w2(32'h3bd815e0),
	.w3(32'hbc1159da),
	.w4(32'hbc79c494),
	.w5(32'h395b95cc),
	.w6(32'hbc0cfde0),
	.w7(32'hbc533774),
	.w8(32'h385b6cd0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb353fe7),
	.w1(32'hbcaac6ec),
	.w2(32'hbc477ba2),
	.w3(32'hbc72e552),
	.w4(32'hbd0adae4),
	.w5(32'hbc854128),
	.w6(32'hbc3257fa),
	.w7(32'hbce19f77),
	.w8(32'hbbd31550),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5382d),
	.w1(32'h39a6cc32),
	.w2(32'hbb2aa16f),
	.w3(32'h3ae7a277),
	.w4(32'hba4f63c6),
	.w5(32'h3c005c1c),
	.w6(32'hb9411731),
	.w7(32'hbb5d4f90),
	.w8(32'h3bfe637a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cace8),
	.w1(32'h3c92e56e),
	.w2(32'h3c34d1ed),
	.w3(32'h3c50f469),
	.w4(32'h3c557e62),
	.w5(32'hbb31cbb6),
	.w6(32'h3ca7121c),
	.w7(32'h3c111c28),
	.w8(32'hbb8ca1da),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73aab1),
	.w1(32'hbb0a6219),
	.w2(32'hbbad1656),
	.w3(32'h3a431f70),
	.w4(32'h3a0cd1a4),
	.w5(32'hbb7404e8),
	.w6(32'hb9b2ab1f),
	.w7(32'hbbc9c0d9),
	.w8(32'hba2c700f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c1b99),
	.w1(32'hb96e1ef2),
	.w2(32'hbac27984),
	.w3(32'hbb161541),
	.w4(32'hbbba93c0),
	.w5(32'hbb271be2),
	.w6(32'h3ab17fe4),
	.w7(32'hba3556ae),
	.w8(32'hbb575784),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806209),
	.w1(32'hbbd0d130),
	.w2(32'h3b30dce9),
	.w3(32'h3b56edd8),
	.w4(32'hbb0c4bc4),
	.w5(32'hbbd9c7a4),
	.w6(32'h3b8ea0d7),
	.w7(32'hbc5b0adb),
	.w8(32'hbbc9a5ca),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb0444),
	.w1(32'h39958820),
	.w2(32'h3ba084d5),
	.w3(32'h3b2d7755),
	.w4(32'h3b41f3b2),
	.w5(32'h3c124501),
	.w6(32'h3bd7b3f2),
	.w7(32'h3a842f46),
	.w8(32'h3b72cf18),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ffd45),
	.w1(32'h3bc72802),
	.w2(32'h3b66f83a),
	.w3(32'h3c1f0730),
	.w4(32'hbac7a8b7),
	.w5(32'h3bb66d4b),
	.w6(32'h3b3164a8),
	.w7(32'hbb9a7ec8),
	.w8(32'h3b81a2c6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0700d0),
	.w1(32'h3bc478ea),
	.w2(32'h3b2e8f3e),
	.w3(32'h3c30e15b),
	.w4(32'hb83a5f73),
	.w5(32'h3be887af),
	.w6(32'h3c4d1736),
	.w7(32'hbabbfc06),
	.w8(32'h3b215dc0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bb69c),
	.w1(32'hbbb5e0e9),
	.w2(32'hbc692651),
	.w3(32'h3c45ac24),
	.w4(32'h3aa1a28a),
	.w5(32'hbbd4b601),
	.w6(32'hbb9e0237),
	.w7(32'hbcabd8df),
	.w8(32'hbc8d4b01),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e8ec),
	.w1(32'h3b503798),
	.w2(32'hba4bce41),
	.w3(32'hbaee80eb),
	.w4(32'hbb59ace3),
	.w5(32'h39980180),
	.w6(32'hbb8b47c9),
	.w7(32'hbb34dc07),
	.w8(32'hbb104f16),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae72cb8),
	.w1(32'hbad1181b),
	.w2(32'hbbb12ba5),
	.w3(32'h3977bb3c),
	.w4(32'hbb199a03),
	.w5(32'hbb1584dc),
	.w6(32'hbba0b3e6),
	.w7(32'hbba2770a),
	.w8(32'hbb9daab7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29e054),
	.w1(32'h3c099873),
	.w2(32'hbbca05bd),
	.w3(32'h3ba72726),
	.w4(32'hbb606081),
	.w5(32'hbb5ea027),
	.w6(32'h3c81f6a5),
	.w7(32'h3a24f522),
	.w8(32'hbab70859),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f43ef),
	.w1(32'hbb392b62),
	.w2(32'hbb1cd0c7),
	.w3(32'hba0c49b9),
	.w4(32'hbb32081c),
	.w5(32'h3ade796b),
	.w6(32'hbab2f4e4),
	.w7(32'hbb91b2df),
	.w8(32'h3c36d2b8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbad584),
	.w1(32'h3c249c50),
	.w2(32'h3cb0dc2f),
	.w3(32'h3c8ae7aa),
	.w4(32'h3cfb1008),
	.w5(32'hbad11beb),
	.w6(32'h3d177d56),
	.w7(32'h3d0c0db5),
	.w8(32'hbb79002b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa842),
	.w1(32'hbbb867a8),
	.w2(32'hbc2c5158),
	.w3(32'h3c0a40a3),
	.w4(32'hbb246e3e),
	.w5(32'hbc28b927),
	.w6(32'h3be605c6),
	.w7(32'hbc3a743c),
	.w8(32'hbc9c9ded),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93e241),
	.w1(32'hbc3f96b7),
	.w2(32'hbbedcdaa),
	.w3(32'hbc809b39),
	.w4(32'hbb4f8164),
	.w5(32'hbb27693f),
	.w6(32'hbc57b2c5),
	.w7(32'hbbdcf168),
	.w8(32'hbbc9ff16),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6b95e),
	.w1(32'hbc190732),
	.w2(32'hbb01998c),
	.w3(32'hbba6daed),
	.w4(32'hbbdaf9ed),
	.w5(32'h3c1eb13e),
	.w6(32'h3c0dfd18),
	.w7(32'hbbc60645),
	.w8(32'h3b157e49),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147355),
	.w1(32'h3c1e4590),
	.w2(32'h3c2298f2),
	.w3(32'h3c493c94),
	.w4(32'h3c2c804e),
	.w5(32'hbbe2b08d),
	.w6(32'h3c7f229b),
	.w7(32'h3bf2b990),
	.w8(32'hbb3aa8fe),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44f959),
	.w1(32'h39dddc1d),
	.w2(32'h3b4420a0),
	.w3(32'h3afd9f77),
	.w4(32'h3b9e1af1),
	.w5(32'hbb621d33),
	.w6(32'h3c4e6a9d),
	.w7(32'h3ba5ba5a),
	.w8(32'hbbb3c1ca),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d35d6),
	.w1(32'hbb2f30ed),
	.w2(32'hbba67879),
	.w3(32'hb9d8cf43),
	.w4(32'hbb87700a),
	.w5(32'h3a606e56),
	.w6(32'hbbb36ef1),
	.w7(32'hbbf94765),
	.w8(32'h3ac50a7f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c5f1b),
	.w1(32'hba151931),
	.w2(32'hbbf106f6),
	.w3(32'hbb78b92d),
	.w4(32'hbbebdd1d),
	.w5(32'hbb560878),
	.w6(32'hbc0b32eb),
	.w7(32'hbbf9138f),
	.w8(32'hbb46e201),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4e92c),
	.w1(32'hbaefe6a1),
	.w2(32'hb8713467),
	.w3(32'h3b8c4f1b),
	.w4(32'hbb3e4543),
	.w5(32'h3b2348f2),
	.w6(32'h3b526a0b),
	.w7(32'hbbf6f918),
	.w8(32'h39c6a8c4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b376f),
	.w1(32'hbb942596),
	.w2(32'h3abdc992),
	.w3(32'hbb078687),
	.w4(32'hbaa624d0),
	.w5(32'h3bbe3195),
	.w6(32'hbb1c5343),
	.w7(32'hbc86cbf7),
	.w8(32'h3bce24a0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c0bf),
	.w1(32'hbc11085e),
	.w2(32'hb9eb6ca5),
	.w3(32'hbb2f3113),
	.w4(32'h3c75812a),
	.w5(32'hbbc0aeb9),
	.w6(32'hb89d4290),
	.w7(32'h3b36211b),
	.w8(32'hbc57b64c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c6fcc),
	.w1(32'h3b18043c),
	.w2(32'h3bb76713),
	.w3(32'h3b29ea28),
	.w4(32'hbabf2bd0),
	.w5(32'hbc14fb02),
	.w6(32'h3c422369),
	.w7(32'h3a5d309e),
	.w8(32'hbc2df8fb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fdd44),
	.w1(32'hbc9dde12),
	.w2(32'h3c345337),
	.w3(32'hbcbacf16),
	.w4(32'h3c8575df),
	.w5(32'h3a74af53),
	.w6(32'hbc7f91ba),
	.w7(32'h3c185e63),
	.w8(32'h3bbf8a8f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d3734),
	.w1(32'h3baec02c),
	.w2(32'h3be211f9),
	.w3(32'h3b88e44a),
	.w4(32'h3c8cc7c9),
	.w5(32'hbb4a25da),
	.w6(32'h3c4c79d2),
	.w7(32'h3c88f245),
	.w8(32'hbad2c14a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a5a30),
	.w1(32'hbbc9401b),
	.w2(32'hbc228ee1),
	.w3(32'h3be64067),
	.w4(32'h3a2f77cf),
	.w5(32'h3b8586da),
	.w6(32'h3b65950a),
	.w7(32'hbc75e5ea),
	.w8(32'hbbf7b8be),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3836c4),
	.w1(32'h3bcef187),
	.w2(32'h3c2593be),
	.w3(32'h3c2b14d8),
	.w4(32'hbc3997f6),
	.w5(32'hbc20c3a6),
	.w6(32'h3a3f95ef),
	.w7(32'hbbf6634a),
	.w8(32'hbc10a577),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad0b7),
	.w1(32'hbcababa1),
	.w2(32'h3c37a76a),
	.w3(32'hbc2b2e95),
	.w4(32'hbaf4280e),
	.w5(32'hbae99116),
	.w6(32'hbc276655),
	.w7(32'hbc1217e3),
	.w8(32'hbb9b66d1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c433),
	.w1(32'h3a9b416b),
	.w2(32'h3c5fb8c1),
	.w3(32'hba0001ec),
	.w4(32'hbb00076a),
	.w5(32'h3c01722c),
	.w6(32'hbc321ebc),
	.w7(32'hbbe35cce),
	.w8(32'h3c0b6ef5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4167c5),
	.w1(32'h3b87d616),
	.w2(32'h3badb395),
	.w3(32'h3b809d73),
	.w4(32'h3aa7607f),
	.w5(32'hbbcfce3c),
	.w6(32'h3b9f7947),
	.w7(32'h3bbb2c4a),
	.w8(32'hbc0d349d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e73d5),
	.w1(32'hbb4ec08f),
	.w2(32'hb93a9b83),
	.w3(32'hbc1b9e51),
	.w4(32'h3b865aa6),
	.w5(32'hbb939adb),
	.w6(32'hbb4ef2a6),
	.w7(32'h3b8a8208),
	.w8(32'hba3490e7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f28aa1),
	.w1(32'hbb6fc069),
	.w2(32'hbb15581c),
	.w3(32'hbb2163a1),
	.w4(32'hb98735b4),
	.w5(32'h3984dfcf),
	.w6(32'hbb9f28c2),
	.w7(32'hbb9105ea),
	.w8(32'h3b5b8bae),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29467c),
	.w1(32'hbb19f83a),
	.w2(32'hbbdd876a),
	.w3(32'h39f16a7e),
	.w4(32'hba8dcae1),
	.w5(32'h3ac4add6),
	.w6(32'h3b3a2550),
	.w7(32'hbbc75d07),
	.w8(32'h3ac210b0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92688e),
	.w1(32'hbaa363e6),
	.w2(32'h3b56e16c),
	.w3(32'h397641e2),
	.w4(32'h3ac442ca),
	.w5(32'hbbad0cb9),
	.w6(32'h3b7879aa),
	.w7(32'h3abbf968),
	.w8(32'hbb15a9d4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca0b32),
	.w1(32'h3b6f7452),
	.w2(32'hbbe61b31),
	.w3(32'h3ba8bda1),
	.w4(32'hbb3b6f5f),
	.w5(32'hbc3cf789),
	.w6(32'h3b1a1542),
	.w7(32'hbbd965dc),
	.w8(32'hbc8a988c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c448675),
	.w1(32'h3ba12420),
	.w2(32'hbc10ac10),
	.w3(32'h3b4220e0),
	.w4(32'hbb958f19),
	.w5(32'h3b07a4f7),
	.w6(32'h3c3845db),
	.w7(32'hbbd4374e),
	.w8(32'hbbfe53ba),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af27701),
	.w1(32'h3b9866f7),
	.w2(32'h3b803b82),
	.w3(32'h3bf110b8),
	.w4(32'h3b3e4213),
	.w5(32'h3be255d9),
	.w6(32'h3c1ad093),
	.w7(32'h3ab20a6f),
	.w8(32'h3bfd1f66),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa96f5e),
	.w1(32'h3a848709),
	.w2(32'h3b60a519),
	.w3(32'h3b2af942),
	.w4(32'hbb15adb6),
	.w5(32'h3c1f7d93),
	.w6(32'hbb424133),
	.w7(32'hbb9105e2),
	.w8(32'h3bb70dd1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d944a),
	.w1(32'hbb5e6ca9),
	.w2(32'hbc189068),
	.w3(32'h3971be8a),
	.w4(32'hbb825873),
	.w5(32'hbc015a5f),
	.w6(32'h3aa3c54a),
	.w7(32'hbc31b6ee),
	.w8(32'hbbfc5159),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e297),
	.w1(32'h3b6f4888),
	.w2(32'h3b99bd66),
	.w3(32'h3a9d766f),
	.w4(32'h3b2581c1),
	.w5(32'hbb32868c),
	.w6(32'hbb3da870),
	.w7(32'hbb23b09f),
	.w8(32'hbad438e7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6c91),
	.w1(32'hbb209f47),
	.w2(32'hbc256af7),
	.w3(32'hbadadac1),
	.w4(32'hbba96d3e),
	.w5(32'h3bf342c1),
	.w6(32'hbbde8bc6),
	.w7(32'hbc2f481d),
	.w8(32'hbc68753f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52ca3a),
	.w1(32'hbc6613a7),
	.w2(32'h3c592b9e),
	.w3(32'hbc2fe666),
	.w4(32'h3bb48757),
	.w5(32'hbbdc26d5),
	.w6(32'hbc862bd5),
	.w7(32'h3bab30e3),
	.w8(32'h3a65f1e3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada3b50),
	.w1(32'h38b774fd),
	.w2(32'hbb7ae918),
	.w3(32'h3b0c5461),
	.w4(32'hbb9c3860),
	.w5(32'h3c8996b2),
	.w6(32'h3c103500),
	.w7(32'hbbbdc33f),
	.w8(32'h3c343b32),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c203e4b),
	.w1(32'h3a97a615),
	.w2(32'h3c4917eb),
	.w3(32'h3b8957b4),
	.w4(32'h3c47b69b),
	.w5(32'h3a508b67),
	.w6(32'hbb34d3ea),
	.w7(32'h3c3745fa),
	.w8(32'h3aa20bd4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3e95b),
	.w1(32'hbc0a21ac),
	.w2(32'hbb884bee),
	.w3(32'hbb9b6e20),
	.w4(32'hbbf8a39f),
	.w5(32'hbb7b9301),
	.w6(32'hba27a6c3),
	.w7(32'hbb219e94),
	.w8(32'hbb88b998),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ff5c),
	.w1(32'hbb4441be),
	.w2(32'h3b74e9eb),
	.w3(32'h3a5594df),
	.w4(32'hb691685d),
	.w5(32'hbc224f99),
	.w6(32'h3b6ba9aa),
	.w7(32'hbb8b5b28),
	.w8(32'hbc6c01b4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b650a),
	.w1(32'hbc15f12e),
	.w2(32'hbbca8850),
	.w3(32'hbc519dec),
	.w4(32'hbc81a028),
	.w5(32'h3b54e474),
	.w6(32'hbc4a90e6),
	.w7(32'hbc2b28e0),
	.w8(32'h3b0f6ec5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98a8a6),
	.w1(32'h3be3f0a8),
	.w2(32'h3c157c3a),
	.w3(32'h3be83431),
	.w4(32'h3b9b8a2c),
	.w5(32'h3c687878),
	.w6(32'h3a34bc1b),
	.w7(32'h3b324f8b),
	.w8(32'h3bf208f2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc8154),
	.w1(32'h3ad3f652),
	.w2(32'hbc09ff7e),
	.w3(32'h3bcc66e2),
	.w4(32'h3a5ab653),
	.w5(32'h3ba0a7bb),
	.w6(32'h3c2daf4a),
	.w7(32'hbc2d033c),
	.w8(32'hbbc22890),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bec52),
	.w1(32'hbb5b9592),
	.w2(32'hbc053b98),
	.w3(32'hbbb57803),
	.w4(32'hbc1a988a),
	.w5(32'hbc0bf22c),
	.w6(32'hbbcb25e1),
	.w7(32'hbc3db4a9),
	.w8(32'hbb640862),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f64ce),
	.w1(32'hbbb5fc1f),
	.w2(32'hbbe8b732),
	.w3(32'h3c55b96f),
	.w4(32'h3b341bd5),
	.w5(32'hbb109b63),
	.w6(32'h3cb2a1f0),
	.w7(32'hbba52ba8),
	.w8(32'hbc825e5b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd212c9),
	.w1(32'h3ab22215),
	.w2(32'hba16baf5),
	.w3(32'hbad1d61a),
	.w4(32'hbc6e685a),
	.w5(32'h3ae96ff3),
	.w6(32'hbb43b0ea),
	.w7(32'hbc7bf9d2),
	.w8(32'h3a5c6164),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb8ba9),
	.w1(32'hbab60be2),
	.w2(32'h3c6a3b36),
	.w3(32'h3c0e2be6),
	.w4(32'h3b92d5fb),
	.w5(32'h3c0dd09c),
	.w6(32'h3c377dcd),
	.w7(32'hba885a08),
	.w8(32'h3ba9a3fb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827fa6),
	.w1(32'hbbe097cf),
	.w2(32'hbba02252),
	.w3(32'hbba1c398),
	.w4(32'hb914fd15),
	.w5(32'h3a9f57b3),
	.w6(32'hbb0550a0),
	.w7(32'hbb8dc878),
	.w8(32'h3affa8af),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9dfe7),
	.w1(32'hbbd1ff38),
	.w2(32'h3b93bbd9),
	.w3(32'hbc40fe24),
	.w4(32'hbc504ce0),
	.w5(32'h3b8c3c07),
	.w6(32'hbba06058),
	.w7(32'hbbdbdd70),
	.w8(32'h3c182b12),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09910c),
	.w1(32'h3a1805dc),
	.w2(32'hbb38b520),
	.w3(32'h3b0a779d),
	.w4(32'hbb6c0eb7),
	.w5(32'h3c026306),
	.w6(32'hbb5a1c9a),
	.w7(32'hbae45463),
	.w8(32'h3c0463e8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94085a),
	.w1(32'h3b6457c7),
	.w2(32'h3acbb2b2),
	.w3(32'h3c96d425),
	.w4(32'h3bfd367a),
	.w5(32'h3a417045),
	.w6(32'h3cc81805),
	.w7(32'hba3cec86),
	.w8(32'hbb138fa7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b46a5),
	.w1(32'hbbb182c9),
	.w2(32'hbc9ebe16),
	.w3(32'h3a9b9c4c),
	.w4(32'hbbcccb1d),
	.w5(32'hbbf30262),
	.w6(32'h3addbef5),
	.w7(32'hbc9541bf),
	.w8(32'hbc81ec67),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8b6f2),
	.w1(32'h3c0ba665),
	.w2(32'h3c71756f),
	.w3(32'h3c3bd602),
	.w4(32'h3c0dff84),
	.w5(32'h3c4e4299),
	.w6(32'h3c206b7c),
	.w7(32'h3c717daa),
	.w8(32'hbbe74348),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baed731),
	.w1(32'hbabb272b),
	.w2(32'h3b967891),
	.w3(32'hbba6f1e3),
	.w4(32'hbbe247c3),
	.w5(32'h3b609195),
	.w6(32'h3ad17d8f),
	.w7(32'h3ac1fb2f),
	.w8(32'h3bff7140),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0274f3),
	.w1(32'h3baa4d26),
	.w2(32'h3c34ae8a),
	.w3(32'h39f93796),
	.w4(32'h3b0ac9d0),
	.w5(32'h3bf55aca),
	.w6(32'h3adc6a44),
	.w7(32'hba1d1063),
	.w8(32'h3ba52336),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c490e43),
	.w1(32'hbc160b1c),
	.w2(32'hbc2d57c5),
	.w3(32'h3b9d7636),
	.w4(32'hbbea7d52),
	.w5(32'hbc0bd0d1),
	.w6(32'h3b984549),
	.w7(32'hbc80ad0a),
	.w8(32'hbcb7aba9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cc520),
	.w1(32'hba326710),
	.w2(32'hba2c49a9),
	.w3(32'hb90fc521),
	.w4(32'hba6b4d47),
	.w5(32'hb98ba0f4),
	.w6(32'hb82d56e5),
	.w7(32'h39a90edd),
	.w8(32'h39c0e4bb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351267),
	.w1(32'h3c57cc5d),
	.w2(32'h3c595982),
	.w3(32'h3c04d850),
	.w4(32'h3b47217e),
	.w5(32'h3c897572),
	.w6(32'h3c104134),
	.w7(32'h3be2592d),
	.w8(32'h3b084b99),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341d68),
	.w1(32'hbbb22635),
	.w2(32'hbc3caf0b),
	.w3(32'hbbaa8e4b),
	.w4(32'hbbd20194),
	.w5(32'hbc224fe7),
	.w6(32'hbb2e87d6),
	.w7(32'hbbde51c9),
	.w8(32'hbc5130eb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9732cd2),
	.w1(32'hb89245a4),
	.w2(32'h3930b83f),
	.w3(32'hb9846890),
	.w4(32'h36df40ec),
	.w5(32'h3978eaaf),
	.w6(32'hb88a1714),
	.w7(32'h38e4ff2e),
	.w8(32'h39d7603b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb837866e),
	.w1(32'h3aad5b2f),
	.w2(32'h3ba94c39),
	.w3(32'hb9c502ba),
	.w4(32'h3b971204),
	.w5(32'h3bae684c),
	.w6(32'hb7930365),
	.w7(32'h3a7fac4d),
	.w8(32'h3b77dcc9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc169be),
	.w1(32'h3a2a7612),
	.w2(32'h3a48e0ca),
	.w3(32'h3b87c7d8),
	.w4(32'h38971199),
	.w5(32'h386ee3db),
	.w6(32'h3b0c6d4a),
	.w7(32'hbb40b32b),
	.w8(32'hbb50ea99),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab088e9),
	.w1(32'h3abdc9ac),
	.w2(32'h3b996d4b),
	.w3(32'hb9cad6e5),
	.w4(32'hba255804),
	.w5(32'h3b1a6ab1),
	.w6(32'h3ac31a8e),
	.w7(32'hbb06dace),
	.w8(32'h3a033d04),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dfb09),
	.w1(32'hbc0da412),
	.w2(32'hbbb17413),
	.w3(32'hbbad65eb),
	.w4(32'hbc2139ef),
	.w5(32'hbc06cd81),
	.w6(32'hbb5775b1),
	.w7(32'hbc181139),
	.w8(32'hbb1bcf7e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bb5f4),
	.w1(32'h3b249b6f),
	.w2(32'h3bd72fa7),
	.w3(32'h3aeb5f5c),
	.w4(32'h3ab5e85b),
	.w5(32'h3bc161d1),
	.w6(32'h3b1b72cb),
	.w7(32'h3b38f562),
	.w8(32'h3bba119d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be95545),
	.w1(32'h3baa4555),
	.w2(32'h3a41d4be),
	.w3(32'h3bbbda3f),
	.w4(32'hb9c25262),
	.w5(32'hbb13e78a),
	.w6(32'h3b9f2932),
	.w7(32'hb9d38f3c),
	.w8(32'hb9d68447),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82a436),
	.w1(32'hb889c13a),
	.w2(32'h3c33183c),
	.w3(32'h3acbbfeb),
	.w4(32'h3bdcaea0),
	.w5(32'h3c5d5f94),
	.w6(32'h3b939993),
	.w7(32'h3b9d7e54),
	.w8(32'h3c4aae7b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45ed95),
	.w1(32'h3984e752),
	.w2(32'h3ab0945d),
	.w3(32'h3b1a3129),
	.w4(32'h393842b5),
	.w5(32'h3a6d592b),
	.w6(32'h3b1344bf),
	.w7(32'hba36bdf2),
	.w8(32'hba39c1b0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39137dca),
	.w1(32'h394d8702),
	.w2(32'h391efd3d),
	.w3(32'h3833671f),
	.w4(32'h3904e895),
	.w5(32'h38c5a769),
	.w6(32'hb8889661),
	.w7(32'h388e958e),
	.w8(32'h38c8c91a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb07a4),
	.w1(32'h3abb6f89),
	.w2(32'h3ab83544),
	.w3(32'h38cfc54e),
	.w4(32'h3abf7366),
	.w5(32'h3aa64a42),
	.w6(32'h3a0c89ef),
	.w7(32'h3a92c515),
	.w8(32'h3a362f2e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38027421),
	.w1(32'hb8651e95),
	.w2(32'hb602adb1),
	.w3(32'h384b7119),
	.w4(32'hb82b2f77),
	.w5(32'hb8cae427),
	.w6(32'h38413623),
	.w7(32'hb7d41cb0),
	.w8(32'hb8732e8a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8caff30),
	.w1(32'hb679f68b),
	.w2(32'hb8a0135e),
	.w3(32'hb9535493),
	.w4(32'hb85633bc),
	.w5(32'hb91e6b26),
	.w6(32'hb9844748),
	.w7(32'hb9334c88),
	.w8(32'hb933c748),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6330c8),
	.w1(32'h3aa49341),
	.w2(32'h3b62b06d),
	.w3(32'h3ae3c0fc),
	.w4(32'hb8ed3902),
	.w5(32'h3a92dc7a),
	.w6(32'h3b073548),
	.w7(32'hbac467db),
	.w8(32'hba1f31fa),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ca033),
	.w1(32'h3811e63d),
	.w2(32'h388ccd89),
	.w3(32'h38fe7b9f),
	.w4(32'h38460e2b),
	.w5(32'h39d0a10b),
	.w6(32'h3984085b),
	.w7(32'h381ba322),
	.w8(32'h3997f6bc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d4547),
	.w1(32'hbb932b8e),
	.w2(32'hbbf7e294),
	.w3(32'h3b1aaef8),
	.w4(32'hbb7b2a75),
	.w5(32'hbb6ded9c),
	.w6(32'hbab9f15a),
	.w7(32'hbc1afed9),
	.w8(32'hbc0d5b76),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e7d0f),
	.w1(32'h3bac2ef8),
	.w2(32'h3c6c6e3b),
	.w3(32'h3836f503),
	.w4(32'h39f857b4),
	.w5(32'h3c3179db),
	.w6(32'h3a564005),
	.w7(32'h3b18744b),
	.w8(32'h3c5ceb6b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962dc64),
	.w1(32'h379ce68e),
	.w2(32'h388873ed),
	.w3(32'hb91798d2),
	.w4(32'h372ac1af),
	.w5(32'h37fdfc6b),
	.w6(32'hb9382c2e),
	.w7(32'hb80a48c5),
	.w8(32'h38899988),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868f333),
	.w1(32'h38755be6),
	.w2(32'h389520f6),
	.w3(32'hb9a3b0bb),
	.w4(32'hb89a3f9d),
	.w5(32'hb913ea0d),
	.w6(32'hb90f75da),
	.w7(32'h38a500ae),
	.w8(32'h395af879),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8982aae),
	.w1(32'hb8526bb5),
	.w2(32'hb76a2ee7),
	.w3(32'hb8c66a54),
	.w4(32'hb8c516fb),
	.w5(32'hb7cf7e22),
	.w6(32'hb8900fe5),
	.w7(32'hb8957a9d),
	.w8(32'hb82fedcf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a282c2c),
	.w1(32'h398af63a),
	.w2(32'h39d6d08f),
	.w3(32'h39a897c1),
	.w4(32'hb8ab48f0),
	.w5(32'h38c537b2),
	.w6(32'h3a18b458),
	.w7(32'h39dd74a6),
	.w8(32'h3a393772),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d6a72),
	.w1(32'hbbd6cad0),
	.w2(32'hbbdc9e4b),
	.w3(32'hb91961b5),
	.w4(32'hbbbacfd3),
	.w5(32'hbc550ff5),
	.w6(32'h3a855617),
	.w7(32'hbc149d84),
	.w8(32'hbb955f77),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43ef0b),
	.w1(32'hbb4b767d),
	.w2(32'hbb46f2b5),
	.w3(32'h3b251557),
	.w4(32'hbb315fbd),
	.w5(32'hbaea5af8),
	.w6(32'h3b5258d1),
	.w7(32'hbc0ae181),
	.w8(32'hbb8f1965),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1616fd),
	.w1(32'hbaf62a30),
	.w2(32'hbaf88002),
	.w3(32'h39e0a35d),
	.w4(32'hba2194e5),
	.w5(32'hba893ee7),
	.w6(32'hb9bb72bb),
	.w7(32'hbb148cd0),
	.w8(32'hbb1e5313),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d6949),
	.w1(32'h3a2fcc47),
	.w2(32'h3b3479c9),
	.w3(32'h395e4468),
	.w4(32'hbac65286),
	.w5(32'h3a73f510),
	.w6(32'hbaffebca),
	.w7(32'hba4a9489),
	.w8(32'h3a8f95f0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b9172),
	.w1(32'h3a618e1c),
	.w2(32'h3aad358b),
	.w3(32'h3a2de720),
	.w4(32'h39cf6910),
	.w5(32'h3a651050),
	.w6(32'h3a3aa35c),
	.w7(32'h39688cf5),
	.w8(32'h3a37bbff),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c8f78),
	.w1(32'h3aef7828),
	.w2(32'h3b7c6b25),
	.w3(32'h3b694f60),
	.w4(32'h3878d148),
	.w5(32'h3b89af38),
	.w6(32'h3b51ae97),
	.w7(32'hb9b27a8d),
	.w8(32'h3b501b57),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f6366),
	.w1(32'h3aecb767),
	.w2(32'h3c08067f),
	.w3(32'hba6d669c),
	.w4(32'h3b11bf23),
	.w5(32'h3bf19b7e),
	.w6(32'h3b31859b),
	.w7(32'h3b1a5c02),
	.w8(32'h3bfdfc14),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d33cc),
	.w1(32'hbbcaf895),
	.w2(32'hbc53d1f9),
	.w3(32'h3ba0ac92),
	.w4(32'hba53e1e7),
	.w5(32'hbb9ffc1f),
	.w6(32'h39e679ce),
	.w7(32'hbc7722cf),
	.w8(32'hbc5a34bf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a973),
	.w1(32'h3b19ae0c),
	.w2(32'h3bebe94b),
	.w3(32'h3a29f8d6),
	.w4(32'h3aa21d9d),
	.w5(32'h3ba850e6),
	.w6(32'h3b250647),
	.w7(32'h3b2e2a46),
	.w8(32'h3ba6d8db),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be83467),
	.w1(32'h39f2ac98),
	.w2(32'h3aa95407),
	.w3(32'h3bac398a),
	.w4(32'h3b2de35d),
	.w5(32'h3b31fd3d),
	.w6(32'h3b31f96b),
	.w7(32'hbaa08120),
	.w8(32'h3a3d1a7e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809be9),
	.w1(32'hbc16c5b5),
	.w2(32'hbc420aba),
	.w3(32'h3ba01ced),
	.w4(32'hbb6a3f0c),
	.w5(32'hbba57b6e),
	.w6(32'h3a82c43b),
	.w7(32'hbc499dba),
	.w8(32'hbc354879),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4f254),
	.w1(32'h3c155636),
	.w2(32'h3c233cdc),
	.w3(32'h3b99f282),
	.w4(32'h3bdb0c7a),
	.w5(32'h3ba7f911),
	.w6(32'h3bc640a6),
	.w7(32'h3bdb16c6),
	.w8(32'h3b840cd7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0b9f6),
	.w1(32'h3aff584c),
	.w2(32'h3a8da812),
	.w3(32'h3b9b2375),
	.w4(32'h3b106e33),
	.w5(32'h3b6d0154),
	.w6(32'h3b5cabec),
	.w7(32'hbafa333f),
	.w8(32'hbb392265),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2074d),
	.w1(32'h3a608f47),
	.w2(32'h3a908fb2),
	.w3(32'h3a9b0bd6),
	.w4(32'h39b06498),
	.w5(32'h39d51287),
	.w6(32'h3aab4198),
	.w7(32'h3983de18),
	.w8(32'h392ce8b8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ddd7),
	.w1(32'hbbb075f0),
	.w2(32'h3b54ae4f),
	.w3(32'hbb7e7761),
	.w4(32'hbc5d2deb),
	.w5(32'hbafec377),
	.w6(32'hba38488e),
	.w7(32'hbbff451f),
	.w8(32'h3b8f8321),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd4af9),
	.w1(32'h39cbe24a),
	.w2(32'hb949e308),
	.w3(32'h391c9aff),
	.w4(32'hbab524d0),
	.w5(32'hb9a53b9f),
	.w6(32'hba287441),
	.w7(32'hbb46e702),
	.w8(32'hbb01edba),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb228b),
	.w1(32'hb9695d24),
	.w2(32'hb9596259),
	.w3(32'hb8d41e17),
	.w4(32'hb9b954f9),
	.w5(32'hb9352f88),
	.w6(32'hb9b1f0dc),
	.w7(32'hb9f642d8),
	.w8(32'hb919b18e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8372c66),
	.w1(32'h37162cde),
	.w2(32'hb90dadad),
	.w3(32'hb885dd80),
	.w4(32'h38958a1f),
	.w5(32'hb7552f47),
	.w6(32'hb89003db),
	.w7(32'h38170107),
	.w8(32'hb8407062),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b482757),
	.w1(32'h3a1e82b8),
	.w2(32'hba409c59),
	.w3(32'h3a802572),
	.w4(32'h3aa962f7),
	.w5(32'h394a4ed8),
	.w6(32'h3ab788c9),
	.w7(32'hba489556),
	.w8(32'hbb0a839e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02cc62),
	.w1(32'h3b58ae5e),
	.w2(32'h3b843fee),
	.w3(32'h3a9b4c28),
	.w4(32'h3af1222a),
	.w5(32'h3b39a4c6),
	.w6(32'h3b43cafe),
	.w7(32'h3b063aa0),
	.w8(32'h385b3b79),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3f65f),
	.w1(32'hba662f9d),
	.w2(32'h3acca517),
	.w3(32'h3b8cb2c4),
	.w4(32'hbac8795e),
	.w5(32'hb9b57cda),
	.w6(32'h3b407da5),
	.w7(32'hbb5adfb4),
	.w8(32'hbb1ff4ec),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3606c82d),
	.w1(32'h3887d7ea),
	.w2(32'h390d43b6),
	.w3(32'h389b1663),
	.w4(32'h3906d303),
	.w5(32'h39031c40),
	.w6(32'h378b2614),
	.w7(32'h37ec6604),
	.w8(32'h3856cef7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b263),
	.w1(32'hb8453481),
	.w2(32'hb89bad8c),
	.w3(32'h3b9a6ee0),
	.w4(32'hba26fc58),
	.w5(32'h3aad0b32),
	.w6(32'h3b215eac),
	.w7(32'hbba13c3c),
	.w8(32'hbb5f3fbe),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d75d),
	.w1(32'h3ad29be2),
	.w2(32'h3b72356f),
	.w3(32'h3b0220bb),
	.w4(32'h3a845304),
	.w5(32'h3b142817),
	.w6(32'h3b3319eb),
	.w7(32'h3a9db466),
	.w8(32'h3ac76441),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb4855),
	.w1(32'hbbdee80c),
	.w2(32'hbbe31b00),
	.w3(32'h3bf1d745),
	.w4(32'hbb13b8c1),
	.w5(32'hbb12c9d2),
	.w6(32'hbad2ac39),
	.w7(32'hbc6a5af6),
	.w8(32'hbc26edac),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32a7c2),
	.w1(32'hbbfe0412),
	.w2(32'hbb2efdf3),
	.w3(32'hbb7788cb),
	.w4(32'hbc7df697),
	.w5(32'hbc5c0df0),
	.w6(32'hbb7355d7),
	.w7(32'hbc8a80d3),
	.w8(32'hbbf676d2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80d5274),
	.w1(32'h3aee0d9f),
	.w2(32'h3b3e05a0),
	.w3(32'hb891c995),
	.w4(32'h3a41618e),
	.w5(32'h3b53f02d),
	.w6(32'h3a9d5761),
	.w7(32'h3a9ba06a),
	.w8(32'h3b716de0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26e7e4),
	.w1(32'h3a22fb90),
	.w2(32'h3a004eb9),
	.w3(32'hb8fd8810),
	.w4(32'h39fe0811),
	.w5(32'h383c720d),
	.w6(32'h3a1d150e),
	.w7(32'h3a3cb7e9),
	.w8(32'h3a705f0f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2c469),
	.w1(32'h3b3e3c0e),
	.w2(32'h3b59dba3),
	.w3(32'h3b454a04),
	.w4(32'h3ad60cd0),
	.w5(32'h3b03a0d1),
	.w6(32'h3b279cec),
	.w7(32'hb9f78aa8),
	.w8(32'h3a31e29c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5effe3),
	.w1(32'h3a81627b),
	.w2(32'h3b1a2318),
	.w3(32'h3a5e5b1b),
	.w4(32'h39006e5a),
	.w5(32'h3b098cbe),
	.w6(32'h3a8cbd11),
	.w7(32'hba25252e),
	.w8(32'h3b55b695),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8291b),
	.w1(32'hb9d6b552),
	.w2(32'h3b5cedb0),
	.w3(32'hbace5d3e),
	.w4(32'hbb0c4c28),
	.w5(32'h3b148c38),
	.w6(32'hba72f569),
	.w7(32'hbad404a4),
	.w8(32'h3b1eba8f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae46a4d),
	.w1(32'hbb17e9fa),
	.w2(32'hbb69dbed),
	.w3(32'h3ad29096),
	.w4(32'hba83328c),
	.w5(32'hbb279611),
	.w6(32'hba5ea3b1),
	.w7(32'hbb8a3bd1),
	.w8(32'hbb989448),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb4114),
	.w1(32'hba0dd8dd),
	.w2(32'h377993fd),
	.w3(32'hb9c2197b),
	.w4(32'hb99901b8),
	.w5(32'hb9157e37),
	.w6(32'hb98f9511),
	.w7(32'hb8fe1be3),
	.w8(32'h38e39f92),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5b45),
	.w1(32'hbb1975e3),
	.w2(32'hbb3944ac),
	.w3(32'h3ae449b3),
	.w4(32'hbb1bf4fb),
	.w5(32'hbabf75bd),
	.w6(32'h3a508c3f),
	.w7(32'hbbc124aa),
	.w8(32'hbb4b4a72),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e9d7),
	.w1(32'hbb4d4876),
	.w2(32'hbba6ab9a),
	.w3(32'h384430ce),
	.w4(32'hbb37e716),
	.w5(32'hbb8c37b9),
	.w6(32'h3aa9b4e8),
	.w7(32'hbb07e427),
	.w8(32'hbb7f875f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd7d3),
	.w1(32'h399e1f8d),
	.w2(32'h3b8784b0),
	.w3(32'hbb1e8d02),
	.w4(32'hbb2b0eb8),
	.w5(32'h39db3d50),
	.w6(32'hbb0421a8),
	.w7(32'hbb8e4ddd),
	.w8(32'h3a18ac54),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989e602),
	.w1(32'hb8a7020e),
	.w2(32'hb8846d05),
	.w3(32'h3a00b305),
	.w4(32'hb8158aa2),
	.w5(32'hb851f143),
	.w6(32'h37269d84),
	.w7(32'hb92df79f),
	.w8(32'hb93335df),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05f651),
	.w1(32'hbb138307),
	.w2(32'hbb3c4afb),
	.w3(32'h3ad135a4),
	.w4(32'hbba425d9),
	.w5(32'hbb6fbc39),
	.w6(32'hba00624a),
	.w7(32'hbb9b80f4),
	.w8(32'hbacd5ceb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3823bf52),
	.w1(32'h38015b39),
	.w2(32'h38aa7cbc),
	.w3(32'h36708540),
	.w4(32'h3866aa73),
	.w5(32'h380cfc49),
	.w6(32'h38944c6a),
	.w7(32'h38f3f92d),
	.w8(32'h38a2bed2),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fff75),
	.w1(32'hb9cfd06e),
	.w2(32'hb939902d),
	.w3(32'hb9980f7b),
	.w4(32'hb97c08b4),
	.w5(32'h398b9729),
	.w6(32'hb9660947),
	.w7(32'hb99fee4a),
	.w8(32'h3945604f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ab68),
	.w1(32'h3a82e7cd),
	.w2(32'h3b9745f8),
	.w3(32'hba292883),
	.w4(32'hba320264),
	.w5(32'h3b8f552a),
	.w6(32'h3a806a5b),
	.w7(32'hb82d0a37),
	.w8(32'h3b82289c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f8fb9),
	.w1(32'h3a066ae5),
	.w2(32'hbb852a0e),
	.w3(32'h3c09458a),
	.w4(32'hbbda59fc),
	.w5(32'hbbac99f7),
	.w6(32'h3bb78085),
	.w7(32'hbc027bb0),
	.w8(32'hbc245843),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ad5e1),
	.w1(32'hbabb97b8),
	.w2(32'hba1a5560),
	.w3(32'hb9ae3795),
	.w4(32'hbb121676),
	.w5(32'hbaae6ac5),
	.w6(32'h397ed57c),
	.w7(32'hbaf3cbc6),
	.w8(32'hba0465cd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a711782),
	.w1(32'hb920fa50),
	.w2(32'h3bc237dc),
	.w3(32'hba33ebda),
	.w4(32'hbb249f0a),
	.w5(32'h3b390fab),
	.w6(32'h3a3875a0),
	.w7(32'hba8192d4),
	.w8(32'h3b82739a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba040f25),
	.w1(32'hba84e555),
	.w2(32'hbb2f3338),
	.w3(32'hbb055aba),
	.w4(32'hbb077c37),
	.w5(32'hbb1253e6),
	.w6(32'hbab8d101),
	.w7(32'hbaccf563),
	.w8(32'hb80d9f1b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8c097),
	.w1(32'hbbb62f57),
	.w2(32'h3b3386e4),
	.w3(32'h3b07e02e),
	.w4(32'hbb7ae0a0),
	.w5(32'h3926e858),
	.w6(32'hbb87a5be),
	.w7(32'hbc62ca30),
	.w8(32'h37ba6d47),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a18fc),
	.w1(32'hba620069),
	.w2(32'h3ad11d96),
	.w3(32'h3b662437),
	.w4(32'hb8e12926),
	.w5(32'h3b5b53ed),
	.w6(32'h3bc95957),
	.w7(32'hbaaf9ec8),
	.w8(32'h3aa21954),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7503e8),
	.w1(32'hbb634ec1),
	.w2(32'hbb286d3d),
	.w3(32'h3b6ea6c1),
	.w4(32'hbaa2a2ab),
	.w5(32'hb959b01d),
	.w6(32'h3af406b0),
	.w7(32'hbbf807f9),
	.w8(32'hbb85d2ce),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966ea39),
	.w1(32'hb95f562e),
	.w2(32'hb9607184),
	.w3(32'h37d6931e),
	.w4(32'hba0f16bb),
	.w5(32'hba0604e0),
	.w6(32'hb991e8c3),
	.w7(32'hba2fb00c),
	.w8(32'hba527fc9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3eac4),
	.w1(32'hbb6dedc1),
	.w2(32'h3985e3cb),
	.w3(32'h3a8bdac1),
	.w4(32'hba9de300),
	.w5(32'h3b16a030),
	.w6(32'h3ae9c672),
	.w7(32'hbb63b5a7),
	.w8(32'h3a69252a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2f980),
	.w1(32'hb7d5309e),
	.w2(32'hb7ce30fd),
	.w3(32'hb8b36939),
	.w4(32'hb41a6b01),
	.w5(32'hb85e5eef),
	.w6(32'hb8667f70),
	.w7(32'hb746cc29),
	.w8(32'hb84da9a0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ea7b7),
	.w1(32'hba460c6e),
	.w2(32'hb9b3b7b3),
	.w3(32'hb8fc5b99),
	.w4(32'hbad1449d),
	.w5(32'hba3b0a82),
	.w6(32'h3a45dfa5),
	.w7(32'hbad3865d),
	.w8(32'hba5de3f7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f4781),
	.w1(32'h392ec323),
	.w2(32'h3a8c9eab),
	.w3(32'hb8dc9b36),
	.w4(32'h39c2857b),
	.w5(32'h3a064df9),
	.w6(32'hba0c99e1),
	.w7(32'hb91631b7),
	.w8(32'h3affeb25),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8448ba),
	.w1(32'hba528a2c),
	.w2(32'h3bf673ee),
	.w3(32'h3b6a263b),
	.w4(32'h3b772bed),
	.w5(32'h3c15658a),
	.w6(32'h3b231c6c),
	.w7(32'hb9bf5b4f),
	.w8(32'h3bd09935),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a4381),
	.w1(32'h3863fb6c),
	.w2(32'h38325a0e),
	.w3(32'hb75c4f3a),
	.w4(32'h38be28ab),
	.w5(32'h3802498a),
	.w6(32'hb7e088f6),
	.w7(32'h383b5f69),
	.w8(32'h37f5ba97),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3802187a),
	.w1(32'h3817f2a5),
	.w2(32'h38cf403f),
	.w3(32'h36f99744),
	.w4(32'h38cef954),
	.w5(32'h395c898f),
	.w6(32'h37784cec),
	.w7(32'h39034116),
	.w8(32'h39627fe5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5c815),
	.w1(32'h3aa228d6),
	.w2(32'h3b48a2c3),
	.w3(32'h38978246),
	.w4(32'h39b6ec8e),
	.w5(32'h3ace976b),
	.w6(32'hba2ca674),
	.w7(32'hbb4f9eda),
	.w8(32'hb90e5a84),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb0618),
	.w1(32'hbc03e7c5),
	.w2(32'hbbb4fe0c),
	.w3(32'h39e606c5),
	.w4(32'hba078ba7),
	.w5(32'hbbbfc151),
	.w6(32'h3b9940bf),
	.w7(32'hbbc50c10),
	.w8(32'hbc2d270b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac8787),
	.w1(32'h3b109560),
	.w2(32'hbb8f102e),
	.w3(32'hbb26d4b8),
	.w4(32'hbad33a37),
	.w5(32'hbba8a7b3),
	.w6(32'hbb84573e),
	.w7(32'hbb2862ba),
	.w8(32'hbc78b205),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2c6ce),
	.w1(32'hb95ed036),
	.w2(32'h384a070b),
	.w3(32'h396acd73),
	.w4(32'h39a7613a),
	.w5(32'h39d86eb2),
	.w6(32'h39c7e22a),
	.w7(32'h393bae1e),
	.w8(32'h3a272f2c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24a314),
	.w1(32'hbbd57f6e),
	.w2(32'hbb14c5c5),
	.w3(32'h3bc8c7a0),
	.w4(32'hbb4e6b8b),
	.w5(32'hbb4c2318),
	.w6(32'h3b386acd),
	.w7(32'hbc5f7455),
	.w8(32'hbba62abf),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d2cd),
	.w1(32'hba953e8f),
	.w2(32'h3bb4d44b),
	.w3(32'h3b819020),
	.w4(32'hbaa54245),
	.w5(32'h3bc5854b),
	.w6(32'h3ba09944),
	.w7(32'hbbd87e0e),
	.w8(32'h3bd6fa0d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b364c33),
	.w1(32'hba7c3ddc),
	.w2(32'hbc06233e),
	.w3(32'hb937dfb8),
	.w4(32'hbb41d955),
	.w5(32'hbb8588c5),
	.w6(32'h39cbd592),
	.w7(32'hbb97b469),
	.w8(32'hbbdd70e4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89547dc),
	.w1(32'hb75661b0),
	.w2(32'hb80d03c8),
	.w3(32'hb8cd8ce2),
	.w4(32'hb7c3cdda),
	.w5(32'hb826bd27),
	.w6(32'hb8adc207),
	.w7(32'h387d072e),
	.w8(32'h382ae6a6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5915a),
	.w1(32'h38cd14fb),
	.w2(32'h3982aa89),
	.w3(32'hb8daac3a),
	.w4(32'hb8735161),
	.w5(32'h39a024fe),
	.w6(32'hb9367fc9),
	.w7(32'h38f4ca8e),
	.w8(32'h3a04f19b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923ef8a),
	.w1(32'hb811f486),
	.w2(32'hb7db3759),
	.w3(32'hb8c5cd57),
	.w4(32'hb816eb90),
	.w5(32'hb84a07f2),
	.w6(32'hb883814a),
	.w7(32'hb8025fe6),
	.w8(32'hb806afab),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b8ba),
	.w1(32'hbb80d722),
	.w2(32'hbc2cf16d),
	.w3(32'hba8d1448),
	.w4(32'hbb96c92c),
	.w5(32'hbbbdabc5),
	.w6(32'h3801b762),
	.w7(32'hbbeb79b6),
	.w8(32'hbc1abfef),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdd0c5),
	.w1(32'h3a6bd550),
	.w2(32'hb910e3b3),
	.w3(32'h3b6e68d2),
	.w4(32'hbb147f61),
	.w5(32'hbb65c14a),
	.w6(32'h3b581b2d),
	.w7(32'hbac27a7e),
	.w8(32'hbaf29433),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f65f),
	.w1(32'h3be51f90),
	.w2(32'h3c5d8fc5),
	.w3(32'h3b619601),
	.w4(32'h3b42dce7),
	.w5(32'h3c087f51),
	.w6(32'h3b86a275),
	.w7(32'h3b8c16cc),
	.w8(32'h3bc2e700),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a037f11),
	.w1(32'hb90a9f5c),
	.w2(32'h3a3e87ff),
	.w3(32'h3a2a84fb),
	.w4(32'hb9bf5e0f),
	.w5(32'hb99ae829),
	.w6(32'h3a23699a),
	.w7(32'hb9e4b2f4),
	.w8(32'h3a37a397),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd9e9b),
	.w1(32'hbae5ba73),
	.w2(32'hbb66a17b),
	.w3(32'h3b9136fd),
	.w4(32'hbb0a1038),
	.w5(32'hbb12c98c),
	.w6(32'h3acf619d),
	.w7(32'hbbe6c5e2),
	.w8(32'hbbc90e78),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51af89),
	.w1(32'h3b7772d2),
	.w2(32'hb9c4f9b0),
	.w3(32'h3a81195d),
	.w4(32'h3b2f8214),
	.w5(32'hbb223b02),
	.w6(32'h3aa33f3d),
	.w7(32'h3ae0ac6c),
	.w8(32'hbbb7a5ef),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db85ec),
	.w1(32'h38023abe),
	.w2(32'h374f311a),
	.w3(32'hb87236ac),
	.w4(32'h3884c204),
	.w5(32'hb7c4000c),
	.w6(32'hb89c1c8f),
	.w7(32'h376a962c),
	.w8(32'hb8863739),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1cf86),
	.w1(32'h3afb1516),
	.w2(32'h3ba322dc),
	.w3(32'hbb4c3fc8),
	.w4(32'h3b2267a5),
	.w5(32'h3bbd178c),
	.w6(32'hba0ab790),
	.w7(32'h3b1818e6),
	.w8(32'h3b0d6730),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978e0a0),
	.w1(32'h38643f3c),
	.w2(32'hb8228363),
	.w3(32'hb95a52b8),
	.w4(32'h38d7cd3a),
	.w5(32'hb800f11b),
	.w6(32'hb982976d),
	.w7(32'hb3f05ef0),
	.w8(32'hb859f065),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e76a),
	.w1(32'hba905e8b),
	.w2(32'hba7e992f),
	.w3(32'h3b2237a7),
	.w4(32'hbacd0eae),
	.w5(32'hbb163716),
	.w6(32'h3aff62e3),
	.w7(32'hbb771d7f),
	.w8(32'hbb4f3f38),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f358),
	.w1(32'h3b1d9a72),
	.w2(32'h3bde6438),
	.w3(32'h3b65b82f),
	.w4(32'h3a94c6be),
	.w5(32'h3b861342),
	.w6(32'h3b575458),
	.w7(32'hbaaf3b16),
	.w8(32'h3b56f441),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840dbd),
	.w1(32'h3b207d9a),
	.w2(32'h3b747d54),
	.w3(32'h3b0e37c7),
	.w4(32'h3a7beeb0),
	.w5(32'h3ac7f774),
	.w6(32'h3b166bf3),
	.w7(32'h38d3c83c),
	.w8(32'h3a196887),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fb98e),
	.w1(32'hb93fa618),
	.w2(32'hba698de8),
	.w3(32'h39f70500),
	.w4(32'hb9ad6fb2),
	.w5(32'hba417cb3),
	.w6(32'h3a0e766c),
	.w7(32'hb95affd8),
	.w8(32'h38567401),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34d214),
	.w1(32'h3b97edca),
	.w2(32'h3c380272),
	.w3(32'h3ae0f319),
	.w4(32'h3b309542),
	.w5(32'h3c1a4fe7),
	.w6(32'h3b6346f7),
	.w7(32'h3b6cf686),
	.w8(32'h3c055031),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e244),
	.w1(32'h3adf57e1),
	.w2(32'h3b2e7364),
	.w3(32'h3b6d5364),
	.w4(32'h3b1e7bbf),
	.w5(32'h3ba6bbe8),
	.w6(32'h3b75f4e1),
	.w7(32'hba8e32d9),
	.w8(32'h39303b7a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0182f),
	.w1(32'hbaa8b316),
	.w2(32'h38ca0cfb),
	.w3(32'h3ba75b0d),
	.w4(32'hbb005b7f),
	.w5(32'hba4c9958),
	.w6(32'h3b6fc2e4),
	.w7(32'hbb366b14),
	.w8(32'hbadfe2ad),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d19c9),
	.w1(32'hb98b37ad),
	.w2(32'hb9dbf05f),
	.w3(32'hb98fd55d),
	.w4(32'hb9dc75ff),
	.w5(32'hb9d3fa23),
	.w6(32'hba02c764),
	.w7(32'hba0d2734),
	.w8(32'hb99c1f9f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14fd70),
	.w1(32'hb974f6c8),
	.w2(32'hb8d8c0d3),
	.w3(32'hb9726790),
	.w4(32'hb95ea7a2),
	.w5(32'h395b8ca4),
	.w6(32'hb9d3dfff),
	.w7(32'h3705f4bd),
	.w8(32'h396695d6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a4b57),
	.w1(32'h38ef866e),
	.w2(32'hbb070d1d),
	.w3(32'h3c181ed4),
	.w4(32'hbbfc0a6f),
	.w5(32'hbc430732),
	.w6(32'h3b999975),
	.w7(32'hbb835b31),
	.w8(32'hbc1425b5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03f375),
	.w1(32'hbac01dc4),
	.w2(32'h3afbd08e),
	.w3(32'h3b79577e),
	.w4(32'hbbd3c615),
	.w5(32'hbb6f3430),
	.w6(32'h3b1f9a35),
	.w7(32'hbc152889),
	.w8(32'hbbb06331),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1683),
	.w1(32'h3bc29500),
	.w2(32'h3c245c59),
	.w3(32'h3baceb5c),
	.w4(32'h3b85c3fc),
	.w5(32'h3bcca744),
	.w6(32'h3bb30f5d),
	.w7(32'h3aa62f5e),
	.w8(32'h3ac65278),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4517f),
	.w1(32'hba2db01c),
	.w2(32'hbc732a09),
	.w3(32'h3b5219e4),
	.w4(32'h3a82330a),
	.w5(32'hbb788768),
	.w6(32'h3bc46791),
	.w7(32'hbc44d0ea),
	.w8(32'hbc4f7b89),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c026f),
	.w1(32'hbb0de111),
	.w2(32'h3990d8dc),
	.w3(32'hba8194c7),
	.w4(32'hba94d37d),
	.w5(32'hba4caefb),
	.w6(32'hbadcaf03),
	.w7(32'hbad88f9c),
	.w8(32'hba246107),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89223a),
	.w1(32'hb978802c),
	.w2(32'h3aa20cfa),
	.w3(32'hb9ecae42),
	.w4(32'hba75e6d8),
	.w5(32'h3a9aa8eb),
	.w6(32'h3a1791c8),
	.w7(32'hb988a4ad),
	.w8(32'h3b1b4033),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ef00),
	.w1(32'hbb475b54),
	.w2(32'hbcc43f95),
	.w3(32'hba782667),
	.w4(32'hbc262254),
	.w5(32'hbca17483),
	.w6(32'h387c3302),
	.w7(32'hbbd35074),
	.w8(32'hbcddb0b7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fb93f),
	.w1(32'hbbdb5a8c),
	.w2(32'hbbcbf96f),
	.w3(32'h3bcae873),
	.w4(32'hbb20859c),
	.w5(32'hbb892369),
	.w6(32'h3931ce9b),
	.w7(32'hbc474538),
	.w8(32'hbbd25134),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4220aa),
	.w1(32'hbbae806c),
	.w2(32'hbb8fbe7a),
	.w3(32'h3be32bbb),
	.w4(32'hbb026d55),
	.w5(32'hbb197f92),
	.w6(32'h3b587240),
	.w7(32'hbc0b7295),
	.w8(32'hbc6527b8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3ad5b),
	.w1(32'hbaac5c8b),
	.w2(32'h3b6388c8),
	.w3(32'hbb10236f),
	.w4(32'hbbb2df83),
	.w5(32'h3886adb2),
	.w6(32'hbb1d1b46),
	.w7(32'hbb873dd5),
	.w8(32'hb89c2187),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a3f75),
	.w1(32'hba80b91f),
	.w2(32'h3bfc0c7e),
	.w3(32'hbac2d7a5),
	.w4(32'hbb3197e3),
	.w5(32'h3bb9bf31),
	.w6(32'h37605372),
	.w7(32'hbb011cb1),
	.w8(32'h3bb7450d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892245e),
	.w1(32'hb787bf1c),
	.w2(32'hb7cd8fb1),
	.w3(32'hb834a49a),
	.w4(32'h36514550),
	.w5(32'hb83fd795),
	.w6(32'hb87b392d),
	.w7(32'hb7e5182c),
	.w8(32'hb837bbc5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892871b),
	.w1(32'hb7a76f51),
	.w2(32'hb8142aaf),
	.w3(32'hb8524d1d),
	.w4(32'hb78bd01c),
	.w5(32'hb843da43),
	.w6(32'hb8a86bca),
	.w7(32'hb7a6aba5),
	.w8(32'hb8412765),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53df1a),
	.w1(32'hbad78997),
	.w2(32'hbab21920),
	.w3(32'hb9643540),
	.w4(32'hbb0cd75f),
	.w5(32'hbb657745),
	.w6(32'h3a34d66d),
	.w7(32'hbaf332cb),
	.w8(32'hbaa0fe03),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d34d73),
	.w1(32'hb773447e),
	.w2(32'hb7b4f92d),
	.w3(32'hb8d7a4f6),
	.w4(32'hb77515c5),
	.w5(32'hb9b527ed),
	.w6(32'hb8bb2add),
	.w7(32'hb75e2dcf),
	.w8(32'h375677c3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fb9bd),
	.w1(32'hbbbba3d8),
	.w2(32'hbbf092cc),
	.w3(32'hbb2a34ba),
	.w4(32'hbbed3b1d),
	.w5(32'hbbc90502),
	.w6(32'h3992705a),
	.w7(32'hbb8df2ea),
	.w8(32'hbbc9b75d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bba8d),
	.w1(32'hbb28cc9c),
	.w2(32'h3bea6e76),
	.w3(32'h3aa6ed19),
	.w4(32'hbb263d1b),
	.w5(32'h3a25c9ec),
	.w6(32'h3a1d6d60),
	.w7(32'hbb994888),
	.w8(32'h3ae7cbb3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd2be6),
	.w1(32'h3b00433a),
	.w2(32'h3ae40385),
	.w3(32'h3b3d2a5b),
	.w4(32'h395b0573),
	.w5(32'h3ac211bd),
	.w6(32'h3acb081b),
	.w7(32'hb995fdb1),
	.w8(32'h3a92a7fb),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23ccb0),
	.w1(32'h39dfebe7),
	.w2(32'h3a8b9332),
	.w3(32'h39de6275),
	.w4(32'hb9a9d48a),
	.w5(32'h3a0bf977),
	.w6(32'h357d2ebd),
	.w7(32'hb8ba3beb),
	.w8(32'h39a80f85),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b6a36),
	.w1(32'hbc22237b),
	.w2(32'hbc10e98b),
	.w3(32'h3bd9b24a),
	.w4(32'hbba49f78),
	.w5(32'hbbfec1bf),
	.w6(32'h3b0513d9),
	.w7(32'hbc83ac17),
	.w8(32'hbcb174a9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e46f08),
	.w1(32'hbb32d15a),
	.w2(32'hbb98f980),
	.w3(32'h3b2d7396),
	.w4(32'hba8b76df),
	.w5(32'h3a0a2d35),
	.w6(32'hb9ceab2b),
	.w7(32'hbbbec3f4),
	.w8(32'hbb32db1e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa65d6a),
	.w1(32'hba60a677),
	.w2(32'h38f5e53a),
	.w3(32'h3a6d62b5),
	.w4(32'h3845a1be),
	.w5(32'hba4a35d5),
	.w6(32'hb9e0e675),
	.w7(32'h36af0f3b),
	.w8(32'hba2bebe5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cbfc5),
	.w1(32'hbbc2fbb3),
	.w2(32'hbc2001e4),
	.w3(32'h3b1efc51),
	.w4(32'hbb90c279),
	.w5(32'hbb82c955),
	.w6(32'h39b4a889),
	.w7(32'hbc0e7a4a),
	.w8(32'hbbbc086c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e4725),
	.w1(32'hb9abaf51),
	.w2(32'hb9f140af),
	.w3(32'hba0bc409),
	.w4(32'hba9c94b0),
	.w5(32'hba5ffdd2),
	.w6(32'h39bac648),
	.w7(32'hba5a465b),
	.w8(32'hba85a827),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39deb867),
	.w1(32'hb9df95bf),
	.w2(32'hb9a9cffa),
	.w3(32'hba867945),
	.w4(32'hba2e5398),
	.w5(32'hb99f023e),
	.w6(32'hba80bf60),
	.w7(32'hba191883),
	.w8(32'h3829078d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a509608),
	.w1(32'h3a42847e),
	.w2(32'h3ab7c19f),
	.w3(32'h3a4acb48),
	.w4(32'h3a9d439b),
	.w5(32'hba6f8bb6),
	.w6(32'h3a2ac6ff),
	.w7(32'h3a8d5137),
	.w8(32'hba6a8b10),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d37f2),
	.w1(32'hbad1b3a2),
	.w2(32'hb927a9bb),
	.w3(32'hba9f0075),
	.w4(32'hb96ac0a9),
	.w5(32'hba8b7f74),
	.w6(32'hbadcc15e),
	.w7(32'hba09ef1d),
	.w8(32'hb9dbdcf0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94b97),
	.w1(32'hbb57a028),
	.w2(32'hbafc25e5),
	.w3(32'hbb436c89),
	.w4(32'hbb9859ca),
	.w5(32'hbaa52a1e),
	.w6(32'hbafb8d69),
	.w7(32'hbb69bf44),
	.w8(32'hbb035959),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e6a40),
	.w1(32'hbc02a675),
	.w2(32'hbb5896f0),
	.w3(32'h3b0b6520),
	.w4(32'hbaf024ff),
	.w5(32'hba89e220),
	.w6(32'h3b30ef0f),
	.w7(32'hbc46cc80),
	.w8(32'hbbe09787),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f906c),
	.w1(32'hbb58dfe1),
	.w2(32'hbb97ab33),
	.w3(32'h3b7adf8e),
	.w4(32'hbade3201),
	.w5(32'h3925a22a),
	.w6(32'h3b5423a6),
	.w7(32'hbbea0add),
	.w8(32'hbb751855),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d50f0),
	.w1(32'hbbd8cac6),
	.w2(32'hbbca9edb),
	.w3(32'h3adc71f8),
	.w4(32'hbb9b8d41),
	.w5(32'hbbc2922d),
	.w6(32'hbb193ee5),
	.w7(32'hbc2d414a),
	.w8(32'hbc14c993),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97593f),
	.w1(32'hba221fc5),
	.w2(32'hba086bf3),
	.w3(32'hb9febbf7),
	.w4(32'hb994887f),
	.w5(32'h3a2f6d03),
	.w6(32'hba57d84d),
	.w7(32'hb9b83c29),
	.w8(32'h393a4b26),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976f725),
	.w1(32'h382daa5e),
	.w2(32'h3a3c4387),
	.w3(32'h39d35eff),
	.w4(32'h3a18c00b),
	.w5(32'h3a823379),
	.w6(32'h3a100ce9),
	.w7(32'h3989086a),
	.w8(32'h3a6891ee),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfad47),
	.w1(32'h3a5aa078),
	.w2(32'hb7b26969),
	.w3(32'h3a3da18e),
	.w4(32'h3985ba28),
	.w5(32'hb9d2aad7),
	.w6(32'h3a4cbd3a),
	.w7(32'hb939a33f),
	.w8(32'hb9e9b350),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbc97e),
	.w1(32'h3843b54f),
	.w2(32'h3abbd727),
	.w3(32'h39f0a773),
	.w4(32'h3a570985),
	.w5(32'h39e18d4b),
	.w6(32'hb81098ae),
	.w7(32'h3a5b5bc0),
	.w8(32'h3a9f4fc4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa76e6e),
	.w1(32'hb99eb468),
	.w2(32'h3c05cc78),
	.w3(32'h3b542117),
	.w4(32'h3b07308f),
	.w5(32'h3be3e059),
	.w6(32'h3b1e0cd5),
	.w7(32'hbac7adb5),
	.w8(32'h3b6fbd64),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa94263),
	.w1(32'hbab0e7f6),
	.w2(32'hba6dd96b),
	.w3(32'hbacb1f6d),
	.w4(32'hba35e100),
	.w5(32'hb9f7def9),
	.w6(32'hbb209b03),
	.w7(32'hba8939c1),
	.w8(32'hba88e963),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c793d),
	.w1(32'hb77e1924),
	.w2(32'hb91b15c4),
	.w3(32'hb6b8e62f),
	.w4(32'hba1e489d),
	.w5(32'hbaa193c2),
	.w6(32'h38f3379a),
	.w7(32'hba089dc7),
	.w8(32'hba403720),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad30886),
	.w1(32'h3a53bbca),
	.w2(32'h3b661a96),
	.w3(32'hbab6d4b1),
	.w4(32'h3b04cf3c),
	.w5(32'h3b509522),
	.w6(32'hba8668ac),
	.w7(32'h3adb6c6a),
	.w8(32'h3aae94ff),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a022a3a),
	.w1(32'hb9d029d4),
	.w2(32'hb94b7ca7),
	.w3(32'h3aa10df2),
	.w4(32'h39d31844),
	.w5(32'hba2a5376),
	.w6(32'h38387ba5),
	.w7(32'h38f53b38),
	.w8(32'hb9c62526),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89534f),
	.w1(32'hbaceddcf),
	.w2(32'hbaf49a92),
	.w3(32'h39979b97),
	.w4(32'hbaed1394),
	.w5(32'hba36e660),
	.w6(32'hbaa43df1),
	.w7(32'hbb30c3d6),
	.w8(32'hbabbc996),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba795750),
	.w1(32'hba254a60),
	.w2(32'h3a0a3559),
	.w3(32'h381d6833),
	.w4(32'h38f91f24),
	.w5(32'h3a35c1fb),
	.w6(32'hb887bf9a),
	.w7(32'h39b2d1d7),
	.w8(32'hb95841b8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef230),
	.w1(32'hbbbef829),
	.w2(32'h3c2d4598),
	.w3(32'h3910132c),
	.w4(32'h3b49e337),
	.w5(32'h3c6341a5),
	.w6(32'hb9f546a1),
	.w7(32'hbbe5cdd0),
	.w8(32'h3c3ef70c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820395),
	.w1(32'hba65ef43),
	.w2(32'hba2787d9),
	.w3(32'hba2746db),
	.w4(32'hba25c58f),
	.w5(32'h3a3eab0f),
	.w6(32'hba1950c9),
	.w7(32'hba139bc4),
	.w8(32'h39e47100),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7c7a),
	.w1(32'h3b717128),
	.w2(32'h3af677c5),
	.w3(32'h3bb36037),
	.w4(32'hb93eb0a2),
	.w5(32'h3a5ddd2d),
	.w6(32'h3b94bd54),
	.w7(32'h3998f890),
	.w8(32'hbb236d00),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule