module layer_10_featuremap_311(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36230fde),
	.w1(32'h36d60348),
	.w2(32'h364f1f86),
	.w3(32'hb690e78d),
	.w4(32'h35a9ee5e),
	.w5(32'hb613742e),
	.w6(32'hb7047330),
	.w7(32'hb5ae12c7),
	.w8(32'hb680e4fb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3651badb),
	.w1(32'hb80228b8),
	.w2(32'hb90b2054),
	.w3(32'h3a1b808d),
	.w4(32'hb8c11a08),
	.w5(32'hb9558aa4),
	.w6(32'h3a7ff7e9),
	.w7(32'h39d7dc85),
	.w8(32'h3a2d7659),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb691c7e3),
	.w1(32'hb67ccfb6),
	.w2(32'hb6ac839f),
	.w3(32'hb683be30),
	.w4(32'hb53f7047),
	.w5(32'hb6113d90),
	.w6(32'h37151bab),
	.w7(32'h36a749df),
	.w8(32'hb5608da7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84c8c8),
	.w1(32'hba934a63),
	.w2(32'hba6c246c),
	.w3(32'hb909e4d3),
	.w4(32'hb960d3f5),
	.w5(32'h38b9aba1),
	.w6(32'hb90f51c3),
	.w7(32'hb814b149),
	.w8(32'h3957521d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38085cf2),
	.w1(32'h38312d6f),
	.w2(32'h384b71b4),
	.w3(32'h380637f7),
	.w4(32'h382a94fc),
	.w5(32'h3819125b),
	.w6(32'hb7789ae5),
	.w7(32'hb786676e),
	.w8(32'h36e16e80),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a84792),
	.w1(32'h33f3dd80),
	.w2(32'h3626a6e5),
	.w3(32'h35a444c2),
	.w4(32'h33b83982),
	.w5(32'h366b11b3),
	.w6(32'h366c5b2e),
	.w7(32'h3640b1e0),
	.w8(32'h36e19824),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae04da8),
	.w1(32'h3ae3c361),
	.w2(32'h3aa626fb),
	.w3(32'hba90b69c),
	.w4(32'h3af208bf),
	.w5(32'h3af4ace9),
	.w6(32'hbb0eac3c),
	.w7(32'h3a2842a7),
	.w8(32'h3ac8ddd1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b575901),
	.w1(32'h3b76a98f),
	.w2(32'h39d51056),
	.w3(32'h3b747480),
	.w4(32'h3b7f7c61),
	.w5(32'h3b02df3b),
	.w6(32'hb97c8072),
	.w7(32'hbafa693c),
	.w8(32'hba8615ed),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7d6e6),
	.w1(32'h353a8aeb),
	.w2(32'h393a36fc),
	.w3(32'hb9d68c4a),
	.w4(32'hb83096a8),
	.w5(32'h392361e3),
	.w6(32'hb9cd0800),
	.w7(32'hb91026f9),
	.w8(32'h38b6caa6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f743da),
	.w1(32'h39e9319a),
	.w2(32'h3a19f45a),
	.w3(32'h3ac4a380),
	.w4(32'h3b0fa934),
	.w5(32'h3ac1fd10),
	.w6(32'h3a6ef9b5),
	.w7(32'h3afc3a6f),
	.w8(32'h3b2c5076),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c8e88),
	.w1(32'h39352532),
	.w2(32'h390de162),
	.w3(32'hb89ea321),
	.w4(32'h393a9323),
	.w5(32'h39411796),
	.w6(32'h381698fe),
	.w7(32'h39395a6c),
	.w8(32'h395f14ce),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2edee4),
	.w1(32'h3a565bda),
	.w2(32'h3aeda5d2),
	.w3(32'hbb43c74e),
	.w4(32'h3a145032),
	.w5(32'h3b37d10d),
	.w6(32'hbb85a4bd),
	.w7(32'hba48b264),
	.w8(32'h3ab80c46),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbc2d0),
	.w1(32'h3a8fdb00),
	.w2(32'h3a054f5f),
	.w3(32'h3a8f3ea6),
	.w4(32'h3b10302d),
	.w5(32'h3ab8479a),
	.w6(32'hba30776e),
	.w7(32'h3ad860a3),
	.w8(32'h3ae11b08),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85f846),
	.w1(32'h3aab60b8),
	.w2(32'h3a3eab48),
	.w3(32'h398414e0),
	.w4(32'h3a3ca4fa),
	.w5(32'h3a26e932),
	.w6(32'hb988b521),
	.w7(32'h3a4d39c3),
	.w8(32'h39dd6f36),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f6a6c),
	.w1(32'hbaa18392),
	.w2(32'hba82222d),
	.w3(32'h3a8ade21),
	.w4(32'h38ab3aed),
	.w5(32'h396709fc),
	.w6(32'h3af8231f),
	.w7(32'h3a35afe9),
	.w8(32'h3a9685cd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d1f01),
	.w1(32'h3a8c715e),
	.w2(32'h3ae1c0ad),
	.w3(32'h3b096b97),
	.w4(32'h3adf3a3e),
	.w5(32'h3a4ee63f),
	.w6(32'h3b08c8d3),
	.w7(32'h3b34f93e),
	.w8(32'h3a880058),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8881efc),
	.w1(32'h37cbecf2),
	.w2(32'h38977dcb),
	.w3(32'hb85d6c35),
	.w4(32'h38a45794),
	.w5(32'h38e633fe),
	.w6(32'h38a76b4f),
	.w7(32'h39231e86),
	.w8(32'h39360756),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb9782),
	.w1(32'h3ab9a734),
	.w2(32'h3b081548),
	.w3(32'h39f48275),
	.w4(32'h3b3e2535),
	.w5(32'h3b5d6089),
	.w6(32'hbb02fc4d),
	.w7(32'hbab9108f),
	.w8(32'hb90335cd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e9a23),
	.w1(32'h3a60269d),
	.w2(32'h3a2b1315),
	.w3(32'h3992db10),
	.w4(32'h3acc6649),
	.w5(32'h3ab47665),
	.w6(32'hba66f4c9),
	.w7(32'hb95f17e2),
	.w8(32'h3a3b5441),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c6e509),
	.w1(32'hb8a3005c),
	.w2(32'hb82cb1e8),
	.w3(32'hb75a736e),
	.w4(32'hb8953146),
	.w5(32'hb7b441e6),
	.w6(32'h37b60c61),
	.w7(32'hb8159500),
	.w8(32'h3731cffe),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b3e92),
	.w1(32'hb7cf97d8),
	.w2(32'hb550fec3),
	.w3(32'hb77f26bf),
	.w4(32'h3570a7d9),
	.w5(32'hb73fb324),
	.w6(32'hb84c91f4),
	.w7(32'hb84356e1),
	.w8(32'hb802aa72),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2f931),
	.w1(32'hba96efae),
	.w2(32'hba137a17),
	.w3(32'hba42eb47),
	.w4(32'hba6cee0d),
	.w5(32'hb92f51a2),
	.w6(32'hb9c82712),
	.w7(32'hba1855a3),
	.w8(32'hb75e98eb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8579e2c),
	.w1(32'hb9b0b0b2),
	.w2(32'h3b6bdceb),
	.w3(32'h39a760aa),
	.w4(32'h3af218ec),
	.w5(32'h3b91ef56),
	.w6(32'hbb46210a),
	.w7(32'hb81b19c3),
	.w8(32'h39024bbf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba211714),
	.w1(32'hb9f038cf),
	.w2(32'hb9ef72b8),
	.w3(32'h3a27ee11),
	.w4(32'h3a330224),
	.w5(32'h399be3b8),
	.w6(32'h3a06fb9a),
	.w7(32'h3a4b8397),
	.w8(32'h3aa9762e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18deca),
	.w1(32'hbb3c6995),
	.w2(32'hbb445409),
	.w3(32'h3a007e94),
	.w4(32'hba95b2e0),
	.w5(32'hbaf0b50c),
	.w6(32'h3ad6e947),
	.w7(32'hb96e6bf6),
	.w8(32'hb945b025),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a89c35),
	.w1(32'hb7422488),
	.w2(32'h3902b6fb),
	.w3(32'h387ca85d),
	.w4(32'h3990ac99),
	.w5(32'h39c151e3),
	.w6(32'h39a18e73),
	.w7(32'h3a126524),
	.w8(32'h3a14afc4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378841c0),
	.w1(32'hb64523de),
	.w2(32'hb7bab603),
	.w3(32'h370ce342),
	.w4(32'hb7861918),
	.w5(32'hb7eb1a42),
	.w6(32'h379b57b5),
	.w7(32'hb794aac3),
	.w8(32'hb8214bdf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3a112),
	.w1(32'hba391df8),
	.w2(32'hb978980a),
	.w3(32'h3a227dcb),
	.w4(32'h3abfb52e),
	.w5(32'hb8331a44),
	.w6(32'h3addd0d4),
	.w7(32'h3b34d436),
	.w8(32'h3aa11f35),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba438d27),
	.w1(32'hb9c0c810),
	.w2(32'hb9821f8b),
	.w3(32'hbaa4cec2),
	.w4(32'hba2ba41f),
	.w5(32'hb915aedc),
	.w6(32'hbaa7540b),
	.w7(32'hba71f186),
	.w8(32'hb9e53056),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cd07b),
	.w1(32'hbb6b7a99),
	.w2(32'hbb90e976),
	.w3(32'hb7c37a8d),
	.w4(32'h3a86cc89),
	.w5(32'hba16bd0e),
	.w6(32'h3b0f0734),
	.w7(32'h3b638350),
	.w8(32'h3b1e1b0d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3776d0a2),
	.w1(32'h3723b007),
	.w2(32'h35fa75eb),
	.w3(32'h37a5b576),
	.w4(32'h3742279f),
	.w5(32'hb6c21b03),
	.w6(32'h3611ddd6),
	.w7(32'h35d45626),
	.w8(32'h372e002b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b83bc5),
	.w1(32'hb6548f98),
	.w2(32'hb7576116),
	.w3(32'hb38f602e),
	.w4(32'h35d5a6d6),
	.w5(32'hb68aa63a),
	.w6(32'h379dbfb6),
	.w7(32'h3795c3eb),
	.w8(32'hb6edc235),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9469bee),
	.w1(32'h398d1eef),
	.w2(32'h39cbc07e),
	.w3(32'h3967f4b7),
	.w4(32'h3a744b88),
	.w5(32'h3a87d786),
	.w6(32'hb9993d0c),
	.w7(32'h398558a8),
	.w8(32'h3a293a49),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3a059),
	.w1(32'hb7fc2c96),
	.w2(32'hb7b1c44e),
	.w3(32'h39850837),
	.w4(32'h38deb70a),
	.w5(32'h38e027cf),
	.w6(32'h39d9a2cb),
	.w7(32'h3987849f),
	.w8(32'h39d6137d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9930945),
	.w1(32'hb8df3e0e),
	.w2(32'hb92bd769),
	.w3(32'hb9bb4e4e),
	.w4(32'h38d450c4),
	.w5(32'h37d536f7),
	.w6(32'hb9aaafbb),
	.w7(32'hb9934903),
	.w8(32'hb60e2a6e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cc92b),
	.w1(32'h3a6e4351),
	.w2(32'h3a9fc6e2),
	.w3(32'hb983faa8),
	.w4(32'h3a7cdb92),
	.w5(32'h3ac938ac),
	.w6(32'hbaec9e09),
	.w7(32'hba44df8c),
	.w8(32'h396b4bb9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88f520),
	.w1(32'hb8e4e0be),
	.w2(32'h3b7293a2),
	.w3(32'h3b548477),
	.w4(32'h3b1e44ec),
	.w5(32'h3bb0c186),
	.w6(32'h3aa3e1d2),
	.w7(32'hb916c491),
	.w8(32'h3b810f94),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38f484),
	.w1(32'hbb9a37ee),
	.w2(32'hbb6a0df6),
	.w3(32'hbaa41cf5),
	.w4(32'hbb8b7e55),
	.w5(32'hbb1b3a8c),
	.w6(32'h3a3b09d8),
	.w7(32'hbb3016e3),
	.w8(32'h395162db),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320420),
	.w1(32'hbb0d403c),
	.w2(32'hbb3ad70e),
	.w3(32'hba0d20d4),
	.w4(32'hb700a769),
	.w5(32'hba06d0df),
	.w6(32'h3a85a6f7),
	.w7(32'hb8335b03),
	.w8(32'h38982515),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f36c8),
	.w1(32'hba569fa8),
	.w2(32'hba37765c),
	.w3(32'h39f8fb18),
	.w4(32'hb9ee5cd8),
	.w5(32'hb9d49150),
	.w6(32'h3a64c3ba),
	.w7(32'h389bc595),
	.w8(32'h381097b3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7321ff8),
	.w1(32'hb5cafcb5),
	.w2(32'hb5d6057f),
	.w3(32'h3601b791),
	.w4(32'h3729e60e),
	.w5(32'h37559888),
	.w6(32'h37ddd6e7),
	.w7(32'h37f62327),
	.w8(32'h378e397c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3778d07d),
	.w1(32'hb7001aa7),
	.w2(32'hb79d3c2b),
	.w3(32'hb788a8da),
	.w4(32'hb887dcb6),
	.w5(32'hb86b5857),
	.w6(32'hb7add461),
	.w7(32'hb893bf55),
	.w8(32'hb8a295fc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b29e24),
	.w1(32'h3a117350),
	.w2(32'h39d769f3),
	.w3(32'hba8efd24),
	.w4(32'hba2b786f),
	.w5(32'hb8b947bf),
	.w6(32'hbabe4929),
	.w7(32'hba84883f),
	.w8(32'hb97ce6ac),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92fe47f),
	.w1(32'h3a9ff318),
	.w2(32'h3b10a86e),
	.w3(32'h3acd20d1),
	.w4(32'h3b0918c4),
	.w5(32'h3af93d78),
	.w6(32'h39944c72),
	.w7(32'h3af02cbe),
	.w8(32'h3abbf98b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba873da9),
	.w1(32'hbabeae5e),
	.w2(32'hbac2e35c),
	.w3(32'h39f2f34e),
	.w4(32'h37e384d7),
	.w5(32'hb97174eb),
	.w6(32'h3aa9adbf),
	.w7(32'h3a9b0d73),
	.w8(32'h3acb6dc6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399149cc),
	.w1(32'hb9e13ea4),
	.w2(32'hbaca9596),
	.w3(32'h3a1139f4),
	.w4(32'h3a0b9043),
	.w5(32'h3909d1de),
	.w6(32'h3981a313),
	.w7(32'h38856e1a),
	.w8(32'h3a01a2c4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8a961),
	.w1(32'hb9b58610),
	.w2(32'h39911fb4),
	.w3(32'h398588d4),
	.w4(32'h37dce782),
	.w5(32'h39a79ffb),
	.w6(32'h393a7652),
	.w7(32'hb8d0df05),
	.w8(32'h39fb68f0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e83f9),
	.w1(32'h3ab5e7b1),
	.w2(32'h3b462adc),
	.w3(32'hba852734),
	.w4(32'h3b2bb8d3),
	.w5(32'h3b9e1901),
	.w6(32'hbb6f5402),
	.w7(32'hbac55553),
	.w8(32'h3a887b10),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836b654),
	.w1(32'hb6e4d3ba),
	.w2(32'hb76765c5),
	.w3(32'h371d724a),
	.w4(32'h37b73953),
	.w5(32'h3796d4ce),
	.w6(32'h380addf5),
	.w7(32'h381f040c),
	.w8(32'h37b42a12),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8daa317),
	.w1(32'h38d4fa14),
	.w2(32'hb8313bdf),
	.w3(32'h3896dd2a),
	.w4(32'h38fa6f2f),
	.w5(32'hb86e7250),
	.w6(32'h3824c094),
	.w7(32'h395d6d9a),
	.w8(32'h39388318),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb815f54b),
	.w1(32'hb62d3da3),
	.w2(32'hb7e3fd0c),
	.w3(32'hb762f83e),
	.w4(32'hb73c67a5),
	.w5(32'hb7605b30),
	.w6(32'hb81dcb56),
	.w7(32'hb7d2d1bd),
	.w8(32'hb70781d2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47870),
	.w1(32'h39f1f911),
	.w2(32'h39234196),
	.w3(32'h3a7232d9),
	.w4(32'h3a462ebf),
	.w5(32'h3a213c90),
	.w6(32'h3a72bbec),
	.w7(32'h3a4d6d3f),
	.w8(32'h391f04db),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883b64e),
	.w1(32'h38e37067),
	.w2(32'hb69e83c2),
	.w3(32'hb728c596),
	.w4(32'h3909ff28),
	.w5(32'h39459b93),
	.w6(32'hba2e01b0),
	.w7(32'hb9e04b76),
	.w8(32'hb9a4b288),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97dc1e2),
	.w1(32'h3ab58b57),
	.w2(32'h3aebcd78),
	.w3(32'h3a177f10),
	.w4(32'h3b3c81be),
	.w5(32'h3b5a42b5),
	.w6(32'hbabba1b3),
	.w7(32'hb956e38a),
	.w8(32'h3afb615f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2f9fb),
	.w1(32'h3920ffd9),
	.w2(32'h39536f3c),
	.w3(32'h381474da),
	.w4(32'h3a1525f2),
	.w5(32'h39e80dcc),
	.w6(32'hb9f32182),
	.w7(32'hb9e7fd08),
	.w8(32'hb86368c6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8090f1a),
	.w1(32'hb81f8dc8),
	.w2(32'hb8168f62),
	.w3(32'hb7a047fd),
	.w4(32'h370bde4f),
	.w5(32'h379f4f10),
	.w6(32'h3920de2a),
	.w7(32'h394fe3c4),
	.w8(32'h3920dba8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4bd5eb4),
	.w1(32'h3694ce5f),
	.w2(32'h372797bf),
	.w3(32'h3658c6db),
	.w4(32'h36a460bc),
	.w5(32'h377424f9),
	.w6(32'h3706949f),
	.w7(32'h37882cce),
	.w8(32'h37c4c86c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9154f8b),
	.w1(32'hb9508002),
	.w2(32'hb87b7e4f),
	.w3(32'h38971351),
	.w4(32'h38fe434c),
	.w5(32'h390478ce),
	.w6(32'h392876a3),
	.w7(32'h3975075a),
	.w8(32'h39892ce1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0950a0),
	.w1(32'hba088e47),
	.w2(32'hb9c9cdc0),
	.w3(32'hb9e7e46c),
	.w4(32'hb9d8a046),
	.w5(32'hb94b68b8),
	.w6(32'hb9d9636b),
	.w7(32'hb9f9be71),
	.w8(32'hb983090e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b81fbb),
	.w1(32'h388e92e2),
	.w2(32'hb73dedf7),
	.w3(32'h394ac00d),
	.w4(32'h39578a81),
	.w5(32'h3985b829),
	.w6(32'hb80b4fda),
	.w7(32'h390798d8),
	.w8(32'h39447c9a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399810b6),
	.w1(32'h3a1e4d49),
	.w2(32'h3a27f8a0),
	.w3(32'h3a0505a9),
	.w4(32'h3a836bf8),
	.w5(32'h3a9b5c0d),
	.w6(32'hba3c642c),
	.w7(32'h389a9262),
	.w8(32'h391f169c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a3ab7),
	.w1(32'h37aee32c),
	.w2(32'h3ac36331),
	.w3(32'h39dfd00a),
	.w4(32'h3a881851),
	.w5(32'h3aa0921d),
	.w6(32'h3955ada5),
	.w7(32'h395923b1),
	.w8(32'h39dbc43b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37012501),
	.w1(32'hb6624f87),
	.w2(32'hb64f02db),
	.w3(32'h37d104e1),
	.w4(32'h378b59e8),
	.w5(32'hb641436d),
	.w6(32'h3521b762),
	.w7(32'hb59d990b),
	.w8(32'h369b652e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb729d1a0),
	.w1(32'hb74e545d),
	.w2(32'hb78014a2),
	.w3(32'hb654680c),
	.w4(32'hb6e5e801),
	.w5(32'hb7174a33),
	.w6(32'h373085f9),
	.w7(32'h36d5b602),
	.w8(32'h360faad7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38106c65),
	.w1(32'h382c49e7),
	.w2(32'h3757d8a6),
	.w3(32'h37f1d193),
	.w4(32'h381ff59a),
	.w5(32'h37affb69),
	.w6(32'h3816be57),
	.w7(32'h3803a6be),
	.w8(32'h3719872d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c8f900),
	.w1(32'hb7734ae4),
	.w2(32'hb7c2a151),
	.w3(32'hb7321df7),
	.w4(32'hb7a0d8d1),
	.w5(32'hb78cbfc3),
	.w6(32'hb7ba5246),
	.w7(32'hb7fe4440),
	.w8(32'hb813a8da),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77bef5),
	.w1(32'hba1f70e7),
	.w2(32'h3a815cb9),
	.w3(32'h3a84e855),
	.w4(32'h3ade2db3),
	.w5(32'h3a26d2fe),
	.w6(32'h3a935473),
	.w7(32'h3a2b83a7),
	.w8(32'h3a985d80),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d69683),
	.w1(32'hb7070214),
	.w2(32'hbaa9a7e8),
	.w3(32'hba552313),
	.w4(32'h3aa8db6c),
	.w5(32'h3ac45a7e),
	.w6(32'hbb5165cc),
	.w7(32'hbb41932b),
	.w8(32'hba609275),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa38059),
	.w1(32'h3af61c92),
	.w2(32'h3b05913d),
	.w3(32'hb78e4dde),
	.w4(32'h3aa3dc29),
	.w5(32'h3b09128a),
	.w6(32'hbb28176d),
	.w7(32'hbacced8b),
	.w8(32'hbac2134f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a67f6),
	.w1(32'hbb8f1278),
	.w2(32'hbb72b136),
	.w3(32'h398a3d4a),
	.w4(32'hba923cdc),
	.w5(32'hbaaef600),
	.w6(32'h3b0e9a45),
	.w7(32'hb5d6173f),
	.w8(32'h3aa0b3cf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c9a52e),
	.w1(32'hb64cd351),
	.w2(32'hb5d12d34),
	.w3(32'hb686f93d),
	.w4(32'hb70df51c),
	.w5(32'hb65a6f5c),
	.w6(32'hb5572297),
	.w7(32'hb5e9a8c6),
	.w8(32'h376375d8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64fc232),
	.w1(32'h35a77bf4),
	.w2(32'hb69d45f3),
	.w3(32'hb622e371),
	.w4(32'hb67bee80),
	.w5(32'hb79ef315),
	.w6(32'h373663cc),
	.w7(32'h36d9f3f2),
	.w8(32'hb762a329),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3726ac4d),
	.w1(32'hb6e3310c),
	.w2(32'hb771144c),
	.w3(32'hb72dc545),
	.w4(32'hb7b0a299),
	.w5(32'hb7b42ca3),
	.w6(32'h363a59a9),
	.w7(32'hb6258ea4),
	.w8(32'hb7aa409b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ce7c5),
	.w1(32'h39faf52a),
	.w2(32'h39d4078f),
	.w3(32'h390a5e76),
	.w4(32'h39d2e493),
	.w5(32'h39f6a405),
	.w6(32'hba295ca3),
	.w7(32'hb9b95054),
	.w8(32'h38be8770),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369e5ec9),
	.w1(32'hb77e2838),
	.w2(32'hb78ae832),
	.w3(32'h36be8510),
	.w4(32'hb752e50c),
	.w5(32'hb75a1212),
	.w6(32'hb6046e83),
	.w7(32'hb74490ab),
	.w8(32'hb732c37c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd2786),
	.w1(32'h3a0cc95b),
	.w2(32'h3a39f335),
	.w3(32'hb31da7e0),
	.w4(32'h3a7a1914),
	.w5(32'h3aea125f),
	.w6(32'hba879f55),
	.w7(32'h38b4e7f3),
	.w8(32'h3a97fc46),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20fb8f),
	.w1(32'h3a8fc525),
	.w2(32'h3a5f292f),
	.w3(32'h3a1b5d28),
	.w4(32'h3ad41c00),
	.w5(32'h3b50b671),
	.w6(32'hbaf35448),
	.w7(32'hb8ad2678),
	.w8(32'h3a5cb23f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba061ccc),
	.w1(32'hba37cc90),
	.w2(32'hba34f559),
	.w3(32'h3a2340b8),
	.w4(32'h396dae0a),
	.w5(32'h3696386b),
	.w6(32'h3ac31704),
	.w7(32'h3a815b34),
	.w8(32'h3a906cb8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39beb00b),
	.w1(32'h399e8aac),
	.w2(32'h39e00b10),
	.w3(32'h3a872f9e),
	.w4(32'h3a84929b),
	.w5(32'h3a3ffd4f),
	.w6(32'h39dfb80d),
	.w7(32'h39b670fc),
	.w8(32'h3a067068),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d96613),
	.w1(32'h39b43ccd),
	.w2(32'h396fbad0),
	.w3(32'h394ca4f9),
	.w4(32'h3a8cd924),
	.w5(32'h3a6abdc8),
	.w6(32'hb9fd2ced),
	.w7(32'h39a7b165),
	.w8(32'h3a82434d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fd0e7),
	.w1(32'hb95235c4),
	.w2(32'hb8fbd852),
	.w3(32'h394444e2),
	.w4(32'h39ce025f),
	.w5(32'h38a02c05),
	.w6(32'h3a3de086),
	.w7(32'h3a822292),
	.w8(32'h3a8058af),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397bc03a),
	.w1(32'h3a497ec8),
	.w2(32'h3a886ef2),
	.w3(32'h3898cb9d),
	.w4(32'h3a9fa69e),
	.w5(32'h3aee3924),
	.w6(32'hba6914f2),
	.w7(32'h389a17b2),
	.w8(32'h3a59e5c8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3796a894),
	.w1(32'h3712ff02),
	.w2(32'hb679c9a2),
	.w3(32'h371f52b9),
	.w4(32'h361cd9fe),
	.w5(32'hb6c81dab),
	.w6(32'h364e22ae),
	.w7(32'hb6b371b9),
	.w8(32'hb67f5a81),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35117b96),
	.w1(32'h379912a1),
	.w2(32'h37cd9d07),
	.w3(32'h35c1f731),
	.w4(32'h37c66a40),
	.w5(32'h37a619c4),
	.w6(32'h37414e94),
	.w7(32'h37da972c),
	.w8(32'h37cf420d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38258393),
	.w1(32'h37945930),
	.w2(32'h37012b67),
	.w3(32'h386a65fe),
	.w4(32'h37473023),
	.w5(32'hb7e254c3),
	.w6(32'h3880d799),
	.w7(32'hb5f7758a),
	.w8(32'h36af2546),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff0a9c),
	.w1(32'hb996e3bf),
	.w2(32'hb9d14712),
	.w3(32'h38c78902),
	.w4(32'h3704bfff),
	.w5(32'hb8826e78),
	.w6(32'h39a4d56a),
	.w7(32'h3946b8d0),
	.w8(32'h38f79f42),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3893ba25),
	.w1(32'hb9ce3bd0),
	.w2(32'h3a0f9331),
	.w3(32'h3a814938),
	.w4(32'hba11f2d8),
	.w5(32'h391ad662),
	.w6(32'h3abb68af),
	.w7(32'h3981a3cf),
	.w8(32'h3a000cfc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdb206),
	.w1(32'hba24381d),
	.w2(32'hb9c92fb7),
	.w3(32'hb8f24000),
	.w4(32'hb952687e),
	.w5(32'h374916fd),
	.w6(32'hb9a5dc1e),
	.w7(32'hb99d4716),
	.w8(32'hb8c8d647),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbf7db),
	.w1(32'hb9871afc),
	.w2(32'hba9dc62a),
	.w3(32'h395aec94),
	.w4(32'hb92666d6),
	.w5(32'hba576b0a),
	.w6(32'h39b7cb4c),
	.w7(32'hb72032d5),
	.w8(32'h38f03643),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac42818),
	.w1(32'hb7fba08b),
	.w2(32'h3ab87ba6),
	.w3(32'hbac54e45),
	.w4(32'h3a8c1f38),
	.w5(32'h3b2cfddb),
	.w6(32'hbb54b14e),
	.w7(32'hbafd6de5),
	.w8(32'hb89ebe42),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0df3a),
	.w1(32'hbb00df1b),
	.w2(32'hbace31fd),
	.w3(32'hb91774fe),
	.w4(32'hba31864d),
	.w5(32'hb9c96c49),
	.w6(32'h3a258eef),
	.w7(32'hb9262c54),
	.w8(32'h395fd2bf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf65d29),
	.w1(32'hba5907b9),
	.w2(32'h3ad8f28f),
	.w3(32'h38a726f8),
	.w4(32'h37e9ec26),
	.w5(32'h3ab1b232),
	.w6(32'hbb2517e8),
	.w7(32'h39bdf5ca),
	.w8(32'h3b322e77),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9a393),
	.w1(32'hbaa9f9d5),
	.w2(32'hba7eb8fb),
	.w3(32'h3a0b3a3c),
	.w4(32'hba62ec3e),
	.w5(32'hb9ead74b),
	.w6(32'h3abea55c),
	.w7(32'hb99e9d9d),
	.w8(32'h394ed695),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9214da),
	.w1(32'hb91170ca),
	.w2(32'h3937603b),
	.w3(32'h3a66eafe),
	.w4(32'h3a5186c4),
	.w5(32'hb89926f6),
	.w6(32'hba0f21f5),
	.w7(32'h383ce1f8),
	.w8(32'hb96cb753),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dc727),
	.w1(32'h3935cde2),
	.w2(32'h3a100bf2),
	.w3(32'h38d044f1),
	.w4(32'h3a7dd3bc),
	.w5(32'h39d5102c),
	.w6(32'h3a4f4d2e),
	.w7(32'h3b08b003),
	.w8(32'h3b00ca58),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba086513),
	.w1(32'hbad1503a),
	.w2(32'hbb0a451b),
	.w3(32'h3a8ced6b),
	.w4(32'hb91af204),
	.w5(32'hb9fbc85f),
	.w6(32'h3b23097f),
	.w7(32'h3ae1c308),
	.w8(32'h3a89bb2a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ce293),
	.w1(32'hb9845498),
	.w2(32'hb8f26e9e),
	.w3(32'hb9227324),
	.w4(32'hb967b592),
	.w5(32'hb8cc0e84),
	.w6(32'hb900cba1),
	.w7(32'hb8c3e862),
	.w8(32'hb72c640d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c10496),
	.w1(32'h3a1bae34),
	.w2(32'h3a1ceef9),
	.w3(32'h3a14ab15),
	.w4(32'h3aecb673),
	.w5(32'h3a5171e6),
	.w6(32'hbaab440a),
	.w7(32'h3909372b),
	.w8(32'h3a3ebbb7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb7185),
	.w1(32'h3ae4695d),
	.w2(32'h3b361ef4),
	.w3(32'h3a8dd538),
	.w4(32'h3ab0f0ab),
	.w5(32'h3a7ea0f0),
	.w6(32'hb9407875),
	.w7(32'h3aa776f8),
	.w8(32'h3b105415),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4edb7b),
	.w1(32'h3aca1dfd),
	.w2(32'h3bda85bb),
	.w3(32'hb9f69b60),
	.w4(32'hbad3906e),
	.w5(32'h38e00b6d),
	.w6(32'hbb7831fa),
	.w7(32'hbb70b6ef),
	.w8(32'hbb4653e1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1c7d2),
	.w1(32'hbbccc8c7),
	.w2(32'hbbd0bb1d),
	.w3(32'hbb8b6abf),
	.w4(32'hbc00a171),
	.w5(32'h3b3b989d),
	.w6(32'hbb445ca9),
	.w7(32'hbbf1d4db),
	.w8(32'h3b0e6580),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ad501),
	.w1(32'hbabebafb),
	.w2(32'h394c80c5),
	.w3(32'h3a460f12),
	.w4(32'hbb2dc966),
	.w5(32'h3addb49e),
	.w6(32'h3a5f2101),
	.w7(32'h3b221d00),
	.w8(32'h3b580b4c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7f172),
	.w1(32'hbadbdae5),
	.w2(32'h3a8f9f95),
	.w3(32'h3b201b63),
	.w4(32'h3b08131e),
	.w5(32'hbb604ad9),
	.w6(32'hbab7635f),
	.w7(32'h3a3d482f),
	.w8(32'hbb68c8e2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba33d6c),
	.w1(32'hb9325fb4),
	.w2(32'hbb42b6a6),
	.w3(32'hba822068),
	.w4(32'hbb92e538),
	.w5(32'h3ae63f27),
	.w6(32'hbb4e858c),
	.w7(32'hbb88d130),
	.w8(32'h3a3e89cb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ea2f73),
	.w1(32'h39395ef1),
	.w2(32'h3a60b6d7),
	.w3(32'h3b0a9446),
	.w4(32'hba5a9f0c),
	.w5(32'h3b407036),
	.w6(32'h3a447427),
	.w7(32'hb9e81c22),
	.w8(32'h3b3eeb70),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee20ec),
	.w1(32'hbb8bb38d),
	.w2(32'hba616863),
	.w3(32'hbb8d186d),
	.w4(32'hbb7f1c23),
	.w5(32'hb9e6fc20),
	.w6(32'hbbbef1cc),
	.w7(32'hbb947469),
	.w8(32'h3b84eff6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a716bc9),
	.w1(32'hbb3885ef),
	.w2(32'hbb08f603),
	.w3(32'h3b2270da),
	.w4(32'hbb1a25d2),
	.w5(32'h3a2c9f2e),
	.w6(32'h3ab6ebbc),
	.w7(32'hbba60107),
	.w8(32'hb98ac7e9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a200f9f),
	.w1(32'hb990b676),
	.w2(32'hb9e29716),
	.w3(32'hba840fc0),
	.w4(32'hb98649aa),
	.w5(32'hba76284f),
	.w6(32'hbb50bb17),
	.w7(32'hbb53a7d2),
	.w8(32'hba418ceb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e4760),
	.w1(32'h3ab177bf),
	.w2(32'h3ab31729),
	.w3(32'h3ac0c036),
	.w4(32'h3abae247),
	.w5(32'h3b8ae481),
	.w6(32'hb89dc523),
	.w7(32'h39a7fc67),
	.w8(32'h3b9921d6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f60f9),
	.w1(32'hbaf2e750),
	.w2(32'hbab915bf),
	.w3(32'hb9704dbb),
	.w4(32'hb98c073d),
	.w5(32'h3b8a3da2),
	.w6(32'hb986f34e),
	.w7(32'hbaff1031),
	.w8(32'h3b2038f4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a887ef5),
	.w1(32'hbaefb1a6),
	.w2(32'h3bb740de),
	.w3(32'h3b14a9e7),
	.w4(32'h3ab8507d),
	.w5(32'h3b0728f0),
	.w6(32'h39bf0264),
	.w7(32'h3b4fe371),
	.w8(32'hb90e766e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19fd8d),
	.w1(32'hb9e0adc6),
	.w2(32'h3a325e6f),
	.w3(32'hba509097),
	.w4(32'hbb2ff5e1),
	.w5(32'h3bc5d66f),
	.w6(32'hb7d70500),
	.w7(32'hba9bde72),
	.w8(32'h3bfef841),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ed635),
	.w1(32'h3ab971c1),
	.w2(32'hb6dcf170),
	.w3(32'h3b43e90d),
	.w4(32'h3b949911),
	.w5(32'h39edffef),
	.w6(32'h3b4eaa2a),
	.w7(32'hb705d69f),
	.w8(32'hbb1ecd57),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d1204),
	.w1(32'hbb33bb6e),
	.w2(32'hbb2825f4),
	.w3(32'h3b18351d),
	.w4(32'h3b347f4a),
	.w5(32'h3a842872),
	.w6(32'hbabd3ee8),
	.w7(32'hba9a11b7),
	.w8(32'h3add93dc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a6634d),
	.w1(32'hb9214ba1),
	.w2(32'h3b1dd1b8),
	.w3(32'h3a93404e),
	.w4(32'h3b7ead29),
	.w5(32'h3a229cea),
	.w6(32'h3a2128c6),
	.w7(32'h3b883640),
	.w8(32'hba8ef818),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac743f5),
	.w1(32'h3a060f87),
	.w2(32'h3b51a269),
	.w3(32'hbacec6f7),
	.w4(32'hbb3204a6),
	.w5(32'h3abddd88),
	.w6(32'hbad3b785),
	.w7(32'hb884f023),
	.w8(32'h3ab7ca8a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922b414),
	.w1(32'h3b8a5963),
	.w2(32'h3b024d4b),
	.w3(32'h3b845f01),
	.w4(32'h3be89eb7),
	.w5(32'h391badf2),
	.w6(32'h3b9168c1),
	.w7(32'h3b96c852),
	.w8(32'h3b2af2d7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b033d),
	.w1(32'h3b5e9af7),
	.w2(32'h3a484c4e),
	.w3(32'hba8657ae),
	.w4(32'hba1a8cdf),
	.w5(32'hbafbe155),
	.w6(32'h3b803b43),
	.w7(32'h3a40d0d0),
	.w8(32'hbae902b4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad298f),
	.w1(32'hbae3cee7),
	.w2(32'hbb34f019),
	.w3(32'hbb0ab343),
	.w4(32'hbb22342e),
	.w5(32'hbc16d422),
	.w6(32'hbb3ba105),
	.w7(32'hbb48bda4),
	.w8(32'hbc1ea0ba),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf21f1d),
	.w1(32'hbbe43769),
	.w2(32'hbc0838db),
	.w3(32'hbbbc27a7),
	.w4(32'hbbe06f95),
	.w5(32'h3ae2d4b8),
	.w6(32'hbc02d827),
	.w7(32'hbbe549cf),
	.w8(32'h3a89a764),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad33ac9),
	.w1(32'h39392243),
	.w2(32'h3ac00b8a),
	.w3(32'h3b6a5c8a),
	.w4(32'h3aa3059e),
	.w5(32'h3b897fb2),
	.w6(32'h3a5efed1),
	.w7(32'h3a86a4c8),
	.w8(32'hb9d46242),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f4fa7),
	.w1(32'hbbc7954a),
	.w2(32'h3ab29d34),
	.w3(32'hbba0485f),
	.w4(32'hbb404261),
	.w5(32'hbc025ba8),
	.w6(32'hbbff60f2),
	.w7(32'hb96d0de8),
	.w8(32'hb8fca878),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a243b),
	.w1(32'h3ada21ab),
	.w2(32'h3bb2ba1e),
	.w3(32'hbc071e0f),
	.w4(32'hbbe913ee),
	.w5(32'h3a3775fc),
	.w6(32'hbbb584f8),
	.w7(32'hbac2c25a),
	.w8(32'h3b43774e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de9996),
	.w1(32'hbb39812d),
	.w2(32'h3a048e0d),
	.w3(32'hbb738e2a),
	.w4(32'h3b6bdf57),
	.w5(32'hbb1f94dc),
	.w6(32'hbb446cd5),
	.w7(32'h3b6fc8d7),
	.w8(32'hbb1c569f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e18b),
	.w1(32'hb9cd63fe),
	.w2(32'h3a8fb05c),
	.w3(32'hbbbefd8b),
	.w4(32'hbb836fe0),
	.w5(32'hba1e7ec3),
	.w6(32'hbbc958e3),
	.w7(32'hbb489ddb),
	.w8(32'hbaf4ff0c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e5db4),
	.w1(32'h39bd0f3d),
	.w2(32'hba4a0b38),
	.w3(32'hb8e4b7e7),
	.w4(32'hba3bba8d),
	.w5(32'hbb0c3f0f),
	.w6(32'hbae58af2),
	.w7(32'hbb130f8f),
	.w8(32'h3642cd08),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17fcf1),
	.w1(32'h398b3197),
	.w2(32'hbaad6707),
	.w3(32'hbb1fc689),
	.w4(32'hba8ff5ad),
	.w5(32'h39edf1ea),
	.w6(32'hbb95296f),
	.w7(32'hbb05b5ce),
	.w8(32'hbb031d2d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b6754),
	.w1(32'h3a93cc90),
	.w2(32'hb97e4fac),
	.w3(32'hb9868eaa),
	.w4(32'h3ad2e6c5),
	.w5(32'h3c000d66),
	.w6(32'hbb96ffe1),
	.w7(32'hbb359fae),
	.w8(32'h3bbacb13),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d63a3),
	.w1(32'hbb8a9b7f),
	.w2(32'hbb62334c),
	.w3(32'h3b6c17c8),
	.w4(32'h393aa165),
	.w5(32'h3a8eaf8c),
	.w6(32'hbb9d0ee9),
	.w7(32'hbb8b29b5),
	.w8(32'h3bbec7db),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93d0cf),
	.w1(32'h3b7d9078),
	.w2(32'h3b3050fa),
	.w3(32'hba3675cd),
	.w4(32'h3bb85e9c),
	.w5(32'h3b90fe30),
	.w6(32'h3b31c799),
	.w7(32'h3b730642),
	.w8(32'h3b304617),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addef0c),
	.w1(32'h3a584285),
	.w2(32'hbab11953),
	.w3(32'h3b0ae0bf),
	.w4(32'hbb0adabe),
	.w5(32'hbacf3200),
	.w6(32'hba64656c),
	.w7(32'hbb8ca51b),
	.w8(32'hba1a822c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128c82),
	.w1(32'hbb10d031),
	.w2(32'hbb0a4fe8),
	.w3(32'hbaa33c99),
	.w4(32'hbb615232),
	.w5(32'hbb83e123),
	.w6(32'hba83ff49),
	.w7(32'hbb1910f2),
	.w8(32'hbb1d13ce),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12b4a1),
	.w1(32'hbb170f64),
	.w2(32'hbc03c45b),
	.w3(32'hbb093230),
	.w4(32'hbbb53ae4),
	.w5(32'h3b546746),
	.w6(32'hbbd52bb8),
	.w7(32'hbc20f3ad),
	.w8(32'h3b4a0763),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeadf0),
	.w1(32'h3a8563eb),
	.w2(32'h3a8903b5),
	.w3(32'h3adc320f),
	.w4(32'hb9063412),
	.w5(32'h3aca83a8),
	.w6(32'h3aa27152),
	.w7(32'hba7a0251),
	.w8(32'h3b37373f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb5a36),
	.w1(32'h3b0dac8b),
	.w2(32'hb99b60ed),
	.w3(32'h3b2a3e41),
	.w4(32'h3b8eab09),
	.w5(32'h3c1a95af),
	.w6(32'hba8a5845),
	.w7(32'h3993a0e9),
	.w8(32'h3b5eaa66),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb2d2),
	.w1(32'hbb2e6b24),
	.w2(32'h3b10cbad),
	.w3(32'h3c182049),
	.w4(32'h3b9ff282),
	.w5(32'h3bb59b4b),
	.w6(32'h3b4674bb),
	.w7(32'h3b635cb7),
	.w8(32'h3bcd9bc0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b730775),
	.w1(32'h3b19f4cf),
	.w2(32'h3b8d8325),
	.w3(32'h3b2f420c),
	.w4(32'h3b929d28),
	.w5(32'h39f377cb),
	.w6(32'h3af57939),
	.w7(32'h3b048dc5),
	.w8(32'h3a674b1d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefe0cd),
	.w1(32'h3a7c5d23),
	.w2(32'hbaaf64f3),
	.w3(32'hbac4b894),
	.w4(32'hba8236a1),
	.w5(32'h3b5dfc68),
	.w6(32'hbb1f78f8),
	.w7(32'hbb12d3f6),
	.w8(32'h3b68d988),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a293ec0),
	.w1(32'hbaadf3a1),
	.w2(32'hbb0cab30),
	.w3(32'h3a9de72a),
	.w4(32'hbb0e0e0f),
	.w5(32'h3b64ba37),
	.w6(32'hba4857dd),
	.w7(32'hbb76de73),
	.w8(32'h3b3e12a6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc70da),
	.w1(32'hbb26f260),
	.w2(32'hbb4d0799),
	.w3(32'h3b7a7000),
	.w4(32'h3b1618d0),
	.w5(32'h3a610398),
	.w6(32'h3aca89ae),
	.w7(32'hbac3b718),
	.w8(32'h3af5db7b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba092993),
	.w1(32'hbbdfac20),
	.w2(32'h3a8a6aaf),
	.w3(32'hbb93ff39),
	.w4(32'hbac189bb),
	.w5(32'h3a55cb82),
	.w6(32'hbc00834a),
	.w7(32'hbb95230f),
	.w8(32'h3997041f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e290b),
	.w1(32'hbb8bf044),
	.w2(32'hbb693437),
	.w3(32'h3af60067),
	.w4(32'hba3b6ea1),
	.w5(32'h3b813203),
	.w6(32'h3b3bb010),
	.w7(32'h3b0a93ab),
	.w8(32'h3b639b53),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0a780),
	.w1(32'hba5dac5c),
	.w2(32'h3b26af6b),
	.w3(32'h3ae679da),
	.w4(32'h3a23a3cd),
	.w5(32'h3ac3d454),
	.w6(32'h3a1b6a9f),
	.w7(32'h3b0c325d),
	.w8(32'h3b8e8a40),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd59a5),
	.w1(32'h3c04a9e7),
	.w2(32'h3b8d2099),
	.w3(32'h3c09c161),
	.w4(32'h3bab2af4),
	.w5(32'h3b3691b6),
	.w6(32'h3be68884),
	.w7(32'h3bdb404c),
	.w8(32'h3b254d27),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ef43),
	.w1(32'hbb50bbf8),
	.w2(32'hbad7534e),
	.w3(32'hbb056c35),
	.w4(32'h39f208ea),
	.w5(32'h37b7b400),
	.w6(32'hbbb99a70),
	.w7(32'hbb851587),
	.w8(32'h3a48a899),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3ce11),
	.w1(32'hbb1ebd73),
	.w2(32'hbb43a341),
	.w3(32'hbb0c1136),
	.w4(32'hbb5c9a64),
	.w5(32'hbafdaf17),
	.w6(32'hbb4c6f92),
	.w7(32'hbb82ea36),
	.w8(32'hbac7b55d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e96613),
	.w1(32'h3a46ffc3),
	.w2(32'h3a83641c),
	.w3(32'hba4b593f),
	.w4(32'hbb15a136),
	.w5(32'hba488ff1),
	.w6(32'hb98b3bb0),
	.w7(32'h39c40dad),
	.w8(32'h3b09e9a8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf80c5f),
	.w1(32'h3a26e6c0),
	.w2(32'hbaf0e491),
	.w3(32'h3a79aea1),
	.w4(32'h3a44f421),
	.w5(32'hbb946ca0),
	.w6(32'h39fc251c),
	.w7(32'hbb0a81df),
	.w8(32'hbb42b99e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d47e1a),
	.w1(32'h3c079404),
	.w2(32'h3bb900a1),
	.w3(32'h3b952064),
	.w4(32'h3bc54107),
	.w5(32'h3a8d01b4),
	.w6(32'h3b95c41b),
	.w7(32'h3bfa2752),
	.w8(32'h390ef842),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ee672),
	.w1(32'h3b3595f0),
	.w2(32'h3abb4da3),
	.w3(32'h3ba2ea08),
	.w4(32'h3bf53e5d),
	.w5(32'h3b529536),
	.w6(32'h3b93d305),
	.w7(32'h3ba4403e),
	.w8(32'h3b95efbb),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63ff91),
	.w1(32'hbb11e524),
	.w2(32'hbb8065eb),
	.w3(32'h3b825741),
	.w4(32'h3af64720),
	.w5(32'h3b8f702d),
	.w6(32'h3aff73cc),
	.w7(32'hbaa9e458),
	.w8(32'h3b77e91f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb50dd),
	.w1(32'h3b450d8f),
	.w2(32'h3bb9e6e4),
	.w3(32'h3c1615a0),
	.w4(32'h3b9b46ff),
	.w5(32'h3a9c0920),
	.w6(32'h3b2a7868),
	.w7(32'h3b7283ac),
	.w8(32'h3aa29422),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ea3a1),
	.w1(32'hbad0265e),
	.w2(32'hbaf6d3ca),
	.w3(32'hbb1b5131),
	.w4(32'hbb818f2d),
	.w5(32'hbb1e08cd),
	.w6(32'hbb5c2181),
	.w7(32'h39f5da5d),
	.w8(32'hbb8578d4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad93c2),
	.w1(32'hbb327ee9),
	.w2(32'hba1f07f0),
	.w3(32'hba98b98b),
	.w4(32'h39cdc089),
	.w5(32'hbb0cb62b),
	.w6(32'hbba11af7),
	.w7(32'hb9fa912c),
	.w8(32'hbad004a3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba481bac),
	.w1(32'hbaaef422),
	.w2(32'hbac69b73),
	.w3(32'hba39f77f),
	.w4(32'hba8376a5),
	.w5(32'h3b94e364),
	.w6(32'hba9b0304),
	.w7(32'hbb10088c),
	.w8(32'h3bcdacf7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1d5a),
	.w1(32'h39a59cc0),
	.w2(32'hb975cfbd),
	.w3(32'h39032934),
	.w4(32'h3a245a6d),
	.w5(32'hbaffac80),
	.w6(32'hba95c492),
	.w7(32'hbacf55d7),
	.w8(32'h3ad3b869),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac400ab),
	.w1(32'hb97e9b54),
	.w2(32'h3a41adfa),
	.w3(32'hbab02f99),
	.w4(32'hba1569fa),
	.w5(32'hbaac8a15),
	.w6(32'h3aa1d9f3),
	.w7(32'h3a93fb86),
	.w8(32'hbaec5270),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507bc4),
	.w1(32'hbbc5b66d),
	.w2(32'h378db259),
	.w3(32'hbbb75f36),
	.w4(32'hbaf60ae0),
	.w5(32'h3acee97f),
	.w6(32'hbbc20fd7),
	.w7(32'h3a4d426d),
	.w8(32'hbaaa6f82),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaf4f6),
	.w1(32'h3a179309),
	.w2(32'h3b8081aa),
	.w3(32'hbb83ef57),
	.w4(32'hbb670b2a),
	.w5(32'hbac3a80a),
	.w6(32'hbba259df),
	.w7(32'h3bbaff33),
	.w8(32'hba3cea2a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c5b3),
	.w1(32'hbb3bc853),
	.w2(32'hbaa2f9aa),
	.w3(32'h3a348ce5),
	.w4(32'h3b5b8c70),
	.w5(32'hbaaed938),
	.w6(32'hbaa5b062),
	.w7(32'hbabd6d2c),
	.w8(32'hbaf77c26),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69253c),
	.w1(32'hba0f3980),
	.w2(32'h3b52f0be),
	.w3(32'hbb71239b),
	.w4(32'hbaa1a997),
	.w5(32'h3b3ad24a),
	.w6(32'hbbbb7496),
	.w7(32'h3ae9ac0c),
	.w8(32'h3b682026),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b8b3),
	.w1(32'hbacb7e52),
	.w2(32'hbb6d7d5b),
	.w3(32'hbaac551f),
	.w4(32'hbba4e094),
	.w5(32'hbb8133dd),
	.w6(32'hbb007c2f),
	.w7(32'hbba9b764),
	.w8(32'h3a7efd58),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc810ba),
	.w1(32'h396cae3e),
	.w2(32'hbb19d2af),
	.w3(32'hbbb82ac7),
	.w4(32'hbb2b8889),
	.w5(32'h3b241be5),
	.w6(32'hbb297956),
	.w7(32'hba7b74a3),
	.w8(32'h3aaa4d87),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7467a),
	.w1(32'h3a5092c4),
	.w2(32'h38f91f05),
	.w3(32'h3aaa0974),
	.w4(32'hba43e2e9),
	.w5(32'h39f5e8e9),
	.w6(32'hb99556fe),
	.w7(32'hba0daf3d),
	.w8(32'hba6399fa),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc1ebd),
	.w1(32'h3ae5ea24),
	.w2(32'hbaa7b55d),
	.w3(32'hbb384578),
	.w4(32'hba8c0b6d),
	.w5(32'h39c4a035),
	.w6(32'hbb315a4d),
	.w7(32'h3921abfc),
	.w8(32'hbadea291),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8b339),
	.w1(32'h3ae5243b),
	.w2(32'h3aeff451),
	.w3(32'h3ae3ead9),
	.w4(32'h3afc0d59),
	.w5(32'h3bb47711),
	.w6(32'h3b4c7cf1),
	.w7(32'h3b49fb9d),
	.w8(32'h3b6ef707),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a234),
	.w1(32'hbae740e3),
	.w2(32'hbb1ac96d),
	.w3(32'h3aedaf71),
	.w4(32'h3b8ac2eb),
	.w5(32'h3be1e825),
	.w6(32'h3aedc638),
	.w7(32'h3b5bdf6a),
	.w8(32'h3be93fae),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3cb32),
	.w1(32'h3b68aefa),
	.w2(32'hba63b568),
	.w3(32'h3c057c2d),
	.w4(32'h3ae0993f),
	.w5(32'h3a25be09),
	.w6(32'h3c1b603f),
	.w7(32'h3aaa8e7e),
	.w8(32'h3b106232),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ddb1a),
	.w1(32'hbb1df271),
	.w2(32'hba3fe904),
	.w3(32'hbb04401e),
	.w4(32'h3a87ff6e),
	.w5(32'hbad9304e),
	.w6(32'hbaef6031),
	.w7(32'hba88ae41),
	.w8(32'hbb874143),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab480),
	.w1(32'hbb81b949),
	.w2(32'hbba76f44),
	.w3(32'hbb27235c),
	.w4(32'hbb3f1d19),
	.w5(32'hbbcfd6a8),
	.w6(32'hbbdeb840),
	.w7(32'hbbb0542d),
	.w8(32'hbbac1fc6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76da1a),
	.w1(32'hbaa6f5e8),
	.w2(32'hbaf2d198),
	.w3(32'hbb271034),
	.w4(32'hbb8091bc),
	.w5(32'h3a9f5d56),
	.w6(32'h3a427e89),
	.w7(32'hbb1d5d76),
	.w8(32'h3b74b128),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39bb65),
	.w1(32'hbb351e1f),
	.w2(32'hbb0b04a7),
	.w3(32'hbb8c5ede),
	.w4(32'hbb63443b),
	.w5(32'hbb9ef73a),
	.w6(32'hbbb8a04b),
	.w7(32'hbbdb577d),
	.w8(32'hbb858d15),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2190),
	.w1(32'hbb58b796),
	.w2(32'hbb86d8e6),
	.w3(32'hbb446c74),
	.w4(32'hbb62af07),
	.w5(32'h3b6f3c55),
	.w6(32'hbb8d0ca5),
	.w7(32'hbb7709d9),
	.w8(32'hb8ecce9f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b115f82),
	.w1(32'hb91380dd),
	.w2(32'h3b2fbf29),
	.w3(32'hba1836c0),
	.w4(32'h39c7b427),
	.w5(32'hbacc2d65),
	.w6(32'hbbfef633),
	.w7(32'hbb482542),
	.w8(32'hbb549647),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2969b),
	.w1(32'h39582d6f),
	.w2(32'hba90171b),
	.w3(32'h3a8553d7),
	.w4(32'h3aa30934),
	.w5(32'h3bb5fe82),
	.w6(32'hbb1f801b),
	.w7(32'hbab11b37),
	.w8(32'h3b8c038c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b337b16),
	.w1(32'h3b2f48aa),
	.w2(32'h3ba88395),
	.w3(32'h3afee829),
	.w4(32'h3bf938ce),
	.w5(32'h3aa7bc97),
	.w6(32'h3b801d8e),
	.w7(32'h3be08877),
	.w8(32'hbaba5170),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15667b),
	.w1(32'hbb8b7b10),
	.w2(32'hb9ad49d3),
	.w3(32'hbb75e2ef),
	.w4(32'hbb1fe1ff),
	.w5(32'h3b0578b4),
	.w6(32'hbbe2518a),
	.w7(32'hbb4b1528),
	.w8(32'h3a85a761),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2dcbc),
	.w1(32'h3b77cb60),
	.w2(32'h3b072221),
	.w3(32'h3ba65975),
	.w4(32'h3bdc1fc2),
	.w5(32'hbaf7db20),
	.w6(32'h3b507e02),
	.w7(32'h3bbaff48),
	.w8(32'hbb4ed8bb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03a9e2),
	.w1(32'h3ab34598),
	.w2(32'hb9a64dcc),
	.w3(32'h3b189ae1),
	.w4(32'h39bc5e7d),
	.w5(32'hbaa57c5a),
	.w6(32'hb998e83f),
	.w7(32'hba11c465),
	.w8(32'h3a670c78),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8588f1),
	.w1(32'h3ad8b6f2),
	.w2(32'h38d5b15b),
	.w3(32'hbaac8dbc),
	.w4(32'h3a3b7699),
	.w5(32'h388589a9),
	.w6(32'hb8dd0667),
	.w7(32'hb8b17749),
	.w8(32'hba4cdb91),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3af88),
	.w1(32'hbb97c381),
	.w2(32'hbb25cb4d),
	.w3(32'h3abbb1de),
	.w4(32'hba97262d),
	.w5(32'h3b59f429),
	.w6(32'hb9faf277),
	.w7(32'hbb008b4d),
	.w8(32'h39ba87ed),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3c8a),
	.w1(32'h3b238fe1),
	.w2(32'hba58abae),
	.w3(32'h3bb972d2),
	.w4(32'hba094d2a),
	.w5(32'hbb016c6c),
	.w6(32'h3b8b1da9),
	.w7(32'h3b062a98),
	.w8(32'h39ee86d4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eeeeab),
	.w1(32'h3aaffe75),
	.w2(32'hbab6643b),
	.w3(32'h3920c70c),
	.w4(32'hb9c8e555),
	.w5(32'hbb57757e),
	.w6(32'hba0b539e),
	.w7(32'hbb169caa),
	.w8(32'h3a16edbd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390fd2),
	.w1(32'h3b0688c6),
	.w2(32'h3aa2c113),
	.w3(32'h3ae95e3e),
	.w4(32'h3b0ea044),
	.w5(32'h3a6809fd),
	.w6(32'h3a6a0740),
	.w7(32'h3aee5eeb),
	.w8(32'h3b0b3e3a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f102),
	.w1(32'h3b70a28b),
	.w2(32'h3b850e77),
	.w3(32'h3ace5173),
	.w4(32'h3b99b217),
	.w5(32'h3ac2b37a),
	.w6(32'h3a8bad09),
	.w7(32'h3b22d40f),
	.w8(32'h39a82e51),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a182ad5),
	.w1(32'hba0baf9a),
	.w2(32'h3a033f57),
	.w3(32'h3b8808ef),
	.w4(32'hba484c8e),
	.w5(32'h3b4edd59),
	.w6(32'h3b23d2b1),
	.w7(32'hb8f372b4),
	.w8(32'h3b24ac35),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937ea29),
	.w1(32'h3b78cfe9),
	.w2(32'h3ab20082),
	.w3(32'h3b9b5452),
	.w4(32'h3bd223a1),
	.w5(32'h3b1cbd57),
	.w6(32'h3b40703b),
	.w7(32'h3ba7c70f),
	.w8(32'hb980edb0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d67e5),
	.w1(32'h3c0a6e44),
	.w2(32'h3b8cb70e),
	.w3(32'h3bd83952),
	.w4(32'h3c0a39d6),
	.w5(32'h3c04aa02),
	.w6(32'h3a680d5d),
	.w7(32'h3b30de72),
	.w8(32'h3b80675e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b965a),
	.w1(32'hbba89922),
	.w2(32'hbaa4c765),
	.w3(32'h3af550a1),
	.w4(32'h3b73e288),
	.w5(32'hba8d196a),
	.w6(32'h3aa54bee),
	.w7(32'h3b71529a),
	.w8(32'h3abfc9f7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ec129),
	.w1(32'h3ab4cae8),
	.w2(32'h3b1efb67),
	.w3(32'hba845a6f),
	.w4(32'h3a748543),
	.w5(32'hba4fc8e0),
	.w6(32'hbbe77e85),
	.w7(32'hba8a3004),
	.w8(32'h3a3d3b01),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97e3da),
	.w1(32'h3a09eb82),
	.w2(32'hba704503),
	.w3(32'hbb190851),
	.w4(32'hbae89a2b),
	.w5(32'hba9202ad),
	.w6(32'hbb41e29f),
	.w7(32'hbb5537f7),
	.w8(32'h3afc698e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fcbf7),
	.w1(32'h3a8e3a40),
	.w2(32'h37f18419),
	.w3(32'hb8f27cf1),
	.w4(32'h3a43bd79),
	.w5(32'hbb71243a),
	.w6(32'h3ac9ed76),
	.w7(32'h3aad6ef5),
	.w8(32'h3aca7ddc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba472c7),
	.w1(32'h3b357a46),
	.w2(32'h3aef2e1c),
	.w3(32'h3aad1428),
	.w4(32'h3bacae7e),
	.w5(32'hbb562a9a),
	.w6(32'h399e3a23),
	.w7(32'h3b55a3e9),
	.w8(32'hba8aace5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb126d5f),
	.w1(32'hba556953),
	.w2(32'hba712988),
	.w3(32'hbb1f9646),
	.w4(32'hb9c7d71f),
	.w5(32'h3bf83310),
	.w6(32'hbb9c34bb),
	.w7(32'hbb480634),
	.w8(32'h3b892e87),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f76d8),
	.w1(32'hbb96fa51),
	.w2(32'h39c35680),
	.w3(32'h3b83ec6e),
	.w4(32'hbb32b3b9),
	.w5(32'hba8e2db9),
	.w6(32'hbb0e3d1f),
	.w7(32'hbb4c7541),
	.w8(32'hbbaf8a9a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fa37a),
	.w1(32'hbb1f1098),
	.w2(32'h3b3675e5),
	.w3(32'hbb86b5bd),
	.w4(32'h3b0d7ea2),
	.w5(32'hba8d862d),
	.w6(32'hbab152a5),
	.w7(32'h3b4adea2),
	.w8(32'hbaea214e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65ec2b),
	.w1(32'h3a27d078),
	.w2(32'h3b083d4d),
	.w3(32'h3b468aa7),
	.w4(32'h3ad979cb),
	.w5(32'h3b24fa60),
	.w6(32'h3a615c10),
	.w7(32'h3aeb3ccf),
	.w8(32'h3acddf32),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214357),
	.w1(32'hbaa8d34f),
	.w2(32'h3aa02899),
	.w3(32'hbb0d8cfc),
	.w4(32'hbb1ad94a),
	.w5(32'hbaa6e03a),
	.w6(32'hbb8b7e05),
	.w7(32'hbb8c4e5c),
	.w8(32'hbabc2087),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb4744),
	.w1(32'h3aababad),
	.w2(32'h3aa514cc),
	.w3(32'hbb1c3f89),
	.w4(32'hbade0653),
	.w5(32'hb914edc2),
	.w6(32'hba376a79),
	.w7(32'h3a4b56af),
	.w8(32'hba995ef3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb667e97),
	.w1(32'h3b4922c4),
	.w2(32'h3a2859c4),
	.w3(32'h3bcc1750),
	.w4(32'h3b9d54a2),
	.w5(32'hba97dfb4),
	.w6(32'h3b5e61a7),
	.w7(32'h3bbe5234),
	.w8(32'h3bc02f81),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39077603),
	.w1(32'h3a8c7857),
	.w2(32'hbb5fc3fd),
	.w3(32'hbab6274c),
	.w4(32'hba65fa8f),
	.w5(32'h3aa72362),
	.w6(32'hbb7f06b5),
	.w7(32'hbac7da2a),
	.w8(32'h3b5ddeeb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae786f6),
	.w1(32'hba6b6c27),
	.w2(32'hbb5c5c05),
	.w3(32'hbadf6fa4),
	.w4(32'hbb29af07),
	.w5(32'h3be7ec57),
	.w6(32'hbac9e68e),
	.w7(32'hbb758f30),
	.w8(32'h3c0c5309),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13258d),
	.w1(32'hbaa62798),
	.w2(32'hb9b9be81),
	.w3(32'h3ae40037),
	.w4(32'hbafaf874),
	.w5(32'hba03242c),
	.w6(32'h399ae64c),
	.w7(32'hbb8982c0),
	.w8(32'hbacbc798),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc144d),
	.w1(32'hbb20b846),
	.w2(32'hbac2777e),
	.w3(32'hbb578e1f),
	.w4(32'hbb89d430),
	.w5(32'hb985f1c4),
	.w6(32'hbb835512),
	.w7(32'hbbc036be),
	.w8(32'hb9c6f190),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cafb3),
	.w1(32'hbb5172db),
	.w2(32'hbb65ca9e),
	.w3(32'hba18b148),
	.w4(32'hbb030fed),
	.w5(32'hbb443366),
	.w6(32'hba6ccea6),
	.w7(32'hbb0bbfac),
	.w8(32'hba5f5dd6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a592f),
	.w1(32'hbaa0e281),
	.w2(32'hbb34ed74),
	.w3(32'hbb2bd208),
	.w4(32'hbb8cde54),
	.w5(32'h3900fad3),
	.w6(32'hbb59c48f),
	.w7(32'hbb9eb7a6),
	.w8(32'hba589433),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f0874),
	.w1(32'hbb09711b),
	.w2(32'h3a2d3831),
	.w3(32'hb929d0fe),
	.w4(32'hbb184ae8),
	.w5(32'h3c0ac135),
	.w6(32'hbae12465),
	.w7(32'hbacc9b0d),
	.w8(32'h3c0b8813),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be65163),
	.w1(32'hb82959d0),
	.w2(32'h3b2004c8),
	.w3(32'h3a329045),
	.w4(32'h3b043b8c),
	.w5(32'h390e2deb),
	.w6(32'hbaf2e8f9),
	.w7(32'hb9cde32b),
	.w8(32'hbae1577a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5d24),
	.w1(32'h3bb5e886),
	.w2(32'h3be2906b),
	.w3(32'h3c00d233),
	.w4(32'h3c077083),
	.w5(32'hb9c86773),
	.w6(32'h3bcda4dd),
	.w7(32'h3c0cd973),
	.w8(32'hbb1026da),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22910e),
	.w1(32'hbb028593),
	.w2(32'hba97326e),
	.w3(32'hbb3c5c3e),
	.w4(32'hbba482b7),
	.w5(32'h3aa4d50c),
	.w6(32'hbb973179),
	.w7(32'hbb83e4b1),
	.w8(32'hb91a74c7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a873),
	.w1(32'hbaad8634),
	.w2(32'h3b72a827),
	.w3(32'h3b3b8f42),
	.w4(32'h3b21b671),
	.w5(32'hbafd2455),
	.w6(32'hba099be3),
	.w7(32'h3b6c44db),
	.w8(32'hbb1f12c8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dbffc),
	.w1(32'hbb678a7c),
	.w2(32'hb929d5cb),
	.w3(32'hbb4ecacd),
	.w4(32'hba175e9a),
	.w5(32'h3a8d5d40),
	.w6(32'hbb827cf7),
	.w7(32'hbb420bc6),
	.w8(32'hb7a6f3fb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fcf94),
	.w1(32'hb98c8a68),
	.w2(32'h3b14ec74),
	.w3(32'h39f90034),
	.w4(32'h3939e074),
	.w5(32'h3af7d918),
	.w6(32'hbb38ca9d),
	.w7(32'hba88a40b),
	.w8(32'hba7d4d59),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba730186),
	.w1(32'hbb209416),
	.w2(32'hba9bfba9),
	.w3(32'hbaa9ca15),
	.w4(32'hbab1cce8),
	.w5(32'hbab362c1),
	.w6(32'hbbf5be32),
	.w7(32'hbbaf9a74),
	.w8(32'hbb986ae4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a8535),
	.w1(32'hbac0cf4c),
	.w2(32'hbbc0e786),
	.w3(32'h3b873982),
	.w4(32'hbb07a9c4),
	.w5(32'hbac4d3a8),
	.w6(32'hbacc52e7),
	.w7(32'hbb69bf09),
	.w8(32'h3a1eabe2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24f94e),
	.w1(32'hba118fb8),
	.w2(32'hbaf23193),
	.w3(32'hbb1b96cf),
	.w4(32'hba893a5c),
	.w5(32'h3ba87849),
	.w6(32'hbb0bc2db),
	.w7(32'hbb2c1833),
	.w8(32'h3b5cff9c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89875e),
	.w1(32'h3ad5dd4c),
	.w2(32'h3a83799f),
	.w3(32'h3ac83125),
	.w4(32'h3b01dae0),
	.w5(32'hbafc1d59),
	.w6(32'hba94c447),
	.w7(32'hba3cf6b9),
	.w8(32'hbb109941),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e926),
	.w1(32'hbba0bc26),
	.w2(32'h3beaef23),
	.w3(32'hbbe0b3e6),
	.w4(32'h3b21f5d7),
	.w5(32'h3c3a3255),
	.w6(32'hbc0c72be),
	.w7(32'h3ab5a7fc),
	.w8(32'h3c01ca81),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc16a01),
	.w1(32'h390f7a9a),
	.w2(32'h3b46b659),
	.w3(32'hbab8a609),
	.w4(32'hbaf78b5f),
	.w5(32'h3afa50e5),
	.w6(32'hbb930985),
	.w7(32'hbb24b7a5),
	.w8(32'h386ce8a4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba240de0),
	.w1(32'hbbc2ad06),
	.w2(32'h3b829b32),
	.w3(32'hbbe06286),
	.w4(32'hba5e09cf),
	.w5(32'hb9feecb1),
	.w6(32'hbc0fcea1),
	.w7(32'h3a7dd804),
	.w8(32'hbb070d8f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f0bf),
	.w1(32'hbb6cde4c),
	.w2(32'hbbacafe4),
	.w3(32'hba8efe23),
	.w4(32'hbb5196fd),
	.w5(32'h3a99abc8),
	.w6(32'hbb26d868),
	.w7(32'hbb39b100),
	.w8(32'h3afe4389),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ba4cb),
	.w1(32'hb9c0a669),
	.w2(32'hba7ed1e8),
	.w3(32'h3a24cdeb),
	.w4(32'hba33b5da),
	.w5(32'h3a4e84db),
	.w6(32'h3ae632e7),
	.w7(32'h39e60572),
	.w8(32'h3b39dc8c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5942e),
	.w1(32'h3ab62bac),
	.w2(32'h3b9452a3),
	.w3(32'h3b6bf0cf),
	.w4(32'h3b9512c0),
	.w5(32'h3a315b3b),
	.w6(32'h3a7fc21f),
	.w7(32'h3be22413),
	.w8(32'h3b5f7e52),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12552),
	.w1(32'hbac34588),
	.w2(32'h37ff2b13),
	.w3(32'h3af9b65f),
	.w4(32'h3b07f2fd),
	.w5(32'hbb2695c6),
	.w6(32'h3b2d85a5),
	.w7(32'hba8a173d),
	.w8(32'hbaf8a421),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba215463),
	.w1(32'h3b34ae53),
	.w2(32'hb824241c),
	.w3(32'h3b5d9ef3),
	.w4(32'h3b894757),
	.w5(32'h39df44ae),
	.w6(32'h3b1ba1b5),
	.w7(32'h3a59c5a5),
	.w8(32'hbb896e2c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb702c82),
	.w1(32'h3b01fe77),
	.w2(32'h3bb9d37b),
	.w3(32'hba4cf8c9),
	.w4(32'h3bb95424),
	.w5(32'hb502c421),
	.w6(32'h3a8a8841),
	.w7(32'h3c129ccc),
	.w8(32'hb68c9b23),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2820e7),
	.w1(32'h3a21da74),
	.w2(32'h3a474854),
	.w3(32'hba2c7267),
	.w4(32'h396c827c),
	.w5(32'h3a8ce7a5),
	.w6(32'hbaa653f4),
	.w7(32'hb952a23e),
	.w8(32'h39a61044),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10b454),
	.w1(32'h3938467e),
	.w2(32'h3a01cd51),
	.w3(32'hb9c71086),
	.w4(32'h3a80f740),
	.w5(32'h3ac993c7),
	.w6(32'hbab7f863),
	.w7(32'hb8959a6f),
	.w8(32'h39be7a68),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ee695),
	.w1(32'hb9abf9c3),
	.w2(32'hb96eda45),
	.w3(32'h38d761c9),
	.w4(32'h3920ffb9),
	.w5(32'h38fa2a9d),
	.w6(32'hb9018c86),
	.w7(32'hb981f073),
	.w8(32'hb8d38c17),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59380e7),
	.w1(32'hb6eea17a),
	.w2(32'hb796b371),
	.w3(32'h36a51886),
	.w4(32'hb6ac475d),
	.w5(32'hb72e3942),
	.w6(32'hb6d13fe6),
	.w7(32'hb77af921),
	.w8(32'hb67e335e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362fdde6),
	.w1(32'h39f7d48a),
	.w2(32'h3b16ff69),
	.w3(32'h3916caf6),
	.w4(32'h3ada6256),
	.w5(32'h3b88b747),
	.w6(32'hbb1fee8a),
	.w7(32'hbb0039ed),
	.w8(32'h3a3749ec),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39821f66),
	.w1(32'h3a7251b4),
	.w2(32'h3a258710),
	.w3(32'h39a36d44),
	.w4(32'h3aa661d5),
	.w5(32'h3a947962),
	.w6(32'hba331c04),
	.w7(32'h38fc3c86),
	.w8(32'h39e232ce),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f28c78),
	.w1(32'h3926d31b),
	.w2(32'h3963b2be),
	.w3(32'h39827fea),
	.w4(32'h3984808e),
	.w5(32'h395e3d73),
	.w6(32'h398ef5a7),
	.w7(32'h39821906),
	.w8(32'h391bd44e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba247ee2),
	.w1(32'h397b6e7a),
	.w2(32'h3a30b89e),
	.w3(32'hba6923ae),
	.w4(32'h39df497f),
	.w5(32'h3a8c893b),
	.w6(32'hbadfd7b8),
	.w7(32'hba3420f0),
	.w8(32'h397b3baf),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb637b404),
	.w1(32'hb674b2ee),
	.w2(32'hb7b4c429),
	.w3(32'hb73551e6),
	.w4(32'hb7565917),
	.w5(32'hb7811026),
	.w6(32'hb7f7e066),
	.w7(32'hb7a7d158),
	.w8(32'hb62b1194),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889f266),
	.w1(32'h38d59a96),
	.w2(32'h3941ad2a),
	.w3(32'hb93f03f0),
	.w4(32'h38861f76),
	.w5(32'h38c3f09b),
	.w6(32'hb93a1954),
	.w7(32'h37b2b9c6),
	.w8(32'h3943061d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6786d5f),
	.w1(32'h3642d5e2),
	.w2(32'hb733e4d7),
	.w3(32'hb74814a7),
	.w4(32'hb726516c),
	.w5(32'hb6c9a90e),
	.w6(32'hb6c723b7),
	.w7(32'hb7369031),
	.w8(32'hb60dfeb8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c1af99),
	.w1(32'h3702fe87),
	.w2(32'hb69db96c),
	.w3(32'hb716ec1e),
	.w4(32'h3675d3bc),
	.w5(32'hb6415537),
	.w6(32'hb7408176),
	.w7(32'h3624e074),
	.w8(32'h35477357),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5b0d5),
	.w1(32'hbad4d5f1),
	.w2(32'hba928d9e),
	.w3(32'hb69a7840),
	.w4(32'hba11ee42),
	.w5(32'h36ec7180),
	.w6(32'h3a1de137),
	.w7(32'h393031eb),
	.w8(32'h3a2f819d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f367a4),
	.w1(32'h3a5d0b58),
	.w2(32'h3ac4904d),
	.w3(32'h3b08f4b9),
	.w4(32'h3b21ed40),
	.w5(32'h3acb3f1c),
	.w6(32'h3afb0f23),
	.w7(32'h3b5bf47e),
	.w8(32'h3b317284),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c76a6c),
	.w1(32'h3a142690),
	.w2(32'h39c8b002),
	.w3(32'h37bc0192),
	.w4(32'h3a8e6e2a),
	.w5(32'h3a804b89),
	.w6(32'hba4ab570),
	.w7(32'h38a0147c),
	.w8(32'h3a0ff5a2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dc4c1),
	.w1(32'h39cf90b3),
	.w2(32'h39fc70ce),
	.w3(32'h39950e58),
	.w4(32'h3aafd218),
	.w5(32'h3a417834),
	.w6(32'hba5583bb),
	.w7(32'h3a4287ba),
	.w8(32'h3a907e13),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8377d0f),
	.w1(32'hb88d54b7),
	.w2(32'hb8616920),
	.w3(32'hb780d576),
	.w4(32'h35388bcc),
	.w5(32'hb7b36a60),
	.w6(32'h37b7a696),
	.w7(32'h3866c492),
	.w8(32'h377fdabe),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902dfe1),
	.w1(32'h3959dc39),
	.w2(32'h38adf0c5),
	.w3(32'h37bda9f2),
	.w4(32'h3927462d),
	.w5(32'h38cf2f6d),
	.w6(32'hb8fe667c),
	.w7(32'hb7d5826d),
	.w8(32'h37f02a80),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36db4a7a),
	.w1(32'h36dbd416),
	.w2(32'h36a8decb),
	.w3(32'h3603b36a),
	.w4(32'h36de1b5d),
	.w5(32'h368060df),
	.w6(32'h36c6a86b),
	.w7(32'h372c9a53),
	.w8(32'hb6e27940),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb735edba),
	.w1(32'h36938d8f),
	.w2(32'hb697d17b),
	.w3(32'h35f31067),
	.w4(32'hb6808af5),
	.w5(32'h378ef14b),
	.w6(32'hb77c54f5),
	.w7(32'hb7dcfff8),
	.w8(32'h35b1ee1b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a576235),
	.w1(32'h3a961559),
	.w2(32'h3aa336b3),
	.w3(32'h3ac1fa95),
	.w4(32'h3aceb3e6),
	.w5(32'h3aa683be),
	.w6(32'hb8842703),
	.w7(32'h39ab0ce8),
	.w8(32'h3a21b5a0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb713dac0),
	.w1(32'hb7368a9e),
	.w2(32'hb7b21434),
	.w3(32'hb747c83b),
	.w4(32'hb7ab812d),
	.w5(32'hb805004d),
	.w6(32'hb6fa03fa),
	.w7(32'hb73df703),
	.w8(32'hb7f42f58),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef7a65),
	.w1(32'h38c291b6),
	.w2(32'h398915eb),
	.w3(32'hb912757e),
	.w4(32'hb84497f0),
	.w5(32'h390f849c),
	.w6(32'hb95b836b),
	.w7(32'hb99c8dde),
	.w8(32'hb8eb4a10),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976c791),
	.w1(32'h3943fde7),
	.w2(32'h39d3f491),
	.w3(32'h3917f35b),
	.w4(32'hb80d6c1b),
	.w5(32'h39a77748),
	.w6(32'h395acc8f),
	.w7(32'hb8245e2b),
	.w8(32'hb903da6f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ae2c1c),
	.w1(32'h35532df7),
	.w2(32'hb709a344),
	.w3(32'h372a7747),
	.w4(32'h355c5f02),
	.w5(32'hb6ac18ad),
	.w6(32'h363d0212),
	.w7(32'hb6fb12d1),
	.w8(32'hb529ff28),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e6cdc),
	.w1(32'h39f23e18),
	.w2(32'h39edbe1c),
	.w3(32'h39b312bd),
	.w4(32'h39e40261),
	.w5(32'h3a09af7b),
	.w6(32'hb9fcf2d6),
	.w7(32'hb9452dba),
	.w8(32'hb8f54cc3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39487ddf),
	.w1(32'h3998dc44),
	.w2(32'h395055e9),
	.w3(32'h392c72d2),
	.w4(32'h393d8872),
	.w5(32'h38cd8526),
	.w6(32'h3922136e),
	.w7(32'h39431d0c),
	.w8(32'h38dca221),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9671580),
	.w1(32'h3a3471bb),
	.w2(32'h3b1f15ed),
	.w3(32'h3b08479a),
	.w4(32'h3ad2fbed),
	.w5(32'h3a863eb8),
	.w6(32'h3aea50e4),
	.w7(32'h3ab6e7d4),
	.w8(32'h3a3995e3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72ada4b),
	.w1(32'h37d7c4e6),
	.w2(32'h3774cdc0),
	.w3(32'h375a50fb),
	.w4(32'h37f36ce9),
	.w5(32'h37d98bde),
	.w6(32'hb832d57c),
	.w7(32'hb815173f),
	.w8(32'hb602a0f4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4a8bf),
	.w1(32'hbadac65c),
	.w2(32'hbb2e6f0b),
	.w3(32'hb99da4e7),
	.w4(32'hba320f1e),
	.w5(32'hb8dca710),
	.w6(32'h39b59b40),
	.w7(32'hb8779b12),
	.w8(32'h39eb6a3b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule