module layer_10_featuremap_226(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0293c3),
	.w1(32'h3b94c152),
	.w2(32'hba73f863),
	.w3(32'hb9630b84),
	.w4(32'hbb1ec336),
	.w5(32'hbc1d714a),
	.w6(32'hbd8ac633),
	.w7(32'hba338ac9),
	.w8(32'h3c03fefa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93cbfd),
	.w1(32'h3b0d66e9),
	.w2(32'h3b9f3f53),
	.w3(32'h3b3c20af),
	.w4(32'hbc5e8de1),
	.w5(32'hbb58ea7c),
	.w6(32'h3b36179a),
	.w7(32'h3b78ad07),
	.w8(32'h3beab219),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1911cd),
	.w1(32'hbb4ccbce),
	.w2(32'hbbdf7a32),
	.w3(32'hbb976431),
	.w4(32'h3cf63e8b),
	.w5(32'h3ba67d63),
	.w6(32'h3b044495),
	.w7(32'hbba6775f),
	.w8(32'h3b28b968),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad77a5f),
	.w1(32'h3cc7d30e),
	.w2(32'h3b791b8d),
	.w3(32'hbcae29d8),
	.w4(32'h3c7ba292),
	.w5(32'h3b2084e9),
	.w6(32'h3bc01ca3),
	.w7(32'h3b065bfd),
	.w8(32'h3b133c9a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf215c3),
	.w1(32'hbc4a3ecf),
	.w2(32'hbb7ab3b3),
	.w3(32'hbb869e9a),
	.w4(32'h3c171822),
	.w5(32'hba6b68c7),
	.w6(32'hbc43d6a8),
	.w7(32'h3a29a76f),
	.w8(32'h3cfde813),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbf8ac),
	.w1(32'hbbc28556),
	.w2(32'hbab25be9),
	.w3(32'h3b671e5b),
	.w4(32'hbb1dd3b3),
	.w5(32'hba3cd6ee),
	.w6(32'h3c0b9d7b),
	.w7(32'hbacae0cd),
	.w8(32'h3c35a91d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51150d),
	.w1(32'h3b2ef49e),
	.w2(32'hbb85a5d3),
	.w3(32'hbbb5d789),
	.w4(32'hbb14a7c3),
	.w5(32'h3c41ffe6),
	.w6(32'h3abad6cc),
	.w7(32'hbb66a159),
	.w8(32'hbbd92dd7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdebf3f),
	.w1(32'h3c094348),
	.w2(32'h3ab13e88),
	.w3(32'hbb996962),
	.w4(32'h3a40a400),
	.w5(32'hbb480cb9),
	.w6(32'hbc403b47),
	.w7(32'h3c56ad43),
	.w8(32'hbb8f8dca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bdd67),
	.w1(32'hbc855145),
	.w2(32'h3ba36d4c),
	.w3(32'hbb4c83bd),
	.w4(32'hbb356362),
	.w5(32'h3b1e6737),
	.w6(32'h3ba57715),
	.w7(32'hb9140e4d),
	.w8(32'hbb41bc92),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6822e),
	.w1(32'h3af81e42),
	.w2(32'h3c01fa61),
	.w3(32'hbb6ef622),
	.w4(32'hbbccf869),
	.w5(32'h3b874593),
	.w6(32'h3d10a1fb),
	.w7(32'hbc810870),
	.w8(32'h3bf2ca94),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8077),
	.w1(32'h3c04db3c),
	.w2(32'h390ce685),
	.w3(32'hbc43bb94),
	.w4(32'h3b44661d),
	.w5(32'hbc79e4d7),
	.w6(32'h3c249644),
	.w7(32'hbafe7af3),
	.w8(32'h3afd634e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d9625),
	.w1(32'hbb5a76ed),
	.w2(32'h3c8aeebb),
	.w3(32'hbbd669ac),
	.w4(32'h3c1e2e2b),
	.w5(32'hbb2faa2a),
	.w6(32'hbb0f28cd),
	.w7(32'hb99c80c2),
	.w8(32'h3c444aaa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd3d7c),
	.w1(32'hbbc455cb),
	.w2(32'h3c0601b7),
	.w3(32'hbb83e97c),
	.w4(32'hba9c2b96),
	.w5(32'h3c50f3ed),
	.w6(32'hbbfefe28),
	.w7(32'h3c499e22),
	.w8(32'hba6ea470),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1aa9f),
	.w1(32'h3c1c4561),
	.w2(32'hbbeae166),
	.w3(32'hbbb80233),
	.w4(32'hbb2507c9),
	.w5(32'hbc903732),
	.w6(32'h3c3e34ff),
	.w7(32'h3bb2d703),
	.w8(32'hbb9a3723),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67b736),
	.w1(32'hbbbaf508),
	.w2(32'hbafd7520),
	.w3(32'h3ba20bad),
	.w4(32'h3b7a0666),
	.w5(32'h3c016460),
	.w6(32'hbb792aaf),
	.w7(32'h3b28d1d7),
	.w8(32'h3b9fec82),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41ac12),
	.w1(32'hb99a522c),
	.w2(32'hbbae7058),
	.w3(32'h3c8de3c5),
	.w4(32'h3b9b2f09),
	.w5(32'h3a847abf),
	.w6(32'h3c212f46),
	.w7(32'hbbe0c456),
	.w8(32'hbc8c8a2c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffea48),
	.w1(32'h3bfae7ad),
	.w2(32'hbb70bf6f),
	.w3(32'h3b1cdbaa),
	.w4(32'hba0e966c),
	.w5(32'hbba2e844),
	.w6(32'hba978b5d),
	.w7(32'hbbf5b1a9),
	.w8(32'hbb881d1e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b1cd4),
	.w1(32'h3cb21d20),
	.w2(32'hbcbd6417),
	.w3(32'h3a9051d1),
	.w4(32'hbb8cbe0a),
	.w5(32'h3a667da6),
	.w6(32'hbb2a4bdf),
	.w7(32'h3c1a328a),
	.w8(32'h3af6b4a9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6ee38),
	.w1(32'hbc466b67),
	.w2(32'hbc00fcbb),
	.w3(32'hbb9b81aa),
	.w4(32'h3aeb73f5),
	.w5(32'hbc2b84ad),
	.w6(32'hbc452dff),
	.w7(32'h3b9d2854),
	.w8(32'hbbc32319),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b382681),
	.w1(32'hbaa988e2),
	.w2(32'hbc001c94),
	.w3(32'hbb5ec8af),
	.w4(32'hbb76fbdd),
	.w5(32'hbbef3407),
	.w6(32'h3b538a62),
	.w7(32'hbc2c8451),
	.w8(32'h3bbebb1b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4557a9),
	.w1(32'hbaed81ab),
	.w2(32'hbc77cf81),
	.w3(32'h3bafa8e0),
	.w4(32'hbb55fc88),
	.w5(32'h3b075e5d),
	.w6(32'h3c49af34),
	.w7(32'hbad63379),
	.w8(32'h3c9c952e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8a201),
	.w1(32'hbbc5b51e),
	.w2(32'hbbc43f25),
	.w3(32'h3a246d57),
	.w4(32'h387b478c),
	.w5(32'hbaf23789),
	.w6(32'h396a71e5),
	.w7(32'hb9f19803),
	.w8(32'hbbceedb3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904463),
	.w1(32'hba46f42e),
	.w2(32'h39e28f7d),
	.w3(32'hb901b30b),
	.w4(32'h3b0f02de),
	.w5(32'h3d1dc61f),
	.w6(32'h3899e625),
	.w7(32'hbb97c0e4),
	.w8(32'hba43c7b2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935e93a),
	.w1(32'hbb9f153f),
	.w2(32'hbb20bcb4),
	.w3(32'h3b27292e),
	.w4(32'hba844542),
	.w5(32'h3ad91584),
	.w6(32'h3b43d6fc),
	.w7(32'hbba5fd7f),
	.w8(32'hbab36e82),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49f37a),
	.w1(32'hbbab0fa6),
	.w2(32'hbc062405),
	.w3(32'hbb669b2a),
	.w4(32'hbad05efe),
	.w5(32'h3bb17db6),
	.w6(32'h3aebc04c),
	.w7(32'hbc0ab548),
	.w8(32'h3cce3bce),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d844f),
	.w1(32'h3c438635),
	.w2(32'hbb916a10),
	.w3(32'h3b0dc100),
	.w4(32'h3cac147c),
	.w5(32'h3b525fe9),
	.w6(32'hbb432b9d),
	.w7(32'hbb99f5a3),
	.w8(32'h3a9d3600),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8be8b9),
	.w1(32'h3cb153a4),
	.w2(32'h3bd57cf1),
	.w3(32'h3c04fec8),
	.w4(32'h3b94541e),
	.w5(32'hb9a11d81),
	.w6(32'h3b2b9bd3),
	.w7(32'hbba90d27),
	.w8(32'h39dfb537),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8b427),
	.w1(32'h3c430802),
	.w2(32'hba11e5e5),
	.w3(32'h3b0c4364),
	.w4(32'hba1392c5),
	.w5(32'h3b343518),
	.w6(32'h3c6ac149),
	.w7(32'h3b9965ad),
	.w8(32'h3bd481fe),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77f914),
	.w1(32'h3c42a777),
	.w2(32'hbb64c64f),
	.w3(32'h3a836f1b),
	.w4(32'h3b9281d4),
	.w5(32'h3c796d67),
	.w6(32'hba04ca19),
	.w7(32'hbb4332dc),
	.w8(32'h3c264a55),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7455cd),
	.w1(32'h3bf8c047),
	.w2(32'hbb16af07),
	.w3(32'hbb0b4b63),
	.w4(32'hbbc449f0),
	.w5(32'h3b975b8d),
	.w6(32'h3c301040),
	.w7(32'hbbeb3a78),
	.w8(32'h3c466459),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4754),
	.w1(32'h3a4291b4),
	.w2(32'h383cb9ab),
	.w3(32'hba5f9a0a),
	.w4(32'h3c0a4811),
	.w5(32'h3b6e9b66),
	.w6(32'h3bbe6c12),
	.w7(32'hbb4ba656),
	.w8(32'h3b1905e5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc32f1),
	.w1(32'h3b418d39),
	.w2(32'hba8401b9),
	.w3(32'h3c5deaab),
	.w4(32'h3a94c09f),
	.w5(32'hbc0a368b),
	.w6(32'h3bf58293),
	.w7(32'hba0a2351),
	.w8(32'h3a3910bf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8875f8),
	.w1(32'h3cb0c1c5),
	.w2(32'hbc219c31),
	.w3(32'h3ba8dc6e),
	.w4(32'h3b896496),
	.w5(32'h3ac818ec),
	.w6(32'hbbd927e3),
	.w7(32'h3b7e040c),
	.w8(32'hbab8449c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14984c),
	.w1(32'h3b53477d),
	.w2(32'hb9bdce47),
	.w3(32'h3be69358),
	.w4(32'h3c867c4e),
	.w5(32'hbbc1fc32),
	.w6(32'hb7a7463c),
	.w7(32'h3c584725),
	.w8(32'hba4a9e5c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44b47b),
	.w1(32'hbbaa2396),
	.w2(32'h3b941220),
	.w3(32'h3b6ac998),
	.w4(32'hbadb8c4e),
	.w5(32'h3a9db6f9),
	.w6(32'h3c6c6ed1),
	.w7(32'hbc6be170),
	.w8(32'h3a656d74),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2292e),
	.w1(32'h3b77f54b),
	.w2(32'h3bada52b),
	.w3(32'hbb80fc02),
	.w4(32'hbcaa44c3),
	.w5(32'h3c8653b4),
	.w6(32'hba8cb276),
	.w7(32'hbc08c62d),
	.w8(32'h3c671399),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b8e6),
	.w1(32'h3bfd90d4),
	.w2(32'hbb91f67a),
	.w3(32'h3b8a8093),
	.w4(32'h3bc741d5),
	.w5(32'h3c1833b5),
	.w6(32'h3b90cbf5),
	.w7(32'h3c68ea91),
	.w8(32'hbc846288),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93529e3),
	.w1(32'hb9ff7678),
	.w2(32'h3be0e86e),
	.w3(32'hbb531d3a),
	.w4(32'h3a9d625e),
	.w5(32'h3aafcdef),
	.w6(32'h3aaa1034),
	.w7(32'h3bcd5562),
	.w8(32'h3c33b4c9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b8aa2),
	.w1(32'hbb94fc3a),
	.w2(32'hbb2d19cb),
	.w3(32'hbb929e38),
	.w4(32'h3b84d0cf),
	.w5(32'hba86f1ea),
	.w6(32'hbbf730c8),
	.w7(32'h3b22ec95),
	.w8(32'h3c29c60e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6641e1),
	.w1(32'h3a644b16),
	.w2(32'hbb2d6325),
	.w3(32'h3a889efa),
	.w4(32'h3b25e65c),
	.w5(32'hbc194280),
	.w6(32'hbb7517d6),
	.w7(32'h3afd56a3),
	.w8(32'h3b1fb5b7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a812546),
	.w1(32'h3b947256),
	.w2(32'h3a911f33),
	.w3(32'h3ad1d357),
	.w4(32'hba703d89),
	.w5(32'h3c42dcf6),
	.w6(32'h3ae47f18),
	.w7(32'h3b358cc6),
	.w8(32'hbb0ac063),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b651872),
	.w1(32'hba99d7c0),
	.w2(32'hbc58668d),
	.w3(32'h3ba95472),
	.w4(32'hbade724e),
	.w5(32'h3b1465f5),
	.w6(32'h3b38972b),
	.w7(32'h3c21257a),
	.w8(32'h3c2ca447),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa44449),
	.w1(32'h3b7e5e99),
	.w2(32'hbc2e40e1),
	.w3(32'hb93d4bae),
	.w4(32'hbbf75ecd),
	.w5(32'hbb23ec52),
	.w6(32'hbb4272f0),
	.w7(32'hba0c7de3),
	.w8(32'hba5af21b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ae954),
	.w1(32'hbac52e72),
	.w2(32'hba68ab17),
	.w3(32'h3b0a7d3a),
	.w4(32'h3ae760a4),
	.w5(32'h3aa66d1a),
	.w6(32'hbb74657e),
	.w7(32'hbb86ed9d),
	.w8(32'h3a12197d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c716adb),
	.w1(32'h38d6426e),
	.w2(32'h3b73cc4a),
	.w3(32'h3a23c392),
	.w4(32'h3b701727),
	.w5(32'h3c0765a2),
	.w6(32'hbbdf0b43),
	.w7(32'hbb01a410),
	.w8(32'hba852d2b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c705d2c),
	.w1(32'hba7487d7),
	.w2(32'hbb8b549f),
	.w3(32'h3bf8a2d7),
	.w4(32'h3c04244b),
	.w5(32'hbbabb85a),
	.w6(32'hba1316b2),
	.w7(32'h3b8cae1f),
	.w8(32'hbaa7fcef),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48e7e),
	.w1(32'h3bab79ad),
	.w2(32'h3ba832f3),
	.w3(32'h3b263023),
	.w4(32'hbb32688f),
	.w5(32'hbc45ffbb),
	.w6(32'h3ab5eb42),
	.w7(32'h3af13839),
	.w8(32'hbc2ea0bd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d5d6f),
	.w1(32'h3c7cfe0c),
	.w2(32'h3b961976),
	.w3(32'hbac2f89e),
	.w4(32'hbae368c4),
	.w5(32'hbb6b12bb),
	.w6(32'hbb722d5f),
	.w7(32'h3be99fc1),
	.w8(32'h3b7926b4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50b62),
	.w1(32'h3aa1026c),
	.w2(32'hbb439176),
	.w3(32'h3bccd30f),
	.w4(32'h38d02197),
	.w5(32'h3c0be692),
	.w6(32'hbadb365b),
	.w7(32'hbaaea76f),
	.w8(32'h3a03d0de),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2050d2),
	.w1(32'hbbcc5aaa),
	.w2(32'hbc1c2788),
	.w3(32'hbc01a137),
	.w4(32'h3b93a25b),
	.w5(32'hbb352d3e),
	.w6(32'h3b286ff5),
	.w7(32'h3ad565e5),
	.w8(32'h3bab2eb9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75122f),
	.w1(32'hb9be51ce),
	.w2(32'h3b634c27),
	.w3(32'h3bb71211),
	.w4(32'hbaa28ee1),
	.w5(32'hb7018e23),
	.w6(32'hba3f23c7),
	.w7(32'h3bc7de2d),
	.w8(32'h3964f203),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba20697),
	.w1(32'h3c08f676),
	.w2(32'hbb182cc2),
	.w3(32'hbbdb6849),
	.w4(32'h3bf611b2),
	.w5(32'hbaccc01d),
	.w6(32'hbc3a224b),
	.w7(32'h3badd2d7),
	.w8(32'hbb84b255),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04974a),
	.w1(32'h3c0233b1),
	.w2(32'hbb872fed),
	.w3(32'h3ba288a5),
	.w4(32'hb995921d),
	.w5(32'hbbaa80c4),
	.w6(32'h3a7e133a),
	.w7(32'h3c20a2ac),
	.w8(32'hbb54c6ea),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f8f7c),
	.w1(32'hbc08fd74),
	.w2(32'h3b0465fc),
	.w3(32'hb9e1c6b7),
	.w4(32'hbc001058),
	.w5(32'hbb005a5b),
	.w6(32'hb8eb37ca),
	.w7(32'hbae606a2),
	.w8(32'hbd733a9d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807aa7),
	.w1(32'h3c164c5a),
	.w2(32'h3b67798e),
	.w3(32'hbc2c5780),
	.w4(32'h3d199b10),
	.w5(32'hb9061395),
	.w6(32'h3c7b5efa),
	.w7(32'h3a8ebe63),
	.w8(32'hbb1ebf59),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee00e4),
	.w1(32'h3b68e845),
	.w2(32'h3b8069d8),
	.w3(32'hbae6aef8),
	.w4(32'h3bb19819),
	.w5(32'h3a6c8a86),
	.w6(32'hbafa9c14),
	.w7(32'h3ab7ee3c),
	.w8(32'h3b5bc37b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5a5e8),
	.w1(32'h3ae9d198),
	.w2(32'h3c2a0b66),
	.w3(32'h3b176c53),
	.w4(32'h3ba7e0f8),
	.w5(32'hbbe41805),
	.w6(32'h3aa6cd20),
	.w7(32'hba460477),
	.w8(32'h3bc2499e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13bc3d),
	.w1(32'hbb70ac43),
	.w2(32'h3a20b124),
	.w3(32'hbbe02ad8),
	.w4(32'h3ab0ac00),
	.w5(32'hb92e1262),
	.w6(32'hbb398f05),
	.w7(32'h3a38a4be),
	.w8(32'h3a1454bf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecb777),
	.w1(32'h3c95fa24),
	.w2(32'hbac1ffb7),
	.w3(32'hbb8ae784),
	.w4(32'hbad454a4),
	.w5(32'hbb2d1e0e),
	.w6(32'h3d0328aa),
	.w7(32'hba507024),
	.w8(32'h3c567ed5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b510a),
	.w1(32'h3bb92839),
	.w2(32'hbb5aa1ba),
	.w3(32'hbad6d279),
	.w4(32'h3a20d1a1),
	.w5(32'hbc1781df),
	.w6(32'h3af80a7b),
	.w7(32'h3aed1327),
	.w8(32'hbbd91611),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf55cfd),
	.w1(32'hbafeb4c8),
	.w2(32'h3bf9e4dc),
	.w3(32'hbb8eb483),
	.w4(32'h3bf4bd39),
	.w5(32'h3b9d2bc0),
	.w6(32'h3c142eb3),
	.w7(32'hbc0274a6),
	.w8(32'h3bae801d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c003c17),
	.w1(32'h3afe88de),
	.w2(32'hb89228f5),
	.w3(32'h3c1063d6),
	.w4(32'hbb1f7149),
	.w5(32'h3cbbe219),
	.w6(32'h3cd1f606),
	.w7(32'hbab5c2a0),
	.w8(32'h3b4e220d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01b220),
	.w1(32'h3ad038c6),
	.w2(32'h3cce598c),
	.w3(32'h39d14733),
	.w4(32'hbb53e2df),
	.w5(32'hbad62f81),
	.w6(32'h3b9f4e68),
	.w7(32'h3b2d45ba),
	.w8(32'hb90a63db),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc39097),
	.w1(32'hbc3777d3),
	.w2(32'hbbe75a69),
	.w3(32'h3bffd674),
	.w4(32'hbbacf70a),
	.w5(32'hbc048074),
	.w6(32'hbcce0a77),
	.w7(32'h3b5214d7),
	.w8(32'h3b175deb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf140a9),
	.w1(32'h383a658b),
	.w2(32'hbb14e917),
	.w3(32'h3b8cc412),
	.w4(32'hba9d26bd),
	.w5(32'hbbbaeccd),
	.w6(32'h3ba156a3),
	.w7(32'hbb301505),
	.w8(32'h3a860bc9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b01f9),
	.w1(32'hbbf47f06),
	.w2(32'h3b1a9492),
	.w3(32'h3c1f7f96),
	.w4(32'hbbe2bfb2),
	.w5(32'h3a431205),
	.w6(32'hbc47d3e7),
	.w7(32'hbb88e8c3),
	.w8(32'hbb13d2bf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4287a),
	.w1(32'h3b397a16),
	.w2(32'h397d61b3),
	.w3(32'h3c5d7037),
	.w4(32'h3b721550),
	.w5(32'hb9e7709b),
	.w6(32'h38fd86e3),
	.w7(32'hbc578e65),
	.w8(32'h3ba521a2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c49eb),
	.w1(32'hbb630b7e),
	.w2(32'h3bac0e6b),
	.w3(32'hbb845dbd),
	.w4(32'h3ab0035e),
	.w5(32'hbc0f242d),
	.w6(32'hbb395e43),
	.w7(32'hb9e77394),
	.w8(32'hbb728afc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01e1ce),
	.w1(32'hba3855d9),
	.w2(32'h3a802750),
	.w3(32'hbaf7dcb6),
	.w4(32'hba265da5),
	.w5(32'hbbb73edb),
	.w6(32'h3b7adadf),
	.w7(32'h3acdbff4),
	.w8(32'h3a753810),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc4558),
	.w1(32'hb9a739ec),
	.w2(32'h3b801254),
	.w3(32'h3bd53da4),
	.w4(32'h3c5d7ac4),
	.w5(32'hbb87025c),
	.w6(32'h3c17a907),
	.w7(32'h3c866dc0),
	.w8(32'h380f2265),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06dac4),
	.w1(32'hba7b1689),
	.w2(32'h3c31ac25),
	.w3(32'h3c0b81ff),
	.w4(32'h3b9534c8),
	.w5(32'h3bf58b23),
	.w6(32'h3b0b536e),
	.w7(32'h3bc7331e),
	.w8(32'h3b9eb554),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45534c),
	.w1(32'hbb360d12),
	.w2(32'h3b78254b),
	.w3(32'hbbd2f219),
	.w4(32'h3bad3ab0),
	.w5(32'h3aba3748),
	.w6(32'h3c73582d),
	.w7(32'h39d64c7f),
	.w8(32'h3bfb9406),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc435cab),
	.w1(32'h3ac7cbb8),
	.w2(32'hba073e01),
	.w3(32'h3bb7d0d0),
	.w4(32'h3b391244),
	.w5(32'h3a09544b),
	.w6(32'h3b8dec1c),
	.w7(32'hbbca7c62),
	.w8(32'h3a3d75cb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71c2eb),
	.w1(32'h37b99ded),
	.w2(32'h3ac09551),
	.w3(32'h3bb449e8),
	.w4(32'hba8b1478),
	.w5(32'h3b219851),
	.w6(32'h36a6fa6b),
	.w7(32'h3b8f4a69),
	.w8(32'h3c4f1f0e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9649de),
	.w1(32'h3a51ec65),
	.w2(32'h3795ebd1),
	.w3(32'hbbfb15ad),
	.w4(32'h3b029ad5),
	.w5(32'h3b9fe9b1),
	.w6(32'hbc6b4612),
	.w7(32'hbc76e074),
	.w8(32'h3b8a3f15),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae2b37),
	.w1(32'h3b948a57),
	.w2(32'h3b252c00),
	.w3(32'h3bb171ef),
	.w4(32'h3c8d5832),
	.w5(32'h3ad8a13a),
	.w6(32'h3c1be02c),
	.w7(32'h3c14aa85),
	.w8(32'hbb40b8d9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170b17),
	.w1(32'hbb83af09),
	.w2(32'hbb27e8bd),
	.w3(32'hbb8565c9),
	.w4(32'hbb46a6e5),
	.w5(32'h3c5fde7d),
	.w6(32'h3ac74039),
	.w7(32'h3ad4a31d),
	.w8(32'hbbe85d48),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4938c1),
	.w1(32'hba0dc14f),
	.w2(32'hbbf56375),
	.w3(32'hbbffce3b),
	.w4(32'h37c3bc54),
	.w5(32'hba830e1c),
	.w6(32'h3b7e9b68),
	.w7(32'h3ba72bd6),
	.w8(32'hbbbc711a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c34d1),
	.w1(32'h3a7f11f4),
	.w2(32'h3ac043e5),
	.w3(32'h3ae66871),
	.w4(32'h397c00db),
	.w5(32'h3bb9f795),
	.w6(32'hbb898690),
	.w7(32'hba9e66e3),
	.w8(32'hba2dc848),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6036e),
	.w1(32'h3a005113),
	.w2(32'h3b6fb97c),
	.w3(32'hb9dfd440),
	.w4(32'h3a4c2585),
	.w5(32'h3bd420cb),
	.w6(32'hba135e95),
	.w7(32'h3c025e08),
	.w8(32'h3ad49bee),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab053d3),
	.w1(32'h3bde95ac),
	.w2(32'h3bb613dd),
	.w3(32'h3aa8f74a),
	.w4(32'h3acc3652),
	.w5(32'hbb63f553),
	.w6(32'hb94bdfd5),
	.w7(32'h3b0b19b6),
	.w8(32'hbc04dcee),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b355dd6),
	.w1(32'hbbb6b994),
	.w2(32'h3b261fc0),
	.w3(32'hb87f2622),
	.w4(32'h3c00e097),
	.w5(32'h3bef84a6),
	.w6(32'h3c83fcfa),
	.w7(32'h3b68d454),
	.w8(32'h3bbcbd51),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a47c),
	.w1(32'h3bc13016),
	.w2(32'hbb162429),
	.w3(32'h3b723881),
	.w4(32'h3aa2c3fe),
	.w5(32'h3b6f5f7f),
	.w6(32'h3b997f8a),
	.w7(32'hbbb82802),
	.w8(32'h3cae6338),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb077458),
	.w1(32'h3bdecb5a),
	.w2(32'hbb9c563c),
	.w3(32'h3bed2a9c),
	.w4(32'hbb16861f),
	.w5(32'h3b2f66d4),
	.w6(32'hba9cf462),
	.w7(32'h3bb7b317),
	.w8(32'hbb820f4e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad67d7),
	.w1(32'h3c8658a8),
	.w2(32'hbbd19610),
	.w3(32'hbb40e9e2),
	.w4(32'h3bea7881),
	.w5(32'h3bd92a4f),
	.w6(32'hb9428c6c),
	.w7(32'hbb9c4433),
	.w8(32'h3c25fe3c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9df419),
	.w1(32'h3ba59310),
	.w2(32'hb99eb0ca),
	.w3(32'hb9b57dfd),
	.w4(32'h3aa688e9),
	.w5(32'h38f16361),
	.w6(32'hbc022678),
	.w7(32'hbb3b7a0f),
	.w8(32'h3c148439),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9e15d),
	.w1(32'h3bd8e313),
	.w2(32'hbaaefb6a),
	.w3(32'hbb2da34c),
	.w4(32'hbc684299),
	.w5(32'hbac7b406),
	.w6(32'h3b4c08c9),
	.w7(32'h3c37e2ce),
	.w8(32'h3c3c306e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bbd85),
	.w1(32'hbb5777b0),
	.w2(32'h3b2499e0),
	.w3(32'h3c29af37),
	.w4(32'hbb20a684),
	.w5(32'h3c47e52f),
	.w6(32'h3bc154b5),
	.w7(32'h3c309359),
	.w8(32'hbb0fff9b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1e9a0),
	.w1(32'hbb36972e),
	.w2(32'hbb918255),
	.w3(32'h3c2c5cdc),
	.w4(32'h3a52b4b0),
	.w5(32'h3a9ba19f),
	.w6(32'h3b866a9f),
	.w7(32'hbc07ee4d),
	.w8(32'h3b6c4eaf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c076213),
	.w1(32'h38119768),
	.w2(32'h3b0e5c33),
	.w3(32'h3c3d4e13),
	.w4(32'h3b46f490),
	.w5(32'hbc03d8b7),
	.w6(32'h3cca20de),
	.w7(32'hbc3009cb),
	.w8(32'hbb66b8bf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60c908),
	.w1(32'h3bc8d85c),
	.w2(32'hbbecdb56),
	.w3(32'hba27e189),
	.w4(32'h3ba1fc01),
	.w5(32'h3acbdc94),
	.w6(32'hbb81d379),
	.w7(32'hba41ffe5),
	.w8(32'h3c0b9e0e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3e8fd),
	.w1(32'h3a234cd0),
	.w2(32'hbcfd222f),
	.w3(32'h3c801e41),
	.w4(32'hbbcd936b),
	.w5(32'h3bedcd99),
	.w6(32'hbbaae7ea),
	.w7(32'h3c9c3908),
	.w8(32'hbbcf3f88),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfe8a7),
	.w1(32'h3c8bf54b),
	.w2(32'h3b53c955),
	.w3(32'hba13d3ed),
	.w4(32'h3a702826),
	.w5(32'hba11679a),
	.w6(32'h3c2e159c),
	.w7(32'hba7e7458),
	.w8(32'hbc446207),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3148c),
	.w1(32'h3bb6de18),
	.w2(32'hbc260611),
	.w3(32'hb9ab0d87),
	.w4(32'h3c04c2ca),
	.w5(32'hbc0983c3),
	.w6(32'h3a905f2a),
	.w7(32'hbad8081b),
	.w8(32'hb9c0fd54),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50d76),
	.w1(32'hb814651a),
	.w2(32'h3a225244),
	.w3(32'h3c218422),
	.w4(32'hbaab513e),
	.w5(32'h3bad0612),
	.w6(32'h3a07247c),
	.w7(32'hba11b5ed),
	.w8(32'h3c03149d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc946614),
	.w1(32'hbb42ace5),
	.w2(32'hbb7dd41d),
	.w3(32'h3b1ee9fa),
	.w4(32'hbb363e11),
	.w5(32'h3b9a271f),
	.w6(32'h3b9ae265),
	.w7(32'hbc71ec3a),
	.w8(32'h3bb88319),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b188f04),
	.w1(32'h3b48dcc1),
	.w2(32'hbb2c5a4c),
	.w3(32'hbb4e15f3),
	.w4(32'hbc2c5a2c),
	.w5(32'h3c281f57),
	.w6(32'hbc10b060),
	.w7(32'h36a7adc2),
	.w8(32'hbadaee7f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1ce8b),
	.w1(32'hbbf748bc),
	.w2(32'hbb8bcf4e),
	.w3(32'hbb9a21cb),
	.w4(32'hbaa91a6a),
	.w5(32'h39d52ece),
	.w6(32'hbc87d5b5),
	.w7(32'h3c56df83),
	.w8(32'h3c57dbe9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc532a1),
	.w1(32'h3b1eccff),
	.w2(32'hbbfd1d3f),
	.w3(32'h3b7976f7),
	.w4(32'h3aabbaad),
	.w5(32'hbb5ead43),
	.w6(32'h3b09ccd3),
	.w7(32'hbbc7d9f8),
	.w8(32'h3bc8605c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc935816),
	.w1(32'h3914692a),
	.w2(32'hb9ad5d3b),
	.w3(32'h3b7114db),
	.w4(32'h3abfbb3b),
	.w5(32'hbaf92949),
	.w6(32'h3c2f2737),
	.w7(32'h3b5f65c0),
	.w8(32'hbc02db6e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5f2f3),
	.w1(32'h393023a2),
	.w2(32'hbb844365),
	.w3(32'hbc201b9b),
	.w4(32'hbb0a073c),
	.w5(32'h3b483edb),
	.w6(32'h3bbe8075),
	.w7(32'hba9fb643),
	.w8(32'hbbab9b72),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a349f58),
	.w1(32'h3b30d07a),
	.w2(32'h3c10cfa7),
	.w3(32'h3ae87966),
	.w4(32'hbb44a71a),
	.w5(32'hba87c78a),
	.w6(32'h3bf66f7c),
	.w7(32'h3a95954c),
	.w8(32'h3c2d4ea0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f1a28),
	.w1(32'h3b68dd17),
	.w2(32'hbbe58e9f),
	.w3(32'hba9a32d7),
	.w4(32'h3bc38305),
	.w5(32'h3be0d9e4),
	.w6(32'hba827df6),
	.w7(32'hbc7719c1),
	.w8(32'hbbc15cd2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e0db),
	.w1(32'hbc031588),
	.w2(32'h3b6576c7),
	.w3(32'hbb1f07ce),
	.w4(32'hbbcfc118),
	.w5(32'h399d3924),
	.w6(32'h3bc40cbd),
	.w7(32'h3af8872a),
	.w8(32'h3b4ba99f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e829),
	.w1(32'hba4815c0),
	.w2(32'h3bd53113),
	.w3(32'hbbba93ac),
	.w4(32'hbba82d58),
	.w5(32'h3b7f8bdf),
	.w6(32'hbaf183bb),
	.w7(32'hbb182874),
	.w8(32'h39a3b1b3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba386b9e),
	.w1(32'hbc66e950),
	.w2(32'h3ade299d),
	.w3(32'h3b692fc4),
	.w4(32'hba3a70f0),
	.w5(32'h3b2a6fe6),
	.w6(32'h3c095226),
	.w7(32'hbac4e70c),
	.w8(32'h3a507f1b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94d2d7),
	.w1(32'h3c1bd905),
	.w2(32'h3b013455),
	.w3(32'hbc6042e9),
	.w4(32'hb568fd83),
	.w5(32'hb7244055),
	.w6(32'hbb750a50),
	.w7(32'hbae8da26),
	.w8(32'hb9b08bf2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5e67),
	.w1(32'hbabd46f0),
	.w2(32'hb9056183),
	.w3(32'h3a4d33df),
	.w4(32'h3a4f8417),
	.w5(32'h3b80e82a),
	.w6(32'h3bd278b6),
	.w7(32'hbaf23074),
	.w8(32'hbc0992d0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1010fe),
	.w1(32'hbbca9728),
	.w2(32'h3c4c7ec4),
	.w3(32'hb9a0e924),
	.w4(32'h3c46d726),
	.w5(32'hbbc669e0),
	.w6(32'h3b4f763f),
	.w7(32'hbb5ecc9f),
	.w8(32'h3a7ea0ff),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb098a),
	.w1(32'h3b518c94),
	.w2(32'h3b671a39),
	.w3(32'h3c2f6431),
	.w4(32'h3b080525),
	.w5(32'h3b7b1b72),
	.w6(32'hbb49b9b4),
	.w7(32'h3a6af8c7),
	.w8(32'h3c6c83e3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906be1),
	.w1(32'hbb80ab22),
	.w2(32'h3d0dca91),
	.w3(32'hbadf6503),
	.w4(32'h3b5092ff),
	.w5(32'hbc9a3122),
	.w6(32'hbb5857b5),
	.w7(32'h3ba0e958),
	.w8(32'h3b2b65cd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45ce10),
	.w1(32'h3d0243e9),
	.w2(32'h3ada3742),
	.w3(32'h3bcb32a0),
	.w4(32'h3bad8ccc),
	.w5(32'h3aacf7ee),
	.w6(32'h3c582605),
	.w7(32'h3c5144d2),
	.w8(32'hbc12a9fa),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acad7d6),
	.w1(32'hbb93c60c),
	.w2(32'hbb84d472),
	.w3(32'h38bfb3a4),
	.w4(32'h39bfd986),
	.w5(32'h3c35678f),
	.w6(32'h3a189ea3),
	.w7(32'h3996b770),
	.w8(32'hbb1026f6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1468),
	.w1(32'h3a104930),
	.w2(32'hba8b2e27),
	.w3(32'hbbd5cacc),
	.w4(32'hb9805e28),
	.w5(32'hbb81a71b),
	.w6(32'h3b1a3817),
	.w7(32'h3c4be6c2),
	.w8(32'h3ba22d1e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3ef57),
	.w1(32'hb9a8ea91),
	.w2(32'hbba42933),
	.w3(32'hbaa9eac3),
	.w4(32'h3bae3a45),
	.w5(32'h3a538a72),
	.w6(32'h39d20acf),
	.w7(32'hbcca3e3e),
	.w8(32'h3bcbd27a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf176c),
	.w1(32'h3ba3e50e),
	.w2(32'hbba516fe),
	.w3(32'h3ba06b01),
	.w4(32'hbc04c01a),
	.w5(32'h39e6357a),
	.w6(32'h3b0bda46),
	.w7(32'hbbe30390),
	.w8(32'h3b1f192c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8766ee),
	.w1(32'h3a243eff),
	.w2(32'hbb2fc39e),
	.w3(32'hbbfafa5f),
	.w4(32'hbaf57b6c),
	.w5(32'h3c8430da),
	.w6(32'hbb88758b),
	.w7(32'h3b017f10),
	.w8(32'h3c027fdc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b2dc1),
	.w1(32'h3b6aeb14),
	.w2(32'hbbd0b77e),
	.w3(32'hbbc22d35),
	.w4(32'h3b89f628),
	.w5(32'h3c2da411),
	.w6(32'h3b834e3f),
	.w7(32'h3b939c9c),
	.w8(32'h3c0b00f1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00442b),
	.w1(32'h3ae49336),
	.w2(32'hbc004bec),
	.w3(32'h3c40c638),
	.w4(32'hba9a576c),
	.w5(32'hbb1520b9),
	.w6(32'hbb304487),
	.w7(32'hbaa098f2),
	.w8(32'hbbeddbf4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29a05d),
	.w1(32'h3b297825),
	.w2(32'h3c1f2ac4),
	.w3(32'h3b256115),
	.w4(32'hbb2bc5e0),
	.w5(32'h3b30ce26),
	.w6(32'hba3ede04),
	.w7(32'hbd143904),
	.w8(32'hbc81c95e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5eca0),
	.w1(32'h3c1f58de),
	.w2(32'hbb390fde),
	.w3(32'h3ba4ae6c),
	.w4(32'h3af6fb1d),
	.w5(32'hbac5b5f9),
	.w6(32'hba50a0dc),
	.w7(32'h3c286263),
	.w8(32'hbbc168da),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c157174),
	.w1(32'hbbfc4425),
	.w2(32'h3c085261),
	.w3(32'h3b5e57d2),
	.w4(32'h3ba1033b),
	.w5(32'hba3916d5),
	.w6(32'hbb43b54d),
	.w7(32'hba6dc75f),
	.w8(32'h3bd06d60),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4d981),
	.w1(32'h3a2d6c12),
	.w2(32'hba8e4b3c),
	.w3(32'h3bf9d05d),
	.w4(32'h3c8836e3),
	.w5(32'h3b407605),
	.w6(32'h3bab9e9d),
	.w7(32'h3c5ae395),
	.w8(32'hbc49637b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2db679),
	.w1(32'h3b3a0aea),
	.w2(32'h3b165018),
	.w3(32'h38aa2ee3),
	.w4(32'h3c18d1c1),
	.w5(32'hbac0f30e),
	.w6(32'hb9f66ba3),
	.w7(32'hba130d39),
	.w8(32'h3bdbdf8c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f5f2),
	.w1(32'h3bdf0283),
	.w2(32'h3c3377e5),
	.w3(32'h3bcaef1f),
	.w4(32'hbb60ae0e),
	.w5(32'h3bcaf787),
	.w6(32'h3c47b321),
	.w7(32'h3b0da7a7),
	.w8(32'hbc042c2d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bf32b),
	.w1(32'h381e663f),
	.w2(32'hb89c8444),
	.w3(32'h3abd427c),
	.w4(32'hbb8cd7cc),
	.w5(32'h3c9792d2),
	.w6(32'h3c180266),
	.w7(32'h3a66e25f),
	.w8(32'hbbd28004),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3e80),
	.w1(32'hbb2b30a0),
	.w2(32'hbb15d9d8),
	.w3(32'h3b689fd1),
	.w4(32'hbb7e68cc),
	.w5(32'hbc622149),
	.w6(32'h3b301135),
	.w7(32'hbb6a0834),
	.w8(32'h3bd19aff),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfda836),
	.w1(32'hbb82dd15),
	.w2(32'hbb21032f),
	.w3(32'h3ad89437),
	.w4(32'hbaac2106),
	.w5(32'h3bcfb91f),
	.w6(32'hb9129a62),
	.w7(32'hbaf48d62),
	.w8(32'h3bade47b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89192a),
	.w1(32'h3c2b776e),
	.w2(32'h3b15c592),
	.w3(32'h3b53d486),
	.w4(32'hbc27c86f),
	.w5(32'h3bf6732a),
	.w6(32'hbb80bdfb),
	.w7(32'hbb180b2c),
	.w8(32'h3a498c4b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f67b41),
	.w1(32'h3a57bc35),
	.w2(32'hbab9f6b4),
	.w3(32'hbb49f1c4),
	.w4(32'hbb2f9350),
	.w5(32'hbbe2165f),
	.w6(32'hbba8637b),
	.w7(32'h3a1fc25e),
	.w8(32'hbbeaadb3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf26ab7),
	.w1(32'h3b8b5189),
	.w2(32'h3bf4f10c),
	.w3(32'h3ab77f37),
	.w4(32'hbbb811bb),
	.w5(32'hb97049e8),
	.w6(32'hb8cf6e94),
	.w7(32'h3bfdcd05),
	.w8(32'h3acbc96f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d6d8),
	.w1(32'h3c0e73c1),
	.w2(32'hbb246589),
	.w3(32'h3c13bb50),
	.w4(32'h3c268317),
	.w5(32'hb922a5f0),
	.w6(32'hbb86ab53),
	.w7(32'hb9dd4051),
	.w8(32'hbbce64df),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba266a1b),
	.w1(32'hba8672ee),
	.w2(32'h3aeb461a),
	.w3(32'hb9358d4d),
	.w4(32'hbbebddcc),
	.w5(32'h3c0c84d9),
	.w6(32'h3be39c4a),
	.w7(32'hbbe3f901),
	.w8(32'h3bf5a049),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1116b3),
	.w1(32'h3b65006f),
	.w2(32'hb9257993),
	.w3(32'h3bc76106),
	.w4(32'h3b8e1587),
	.w5(32'h3b254ee9),
	.w6(32'h3b540c3c),
	.w7(32'hbbf2cf56),
	.w8(32'h3be7bfde),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67eb0b),
	.w1(32'h3a9169bb),
	.w2(32'h3a20632d),
	.w3(32'hbb27a12c),
	.w4(32'hba43616c),
	.w5(32'h3c0fc988),
	.w6(32'hbb937e25),
	.w7(32'h3c751be1),
	.w8(32'h39ed5a97),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e40ec),
	.w1(32'hb8698d80),
	.w2(32'hbad1f657),
	.w3(32'hbc661a15),
	.w4(32'hbb8819c5),
	.w5(32'hbbf58498),
	.w6(32'hba6c31d6),
	.w7(32'h3a119077),
	.w8(32'h3aa67795),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba548169),
	.w1(32'hbbc5171a),
	.w2(32'h3bf286f9),
	.w3(32'h3a3907dd),
	.w4(32'h3b52781a),
	.w5(32'h3a1635df),
	.w6(32'h3a8071f6),
	.w7(32'hbcccd37b),
	.w8(32'hbb07a0d3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b710570),
	.w1(32'h3a3066b2),
	.w2(32'hbb0e0cc8),
	.w3(32'h3959396a),
	.w4(32'h3c32bd86),
	.w5(32'hb9c9233a),
	.w6(32'h3b264d7c),
	.w7(32'hbb06ce3e),
	.w8(32'hbb91502a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11603b),
	.w1(32'h3be6926d),
	.w2(32'h3bf87f21),
	.w3(32'hbad3acca),
	.w4(32'h3aab8006),
	.w5(32'h3c9ba160),
	.w6(32'hbb61be1a),
	.w7(32'h3b2a11cc),
	.w8(32'h3badb2dc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace1059),
	.w1(32'hbaedefcd),
	.w2(32'hbb78e2d6),
	.w3(32'hbbb65e93),
	.w4(32'h3b63bb1d),
	.w5(32'h3b973f2e),
	.w6(32'hbbc5fec4),
	.w7(32'h3b27766a),
	.w8(32'hbbb43841),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7e0e3),
	.w1(32'h3ab2f409),
	.w2(32'h3c2f884b),
	.w3(32'hbb671bc9),
	.w4(32'hbabb89e2),
	.w5(32'hbbb987ab),
	.w6(32'h3b60d21c),
	.w7(32'h3b4d46c2),
	.w8(32'hbc1aadc7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52ee79),
	.w1(32'hbc0cfc80),
	.w2(32'h3a487087),
	.w3(32'h39a31855),
	.w4(32'hbbdade40),
	.w5(32'h3b235f5a),
	.w6(32'hbc2b0a31),
	.w7(32'hbc3d022f),
	.w8(32'h3af3e576),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b427b),
	.w1(32'hbb325d4d),
	.w2(32'hbbd4de00),
	.w3(32'h3c8606e5),
	.w4(32'h3b810365),
	.w5(32'hbb140d90),
	.w6(32'hba6f6a9c),
	.w7(32'h3b9b8b99),
	.w8(32'h3c7599c7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1c540),
	.w1(32'h3c500ab1),
	.w2(32'hbbe71ad1),
	.w3(32'h3c85833a),
	.w4(32'h3a127203),
	.w5(32'hbc5d52c0),
	.w6(32'h3bf65db8),
	.w7(32'h3b9f8332),
	.w8(32'h3b5d8b12),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83fe32),
	.w1(32'hba5f82c0),
	.w2(32'h3c23e406),
	.w3(32'hbc17a92e),
	.w4(32'hbb381a89),
	.w5(32'h3b82a612),
	.w6(32'h3c48aca3),
	.w7(32'hbc2491bd),
	.w8(32'h3b34d9fd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73f384),
	.w1(32'hbc061b4b),
	.w2(32'h3aa4bb7d),
	.w3(32'hbb9c322a),
	.w4(32'h3c07fdb1),
	.w5(32'h3c155df2),
	.w6(32'h3c775c0d),
	.w7(32'hbb725645),
	.w8(32'hbb91995b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe69a),
	.w1(32'hbb110e74),
	.w2(32'h39da22f0),
	.w3(32'hbc4a53ee),
	.w4(32'h3b8d5630),
	.w5(32'hbbfe1a25),
	.w6(32'h3ca9774a),
	.w7(32'h3b43ebec),
	.w8(32'h3a1859b5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc744a),
	.w1(32'h3a46b768),
	.w2(32'hba6bb009),
	.w3(32'hbb71979c),
	.w4(32'h39b83027),
	.w5(32'h3af3e8e2),
	.w6(32'h3c64ee37),
	.w7(32'h3984d234),
	.w8(32'hbb45b9cd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c2339),
	.w1(32'hbbaf44fd),
	.w2(32'hbc601d9d),
	.w3(32'h3ba17c97),
	.w4(32'h394b2d9d),
	.w5(32'h3ce71fb3),
	.w6(32'hb8b1b9cb),
	.w7(32'h3cbdfd37),
	.w8(32'hba1f8e02),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c172a1a),
	.w1(32'h3c8b8014),
	.w2(32'hbbbb1b68),
	.w3(32'hbb82a904),
	.w4(32'hbbb70ed6),
	.w5(32'hbc3501cd),
	.w6(32'h3c02f561),
	.w7(32'h3cb8a515),
	.w8(32'hba472b8f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a1ffb),
	.w1(32'h3c8a23ca),
	.w2(32'h3c19ec7e),
	.w3(32'hbc4f8277),
	.w4(32'hb9e8567a),
	.w5(32'h3c196aa7),
	.w6(32'h3aaec67f),
	.w7(32'h3b5f3d6b),
	.w8(32'h3c0b5458),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bceec95),
	.w1(32'hbbab4a1a),
	.w2(32'hbc05fe0d),
	.w3(32'h3b1d439a),
	.w4(32'hbb8cf7e3),
	.w5(32'hbb97e757),
	.w6(32'h3b6f947a),
	.w7(32'h39fa857c),
	.w8(32'h3cb6bc71),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3d6e2),
	.w1(32'h3d101499),
	.w2(32'hba75fb32),
	.w3(32'h39a35efb),
	.w4(32'hbc5a77a2),
	.w5(32'hbbd1b1dd),
	.w6(32'hbb260794),
	.w7(32'hbaac92ad),
	.w8(32'hbaa77d44),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc004126),
	.w1(32'hbba1b77d),
	.w2(32'hba077f48),
	.w3(32'h3c4ae998),
	.w4(32'h3b35f549),
	.w5(32'hba1b40b6),
	.w6(32'hbbb9b8c3),
	.w7(32'h3c6467ad),
	.w8(32'hbbbb167b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa06988),
	.w1(32'h3adb55d8),
	.w2(32'h3c238496),
	.w3(32'hbc8eeb40),
	.w4(32'h3aaedb9a),
	.w5(32'h3ba74146),
	.w6(32'hbb26b266),
	.w7(32'h3c3323d0),
	.w8(32'hba460c99),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b649260),
	.w1(32'h3b1f91b2),
	.w2(32'hbc442312),
	.w3(32'h3c713e64),
	.w4(32'h3b007941),
	.w5(32'hbb86b3b7),
	.w6(32'h3b142696),
	.w7(32'hbbecc926),
	.w8(32'hbb2b6d5c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc1457),
	.w1(32'h3b6d15be),
	.w2(32'h3bd58b57),
	.w3(32'h3b0834ce),
	.w4(32'h3bc982df),
	.w5(32'h3c1baf0b),
	.w6(32'h3c227a7a),
	.w7(32'hbbff891f),
	.w8(32'h3cac85f8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad646),
	.w1(32'hbb95f742),
	.w2(32'hbbcadbc0),
	.w3(32'h394cb8b8),
	.w4(32'h3acff14a),
	.w5(32'hbad8a827),
	.w6(32'h3b415ee0),
	.w7(32'h3a9ec7b4),
	.w8(32'hbc13ac15),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9ce50),
	.w1(32'h3ae9be35),
	.w2(32'hb71950dd),
	.w3(32'hbbc3e19d),
	.w4(32'hbc013b8e),
	.w5(32'h3b478996),
	.w6(32'hbbfd70e8),
	.w7(32'h3a84ee62),
	.w8(32'hbb87dfc1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf6e8b),
	.w1(32'hba41312d),
	.w2(32'hbc0a68d5),
	.w3(32'h3c4c41f0),
	.w4(32'hbb7f3d0c),
	.w5(32'h38c24328),
	.w6(32'hbba639ff),
	.w7(32'h3bb56cfb),
	.w8(32'hbbd1c151),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3797cb),
	.w1(32'hbbf358c6),
	.w2(32'hbbf019a9),
	.w3(32'hbbb7c46e),
	.w4(32'hbb059ee4),
	.w5(32'h3b94c9ba),
	.w6(32'h3a8da5c9),
	.w7(32'hbad86b37),
	.w8(32'h3b994f46),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc45b0),
	.w1(32'h39363c72),
	.w2(32'hbbb5a1df),
	.w3(32'h3c8eb58d),
	.w4(32'h3c647970),
	.w5(32'h3c03cb05),
	.w6(32'h3bd4c2bb),
	.w7(32'hba6feab8),
	.w8(32'h3ba29b19),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc386),
	.w1(32'h38db0dcd),
	.w2(32'hbb8cf421),
	.w3(32'hbbef750c),
	.w4(32'h398d1055),
	.w5(32'hb81a8833),
	.w6(32'h3b54184a),
	.w7(32'hbac68f86),
	.w8(32'h3c1f6fd3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71648a),
	.w1(32'h3b1614ab),
	.w2(32'h3c5ecdb2),
	.w3(32'h3c1f4d4e),
	.w4(32'h3b499a12),
	.w5(32'h395ab960),
	.w6(32'hbb324528),
	.w7(32'h3c345989),
	.w8(32'hbbcad5c7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe40a99),
	.w1(32'h3c3deb82),
	.w2(32'hba8ec0e8),
	.w3(32'hbad3980d),
	.w4(32'h3b5394f5),
	.w5(32'h3a2b6dfc),
	.w6(32'h3bdbd55a),
	.w7(32'h39a25c92),
	.w8(32'h3b81e0dc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc404247),
	.w1(32'hbbf8e5b4),
	.w2(32'hbabae813),
	.w3(32'hbbca9b19),
	.w4(32'h3b9a6449),
	.w5(32'h3c9e0650),
	.w6(32'h3b0e7e65),
	.w7(32'hbb410129),
	.w8(32'hbb97b085),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15a09f),
	.w1(32'h3c770e00),
	.w2(32'hbc8de2f0),
	.w3(32'hbb2aa90c),
	.w4(32'h3a0e67b1),
	.w5(32'h3c30fb22),
	.w6(32'h3bb39005),
	.w7(32'hbc9e7191),
	.w8(32'h3c147005),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77d22a),
	.w1(32'hbc16e080),
	.w2(32'hbc220d87),
	.w3(32'hbb07df02),
	.w4(32'hbb1791c3),
	.w5(32'h3b3cefb0),
	.w6(32'hba4c5bdd),
	.w7(32'hbc41c003),
	.w8(32'h3bb2043b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b168c7d),
	.w1(32'h3c018f5a),
	.w2(32'h3bb6b26a),
	.w3(32'hbb8fa49f),
	.w4(32'h3b3512e2),
	.w5(32'h3b660f20),
	.w6(32'hbc8a1cac),
	.w7(32'h3afbda84),
	.w8(32'hbabd5c67),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ef6e),
	.w1(32'hbc39b243),
	.w2(32'h3aff8494),
	.w3(32'hbb013ebc),
	.w4(32'h3ae80a5f),
	.w5(32'hbbd8795e),
	.w6(32'hbb87627c),
	.w7(32'hbc80bf3d),
	.w8(32'h3c4bb83a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d123502),
	.w1(32'hbb64343c),
	.w2(32'h3bb935a2),
	.w3(32'h3b691be5),
	.w4(32'hbb0d1c96),
	.w5(32'hbb81b601),
	.w6(32'hbb1531e0),
	.w7(32'h3a125e63),
	.w8(32'hbcc97cf9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7bb44),
	.w1(32'hbc16b037),
	.w2(32'hbc5ce2ef),
	.w3(32'hbbdeb753),
	.w4(32'h3ba04d7f),
	.w5(32'h3a7942df),
	.w6(32'hbc0132d1),
	.w7(32'hbbaea008),
	.w8(32'hbb3d5b45),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88149c),
	.w1(32'h3b0937e2),
	.w2(32'h3ba70517),
	.w3(32'hbbd1b4a9),
	.w4(32'hbbef0e7b),
	.w5(32'hb9f374e4),
	.w6(32'hbb8b8a9f),
	.w7(32'hba85596d),
	.w8(32'hbcbfbebf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804053),
	.w1(32'hbbfedfe4),
	.w2(32'hbbb68bba),
	.w3(32'hbc0fd429),
	.w4(32'h3aa99877),
	.w5(32'hb9ff6904),
	.w6(32'h3b99f834),
	.w7(32'hbc32fb42),
	.w8(32'h397b14de),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e75f9),
	.w1(32'hbbc4611f),
	.w2(32'hbb88ce2e),
	.w3(32'h3c952817),
	.w4(32'hbc6fa6d0),
	.w5(32'hbca68245),
	.w6(32'hbbf523cb),
	.w7(32'hbc1037f3),
	.w8(32'hbb5c3d92),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67eb19),
	.w1(32'hbb2e85df),
	.w2(32'hb9a2f035),
	.w3(32'h3bb2fa5b),
	.w4(32'hbacd9f40),
	.w5(32'hba4ccbda),
	.w6(32'hbbbb7344),
	.w7(32'hbcdbebf6),
	.w8(32'h3aeb7a0d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7752e0),
	.w1(32'hba9e229e),
	.w2(32'hbae7a4b5),
	.w3(32'h3b15bb2b),
	.w4(32'hbc5a8bb9),
	.w5(32'h3b83c7af),
	.w6(32'h3ba692af),
	.w7(32'hbb269bd1),
	.w8(32'hbb1113b0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962616),
	.w1(32'h3c344947),
	.w2(32'h3acf71bb),
	.w3(32'h3c2c96de),
	.w4(32'hbc1ba5a2),
	.w5(32'hba416641),
	.w6(32'hbbd4e299),
	.w7(32'hbc43cd4d),
	.w8(32'hbc3e56e4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee71c9),
	.w1(32'h3b1ee343),
	.w2(32'hbbfdb8d3),
	.w3(32'hb953bbf1),
	.w4(32'hb9cefe8b),
	.w5(32'hbbf2720b),
	.w6(32'hbaa7fa6f),
	.w7(32'hb9100c6a),
	.w8(32'hbb409f4c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c634e),
	.w1(32'h3c26cdcd),
	.w2(32'h3cc5301e),
	.w3(32'hbb8f4519),
	.w4(32'hbc03e30c),
	.w5(32'hbbbcc4be),
	.w6(32'hb9bfad83),
	.w7(32'h39a19246),
	.w8(32'h3c980ee5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d05058),
	.w1(32'hbbf98f8c),
	.w2(32'h3b57996c),
	.w3(32'hbbfb99a7),
	.w4(32'hba822c50),
	.w5(32'h3a876024),
	.w6(32'hbb84d729),
	.w7(32'hbb187283),
	.w8(32'hb6e864ad),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae81a04),
	.w1(32'h3c08bf4f),
	.w2(32'h3bab2363),
	.w3(32'hbc926415),
	.w4(32'h3c28182d),
	.w5(32'hbaa7dfe2),
	.w6(32'hbbae516d),
	.w7(32'hbad59c5e),
	.w8(32'h3a630501),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b915e5e),
	.w1(32'h3c1ea13f),
	.w2(32'hbbfb4777),
	.w3(32'h3cd2ec13),
	.w4(32'hbb23f18b),
	.w5(32'h39f2a152),
	.w6(32'hb8da87d7),
	.w7(32'hbb37ce6f),
	.w8(32'h3b4ba908),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf37591),
	.w1(32'h3b7efc78),
	.w2(32'h3c3ada8a),
	.w3(32'hbb925a15),
	.w4(32'h3afc40a8),
	.w5(32'hbc2ab221),
	.w6(32'hbb422a74),
	.w7(32'hbc3e1f1d),
	.w8(32'hbca1ea0f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fdac4),
	.w1(32'h3a73db89),
	.w2(32'hbc950140),
	.w3(32'hbcd426d5),
	.w4(32'hbc3c7f86),
	.w5(32'hbb84de75),
	.w6(32'hbb9502e4),
	.w7(32'hbaf5aa12),
	.w8(32'hbc1e73a2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4ff4b),
	.w1(32'hba059b28),
	.w2(32'hbc0019a7),
	.w3(32'hbbd3fb36),
	.w4(32'hba10de99),
	.w5(32'h3a6ca519),
	.w6(32'hbbd26eac),
	.w7(32'h3b2f5ffb),
	.w8(32'hbb3d010d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75d766),
	.w1(32'h3b081f85),
	.w2(32'hba918741),
	.w3(32'h3a4e43f4),
	.w4(32'hbb463841),
	.w5(32'hbb14fbeb),
	.w6(32'h3bb1a770),
	.w7(32'hbd186b0c),
	.w8(32'hbb0d0a4f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5241f),
	.w1(32'hbc2209b8),
	.w2(32'hbbc2f18c),
	.w3(32'hba501201),
	.w4(32'hbc5338cb),
	.w5(32'hbb3481d7),
	.w6(32'hbc5bdb8f),
	.w7(32'hba47dfb8),
	.w8(32'hbb723c18),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd23213),
	.w1(32'hbc55ddf3),
	.w2(32'h392f454f),
	.w3(32'h3b86b08e),
	.w4(32'hba75ffea),
	.w5(32'h3a4041e8),
	.w6(32'hbd0317d8),
	.w7(32'hbc7ec10b),
	.w8(32'h3afcc330),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b77fc5),
	.w1(32'hbb77fa70),
	.w2(32'hb98ae391),
	.w3(32'hba7048d8),
	.w4(32'h3b7023a2),
	.w5(32'hbb3d251d),
	.w6(32'hbb38f186),
	.w7(32'hbbd81f99),
	.w8(32'hba904b67),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd45b7),
	.w1(32'h3c59a998),
	.w2(32'h3ac33054),
	.w3(32'h3d0c148f),
	.w4(32'h3c062b5f),
	.w5(32'hbbdc4e7f),
	.w6(32'hbb22f0cf),
	.w7(32'hbc1a3163),
	.w8(32'h3bc6dd11),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfff458),
	.w1(32'h3c1dcfc3),
	.w2(32'h3c91f642),
	.w3(32'hbac2fa0e),
	.w4(32'hbb22fb8f),
	.w5(32'hbaf68702),
	.w6(32'h3aff7c5b),
	.w7(32'hbbf2d816),
	.w8(32'h3c2ec82f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caeaa1c),
	.w1(32'hbbceb60c),
	.w2(32'hbba99d14),
	.w3(32'hbb80bd59),
	.w4(32'hbb62699f),
	.w5(32'h3b241ee5),
	.w6(32'hb81b82fa),
	.w7(32'hbbb7d571),
	.w8(32'h389db4d6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941809f),
	.w1(32'hbd64a8a9),
	.w2(32'hbc0bce3a),
	.w3(32'h3bc64757),
	.w4(32'hbbfce737),
	.w5(32'hbb5ed3f8),
	.w6(32'hbae6256a),
	.w7(32'hbc979276),
	.w8(32'h38b88261),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5293ad),
	.w1(32'h3b84c4df),
	.w2(32'hba7ec4b2),
	.w3(32'h3c0125a2),
	.w4(32'hba6a6eed),
	.w5(32'h3c044334),
	.w6(32'h3cbdfaf0),
	.w7(32'h3b120779),
	.w8(32'hb9d3be81),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb14aa),
	.w1(32'h3a0f854b),
	.w2(32'hba8375e7),
	.w3(32'hbd0c43c0),
	.w4(32'h3b078c5e),
	.w5(32'h3a1192a9),
	.w6(32'hbb8de5c0),
	.w7(32'h3cc80d65),
	.w8(32'hbb714aec),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb7da),
	.w1(32'h3c2150b3),
	.w2(32'hbbabf63c),
	.w3(32'h3bfe68d5),
	.w4(32'hbafec71a),
	.w5(32'hbad9412b),
	.w6(32'hbb2afaf4),
	.w7(32'hba44d7b6),
	.w8(32'hbbf035a7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c5d93),
	.w1(32'hbc0d1ab8),
	.w2(32'hbbe7994a),
	.w3(32'hb9b46c6f),
	.w4(32'hbaed29fa),
	.w5(32'hbbd39050),
	.w6(32'hbb497cba),
	.w7(32'h3acd9fd2),
	.w8(32'hbbcbffc8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e88bb),
	.w1(32'hbb904009),
	.w2(32'hbaf9ed84),
	.w3(32'hbb7bb04a),
	.w4(32'h3bff0c99),
	.w5(32'hbaf9bb21),
	.w6(32'hb918011b),
	.w7(32'hb81f0454),
	.w8(32'hbc374f53),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21dde8),
	.w1(32'h3c0f08b7),
	.w2(32'hbabcea9d),
	.w3(32'h3a946a4b),
	.w4(32'h3b558b3b),
	.w5(32'hbb3f92ee),
	.w6(32'h3aa6f967),
	.w7(32'hbb949b77),
	.w8(32'hbab9ee81),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b904be6),
	.w1(32'hbc30e393),
	.w2(32'hbbd64358),
	.w3(32'h39a0d123),
	.w4(32'h3ca373e2),
	.w5(32'hbab4e069),
	.w6(32'hbb1badc6),
	.w7(32'h3c45e6a7),
	.w8(32'h3a9682c0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1228f),
	.w1(32'hba6d22c7),
	.w2(32'hbaf955c1),
	.w3(32'h39fd1ea4),
	.w4(32'hbb04f2de),
	.w5(32'hba60529c),
	.w6(32'hbb2ab280),
	.w7(32'h3b0fb218),
	.w8(32'h3b0768bf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054dd2),
	.w1(32'hbc0374bb),
	.w2(32'hbb046eb1),
	.w3(32'hbbdbe31c),
	.w4(32'h3ca831d7),
	.w5(32'hbab2ca2b),
	.w6(32'hbbad533b),
	.w7(32'hbbcfcf01),
	.w8(32'h3c8d6cab),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a80b),
	.w1(32'h3c154bf4),
	.w2(32'h3b918701),
	.w3(32'h3b23af6f),
	.w4(32'h3cc9b354),
	.w5(32'hbae7b842),
	.w6(32'h3b210778),
	.w7(32'h3ba1e0bc),
	.w8(32'h3a0e1b6a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df250),
	.w1(32'h3b7894b7),
	.w2(32'hbbdfeed0),
	.w3(32'h3abe2cda),
	.w4(32'h3b0e856c),
	.w5(32'h3b63d3a9),
	.w6(32'hbbd9a3ee),
	.w7(32'h3badb540),
	.w8(32'h3c64ab93),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad86c9e),
	.w1(32'hbb8c3ccb),
	.w2(32'hbbf41fb2),
	.w3(32'hbb073375),
	.w4(32'hbc267aca),
	.w5(32'hbba2916a),
	.w6(32'hbb2e25c9),
	.w7(32'h3c1a606e),
	.w8(32'hbb72c13a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b3d1),
	.w1(32'hbb70984f),
	.w2(32'h3c0fb98d),
	.w3(32'h3a91f723),
	.w4(32'hbb1d31e5),
	.w5(32'hba1bd823),
	.w6(32'hbc2c4af7),
	.w7(32'hbaaf8a6a),
	.w8(32'h3a86d037),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba111b02),
	.w1(32'hbb5cc228),
	.w2(32'hbb87915d),
	.w3(32'hbc62dcc5),
	.w4(32'h39fcbd7a),
	.w5(32'h3b0a6d8f),
	.w6(32'h3b8bbb13),
	.w7(32'hbc0d6468),
	.w8(32'hbb4e5d25),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70d61d),
	.w1(32'h3b5b27b5),
	.w2(32'hbbc1c819),
	.w3(32'h3c24e304),
	.w4(32'hb9c6af0b),
	.w5(32'h3ba593de),
	.w6(32'h3c1df756),
	.w7(32'hbbc5e848),
	.w8(32'hbc01bd98),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82b90e),
	.w1(32'h3bad88ee),
	.w2(32'hbbc021aa),
	.w3(32'h3ca42d9e),
	.w4(32'hbc07575e),
	.w5(32'hb8a735cb),
	.w6(32'h3b071b34),
	.w7(32'hbc26a1aa),
	.w8(32'h3a9faafd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4aeb1),
	.w1(32'h3a86d5a0),
	.w2(32'hb5fd1d1c),
	.w3(32'hbaf5a0ae),
	.w4(32'hba973c0b),
	.w5(32'hbc1e4cfa),
	.w6(32'hbb68fc52),
	.w7(32'h3b84af26),
	.w8(32'hbabaed51),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3138c),
	.w1(32'hbbc52e8c),
	.w2(32'h3ca8bebb),
	.w3(32'hbc831729),
	.w4(32'h3af849fe),
	.w5(32'h3c116f49),
	.w6(32'h3b0d9eed),
	.w7(32'hbbbaaaa4),
	.w8(32'h3c40062f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fba01),
	.w1(32'h3c911013),
	.w2(32'hb9d79632),
	.w3(32'h3a90f5fb),
	.w4(32'hba856194),
	.w5(32'hbb97c200),
	.w6(32'hbbc08188),
	.w7(32'h3b3b5ddf),
	.w8(32'h3b92ce37),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b968692),
	.w1(32'hbabcd755),
	.w2(32'hbc00ca02),
	.w3(32'h3995b0c3),
	.w4(32'h3b90dde8),
	.w5(32'hbb0e6408),
	.w6(32'hbc1e1af7),
	.w7(32'h3a99c4c3),
	.w8(32'h3a2fe785),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeed754),
	.w1(32'hbb9c22d2),
	.w2(32'h3a95c2d0),
	.w3(32'h3a9be031),
	.w4(32'hbb566900),
	.w5(32'hbbe45e18),
	.w6(32'hbb1d99ee),
	.w7(32'h39acac8f),
	.w8(32'h3be6560c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6a9f2),
	.w1(32'h3a4b4c7d),
	.w2(32'hbc16dcc9),
	.w3(32'hbc1b9aa3),
	.w4(32'h3b18dfc7),
	.w5(32'hbb437b96),
	.w6(32'h3a962389),
	.w7(32'h36e7e1fb),
	.w8(32'h37fc2c00),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f3c1),
	.w1(32'hbc2d0914),
	.w2(32'hbb3ed7ab),
	.w3(32'h3b975fea),
	.w4(32'hbb854f2e),
	.w5(32'hbb9a10b8),
	.w6(32'hbc1ef3e1),
	.w7(32'h39070224),
	.w8(32'h3988af6a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17592),
	.w1(32'h3ba2a132),
	.w2(32'h3d15fe52),
	.w3(32'h3a8a1e74),
	.w4(32'h3b427a9d),
	.w5(32'hbc096a31),
	.w6(32'hbcaec88d),
	.w7(32'h3b75e446),
	.w8(32'h3c8b139d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e42dd),
	.w1(32'hbb23a929),
	.w2(32'hb9b2bb2e),
	.w3(32'hbb9653ac),
	.w4(32'h39409e56),
	.w5(32'h3b11997d),
	.w6(32'hba41bab2),
	.w7(32'hbb6323a5),
	.w8(32'hba7aaf77),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55a3fc),
	.w1(32'hba355780),
	.w2(32'hbb07e0fa),
	.w3(32'hbb57d55a),
	.w4(32'hbba28fa9),
	.w5(32'h3b556152),
	.w6(32'h3b0b534b),
	.w7(32'hbb2b79a8),
	.w8(32'h3a9a008b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba85b28),
	.w1(32'hbbf30141),
	.w2(32'hb9de34d3),
	.w3(32'hbc30a167),
	.w4(32'hbbf99b51),
	.w5(32'hb947be18),
	.w6(32'hba2cc509),
	.w7(32'hba956475),
	.w8(32'hbad9b866),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8050cc),
	.w1(32'hbb2394c2),
	.w2(32'h3bc174bd),
	.w3(32'hb9689cd6),
	.w4(32'h38d1a3de),
	.w5(32'h3bae9f1b),
	.w6(32'h3b86b51b),
	.w7(32'hbb39759f),
	.w8(32'h3c0266d7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1b117),
	.w1(32'hbb3fdd80),
	.w2(32'h39ec91be),
	.w3(32'hbab43ae9),
	.w4(32'hbad0e342),
	.w5(32'hbbde3efd),
	.w6(32'hbbb53de2),
	.w7(32'hbad67d03),
	.w8(32'h3b1bbc58),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85d00e),
	.w1(32'hbb2eacfb),
	.w2(32'hbb1b5836),
	.w3(32'hbbfca8c4),
	.w4(32'h3c6fed6c),
	.w5(32'h3b83bf25),
	.w6(32'h3b6c87c0),
	.w7(32'hbc46ebfb),
	.w8(32'hbb9618c3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bbaba),
	.w1(32'hbb859ede),
	.w2(32'hbbd2d69e),
	.w3(32'hbb982fee),
	.w4(32'hbb3ce5e7),
	.w5(32'hbc0aa135),
	.w6(32'hbc3ae641),
	.w7(32'h3ba0a343),
	.w8(32'hbbfdfbd2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b226a),
	.w1(32'hbb8f19b2),
	.w2(32'hba270d58),
	.w3(32'h3c2b94ee),
	.w4(32'hbb1b00ea),
	.w5(32'hbc497dbc),
	.w6(32'h3b6df791),
	.w7(32'h3a9d6f13),
	.w8(32'hbb51e617),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31dd58),
	.w1(32'hbbb562aa),
	.w2(32'hbbae8b0f),
	.w3(32'hbb11aa39),
	.w4(32'hbc0ba098),
	.w5(32'hbc333ad4),
	.w6(32'hbb74d013),
	.w7(32'hb9dda860),
	.w8(32'h3b8d0683),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195eff),
	.w1(32'hbbe95e40),
	.w2(32'hbb96e053),
	.w3(32'hb9bcad91),
	.w4(32'hba59085e),
	.w5(32'h3bc5f750),
	.w6(32'h3b925714),
	.w7(32'hbbdb66cd),
	.w8(32'hbb36e9b1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcc45e),
	.w1(32'h3d411a22),
	.w2(32'hbba9abee),
	.w3(32'hbb9f4750),
	.w4(32'hbba0b981),
	.w5(32'hbb03b0d3),
	.w6(32'hbb2acdf2),
	.w7(32'hbb8643f6),
	.w8(32'h3b17b6a7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb975d14),
	.w1(32'hbbb5fde0),
	.w2(32'h3ad870bf),
	.w3(32'hbc007c39),
	.w4(32'hbc57cbc8),
	.w5(32'hb901bfec),
	.w6(32'h3a9362f5),
	.w7(32'hbac1d09b),
	.w8(32'hba3309c0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e1dbc),
	.w1(32'hbbc91765),
	.w2(32'hbbca8809),
	.w3(32'hbb592d6b),
	.w4(32'hbc234507),
	.w5(32'hbc481023),
	.w6(32'hbc85cb62),
	.w7(32'hbc1c56b8),
	.w8(32'hbc0edae5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0329ef),
	.w1(32'hbba0efa8),
	.w2(32'hbc1c9fa1),
	.w3(32'hbc283913),
	.w4(32'h3b666a25),
	.w5(32'h3b6b46a1),
	.w6(32'hbbf98696),
	.w7(32'h3bab7eab),
	.w8(32'hbc2abab7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b7d7a),
	.w1(32'h3ba3dff6),
	.w2(32'hbc11cbf0),
	.w3(32'h3b8e57a2),
	.w4(32'h3abe7619),
	.w5(32'h3b1e2c24),
	.w6(32'hbb55b9a8),
	.w7(32'hbc0983e0),
	.w8(32'hbbf3962e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57d979),
	.w1(32'h3ba63fed),
	.w2(32'hbae6a49f),
	.w3(32'hbbbc1575),
	.w4(32'hbbf3f431),
	.w5(32'h3c31dae2),
	.w6(32'hbb8f463c),
	.w7(32'hba3b8e44),
	.w8(32'hbb0a039d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b401d2a),
	.w1(32'h3b9e7c33),
	.w2(32'hbb941ef7),
	.w3(32'hbc3281bc),
	.w4(32'h3bdebcf7),
	.w5(32'hbaf6a2af),
	.w6(32'hbb89f61b),
	.w7(32'h3b6ba725),
	.w8(32'hbae11a81),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5991c4),
	.w1(32'h3af22eaa),
	.w2(32'hbc3d6c54),
	.w3(32'hb998af56),
	.w4(32'hbc602fd4),
	.w5(32'h38c039e1),
	.w6(32'hbc00cdae),
	.w7(32'hbb0e8206),
	.w8(32'h3bbc9284),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6d36c),
	.w1(32'h3b91e806),
	.w2(32'hbb968f11),
	.w3(32'hbc44fbb7),
	.w4(32'hbb25d35a),
	.w5(32'hbbf378c5),
	.w6(32'h3af969b9),
	.w7(32'hba46b676),
	.w8(32'hb9ac12c4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560b6f),
	.w1(32'hbbd1ffed),
	.w2(32'hbc652a7b),
	.w3(32'hbc1e33cb),
	.w4(32'hbc352b34),
	.w5(32'h3af57b94),
	.w6(32'hbc9ee6c7),
	.w7(32'hbb2c0d44),
	.w8(32'hbb2b0f9c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5438e),
	.w1(32'h3bad8660),
	.w2(32'h3a5da193),
	.w3(32'hbb7136b3),
	.w4(32'hbc031044),
	.w5(32'hbb2e50aa),
	.w6(32'hbb82194e),
	.w7(32'hbba017ea),
	.w8(32'h3afb31ba),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192630),
	.w1(32'hbabd10ff),
	.w2(32'hba6ed7fd),
	.w3(32'h3a6c2e16),
	.w4(32'hbcbb8320),
	.w5(32'h3c43b091),
	.w6(32'hbbbb8094),
	.w7(32'hbce31fc0),
	.w8(32'hbc693db2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24457e),
	.w1(32'hb9074316),
	.w2(32'hbb036cb9),
	.w3(32'hbb6c072e),
	.w4(32'hbb9b13ad),
	.w5(32'hbb5c2b6b),
	.w6(32'hbc19b13c),
	.w7(32'h3c0967d3),
	.w8(32'h3baba77d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75267a),
	.w1(32'hbb3c42b0),
	.w2(32'hbb8143cf),
	.w3(32'h3ba1427b),
	.w4(32'hbbd570ab),
	.w5(32'hbc40f228),
	.w6(32'hbbbd73e8),
	.w7(32'hbc4d693a),
	.w8(32'hbc3b3dcb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d9ae),
	.w1(32'hbbd00053),
	.w2(32'h3c1b0793),
	.w3(32'hbc1b7eb5),
	.w4(32'h3980dfc2),
	.w5(32'hbba28ffa),
	.w6(32'hbbc1e591),
	.w7(32'hbc682528),
	.w8(32'hbc0468ab),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3511b),
	.w1(32'hbbca716c),
	.w2(32'h3bd3cf64),
	.w3(32'hbb19fe3f),
	.w4(32'h3a5f9bc4),
	.w5(32'hbb3107ca),
	.w6(32'h3b49efce),
	.w7(32'h3acea3a2),
	.w8(32'hb9c2254b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e2289d),
	.w1(32'hbb1577e7),
	.w2(32'hbc46c6ca),
	.w3(32'hbb4fca00),
	.w4(32'h3a4ac5c4),
	.w5(32'hbba6b1e9),
	.w6(32'h390f365c),
	.w7(32'hbc038471),
	.w8(32'hbb66b49d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf5202),
	.w1(32'hb9a63f46),
	.w2(32'h3bb8bfaf),
	.w3(32'h3a59e755),
	.w4(32'hb9904f7c),
	.w5(32'h3a9d3466),
	.w6(32'hbc00ed94),
	.w7(32'h3b8baa50),
	.w8(32'hbc725ed5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68dda7),
	.w1(32'hbc2f45ff),
	.w2(32'hbc542f70),
	.w3(32'h3b27ecc5),
	.w4(32'hba726893),
	.w5(32'hbb7378cd),
	.w6(32'hbbeb4032),
	.w7(32'hbb327709),
	.w8(32'hbc220ff7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b04a2),
	.w1(32'hbbeca9b0),
	.w2(32'hbac16253),
	.w3(32'h3a5e6044),
	.w4(32'hbbd9e935),
	.w5(32'hbbaa80d0),
	.w6(32'h3c16c5bc),
	.w7(32'hbc6bff4b),
	.w8(32'hbc0d866f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4256e),
	.w1(32'hbc52cf3c),
	.w2(32'hbabb454c),
	.w3(32'hbaeec0d1),
	.w4(32'hbc1ff3c6),
	.w5(32'hbba3f719),
	.w6(32'h3b8f9e69),
	.w7(32'hbc531284),
	.w8(32'hba5a020d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4b32c),
	.w1(32'hbb25d919),
	.w2(32'hbc2ed03d),
	.w3(32'h365c1b4c),
	.w4(32'hb9775de2),
	.w5(32'h3a886485),
	.w6(32'hbadc2415),
	.w7(32'hbb496a7b),
	.w8(32'hb9a38f8a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89846c),
	.w1(32'hbb1fdae3),
	.w2(32'hbb467a00),
	.w3(32'hbc11bac9),
	.w4(32'hbb513ad2),
	.w5(32'hbc0d48ed),
	.w6(32'h3aaf69d4),
	.w7(32'hbb15fe85),
	.w8(32'hbca8cdd8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0446e8),
	.w1(32'hbb691094),
	.w2(32'hbb9439c9),
	.w3(32'hbc18e73f),
	.w4(32'hbbc0f674),
	.w5(32'hbbf93973),
	.w6(32'h3a029e79),
	.w7(32'h3bb9f6c4),
	.w8(32'h3a9167fb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1629db),
	.w1(32'hbc55b9bd),
	.w2(32'hbbd85e73),
	.w3(32'hbbf8d90d),
	.w4(32'hbc057cf8),
	.w5(32'h3bfe670d),
	.w6(32'hbb85577d),
	.w7(32'hbc6f28e6),
	.w8(32'hbc582e19),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd11d1a),
	.w1(32'hbaa49b8c),
	.w2(32'hbc04fc96),
	.w3(32'h3abbcdc8),
	.w4(32'hbb56a7b2),
	.w5(32'hbaedbe87),
	.w6(32'h3b8f7e53),
	.w7(32'hbcaed09f),
	.w8(32'hba848e0b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8f6eb),
	.w1(32'hbb295b73),
	.w2(32'hbbf1e859),
	.w3(32'h3a17157d),
	.w4(32'hbbc33f93),
	.w5(32'h3a7b4bec),
	.w6(32'hbb2c61fc),
	.w7(32'hbbeac313),
	.w8(32'h3bbd8d56),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b2da),
	.w1(32'hbbbccba8),
	.w2(32'hb9c98980),
	.w3(32'hbb30dc92),
	.w4(32'h3a107261),
	.w5(32'hbb873535),
	.w6(32'hbc1fd5d7),
	.w7(32'h3af5e982),
	.w8(32'hb9f48d3e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule