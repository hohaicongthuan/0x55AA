module layer_10_featuremap_385(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942126b),
	.w1(32'h3a1ff31d),
	.w2(32'h3965c750),
	.w3(32'h39c0e0e0),
	.w4(32'h3a25c622),
	.w5(32'h393c2845),
	.w6(32'h3a8e9506),
	.w7(32'hb71703ea),
	.w8(32'hb938789b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b797dc),
	.w1(32'hba28e6a5),
	.w2(32'hba59a361),
	.w3(32'hb9766d32),
	.w4(32'hba41769c),
	.w5(32'hba0fe252),
	.w6(32'hb9f7ca8e),
	.w7(32'hba617bd3),
	.w8(32'hba1c0a7a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0edce2),
	.w1(32'hb9d40823),
	.w2(32'hba89e2ce),
	.w3(32'h3a12498b),
	.w4(32'hba80a4c6),
	.w5(32'hba3b6b41),
	.w6(32'h38c2bbbc),
	.w7(32'hba4e4c58),
	.w8(32'hbac13191),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2357d),
	.w1(32'h39a172f6),
	.w2(32'h389773fe),
	.w3(32'hb9f8e542),
	.w4(32'h38204093),
	.w5(32'hb9bf6a96),
	.w6(32'hba2867fd),
	.w7(32'hba078a38),
	.w8(32'hb8a00def),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959fd5b),
	.w1(32'hb980bf7d),
	.w2(32'h385d778b),
	.w3(32'hb982bb95),
	.w4(32'hba264ea6),
	.w5(32'hb98dc4c2),
	.w6(32'hb5ccb210),
	.w7(32'hba43e375),
	.w8(32'hba4e76ad),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6538c),
	.w1(32'hb952d025),
	.w2(32'hb91f64ca),
	.w3(32'hb70df38b),
	.w4(32'h38b3ba8a),
	.w5(32'hb9a8edde),
	.w6(32'hb9e2abbf),
	.w7(32'hb9a49c92),
	.w8(32'hb8e07bc9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a704e9),
	.w1(32'h3a815a42),
	.w2(32'h3a35e9af),
	.w3(32'h399064a6),
	.w4(32'hb95d9de1),
	.w5(32'hb74c8973),
	.w6(32'h39b17e93),
	.w7(32'h39b04a7d),
	.w8(32'h3920431a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a45d11),
	.w1(32'h3a3906a5),
	.w2(32'h3a36d6d3),
	.w3(32'hba3a4769),
	.w4(32'h3a4e9699),
	.w5(32'h3a12d68b),
	.w6(32'hb906711e),
	.w7(32'hb9a81a01),
	.w8(32'hb9b93229),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a767cc9),
	.w1(32'hb9865c68),
	.w2(32'hba03d632),
	.w3(32'h3a994380),
	.w4(32'hba270ce1),
	.w5(32'hb9d7e44f),
	.w6(32'hb9b8c8b9),
	.w7(32'hba71c6c0),
	.w8(32'hb9890e83),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33fd74),
	.w1(32'h3a8d29c1),
	.w2(32'h3a58348d),
	.w3(32'hba0a241d),
	.w4(32'hba1a97be),
	.w5(32'hba249534),
	.w6(32'hb9834c72),
	.w7(32'hb99cf7d5),
	.w8(32'hba581bf8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a608222),
	.w1(32'hb9d92ea5),
	.w2(32'h396c2679),
	.w3(32'hba27071e),
	.w4(32'hb9fa015c),
	.w5(32'hb9a6d88d),
	.w6(32'hba903888),
	.w7(32'h3a2a2953),
	.w8(32'hb919dfce),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a97a9),
	.w1(32'h39353c80),
	.w2(32'h3a656e3f),
	.w3(32'h3860fa5c),
	.w4(32'h3a801772),
	.w5(32'h3abc3506),
	.w6(32'h39889225),
	.w7(32'h3a5e91b1),
	.w8(32'h3a6e54ee),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a867e),
	.w1(32'h3a07f540),
	.w2(32'h39a00117),
	.w3(32'h3aa3d751),
	.w4(32'h3a44f71b),
	.w5(32'h3a1a753e),
	.w6(32'h3a6b764b),
	.w7(32'h39fbc028),
	.w8(32'h3a0473d4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3d2af),
	.w1(32'hb9744e9f),
	.w2(32'hb8aa4b92),
	.w3(32'h3a69b8cc),
	.w4(32'hba83f6d5),
	.w5(32'h3920e015),
	.w6(32'h3a33f40f),
	.w7(32'h392b2b95),
	.w8(32'hb90c4f5e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990f82c),
	.w1(32'hba3bcbd0),
	.w2(32'hb9d0620a),
	.w3(32'hb9858d6b),
	.w4(32'hbad0cf5a),
	.w5(32'hb9fd8bba),
	.w6(32'h39e7e506),
	.w7(32'hba66b957),
	.w8(32'hbab77d78),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca876e),
	.w1(32'hba49be7a),
	.w2(32'hb9e6efc8),
	.w3(32'hba9153c4),
	.w4(32'hba33e9b7),
	.w5(32'hb98d7a21),
	.w6(32'hba51a26f),
	.w7(32'hba2a81e9),
	.w8(32'hba22e378),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17dd81),
	.w1(32'h396193f9),
	.w2(32'h3a4e190c),
	.w3(32'hb9d0e48a),
	.w4(32'h3a0195f7),
	.w5(32'h3a9603aa),
	.w6(32'hb9cac8bd),
	.w7(32'h3a5e0fbc),
	.w8(32'h3a88600c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b1ebf6),
	.w1(32'h3a064fc4),
	.w2(32'hb901b475),
	.w3(32'h3a631aa6),
	.w4(32'h3a260e4e),
	.w5(32'h39dd49f0),
	.w6(32'h3a16a4ca),
	.w7(32'h3835c4ff),
	.w8(32'h3a0e682c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cddf40),
	.w1(32'hba152e38),
	.w2(32'h39130d2c),
	.w3(32'h39afb772),
	.w4(32'hb956a0bf),
	.w5(32'h39105ca5),
	.w6(32'h39806800),
	.w7(32'hb9b5e595),
	.w8(32'hb959e5f1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8126c92),
	.w1(32'hb9ba319f),
	.w2(32'h380cfc9e),
	.w3(32'hb87ff066),
	.w4(32'h38509450),
	.w5(32'h3a8a362d),
	.w6(32'hb98fee06),
	.w7(32'h3a830936),
	.w8(32'h38762a21),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c39158),
	.w1(32'hb90e86a4),
	.w2(32'hb9bfa0ba),
	.w3(32'h3a4b6711),
	.w4(32'hb9051959),
	.w5(32'hb9ced9c2),
	.w6(32'h3a8ea3bf),
	.w7(32'hba5e53fe),
	.w8(32'hba269eed),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a4a61),
	.w1(32'hba597e84),
	.w2(32'hba390b03),
	.w3(32'h39053120),
	.w4(32'hba4e7860),
	.w5(32'hba4ee0bc),
	.w6(32'hb9892b8f),
	.w7(32'hba984d70),
	.w8(32'hbabef6d6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ba5c0),
	.w1(32'h39b21037),
	.w2(32'h3a344b2c),
	.w3(32'hba9da5ed),
	.w4(32'h3a17a83d),
	.w5(32'h3a89056d),
	.w6(32'hba4734c2),
	.w7(32'h3a959c1d),
	.w8(32'h3a63f70a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a993d2b),
	.w1(32'hb8c8221d),
	.w2(32'hba0a79d5),
	.w3(32'h3a9618bc),
	.w4(32'hb9fe746e),
	.w5(32'hba8f658b),
	.w6(32'h3a2874ae),
	.w7(32'hb8a91bb4),
	.w8(32'hb9a5840c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8f0a0),
	.w1(32'hba1bad6e),
	.w2(32'h39481387),
	.w3(32'hb9a8807f),
	.w4(32'hb9faf8e5),
	.w5(32'h3a218a41),
	.w6(32'hb8ac1992),
	.w7(32'h393a69b9),
	.w8(32'hba77b745),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba818050),
	.w1(32'h3a5e1766),
	.w2(32'h3a334ea2),
	.w3(32'hb9e8b43e),
	.w4(32'h3a839e89),
	.w5(32'h391cbd91),
	.w6(32'hba806c0e),
	.w7(32'h3a552848),
	.w8(32'h39f739c0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7181ed),
	.w1(32'h3a799b93),
	.w2(32'h3986c954),
	.w3(32'h3a5f2b96),
	.w4(32'h39bab445),
	.w5(32'h38078717),
	.w6(32'h38f74415),
	.w7(32'h3a04db10),
	.w8(32'h3a865512),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39989518),
	.w1(32'h39c637ac),
	.w2(32'h3a0c2dbb),
	.w3(32'h398d9946),
	.w4(32'h39252bbd),
	.w5(32'h3938dd87),
	.w6(32'h3a9dd1dc),
	.w7(32'h393cbf25),
	.w8(32'hb9c234a1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9970978),
	.w1(32'h391a6236),
	.w2(32'hb8d493dc),
	.w3(32'hba1e604a),
	.w4(32'hb89ab22d),
	.w5(32'h3a31c10e),
	.w6(32'hba291463),
	.w7(32'h3a1a8574),
	.w8(32'h39f6bf76),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e9533),
	.w1(32'h38da883e),
	.w2(32'hb9d94c7f),
	.w3(32'h39cbc7d7),
	.w4(32'h388b42c4),
	.w5(32'hb93d440a),
	.w6(32'h39e11523),
	.w7(32'h3800fe6b),
	.w8(32'h38fe5f64),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00b35d),
	.w1(32'hb931bf31),
	.w2(32'h3a0dd104),
	.w3(32'h39a4f8f1),
	.w4(32'hba14f452),
	.w5(32'hb92fd126),
	.w6(32'h39f02d4a),
	.w7(32'h38427e38),
	.w8(32'h38a4176f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f550c),
	.w1(32'hb9cbbc9c),
	.w2(32'hba14c08c),
	.w3(32'hb95e1467),
	.w4(32'hba05b7b1),
	.w5(32'hb9f80312),
	.w6(32'hb9d1f101),
	.w7(32'hb9ca9a53),
	.w8(32'hba51985d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80370c9),
	.w1(32'h3a0471c6),
	.w2(32'h3a075344),
	.w3(32'h3953e167),
	.w4(32'h394a41b5),
	.w5(32'h3a5623ac),
	.w6(32'hb8aa8f9a),
	.w7(32'h3a15abcb),
	.w8(32'h3a21b982),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1bab7),
	.w1(32'h3a7d2b9a),
	.w2(32'h3a9f755c),
	.w3(32'hb9b48706),
	.w4(32'h3a44de56),
	.w5(32'h39a14c1b),
	.w6(32'hb7f0dafd),
	.w7(32'h3a4637bc),
	.w8(32'h3a05e553),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2201e4),
	.w1(32'hb9883058),
	.w2(32'hb88741aa),
	.w3(32'hb9af7d44),
	.w4(32'h39f8af07),
	.w5(32'h39464fe1),
	.w6(32'hba27cc9f),
	.w7(32'h3a38b2a3),
	.w8(32'h3a37fb4d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd26ba),
	.w1(32'h3713aa77),
	.w2(32'hb999a207),
	.w3(32'h39ef6e5d),
	.w4(32'h39983fb5),
	.w5(32'hb6b9074e),
	.w6(32'h3a7b3683),
	.w7(32'hb86e92ed),
	.w8(32'h3a18f947),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e4b84),
	.w1(32'h39df7eda),
	.w2(32'h3a0c83f5),
	.w3(32'h3a2249ec),
	.w4(32'hb9653610),
	.w5(32'hb85152d6),
	.w6(32'h3a2c26a4),
	.w7(32'hb89fac6f),
	.w8(32'hba1a5c47),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971d189),
	.w1(32'h3988f116),
	.w2(32'h399e3638),
	.w3(32'h36e74d06),
	.w4(32'hb9df2da6),
	.w5(32'hb8246e2c),
	.w6(32'h378cf13c),
	.w7(32'hba09ac9a),
	.w8(32'hb99c70be),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b88d6),
	.w1(32'h39e9ef8d),
	.w2(32'h3a1eba06),
	.w3(32'h3a692ddf),
	.w4(32'h3a0f9b5a),
	.w5(32'h3a063dad),
	.w6(32'hb8384654),
	.w7(32'h3a52c9c8),
	.w8(32'hb9d6e369),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9dc65),
	.w1(32'h398e1a1c),
	.w2(32'h39d515ef),
	.w3(32'hb9878c6c),
	.w4(32'h3a00ba61),
	.w5(32'h396afe09),
	.w6(32'h39c650da),
	.w7(32'h3a27807d),
	.w8(32'h37dfdf6b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a6890),
	.w1(32'h3a86691b),
	.w2(32'h39daa59a),
	.w3(32'h3a65442e),
	.w4(32'hb9af11e6),
	.w5(32'h3a8fc51c),
	.w6(32'hb910fea8),
	.w7(32'hb9e71720),
	.w8(32'h3a76e275),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392658dc),
	.w1(32'hb986363d),
	.w2(32'h3947cbb4),
	.w3(32'h39f0a0b7),
	.w4(32'hb9fe44c5),
	.w5(32'hb94d5f60),
	.w6(32'h39732e08),
	.w7(32'hba2ec3bd),
	.w8(32'hb9c392cc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a49e82),
	.w1(32'h395906f7),
	.w2(32'hb9d19bb1),
	.w3(32'hb96fdd8a),
	.w4(32'h38ea5403),
	.w5(32'hb9d47776),
	.w6(32'h37dc8221),
	.w7(32'h393b767e),
	.w8(32'hb815f569),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac9649),
	.w1(32'h3a5381b5),
	.w2(32'h3a469167),
	.w3(32'hb8a23f49),
	.w4(32'h3a96b18c),
	.w5(32'hb94bcc67),
	.w6(32'h39cc251a),
	.w7(32'h3a53c9cd),
	.w8(32'hb8804529),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea01de),
	.w1(32'h39cc69fb),
	.w2(32'h3a0c04de),
	.w3(32'h39e3e3b2),
	.w4(32'h39da4e66),
	.w5(32'h396eaa3a),
	.w6(32'h38be2509),
	.w7(32'h39e242be),
	.w8(32'h39694f0e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a05b1e),
	.w1(32'hba95e1a0),
	.w2(32'hba7fd0da),
	.w3(32'h38ff4237),
	.w4(32'hbaa3f025),
	.w5(32'hba49ff13),
	.w6(32'hb887b8a4),
	.w7(32'hba9eea01),
	.w8(32'hbac05b39),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88b1bd),
	.w1(32'hba2cce96),
	.w2(32'hb9896c90),
	.w3(32'hba6438d0),
	.w4(32'hba8ca515),
	.w5(32'hb924da9b),
	.w6(32'hba293510),
	.w7(32'h39988f22),
	.w8(32'h3882585f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e93f1),
	.w1(32'h3a16d831),
	.w2(32'hb9662c24),
	.w3(32'hba116a6c),
	.w4(32'h3951140a),
	.w5(32'hb9915804),
	.w6(32'h39fbea3a),
	.w7(32'h39f21a33),
	.w8(32'hb9ab8651),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9af25),
	.w1(32'hbab66e15),
	.w2(32'hba4731db),
	.w3(32'hba76e082),
	.w4(32'hb9c9a0e5),
	.w5(32'hb9ac223d),
	.w6(32'hba33d2fe),
	.w7(32'hb9a2e3c4),
	.w8(32'hb8ea1f98),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43342c),
	.w1(32'hba25e070),
	.w2(32'hb9b101aa),
	.w3(32'h394cda58),
	.w4(32'hb9f684b5),
	.w5(32'hb94deefc),
	.w6(32'h393d019e),
	.w7(32'hba1c807d),
	.w8(32'h36810049),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1330b3),
	.w1(32'h39c307be),
	.w2(32'h3909138a),
	.w3(32'h3a5eb90d),
	.w4(32'h3a627f5e),
	.w5(32'h3986dde4),
	.w6(32'h3a23b2f7),
	.w7(32'h39663be4),
	.w8(32'h3a13474e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed77c8),
	.w1(32'h3a60533a),
	.w2(32'h394b23b4),
	.w3(32'h38f6ea58),
	.w4(32'hb81d1f6f),
	.w5(32'hb74c8bcc),
	.w6(32'hb92cf902),
	.w7(32'h39773841),
	.w8(32'h38b514b6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a433d4f),
	.w1(32'h3990c51e),
	.w2(32'h39c0a4d4),
	.w3(32'h390d2fee),
	.w4(32'h39b78913),
	.w5(32'h39f5a1f8),
	.w6(32'h3a344745),
	.w7(32'h38ebfab7),
	.w8(32'h3a2730dc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39187492),
	.w1(32'h39ad3cdb),
	.w2(32'hb8b09d1a),
	.w3(32'h3a563ebb),
	.w4(32'h39e8c952),
	.w5(32'h390c3b24),
	.w6(32'h3a227e10),
	.w7(32'hb9b4dd86),
	.w8(32'hba457006),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba078027),
	.w1(32'hb86e1d69),
	.w2(32'hb95d3fc1),
	.w3(32'h388249a9),
	.w4(32'h39aa6b8a),
	.w5(32'hba1d3a85),
	.w6(32'hba5fdf9c),
	.w7(32'h3aa09dc2),
	.w8(32'hb961c1be),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa80188),
	.w1(32'hba88e43c),
	.w2(32'hba32c607),
	.w3(32'hb9c84ff6),
	.w4(32'hbaa06f63),
	.w5(32'hba2c6f92),
	.w6(32'hba2456c0),
	.w7(32'hba2c0d1d),
	.w8(32'hba43e67c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8537728),
	.w1(32'hb7589514),
	.w2(32'hb940e446),
	.w3(32'h398f201b),
	.w4(32'hb87f7f1f),
	.w5(32'hb96dab95),
	.w6(32'hb9f09bcf),
	.w7(32'hb9d7bb7b),
	.w8(32'hba168ac6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ee1689),
	.w1(32'hb9dbd63b),
	.w2(32'hb987bb63),
	.w3(32'hba3270e2),
	.w4(32'h39d4e367),
	.w5(32'hba4782e1),
	.w6(32'hba201d46),
	.w7(32'hba6aaab6),
	.w8(32'h381babad),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9af8e),
	.w1(32'h3a3c71fd),
	.w2(32'h3a6c07a8),
	.w3(32'hba57b1af),
	.w4(32'h3a52c28b),
	.w5(32'h399a321e),
	.w6(32'hba03fdaa),
	.w7(32'h3a498ba1),
	.w8(32'h39fd529d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a303cd7),
	.w1(32'hb9ea8d22),
	.w2(32'hb8ae37a1),
	.w3(32'h378a8ef4),
	.w4(32'hb8aaefbd),
	.w5(32'h3ae3bd15),
	.w6(32'h38cf0940),
	.w7(32'h3ad3ccc6),
	.w8(32'hb9c06cc1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f212),
	.w1(32'hba912158),
	.w2(32'hbadfcc4a),
	.w3(32'hb9a593fd),
	.w4(32'hba38ef49),
	.w5(32'hba09d698),
	.w6(32'h3a403416),
	.w7(32'h3984fe6b),
	.w8(32'h373799d3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae04d8e),
	.w1(32'hba32a9cb),
	.w2(32'hb9e49c5a),
	.w3(32'hb98a47e6),
	.w4(32'hba3f69bd),
	.w5(32'hba820890),
	.w6(32'h39459740),
	.w7(32'h386021f9),
	.w8(32'hba978f78),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b9780),
	.w1(32'hb9870844),
	.w2(32'hbab15ee8),
	.w3(32'hb9fe537c),
	.w4(32'hb99db906),
	.w5(32'hba7b0ebc),
	.w6(32'hba0dbaa4),
	.w7(32'hb981814c),
	.w8(32'hba88a90b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba280235),
	.w1(32'h3a00ad9f),
	.w2(32'h3a6c7390),
	.w3(32'hb9b0d300),
	.w4(32'h3a6a4602),
	.w5(32'h3a96f354),
	.w6(32'hba34f312),
	.w7(32'h3a4d5009),
	.w8(32'h3a787244),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dca7c),
	.w1(32'h3a7f1736),
	.w2(32'h3a844706),
	.w3(32'h3a2e8e00),
	.w4(32'h3a91110c),
	.w5(32'h3a54c81f),
	.w6(32'h3a20b459),
	.w7(32'h3a55a2d6),
	.w8(32'h3a93ec3b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a0d3b),
	.w1(32'hb991db7d),
	.w2(32'hb7ac8903),
	.w3(32'h3ac3e8e3),
	.w4(32'h375e872c),
	.w5(32'h3997a657),
	.w6(32'h3a7bbab3),
	.w7(32'hb7854f85),
	.w8(32'h39891797),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38642e51),
	.w1(32'hb9cf48e5),
	.w2(32'hb88b781f),
	.w3(32'h3a383afa),
	.w4(32'hb9a33e84),
	.w5(32'hba33b225),
	.w6(32'h3aaf4c65),
	.w7(32'hb9952dde),
	.w8(32'hba0bb23a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e2b3f),
	.w1(32'hbad28746),
	.w2(32'hba90f1cc),
	.w3(32'hba327085),
	.w4(32'hba76878b),
	.w5(32'hba6718f5),
	.w6(32'hb4cd15d6),
	.w7(32'hba839c26),
	.w8(32'hba576164),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65fb6d),
	.w1(32'h39f057aa),
	.w2(32'hba485543),
	.w3(32'hba46df7b),
	.w4(32'h38b04a0f),
	.w5(32'hba8c01a6),
	.w6(32'hbaac9f47),
	.w7(32'h38abce6e),
	.w8(32'hbabcb180),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3850df),
	.w1(32'h3c1a2b03),
	.w2(32'hbc8aa9a7),
	.w3(32'hba957006),
	.w4(32'hbb435564),
	.w5(32'hbb993aea),
	.w6(32'hbac85fd6),
	.w7(32'hbc776d54),
	.w8(32'h3d1e40f7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30c12c),
	.w1(32'hbb5b6428),
	.w2(32'hbb92fa03),
	.w3(32'hbc5e2cb3),
	.w4(32'h3b41d953),
	.w5(32'h3c1d677b),
	.w6(32'h3bf06cd7),
	.w7(32'h3c4d05c8),
	.w8(32'h3cb95ff2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1656),
	.w1(32'h3bd2912e),
	.w2(32'hb8f59e84),
	.w3(32'h3b4695e2),
	.w4(32'h3c299e4a),
	.w5(32'hbb9888e8),
	.w6(32'h3c569428),
	.w7(32'h3ba528a9),
	.w8(32'hbbea7595),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1943ac),
	.w1(32'hbaba4978),
	.w2(32'hbc874fe3),
	.w3(32'h3c2c90ba),
	.w4(32'hbc0671ee),
	.w5(32'hbc021546),
	.w6(32'h3aa02fd2),
	.w7(32'hbb145993),
	.w8(32'h3b72af6e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d9fe1),
	.w1(32'hbb66a06b),
	.w2(32'h3ac7bc4d),
	.w3(32'hbb9d4973),
	.w4(32'hbb832403),
	.w5(32'hb90fdc0b),
	.w6(32'hbbd7aa63),
	.w7(32'hbb489db2),
	.w8(32'hbb0ea395),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10777c),
	.w1(32'hba62b1d8),
	.w2(32'hbbb7ea15),
	.w3(32'hbbf9e662),
	.w4(32'hbcacb73d),
	.w5(32'hbc916ab1),
	.w6(32'hbc1e6a06),
	.w7(32'hbc5cb586),
	.w8(32'hbc65c05b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4945b),
	.w1(32'hbc168a3c),
	.w2(32'hbb11558f),
	.w3(32'hbc919a2f),
	.w4(32'h3bc3dbcb),
	.w5(32'h3cacec43),
	.w6(32'hbbf390e4),
	.w7(32'h3b9a2dc7),
	.w8(32'h3baffa0e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaef8c3),
	.w1(32'h3bc269e3),
	.w2(32'h3c5ec890),
	.w3(32'h3c0c1dd9),
	.w4(32'h3ae541b3),
	.w5(32'hbc19c221),
	.w6(32'hbabed93e),
	.w7(32'hbbb63210),
	.w8(32'hbc15d90e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56b5e6),
	.w1(32'hbc161d18),
	.w2(32'hbce692d5),
	.w3(32'hba6e5dba),
	.w4(32'hbc6a1b23),
	.w5(32'hbafa6818),
	.w6(32'hbba2f123),
	.w7(32'h3b89aef0),
	.w8(32'h3c948d46),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb1bd4),
	.w1(32'h3b929954),
	.w2(32'h3c299438),
	.w3(32'hbbab8303),
	.w4(32'h3aefab19),
	.w5(32'h3a090a17),
	.w6(32'h3c29a26b),
	.w7(32'hbb26e42b),
	.w8(32'hbc5b37a2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14cce4),
	.w1(32'hbc0f5e14),
	.w2(32'hbb8c0fe5),
	.w3(32'hbacd41b5),
	.w4(32'hbbbba25f),
	.w5(32'h3ba85704),
	.w6(32'hbc67e6dc),
	.w7(32'hbbc72a07),
	.w8(32'h3c433702),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9cd1),
	.w1(32'h3cf43950),
	.w2(32'h3d48d275),
	.w3(32'h3c02226f),
	.w4(32'h3c6cc8dd),
	.w5(32'h3c4f4484),
	.w6(32'h3c5fc1b2),
	.w7(32'hbcb97d91),
	.w8(32'hbd92fcd8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d052aa6),
	.w1(32'h3b6e484a),
	.w2(32'hba45fafa),
	.w3(32'h3c570020),
	.w4(32'h3aac50e5),
	.w5(32'h3c034be5),
	.w6(32'hbd0b0216),
	.w7(32'h3aab2164),
	.w8(32'h3bb5e9e6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be49ad0),
	.w1(32'hbc284884),
	.w2(32'hbb3338a7),
	.w3(32'h3ba5987d),
	.w4(32'h3b59fc8c),
	.w5(32'h3c345b63),
	.w6(32'h3af0ce6e),
	.w7(32'h3ad61650),
	.w8(32'h3bdeb292),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc182794),
	.w1(32'h3b3e3815),
	.w2(32'hbb3c4e05),
	.w3(32'h3adb43d3),
	.w4(32'hbbeb0b52),
	.w5(32'h3b9d8847),
	.w6(32'hbb50875a),
	.w7(32'hbb1794b0),
	.w8(32'h3a8bde3e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafea756),
	.w1(32'hbaf192a2),
	.w2(32'hbbc073d1),
	.w3(32'hbb298caf),
	.w4(32'hbb90e2f8),
	.w5(32'hb9a24620),
	.w6(32'hbc3dd1a4),
	.w7(32'h3bd2ed29),
	.w8(32'h3bb0d5f6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ca0b3),
	.w1(32'hbc19ecb1),
	.w2(32'hbcf7dbdf),
	.w3(32'h3bf30391),
	.w4(32'h3bc4a4ad),
	.w5(32'h3c6d1ca6),
	.w6(32'hb7de2347),
	.w7(32'h3ced88a2),
	.w8(32'h3cc51ec1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b3e42),
	.w1(32'hbc35f582),
	.w2(32'hbbed06ae),
	.w3(32'h3a8a65ec),
	.w4(32'hbbd608e7),
	.w5(32'hba8d5fc3),
	.w6(32'hbc34a401),
	.w7(32'h3be71007),
	.w8(32'h3c96a653),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc858149),
	.w1(32'hbbf6ad9a),
	.w2(32'h3bfbd689),
	.w3(32'h3b2a47eb),
	.w4(32'hbbf424a9),
	.w5(32'h3cd9225c),
	.w6(32'h3c605b29),
	.w7(32'hbc08d861),
	.w8(32'h3c414887),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52330d),
	.w1(32'hbb283990),
	.w2(32'h3adca337),
	.w3(32'h3b80dd06),
	.w4(32'h3a252fb5),
	.w5(32'hbb603c68),
	.w6(32'hbbacffb0),
	.w7(32'h3a76dd9d),
	.w8(32'h3c2ecc37),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ff85e),
	.w1(32'hbbfb8e1f),
	.w2(32'hbc20f16b),
	.w3(32'hbb126c00),
	.w4(32'hbbb72b6f),
	.w5(32'hbc2d2213),
	.w6(32'h3af374fb),
	.w7(32'h3a9d91c8),
	.w8(32'h3c2af314),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc689438),
	.w1(32'hbb3f78d9),
	.w2(32'hbcc2174f),
	.w3(32'hbbb53a36),
	.w4(32'hbb527ab8),
	.w5(32'hbc883e71),
	.w6(32'hbb9a95ed),
	.w7(32'h3a70fbf8),
	.w8(32'h3ccb2ee9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbe563),
	.w1(32'hbb15cd84),
	.w2(32'h3ba3dc53),
	.w3(32'hbc2600e4),
	.w4(32'hbc52bac9),
	.w5(32'h3c021872),
	.w6(32'h3c1fe276),
	.w7(32'hbb0e3710),
	.w8(32'hbb0bf2ab),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fc374),
	.w1(32'h3c12dc7d),
	.w2(32'h3c817e46),
	.w3(32'h3c0cf086),
	.w4(32'hbba0ee48),
	.w5(32'hbaab3328),
	.w6(32'hbbe32d3b),
	.w7(32'hbc607efa),
	.w8(32'hbbedfd73),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3918),
	.w1(32'h3a48219f),
	.w2(32'h3c1d9877),
	.w3(32'h3b527be8),
	.w4(32'h3916ec94),
	.w5(32'h3b70f7f1),
	.w6(32'hbc80cc47),
	.w7(32'hbbee26df),
	.w8(32'hbc5f3e69),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027dbc),
	.w1(32'hb94b475c),
	.w2(32'h3c02727e),
	.w3(32'h3b0cc165),
	.w4(32'hba5e215b),
	.w5(32'h3cae173b),
	.w6(32'hbbed2246),
	.w7(32'hbc29b2b1),
	.w8(32'h3be043c2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46c20e),
	.w1(32'hbc47d4ec),
	.w2(32'hbbaf4861),
	.w3(32'h3a54377f),
	.w4(32'hbaf0968a),
	.w5(32'hbc61ad57),
	.w6(32'h3c47c0e7),
	.w7(32'h3c48d5ad),
	.w8(32'h3c89a215),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28b2ad),
	.w1(32'hbc1db456),
	.w2(32'hbcbf61a5),
	.w3(32'hbc1f3b91),
	.w4(32'hbc1c13d0),
	.w5(32'hb7ac351d),
	.w6(32'h3c298311),
	.w7(32'h3c649faf),
	.w8(32'h3ce2507c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc530805),
	.w1(32'hba89f251),
	.w2(32'hbbc9e52e),
	.w3(32'hba88cf9e),
	.w4(32'hbc34034c),
	.w5(32'hbc37455e),
	.w6(32'h3c3908aa),
	.w7(32'hbba70888),
	.w8(32'h3bf9cce5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2df867),
	.w1(32'h3b8db5a4),
	.w2(32'hbbf3e4fd),
	.w3(32'h3b298128),
	.w4(32'hba516961),
	.w5(32'hbbac6812),
	.w6(32'h3be5899b),
	.w7(32'hbaa81244),
	.w8(32'hba4a1162),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18abb),
	.w1(32'hbb606385),
	.w2(32'hbc3db808),
	.w3(32'h3b870441),
	.w4(32'hbb7f69d1),
	.w5(32'hbc316546),
	.w6(32'h3ac868a5),
	.w7(32'hbc576a08),
	.w8(32'hbbef1b44),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b8042),
	.w1(32'hbb7032ce),
	.w2(32'hb88a74b7),
	.w3(32'hbc52a2cc),
	.w4(32'h3b112f37),
	.w5(32'h3c502b33),
	.w6(32'h3a4954f5),
	.w7(32'h399bc10e),
	.w8(32'h3c21eacc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65fd3f),
	.w1(32'hbbe90b90),
	.w2(32'hbc39b5e0),
	.w3(32'h3bc527b2),
	.w4(32'hbc13e9ce),
	.w5(32'hbc00b14f),
	.w6(32'h3c063bd2),
	.w7(32'h3bee7fa2),
	.w8(32'h3ca200ff),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca957),
	.w1(32'h3a1e87fa),
	.w2(32'hbbb93c3c),
	.w3(32'h3a8a7032),
	.w4(32'h3b4a9f05),
	.w5(32'h3afe2327),
	.w6(32'h3c32d3c5),
	.w7(32'h3b68add8),
	.w8(32'h3c0770ea),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e82b3),
	.w1(32'hbc033406),
	.w2(32'hbc2e9cd0),
	.w3(32'hbc0b3816),
	.w4(32'hbc0d1c16),
	.w5(32'hbc12cfc2),
	.w6(32'hbac1a5dc),
	.w7(32'h3b83968e),
	.w8(32'hbad1a5f3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0e89),
	.w1(32'hbbb3a2b7),
	.w2(32'hbb0b0692),
	.w3(32'hba713e63),
	.w4(32'h3b2f12d3),
	.w5(32'h3c49ebd3),
	.w6(32'hbab34c79),
	.w7(32'h3c6bd4c0),
	.w8(32'h3b20033d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85cc3d),
	.w1(32'hbb835ba3),
	.w2(32'hbb186a6a),
	.w3(32'hba150827),
	.w4(32'h3ad47bc6),
	.w5(32'h3c9fb80b),
	.w6(32'h3ba9a14d),
	.w7(32'h3b998127),
	.w8(32'h3be38f54),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99cbc5),
	.w1(32'hbb99450d),
	.w2(32'hbc016c13),
	.w3(32'h3c200602),
	.w4(32'h3b929b93),
	.w5(32'h39e0309d),
	.w6(32'hb936d5cd),
	.w7(32'h3be43734),
	.w8(32'h3ac61ffe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39990a8a),
	.w1(32'hbc482519),
	.w2(32'hbcd42d1a),
	.w3(32'hba1bc4c0),
	.w4(32'hbc64b484),
	.w5(32'hbbed4886),
	.w6(32'hbb266603),
	.w7(32'hbbdba831),
	.w8(32'h3c2478ef),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69ca11),
	.w1(32'hbc23b00f),
	.w2(32'hbc1d229a),
	.w3(32'h3c215764),
	.w4(32'hbc10d92d),
	.w5(32'h3beff7bc),
	.w6(32'h3cef05d1),
	.w7(32'h3b0b6386),
	.w8(32'hbbdcda08),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18e4a8),
	.w1(32'hbb6b2579),
	.w2(32'hbc1c1783),
	.w3(32'h3b9a10b1),
	.w4(32'hbb8c57de),
	.w5(32'h3bfbaeca),
	.w6(32'hbb893e07),
	.w7(32'h3afacb9d),
	.w8(32'h3c493776),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb92558),
	.w1(32'hbc5b24cc),
	.w2(32'hbca548ba),
	.w3(32'h3bce6370),
	.w4(32'hbc0b117f),
	.w5(32'h3ba642e8),
	.w6(32'h3c16c8a8),
	.w7(32'h3c4adfb1),
	.w8(32'h3a6cd297),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c9f2d),
	.w1(32'hbc3adec1),
	.w2(32'hbd03e8ab),
	.w3(32'hbbabf74f),
	.w4(32'hbc1979b2),
	.w5(32'hbcb4c444),
	.w6(32'hbb3e69cc),
	.w7(32'h3caa5068),
	.w8(32'h3d0c723c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca72000),
	.w1(32'h3a66f369),
	.w2(32'hbb7b31f6),
	.w3(32'hbc6eed02),
	.w4(32'h3b7bd339),
	.w5(32'h3bac3326),
	.w6(32'h3b30ae3e),
	.w7(32'hbada94c8),
	.w8(32'hbb186442),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe23058),
	.w1(32'hbbb49914),
	.w2(32'h3b83da4c),
	.w3(32'hb9e84d19),
	.w4(32'h3af84c4a),
	.w5(32'hbb9b1328),
	.w6(32'hbb07b8ed),
	.w7(32'h3bff899d),
	.w8(32'h3b3fe255),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43a586),
	.w1(32'h3ae19dd0),
	.w2(32'h3b696b5c),
	.w3(32'h3ac67410),
	.w4(32'hbbe76d41),
	.w5(32'h3c5f5a36),
	.w6(32'h3bb4c5d4),
	.w7(32'h3a8fb352),
	.w8(32'h3b8f4ae2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac166f6),
	.w1(32'h395e4e82),
	.w2(32'hbb356ec1),
	.w3(32'h3a71bb01),
	.w4(32'h3c42cf72),
	.w5(32'h3c6631c4),
	.w6(32'hb9333eb4),
	.w7(32'h3c922a94),
	.w8(32'h3c8d0ba3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ff8ac),
	.w1(32'hbb46497d),
	.w2(32'hba47bc72),
	.w3(32'h3bb4d521),
	.w4(32'hbb3a0161),
	.w5(32'hba01aa3d),
	.w6(32'h3b63b5f2),
	.w7(32'h3a80e355),
	.w8(32'h3b831ac7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe08480),
	.w1(32'h3b9479bf),
	.w2(32'h3b764659),
	.w3(32'h3af86286),
	.w4(32'h3bfc5874),
	.w5(32'hbc0aca48),
	.w6(32'h3c3fd822),
	.w7(32'h3ad0c4a1),
	.w8(32'h3bf711dc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c2252),
	.w1(32'h3b3fc85b),
	.w2(32'h3b6ca95f),
	.w3(32'hbbc5d5cb),
	.w4(32'hbb2088cc),
	.w5(32'hbb816569),
	.w6(32'h3be575b9),
	.w7(32'hbbc42bf7),
	.w8(32'hbbd9a89e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993a638),
	.w1(32'hbc24458d),
	.w2(32'hbc54716f),
	.w3(32'hbb6d2df7),
	.w4(32'h39997ae8),
	.w5(32'hbbd173a2),
	.w6(32'hba80ccc3),
	.w7(32'hb9998dd6),
	.w8(32'hbba1bed7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dc2d6),
	.w1(32'h3c615ef0),
	.w2(32'h3ca770d1),
	.w3(32'hb9ed51a8),
	.w4(32'h3b7c91bf),
	.w5(32'h39b572d1),
	.w6(32'h385878ca),
	.w7(32'hbc660c34),
	.w8(32'hbcfa8d10),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb20ddf),
	.w1(32'hbc5bd788),
	.w2(32'hbc7b9b7a),
	.w3(32'hbb2c36d3),
	.w4(32'hbc8fa000),
	.w5(32'hbca6457f),
	.w6(32'hbc6fdb64),
	.w7(32'hbbddfbca),
	.w8(32'h3c19a749),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca61249),
	.w1(32'h3b0d8cfb),
	.w2(32'hbb1234ec),
	.w3(32'hbc36d05d),
	.w4(32'hba8653a2),
	.w5(32'h3c428cbf),
	.w6(32'h3bbb225c),
	.w7(32'h3c10d1e9),
	.w8(32'h3c55595c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf37b33),
	.w1(32'hba68592c),
	.w2(32'h3b8809af),
	.w3(32'hbac886ca),
	.w4(32'hbb7997fd),
	.w5(32'hbc06a42a),
	.w6(32'h3c41a729),
	.w7(32'hbac89e0d),
	.w8(32'hbba5009a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace79d9),
	.w1(32'hbbc06641),
	.w2(32'hbbf27cf5),
	.w3(32'hbbbc3ee1),
	.w4(32'hb8bce3ec),
	.w5(32'h3bd8b254),
	.w6(32'hbbb975e6),
	.w7(32'h3b263234),
	.w8(32'h3b987354),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc75562),
	.w1(32'h3a9adbf7),
	.w2(32'hbb3acf66),
	.w3(32'h3b779fce),
	.w4(32'hbb0f144a),
	.w5(32'hbb22d8d3),
	.w6(32'h3b852cbe),
	.w7(32'h3b7810ac),
	.w8(32'h3c16c94c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf81d74),
	.w1(32'hbcfe7d5e),
	.w2(32'hbd5447ca),
	.w3(32'hbc1f0831),
	.w4(32'hbcd8b2b4),
	.w5(32'hbc93ba86),
	.w6(32'h3a268a88),
	.w7(32'h3b187d21),
	.w8(32'h3d43e58c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ba374),
	.w1(32'h3c6cffbe),
	.w2(32'h3b4862a6),
	.w3(32'hbcb3613e),
	.w4(32'h3be96034),
	.w5(32'hbb92eb90),
	.w6(32'h3ccfc658),
	.w7(32'h3c7118c1),
	.w8(32'h3c2c403a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f2a46),
	.w1(32'h3b2f6950),
	.w2(32'h3babd8d1),
	.w3(32'hbc88ed3d),
	.w4(32'h3b676b6f),
	.w5(32'h3ba901c1),
	.w6(32'hbc96b723),
	.w7(32'hbc03adfa),
	.w8(32'hbc8330dc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b217),
	.w1(32'hbc8eb27f),
	.w2(32'hbca73443),
	.w3(32'h3bbe46c6),
	.w4(32'hbc05edd1),
	.w5(32'hbc361174),
	.w6(32'hba6c5ea6),
	.w7(32'h3b90b8d3),
	.w8(32'h3c98bbc3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf8c2e),
	.w1(32'hbc6b1996),
	.w2(32'hbc288fd9),
	.w3(32'hbb18f020),
	.w4(32'hbc3a888e),
	.w5(32'h3acc543b),
	.w6(32'h3c97564c),
	.w7(32'hbbcafbff),
	.w8(32'h3b21b5af),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f757c),
	.w1(32'hbb7b48ff),
	.w2(32'hbaa889b6),
	.w3(32'hbb04c263),
	.w4(32'h3c085609),
	.w5(32'hbb9e5c15),
	.w6(32'h3a0b0f9c),
	.w7(32'h3b7c40c2),
	.w8(32'h3bc542e9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35976),
	.w1(32'hbbcf002d),
	.w2(32'hbbb1aa4b),
	.w3(32'h3b8debaa),
	.w4(32'hbbdac274),
	.w5(32'hbaa6e4b3),
	.w6(32'h3c0bc736),
	.w7(32'hbbe11f51),
	.w8(32'hbb28060f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb847f6),
	.w1(32'hbb38ed6b),
	.w2(32'hbc0a59bf),
	.w3(32'hbb52a9ad),
	.w4(32'hba7ce9f4),
	.w5(32'hbc3e898f),
	.w6(32'hbb0dc255),
	.w7(32'h3c0231f8),
	.w8(32'h3bad3871),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6275e7),
	.w1(32'h3b4bdc31),
	.w2(32'h3b1fa022),
	.w3(32'hbc554223),
	.w4(32'h3a1005e4),
	.w5(32'h3bd28a46),
	.w6(32'h3c1f3d08),
	.w7(32'h3bff33b9),
	.w8(32'h3b1e5c10),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8e090),
	.w1(32'hb7203eff),
	.w2(32'h3af06830),
	.w3(32'hbb7f3246),
	.w4(32'h3b2b5153),
	.w5(32'hbc154d4d),
	.w6(32'h3a5ba814),
	.w7(32'hbaa357a2),
	.w8(32'h3aeb6529),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f858cc),
	.w1(32'h3ade3d13),
	.w2(32'hbb8919ed),
	.w3(32'h3b1e6835),
	.w4(32'h3b275ea5),
	.w5(32'hbb6b9be5),
	.w6(32'h3c35630a),
	.w7(32'h3babf58f),
	.w8(32'hbbbdc016),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e426),
	.w1(32'hbc1c324d),
	.w2(32'hbc2cf6b0),
	.w3(32'h3a863812),
	.w4(32'hb9c8ed0a),
	.w5(32'h3bfc3238),
	.w6(32'hbc0b40f5),
	.w7(32'h3ba2210b),
	.w8(32'h3ba1708e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc775cf4),
	.w1(32'hbbdbfdd4),
	.w2(32'h37397b22),
	.w3(32'hbb9d8c38),
	.w4(32'hbba76a87),
	.w5(32'h3c0008fa),
	.w6(32'h3b072f78),
	.w7(32'hb9a6ba82),
	.w8(32'h3b84d9bb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaa3e9),
	.w1(32'h3c782874),
	.w2(32'h3cb6df05),
	.w3(32'h3c339803),
	.w4(32'h3bc8134a),
	.w5(32'h3b463191),
	.w6(32'h3c217f9f),
	.w7(32'hbbd6d348),
	.w8(32'hbcb8457c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb82a08),
	.w1(32'hbc4b26bc),
	.w2(32'hbca086fe),
	.w3(32'h38c81c8e),
	.w4(32'hbb90f728),
	.w5(32'hbb81660f),
	.w6(32'hbcae09d4),
	.w7(32'h3c569787),
	.w8(32'h3cad1a6c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc860a6c),
	.w1(32'hbc26f3f5),
	.w2(32'hb8c29613),
	.w3(32'hbc417b70),
	.w4(32'hbc55c2c9),
	.w5(32'h3b16dfea),
	.w6(32'h3c19c2f8),
	.w7(32'hbb5d9bf9),
	.w8(32'h3be7ef42),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b74b3),
	.w1(32'hbbcdfac3),
	.w2(32'hbc60ee8f),
	.w3(32'h39bdee05),
	.w4(32'h3af73e4c),
	.w5(32'h39957d1a),
	.w6(32'hbb813047),
	.w7(32'h3c27719e),
	.w8(32'h3be12aef),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866923),
	.w1(32'h3be8e33b),
	.w2(32'h3b8b2a2c),
	.w3(32'h39d9d1ec),
	.w4(32'h3b5f7cd5),
	.w5(32'h3c32f61e),
	.w6(32'h3b4d71bb),
	.w7(32'hbbcd483c),
	.w8(32'hbb4200ad),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba753f7),
	.w1(32'h3b4d2861),
	.w2(32'hbbadc5b9),
	.w3(32'h3be77e4e),
	.w4(32'hbc6df974),
	.w5(32'hbcb8731c),
	.w6(32'h3a763b0b),
	.w7(32'h3c28c9fb),
	.w8(32'h3a9fb63a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b398a4a),
	.w1(32'h3b8a2901),
	.w2(32'h3c37993f),
	.w3(32'hbc490d2b),
	.w4(32'hbbeecf14),
	.w5(32'hbc868710),
	.w6(32'h3adc130d),
	.w7(32'hbb8773f4),
	.w8(32'hbbed9c38),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c144e94),
	.w1(32'h3a30489b),
	.w2(32'hbbbfe15b),
	.w3(32'hbb8b8644),
	.w4(32'hbbafc994),
	.w5(32'hbc882c41),
	.w6(32'h3b864b59),
	.w7(32'h3b641473),
	.w8(32'h3bea97ba),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943e26),
	.w1(32'hbb326557),
	.w2(32'hba7af1d8),
	.w3(32'hbb8194e6),
	.w4(32'hbb4ca74e),
	.w5(32'h3bd331d0),
	.w6(32'h3b76bdcc),
	.w7(32'hbc767c37),
	.w8(32'hbb2ead9f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a939e),
	.w1(32'h3b73e92c),
	.w2(32'h3bdceb8f),
	.w3(32'hbbced9be),
	.w4(32'hbb48cfdf),
	.w5(32'hb9210bdb),
	.w6(32'h3c131a41),
	.w7(32'hbc330d1e),
	.w8(32'hbb40ef6a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e40a0),
	.w1(32'h3a1ff293),
	.w2(32'hbc980445),
	.w3(32'hbb8a1113),
	.w4(32'hbbec0c3f),
	.w5(32'hbb09320b),
	.w6(32'h3b85221d),
	.w7(32'hbbab69bb),
	.w8(32'h3cc423a1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24bf89),
	.w1(32'hbb9eb85b),
	.w2(32'hbc9b7d80),
	.w3(32'hbbd15f6d),
	.w4(32'hba43c257),
	.w5(32'hba910798),
	.w6(32'h3c44b936),
	.w7(32'h3bd1159b),
	.w8(32'h3c519967),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e4f5f),
	.w1(32'hbc038255),
	.w2(32'hba2345d9),
	.w3(32'hbb64de02),
	.w4(32'hbca519b4),
	.w5(32'hbc25c5ad),
	.w6(32'hbb8ea58d),
	.w7(32'h3a370ea0),
	.w8(32'h3c5bb6aa),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b7233),
	.w1(32'hbca071e5),
	.w2(32'hbd2a1d7f),
	.w3(32'hbc6ebdbd),
	.w4(32'hbc7ad505),
	.w5(32'hbca151a2),
	.w6(32'h3b8d3067),
	.w7(32'h3a90ad3c),
	.w8(32'h3d3cc8be),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9762d7),
	.w1(32'h3b46515f),
	.w2(32'hbbc02610),
	.w3(32'hbc8cb992),
	.w4(32'h3c140e73),
	.w5(32'h3ab15880),
	.w6(32'h3bbe3e17),
	.w7(32'h3c0dbd17),
	.w8(32'h3c4d6ac2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a6b09),
	.w1(32'hbb8ac584),
	.w2(32'hbbdd4754),
	.w3(32'hba4f888d),
	.w4(32'h3aa0e7d0),
	.w5(32'hbce68b20),
	.w6(32'h3c1575c1),
	.w7(32'h3c99d184),
	.w8(32'h3c4f124a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc695791),
	.w1(32'hbc00096e),
	.w2(32'hbc867ca7),
	.w3(32'hbca01ec4),
	.w4(32'hbaaa1132),
	.w5(32'hbc038b26),
	.w6(32'h3c70e995),
	.w7(32'h3be40d9b),
	.w8(32'h3c91265b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc842d7a),
	.w1(32'hbad27672),
	.w2(32'hbbec3a91),
	.w3(32'hbc2f91c7),
	.w4(32'hbabbbdb2),
	.w5(32'hbc20b40b),
	.w6(32'h3bd54c23),
	.w7(32'hb82917bf),
	.w8(32'hbc05baac),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb415a0c),
	.w1(32'h3b93ce56),
	.w2(32'h3beb3a5e),
	.w3(32'hbc1c01fe),
	.w4(32'h3b8c00eb),
	.w5(32'h3b668722),
	.w6(32'hbb47897f),
	.w7(32'hbc112f7a),
	.w8(32'hbc9b0e15),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71578b),
	.w1(32'h3c28d6e2),
	.w2(32'h3c515e47),
	.w3(32'h3a9808aa),
	.w4(32'h3c9c2213),
	.w5(32'h3b3dd146),
	.w6(32'hbc827941),
	.w7(32'h3c37f143),
	.w8(32'hbb52c218),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16f0fa),
	.w1(32'hbb9b85ea),
	.w2(32'hbbd34a78),
	.w3(32'h3b94009f),
	.w4(32'h398dd66a),
	.w5(32'hba62ddf7),
	.w6(32'h3b41c325),
	.w7(32'h3b80b40a),
	.w8(32'hbb804cbb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a1c6),
	.w1(32'hbafba99c),
	.w2(32'hb96733c3),
	.w3(32'h3b08574b),
	.w4(32'hbaabc9cb),
	.w5(32'h3c02d6cb),
	.w6(32'h3b9f0475),
	.w7(32'hb9ae6553),
	.w8(32'hbc3808e0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab679b1),
	.w1(32'hbbd8fc53),
	.w2(32'hbc3321d0),
	.w3(32'h3c1f68a8),
	.w4(32'h3b08cd86),
	.w5(32'h3bfc779a),
	.w6(32'hbbf4855c),
	.w7(32'h3be0c394),
	.w8(32'h3c166557),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670a05),
	.w1(32'h3ab25bba),
	.w2(32'h3bae39fb),
	.w3(32'hbb9ecdde),
	.w4(32'h3b01087e),
	.w5(32'hbc77da6b),
	.w6(32'h3b7e85ac),
	.w7(32'h3bc5240b),
	.w8(32'hbb766294),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b080511),
	.w1(32'h3c8769e7),
	.w2(32'h3c275457),
	.w3(32'hbad6ed0f),
	.w4(32'h39500250),
	.w5(32'hbb33a130),
	.w6(32'hbafe8cf7),
	.w7(32'hbc119027),
	.w8(32'hbc22bf56),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90a805),
	.w1(32'hbc18c9f5),
	.w2(32'h3b056ef6),
	.w3(32'h3b1fe08f),
	.w4(32'hbb3d7b32),
	.w5(32'h3be4c9ea),
	.w6(32'hbba4cdc0),
	.w7(32'hbadd3b22),
	.w8(32'hbb6c3369),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff2a91),
	.w1(32'h3b0ac0e3),
	.w2(32'hb9e3eb68),
	.w3(32'h3bebd0d0),
	.w4(32'hbb80db96),
	.w5(32'hbb041046),
	.w6(32'h3b143f88),
	.w7(32'h3b4b3086),
	.w8(32'hbb872f12),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b403316),
	.w1(32'h39e46cae),
	.w2(32'hbafba049),
	.w3(32'h3b3e6954),
	.w4(32'hbb8f2484),
	.w5(32'hbb2ebeba),
	.w6(32'h3b9bd2fd),
	.w7(32'hba64b8e2),
	.w8(32'h3bf0bf2a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1412),
	.w1(32'hbbeb3203),
	.w2(32'hbbe99f10),
	.w3(32'h3b46a593),
	.w4(32'hbb7888e4),
	.w5(32'hbba4814f),
	.w6(32'h3bef11d6),
	.w7(32'hbb8258d0),
	.w8(32'hbaee919c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068ab1),
	.w1(32'hbbe79311),
	.w2(32'hb9d20550),
	.w3(32'h3a4d92e7),
	.w4(32'h3a986630),
	.w5(32'hbba57a66),
	.w6(32'h3bc5dcec),
	.w7(32'h3a9767b1),
	.w8(32'h3b7f1cbf),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b2b9),
	.w1(32'hbb53a9db),
	.w2(32'hbb5e0bbb),
	.w3(32'h3ab7aa0a),
	.w4(32'h39052f5c),
	.w5(32'hbb8fa37e),
	.w6(32'h3c431521),
	.w7(32'h3b32e31b),
	.w8(32'h3abc874f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae86025),
	.w1(32'hbb58f762),
	.w2(32'h3ae023e5),
	.w3(32'hbab5f0f4),
	.w4(32'h3b7e2022),
	.w5(32'hbc4f648e),
	.w6(32'h3bfcb326),
	.w7(32'h3bde1af7),
	.w8(32'h3b51efac),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f957a),
	.w1(32'h3ba5a12d),
	.w2(32'h3c4013a3),
	.w3(32'hbb942763),
	.w4(32'h3c465d43),
	.w5(32'h39b454d0),
	.w6(32'h3b0682d5),
	.w7(32'h3b59d532),
	.w8(32'hbb9fc095),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa94666),
	.w1(32'hbae63e3d),
	.w2(32'hbb078ecf),
	.w3(32'h39c247b6),
	.w4(32'h3b4653bf),
	.w5(32'h3a7ae2f9),
	.w6(32'hbc3bb4f0),
	.w7(32'h3ba90829),
	.w8(32'hbc19c93d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8410),
	.w1(32'h3c1b18b2),
	.w2(32'h3b84d291),
	.w3(32'hbb67f41b),
	.w4(32'h3c86ce78),
	.w5(32'hbb211235),
	.w6(32'hbab8f0cb),
	.w7(32'h3b60cfc5),
	.w8(32'hbb7b5273),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27414),
	.w1(32'hbc22c4d1),
	.w2(32'hbc325839),
	.w3(32'h3c0472aa),
	.w4(32'hbc1dea2a),
	.w5(32'h3c3f6b37),
	.w6(32'hbb06c8ed),
	.w7(32'h3af7ab31),
	.w8(32'h3cd6b3dd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4db664),
	.w1(32'hba9ccd3a),
	.w2(32'hbc3d74cd),
	.w3(32'h3a156725),
	.w4(32'h3841881e),
	.w5(32'hbb99f8a7),
	.w6(32'h3bcefe3f),
	.w7(32'h3c0b1a09),
	.w8(32'h3c0ea84e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16388d),
	.w1(32'h3c4d6bb2),
	.w2(32'h3c2453b5),
	.w3(32'h3a1a5296),
	.w4(32'hbb523916),
	.w5(32'hba843dab),
	.w6(32'h3bee4127),
	.w7(32'hbb13f516),
	.w8(32'hba68810c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07dd6a),
	.w1(32'h3a67cc19),
	.w2(32'h3c564b48),
	.w3(32'h3b7f5cf2),
	.w4(32'hbaab8e0f),
	.w5(32'h3aac6bec),
	.w6(32'hba850109),
	.w7(32'hbb43473e),
	.w8(32'hbc46a82a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9bc85),
	.w1(32'hba34ca46),
	.w2(32'hbbb85176),
	.w3(32'hbafb980c),
	.w4(32'hbc85a428),
	.w5(32'hbc373729),
	.w6(32'hbc355972),
	.w7(32'hbafdcde7),
	.w8(32'h3c25220d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e557a),
	.w1(32'h3b1c6d03),
	.w2(32'hbb1a040c),
	.w3(32'hbbdd1e25),
	.w4(32'h3c09a5a2),
	.w5(32'h3b80e264),
	.w6(32'h3c8602a8),
	.w7(32'hbb84a48e),
	.w8(32'hbadf2112),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc135a48),
	.w1(32'h3c339bd9),
	.w2(32'h3cb447e0),
	.w3(32'h3be5ed63),
	.w4(32'h3b6f491a),
	.w5(32'hbac719ae),
	.w6(32'h3c57898e),
	.w7(32'hbbfc37df),
	.w8(32'hbc855100),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc12f7),
	.w1(32'hbbe60f74),
	.w2(32'h3af02748),
	.w3(32'hbb04f96a),
	.w4(32'hbb2de42d),
	.w5(32'h3c2f7b30),
	.w6(32'hbc818588),
	.w7(32'hbb44adf3),
	.w8(32'h3b5cceba),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae27ffa),
	.w1(32'hbbd2c78a),
	.w2(32'hbc847486),
	.w3(32'h3c33d4d1),
	.w4(32'hbc0aa6aa),
	.w5(32'hbbcb0e8f),
	.w6(32'h3b2f3b51),
	.w7(32'h3b9fe2d6),
	.w8(32'h3c69eedf),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210131),
	.w1(32'hbc113ed2),
	.w2(32'hbb90e849),
	.w3(32'hbb9cee5b),
	.w4(32'hbb0e182e),
	.w5(32'hbbfa15a6),
	.w6(32'h3af677d5),
	.w7(32'h3c5e3a56),
	.w8(32'h3c2f7125),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8949e3),
	.w1(32'hbb473a16),
	.w2(32'hbc3f2aaf),
	.w3(32'h3baa2f6d),
	.w4(32'hbbf58efd),
	.w5(32'hbc6a8f0c),
	.w6(32'h3c784633),
	.w7(32'h3bab0263),
	.w8(32'hb88b496a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d3ce9),
	.w1(32'hbc96138e),
	.w2(32'hbc94b5cc),
	.w3(32'hbc1d5ff0),
	.w4(32'hbc3238da),
	.w5(32'hbbad350b),
	.w6(32'h3ab22f6a),
	.w7(32'h3ab2f909),
	.w8(32'h3d1bbeb0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4d939),
	.w1(32'hb82d1976),
	.w2(32'hbbfce607),
	.w3(32'hbba3815f),
	.w4(32'h399159c5),
	.w5(32'hbae29bde),
	.w6(32'hbbfd276f),
	.w7(32'hbae916b4),
	.w8(32'h3c5de7c3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed73b6),
	.w1(32'hbcfa16fd),
	.w2(32'hbd087c3a),
	.w3(32'hbb3b7b81),
	.w4(32'hbc99ac60),
	.w5(32'h3ab65c0f),
	.w6(32'hbb080e02),
	.w7(32'hbc54abe8),
	.w8(32'h3ce7fe1b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00a5b),
	.w1(32'h3963794f),
	.w2(32'h3b7ad472),
	.w3(32'h3bdcea6f),
	.w4(32'hbc00e16a),
	.w5(32'hbc8b943b),
	.w6(32'h3ceb9e63),
	.w7(32'hba62be1a),
	.w8(32'h3b825f5a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad25724),
	.w1(32'hbb9049ec),
	.w2(32'hbbda4f44),
	.w3(32'hbba0968b),
	.w4(32'hbb383899),
	.w5(32'hba7a0882),
	.w6(32'h3c754680),
	.w7(32'h3b0beca4),
	.w8(32'hbb678dcd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21ce9),
	.w1(32'hbba90474),
	.w2(32'hbc50dbb4),
	.w3(32'h3b47d1f8),
	.w4(32'hbab50c93),
	.w5(32'hbc523ac9),
	.w6(32'h38dd10e8),
	.w7(32'h3b698d76),
	.w8(32'h3cc026e0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7063e9),
	.w1(32'h3b86b499),
	.w2(32'h3b974b2d),
	.w3(32'hbb4ccf78),
	.w4(32'h3b4089a6),
	.w5(32'h3b9861bf),
	.w6(32'h3ca5a5aa),
	.w7(32'hbbbef016),
	.w8(32'hbbd5de35),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f1df7),
	.w1(32'h3c9f44a9),
	.w2(32'h3cf0be40),
	.w3(32'hbb919d54),
	.w4(32'hb9e21bbd),
	.w5(32'hbbb854e9),
	.w6(32'hbbb2d381),
	.w7(32'hbc0122e7),
	.w8(32'hbcf346a3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c8db8),
	.w1(32'h3bd9633b),
	.w2(32'h3c86320b),
	.w3(32'hbb6d0944),
	.w4(32'hbab5c181),
	.w5(32'hbb75776c),
	.w6(32'hbc1cf0ea),
	.w7(32'hba482a9f),
	.w8(32'hbcb057c4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dce21),
	.w1(32'hbc476719),
	.w2(32'hbc89d3e8),
	.w3(32'h3b848025),
	.w4(32'hba1c1ddb),
	.w5(32'h3c9357df),
	.w6(32'hbc03b9f2),
	.w7(32'h3c07efbd),
	.w8(32'h3bc1d50d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bae7b),
	.w1(32'hbc0c2519),
	.w2(32'hbc8fa53f),
	.w3(32'hbac7e8fe),
	.w4(32'hbbb07904),
	.w5(32'hbc04e122),
	.w6(32'h3ba3b23c),
	.w7(32'h3c23b266),
	.w8(32'h3cc779fb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76608d),
	.w1(32'hbbedb8de),
	.w2(32'hbc447bbf),
	.w3(32'hbb827780),
	.w4(32'hbba1192c),
	.w5(32'hbb0ba2d0),
	.w6(32'h3cc5a9dd),
	.w7(32'h3bdb5074),
	.w8(32'h3c835c0a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308e7b),
	.w1(32'h3a6967ce),
	.w2(32'h3b2b675d),
	.w3(32'hbaf2dd90),
	.w4(32'h3aa1a816),
	.w5(32'h3b9917dc),
	.w6(32'h3a8d636f),
	.w7(32'h3b56543f),
	.w8(32'h3a35f9ab),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e738),
	.w1(32'hba128816),
	.w2(32'h3af83829),
	.w3(32'hbb92b256),
	.w4(32'h3ab8d011),
	.w5(32'h3c04bb5e),
	.w6(32'hbbb793dd),
	.w7(32'h3b601e55),
	.w8(32'h3aed59ef),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b33f),
	.w1(32'hbb386af5),
	.w2(32'hbaa9cda4),
	.w3(32'hba12621c),
	.w4(32'hbb779b89),
	.w5(32'hbbb9b120),
	.w6(32'hbb2190a3),
	.w7(32'hbb04710e),
	.w8(32'h3a0c1421),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09abf3),
	.w1(32'h3b63d81b),
	.w2(32'h3bbcaaf1),
	.w3(32'h3aedffc6),
	.w4(32'h3ae323d9),
	.w5(32'hbaa5f8b2),
	.w6(32'h3bc8266b),
	.w7(32'hba624bbc),
	.w8(32'h39e5f7a3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d47c0),
	.w1(32'hbb00ddbd),
	.w2(32'hba9b675f),
	.w3(32'h3b4a6e85),
	.w4(32'hbb4b10aa),
	.w5(32'hbaadfadb),
	.w6(32'h3b1a1c67),
	.w7(32'hbb1b9c1c),
	.w8(32'h3aaeb7a4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d626),
	.w1(32'h3b69fd82),
	.w2(32'h3b48fcb5),
	.w3(32'hb9305d40),
	.w4(32'hbb3a5b59),
	.w5(32'h3b093671),
	.w6(32'h3b281608),
	.w7(32'hbabe04d1),
	.w8(32'h3a0de1d7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14a782),
	.w1(32'hbbc4bddf),
	.w2(32'hbb0aeb24),
	.w3(32'h3b543a4a),
	.w4(32'hb994ccb6),
	.w5(32'h3a333c34),
	.w6(32'hbb958bf2),
	.w7(32'hbb5a93d9),
	.w8(32'hbb85a221),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb18684),
	.w1(32'hbbf9d051),
	.w2(32'hbc07f895),
	.w3(32'hb98d2aab),
	.w4(32'hbc10a947),
	.w5(32'hbb9bd6d8),
	.w6(32'hba8e6f70),
	.w7(32'hbc159f84),
	.w8(32'hbbe47267),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d8333),
	.w1(32'hbbaddff7),
	.w2(32'h3b1c4ecd),
	.w3(32'hbc1a39ac),
	.w4(32'hb6359152),
	.w5(32'hbac32520),
	.w6(32'hbc02e526),
	.w7(32'hbaf490c5),
	.w8(32'h3a8b06f7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5164e0),
	.w1(32'hbada7749),
	.w2(32'hbaf58387),
	.w3(32'hbbf72220),
	.w4(32'h3aca5a52),
	.w5(32'h3ac6601f),
	.w6(32'hbbcc7d64),
	.w7(32'hbb6874ca),
	.w8(32'h3aa9895d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba321856),
	.w1(32'hb99ca492),
	.w2(32'hb942282f),
	.w3(32'h3aa72cb6),
	.w4(32'h3a146c68),
	.w5(32'h3b721c2b),
	.w6(32'hb9b04901),
	.w7(32'hbaa43b16),
	.w8(32'h3b2bae08),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8201a0),
	.w1(32'h3b2607ce),
	.w2(32'h3b686c33),
	.w3(32'hbba3373f),
	.w4(32'h3bb5ee8d),
	.w5(32'hba242dc7),
	.w6(32'h3ae4fdf6),
	.w7(32'h3b6637ff),
	.w8(32'h3b753aac),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2c423),
	.w1(32'hb9e862af),
	.w2(32'h3b82acd5),
	.w3(32'h3ba2b4c6),
	.w4(32'hb9bf783e),
	.w5(32'h3bad3eec),
	.w6(32'h3bf26874),
	.w7(32'hb9650d93),
	.w8(32'h3b048efc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d123),
	.w1(32'h3944ab1c),
	.w2(32'h3aab2c21),
	.w3(32'h3b1d8286),
	.w4(32'hbab50090),
	.w5(32'h3ab9902e),
	.w6(32'h3b24d215),
	.w7(32'hba8c5707),
	.w8(32'hba699b83),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0557aa),
	.w1(32'h3c1413fe),
	.w2(32'h3c592d1c),
	.w3(32'h3b29105c),
	.w4(32'h3c13a4c1),
	.w5(32'h3caf4e89),
	.w6(32'h3b8d9b08),
	.w7(32'h3c805074),
	.w8(32'h3ce088fd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd91a3d),
	.w1(32'h3a80c5df),
	.w2(32'h3bd8edd1),
	.w3(32'h3cdf864f),
	.w4(32'hba576a81),
	.w5(32'h3b8628f1),
	.w6(32'h3c441e89),
	.w7(32'h3b301b75),
	.w8(32'h3bbc6875),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09e4a9),
	.w1(32'hbab2b1df),
	.w2(32'h39fc2ede),
	.w3(32'h3b884d13),
	.w4(32'hbb17968d),
	.w5(32'h3c3e3df3),
	.w6(32'h3bfce61c),
	.w7(32'h3a969369),
	.w8(32'h3adc848c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8972f),
	.w1(32'hba562946),
	.w2(32'hbb2abd33),
	.w3(32'hbb4d82ba),
	.w4(32'h3b848779),
	.w5(32'hbb46453b),
	.w6(32'h3a18c9f4),
	.w7(32'hbad78dde),
	.w8(32'h3a359813),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e8fbd),
	.w1(32'hba9341fe),
	.w2(32'hbbd87c6f),
	.w3(32'hba616b4d),
	.w4(32'hbac6c4a2),
	.w5(32'hbbf5c3f5),
	.w6(32'h3b221398),
	.w7(32'hbb1b3866),
	.w8(32'h3b3d7a45),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba519eaa),
	.w1(32'hb907decd),
	.w2(32'hbaa7efac),
	.w3(32'h3a427812),
	.w4(32'h390173a0),
	.w5(32'hbb5dbc4e),
	.w6(32'h3b422c9a),
	.w7(32'hbae4f0fc),
	.w8(32'hbb7361fd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5b34f),
	.w1(32'hbab4cb2d),
	.w2(32'h3b097df6),
	.w3(32'h3bed7286),
	.w4(32'h36d1e551),
	.w5(32'h3b1545b6),
	.w6(32'h3abd5fd9),
	.w7(32'hbb0d69af),
	.w8(32'hba67d027),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf268),
	.w1(32'hbb9160ca),
	.w2(32'hb8c72868),
	.w3(32'hbb76424c),
	.w4(32'hbc04badd),
	.w5(32'hbada19e9),
	.w6(32'hbaf19976),
	.w7(32'hbbe0984a),
	.w8(32'hbae18400),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc5701),
	.w1(32'hbaf82d57),
	.w2(32'hbac0413d),
	.w3(32'h3bd63b66),
	.w4(32'hbb4537ce),
	.w5(32'h3ba11f21),
	.w6(32'h3b8c7ed1),
	.w7(32'h3b04d2a3),
	.w8(32'hb971b936),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e84de),
	.w1(32'h3b37730d),
	.w2(32'h39222a38),
	.w3(32'h3b3b69a1),
	.w4(32'h3b27607c),
	.w5(32'h3a4f0a86),
	.w6(32'hbb81bbec),
	.w7(32'h3a9c57c7),
	.w8(32'hba085e8a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26a473),
	.w1(32'hbb060973),
	.w2(32'h3b09a3b9),
	.w3(32'h3ab1b189),
	.w4(32'h3ad66968),
	.w5(32'h3aa1b4f5),
	.w6(32'h3b212a03),
	.w7(32'h3a5a4a5d),
	.w8(32'h38231060),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73fdce),
	.w1(32'hbae9b44f),
	.w2(32'hbb4273be),
	.w3(32'h3b3bb157),
	.w4(32'h3b04458d),
	.w5(32'h3be1159f),
	.w6(32'h3b832c7b),
	.w7(32'h3a1ea227),
	.w8(32'h3c4524b0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2ebca),
	.w1(32'h3a817faa),
	.w2(32'h3aba8737),
	.w3(32'h3c2bf7d3),
	.w4(32'h3a07c35e),
	.w5(32'hbaa17fdf),
	.w6(32'h3b2b4812),
	.w7(32'h39c31a3d),
	.w8(32'h3b6f7035),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54620c),
	.w1(32'hbb3fa021),
	.w2(32'hbaf037cf),
	.w3(32'hb9d31aa6),
	.w4(32'hbb287df6),
	.w5(32'h3c178957),
	.w6(32'h3b64383b),
	.w7(32'h3a9e0c79),
	.w8(32'h3bcea5f1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9fc7b),
	.w1(32'hba0f40ca),
	.w2(32'h3bff6953),
	.w3(32'h3b2fd0c0),
	.w4(32'hbac12100),
	.w5(32'h3bb89f9d),
	.w6(32'h38a3d805),
	.w7(32'h3b27c75d),
	.w8(32'h3bcd5c99),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb826e841),
	.w1(32'h3a35fc23),
	.w2(32'h3b9acd29),
	.w3(32'hbb55636d),
	.w4(32'h3b267a4b),
	.w5(32'hbb0d0b41),
	.w6(32'h3a5e3977),
	.w7(32'h3a6666ab),
	.w8(32'hbbb1ab76),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886649),
	.w1(32'h3ba0bb7f),
	.w2(32'h3acac1b5),
	.w3(32'h39bd9dd2),
	.w4(32'hbb7cb25e),
	.w5(32'h3a80f148),
	.w6(32'hb8a75e5d),
	.w7(32'h39c1f5c2),
	.w8(32'h3b7aada2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2df164),
	.w1(32'hbacbc7af),
	.w2(32'hbac19b70),
	.w3(32'h398f8373),
	.w4(32'h3a8b3f24),
	.w5(32'h3a5cf48b),
	.w6(32'h3bb649ea),
	.w7(32'hbaffb376),
	.w8(32'h3b41a426),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75a293),
	.w1(32'hba599562),
	.w2(32'hbb4bb5da),
	.w3(32'h3bb81659),
	.w4(32'hbb3cd010),
	.w5(32'h3bcb2d8f),
	.w6(32'h3b76991a),
	.w7(32'h3ab26d64),
	.w8(32'h390a6878),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af79a40),
	.w1(32'h3b317fd6),
	.w2(32'h3b29b857),
	.w3(32'hbab71f82),
	.w4(32'hbaac4fd8),
	.w5(32'h39147600),
	.w6(32'h3ae9915e),
	.w7(32'h3a18de23),
	.w8(32'h3b4a6fca),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddc571),
	.w1(32'hbb16dac8),
	.w2(32'hb94016a3),
	.w3(32'h3b44918c),
	.w4(32'hba2f68d0),
	.w5(32'hb81de64e),
	.w6(32'h3abdd892),
	.w7(32'hbaf26346),
	.w8(32'h3aa8177a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f7b5a),
	.w1(32'hbaadcd02),
	.w2(32'hbbaf6df8),
	.w3(32'hbb8b4027),
	.w4(32'hb9a840de),
	.w5(32'hbaad93b1),
	.w6(32'h38e3e152),
	.w7(32'h3ac5b2c2),
	.w8(32'h3b97d511),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed009b),
	.w1(32'hba6ac9eb),
	.w2(32'h3944d08b),
	.w3(32'h3b432a72),
	.w4(32'hb9c49ae7),
	.w5(32'h3a7ab432),
	.w6(32'h3a815094),
	.w7(32'h3a699b08),
	.w8(32'h3a062c0e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85ae09),
	.w1(32'h3ae310b9),
	.w2(32'h3afd8071),
	.w3(32'h3b8ade53),
	.w4(32'hba98fb29),
	.w5(32'h3bbea032),
	.w6(32'h3b4d2423),
	.w7(32'hbaf1cb27),
	.w8(32'hbabebdcb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e89b0),
	.w1(32'h3ab04862),
	.w2(32'hb9598af2),
	.w3(32'hba9ecd97),
	.w4(32'hbb16e49d),
	.w5(32'h3af54de9),
	.w6(32'hbb1e158a),
	.w7(32'h3a48f012),
	.w8(32'h3b7d92f1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb776866),
	.w1(32'hbbcdbe36),
	.w2(32'hbb1b11a5),
	.w3(32'hb95e5cd8),
	.w4(32'hbb8303b8),
	.w5(32'hbb67000f),
	.w6(32'h3a516e2e),
	.w7(32'hbb3237a2),
	.w8(32'hbb68f1c3),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e35e6),
	.w1(32'hbb69cd42),
	.w2(32'hbb366037),
	.w3(32'hbacfa6d4),
	.w4(32'h3a0f8d18),
	.w5(32'hba75c713),
	.w6(32'h3acb4dcc),
	.w7(32'h3b2a4d69),
	.w8(32'h39ad7d02),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1948a4),
	.w1(32'hbb32e58e),
	.w2(32'h3c67959a),
	.w3(32'h3b4957e3),
	.w4(32'h3bd89d68),
	.w5(32'h3bf88d33),
	.w6(32'hb9c8a357),
	.w7(32'h3b05d50a),
	.w8(32'hbbd1aa05),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33e399),
	.w1(32'h3ac705dd),
	.w2(32'h3b9d081e),
	.w3(32'hbb857974),
	.w4(32'h3a55e446),
	.w5(32'h3bb08422),
	.w6(32'hbb2d357f),
	.w7(32'h3b1bdc98),
	.w8(32'h3b35f5bc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc727ca),
	.w1(32'h38c37a3a),
	.w2(32'h38b92cfd),
	.w3(32'hba13708c),
	.w4(32'hbb3255ba),
	.w5(32'hba1f8b9f),
	.w6(32'hba445baa),
	.w7(32'hbac20a5a),
	.w8(32'h3a98cd00),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba996950),
	.w1(32'hbb8bb775),
	.w2(32'hbbbdab78),
	.w3(32'hbb24c162),
	.w4(32'hbb8b5d0c),
	.w5(32'h3a0b31b6),
	.w6(32'hbb51df22),
	.w7(32'hbb7fd27b),
	.w8(32'hbb1ad0da),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc5f89),
	.w1(32'h3ba46df2),
	.w2(32'hbace340f),
	.w3(32'h3aa7d49a),
	.w4(32'h3b208e05),
	.w5(32'hbb1f3123),
	.w6(32'hba53cfb9),
	.w7(32'h3a8d3093),
	.w8(32'h3b0209ec),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae44c5d),
	.w1(32'hbbfeb380),
	.w2(32'hbaac409e),
	.w3(32'hbadcf7d5),
	.w4(32'hbbd85b13),
	.w5(32'h3bf82847),
	.w6(32'h3a0ffcae),
	.w7(32'hbb895c71),
	.w8(32'h3abaef2e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec200),
	.w1(32'hbaad2d0e),
	.w2(32'h3b8deae5),
	.w3(32'h3a879152),
	.w4(32'hbb6ac4bc),
	.w5(32'h3abf39c3),
	.w6(32'h3a0789e5),
	.w7(32'hbb22599a),
	.w8(32'h3a53ebdf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009523),
	.w1(32'hbad734a4),
	.w2(32'h3b25ce71),
	.w3(32'h3bbed2cc),
	.w4(32'h3b05cadc),
	.w5(32'hba379126),
	.w6(32'h387750e1),
	.w7(32'h3a837235),
	.w8(32'hbae1aba8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dadc7),
	.w1(32'h3a242658),
	.w2(32'hbb1f1b21),
	.w3(32'h3ab61b02),
	.w4(32'hbac0ccec),
	.w5(32'hbbb44751),
	.w6(32'h3a4a1b95),
	.w7(32'hbb10eb1c),
	.w8(32'h3a8e0f7b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e83ba),
	.w1(32'hba2fbff0),
	.w2(32'h3aa182b6),
	.w3(32'hbb3613e3),
	.w4(32'hbb513756),
	.w5(32'h3aada207),
	.w6(32'h3afc31eb),
	.w7(32'hba63bd3a),
	.w8(32'h3a87a5eb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16716e),
	.w1(32'hbb73f906),
	.w2(32'hbb8ebc43),
	.w3(32'h3b40d22e),
	.w4(32'hbb9f3248),
	.w5(32'hbb918f5f),
	.w6(32'h3b8df391),
	.w7(32'hbbe3293e),
	.w8(32'hbba0f730),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecc5d0),
	.w1(32'hbbdbb8de),
	.w2(32'hbb7d8532),
	.w3(32'h3b22551a),
	.w4(32'hb98ae476),
	.w5(32'hb9cc235d),
	.w6(32'hbb37152b),
	.w7(32'hbac4fc59),
	.w8(32'hbb2b3c3e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab01064),
	.w1(32'hbb0362f7),
	.w2(32'hbafdda87),
	.w3(32'h3a85270e),
	.w4(32'hba59e6b5),
	.w5(32'h3b324408),
	.w6(32'hbbe1579b),
	.w7(32'hb98f5ac0),
	.w8(32'h3b56229b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4072b5),
	.w1(32'hbb579b1f),
	.w2(32'hbbce2f25),
	.w3(32'h3b2c5b4b),
	.w4(32'hbb07640f),
	.w5(32'hba74eee4),
	.w6(32'hba44c41d),
	.w7(32'hba662b40),
	.w8(32'hbb162df5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf59b70),
	.w1(32'hba21e596),
	.w2(32'h3b93a6d3),
	.w3(32'hbaa6e090),
	.w4(32'h3a0f2d8c),
	.w5(32'hba858f58),
	.w6(32'h3ab2bd96),
	.w7(32'hbb1c4650),
	.w8(32'hbb59d92a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3d75),
	.w1(32'hbb022652),
	.w2(32'hbb144e2b),
	.w3(32'hba888213),
	.w4(32'hb7aa36cf),
	.w5(32'h3b0a5c5d),
	.w6(32'h3b103218),
	.w7(32'h3b03ea1a),
	.w8(32'h3b54cd70),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67ac3b),
	.w1(32'h3bb41113),
	.w2(32'h3b74f712),
	.w3(32'h3b6ea516),
	.w4(32'h3bba293e),
	.w5(32'hbbba3d6d),
	.w6(32'h3b1bbf09),
	.w7(32'h3b66ba61),
	.w8(32'h3a25cd11),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30969f),
	.w1(32'hbbbb1d58),
	.w2(32'hbc1318fb),
	.w3(32'hbc1b7a3d),
	.w4(32'hbbb1e2b7),
	.w5(32'hb801b581),
	.w6(32'hbc15eb9d),
	.w7(32'hbb84f99b),
	.w8(32'h3b93fb29),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule