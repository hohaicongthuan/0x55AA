module layer_10_featuremap_193(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78c8bfa),
	.w1(32'h363ec326),
	.w2(32'hb74af0bc),
	.w3(32'hb7d3b359),
	.w4(32'hb7630cbf),
	.w5(32'hb79b2cf9),
	.w6(32'hb7bb46b7),
	.w7(32'hb7b3f151),
	.w8(32'hb803328b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d012f3),
	.w1(32'hba85d913),
	.w2(32'h3a485029),
	.w3(32'h378add9f),
	.w4(32'hba2f0479),
	.w5(32'h3aa05176),
	.w6(32'h3ae61507),
	.w7(32'h3b607277),
	.w8(32'h3bbc2665),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76a7f8c),
	.w1(32'hb5cf2f4d),
	.w2(32'hb6cedd4a),
	.w3(32'hb7863a47),
	.w4(32'hb696dd1b),
	.w5(32'hb6f8ada7),
	.w6(32'hb780ed44),
	.w7(32'hb6df33af),
	.w8(32'hb75e1cde),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585d71),
	.w1(32'hba349b72),
	.w2(32'hba9d4480),
	.w3(32'h3a4cdd8e),
	.w4(32'h3ab09828),
	.w5(32'h3ab35cb6),
	.w6(32'h39b0172a),
	.w7(32'h3a4beb2a),
	.w8(32'h3a36aea0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a2d95),
	.w1(32'h394b377e),
	.w2(32'h39e4b31e),
	.w3(32'hb94b28d7),
	.w4(32'h383cfa77),
	.w5(32'h399ec13a),
	.w6(32'hb970895e),
	.w7(32'hb8c67890),
	.w8(32'h389cc95c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f6c36e),
	.w1(32'h37679806),
	.w2(32'hb78c08a0),
	.w3(32'hb782412c),
	.w4(32'hb6fa1a29),
	.w5(32'hb8157ae1),
	.w6(32'hb7edca31),
	.w7(32'hb754d8f6),
	.w8(32'hb8480041),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32645a),
	.w1(32'h3b820712),
	.w2(32'h3b71c48e),
	.w3(32'h3b20ba2c),
	.w4(32'h3b8c2a23),
	.w5(32'h3b6daf18),
	.w6(32'h3b72c747),
	.w7(32'h3930d28f),
	.w8(32'h3abb8bb3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d47d9),
	.w1(32'h3b995256),
	.w2(32'hbb8de15e),
	.w3(32'h3c8d8a86),
	.w4(32'h3b774f86),
	.w5(32'hbb6a1a20),
	.w6(32'h3c796dec),
	.w7(32'h3bc29967),
	.w8(32'h390b5751),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a577658),
	.w1(32'hb84e11b7),
	.w2(32'h3966062c),
	.w3(32'h3a21c013),
	.w4(32'hba2d1512),
	.w5(32'hb9baf63a),
	.w6(32'h39d5c329),
	.w7(32'hba3c5645),
	.w8(32'hb9ead536),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7b2f1),
	.w1(32'hba60674c),
	.w2(32'hb92c1405),
	.w3(32'h3be43dd1),
	.w4(32'hbb3a5a3b),
	.w5(32'hbb2cf4c0),
	.w6(32'h3c218553),
	.w7(32'hb88cda7a),
	.w8(32'h3949a1ce),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60dfc4),
	.w1(32'h3a5a322d),
	.w2(32'h3a9a3b20),
	.w3(32'h3a2dd6c6),
	.w4(32'h392bab22),
	.w5(32'h3a38ce93),
	.w6(32'h398ee246),
	.w7(32'h38eb0b0b),
	.w8(32'h3a1f4bb9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284497),
	.w1(32'h3a837bab),
	.w2(32'h3ac114f8),
	.w3(32'h3b75a9ed),
	.w4(32'hbabff26d),
	.w5(32'h3b286e02),
	.w6(32'h3b8a9b0d),
	.w7(32'hbba638f9),
	.w8(32'hba6339a2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd258dc),
	.w1(32'hbb1a4511),
	.w2(32'hbad383c0),
	.w3(32'h3bd3af40),
	.w4(32'hbb1a8c29),
	.w5(32'hbb1838f1),
	.w6(32'h3bdfa130),
	.w7(32'hbac6cd31),
	.w8(32'hba2af50e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b083f36),
	.w1(32'h3ae114d9),
	.w2(32'h3b3f045a),
	.w3(32'h3aaaddc0),
	.w4(32'hbad3dfef),
	.w5(32'hbaab624f),
	.w6(32'h3a64ff13),
	.w7(32'hba3337d6),
	.w8(32'hba015488),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000c96),
	.w1(32'hbb0c1251),
	.w2(32'h39513b9f),
	.w3(32'h39b73741),
	.w4(32'hbb2e2d42),
	.w5(32'hba8bf607),
	.w6(32'h3b315cb1),
	.w7(32'h3b17f069),
	.w8(32'h3b911356),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d9f6a),
	.w1(32'h39bb9eee),
	.w2(32'hbb9151e6),
	.w3(32'h3ba2570f),
	.w4(32'hbb68c372),
	.w5(32'hbb97602c),
	.w6(32'h3bfa1f5f),
	.w7(32'hbac4ae3d),
	.w8(32'h3aa5551a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a056a63),
	.w1(32'hb87bf2a9),
	.w2(32'hb92d9491),
	.w3(32'h39c44e9f),
	.w4(32'hb9de5a6d),
	.w5(32'hb9e49152),
	.w6(32'h393b79d8),
	.w7(32'hb98d5ebe),
	.w8(32'hb9cb1eaf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c181),
	.w1(32'h3aa33fbf),
	.w2(32'hbbca756c),
	.w3(32'h3c34d937),
	.w4(32'hbaf51565),
	.w5(32'hbaa1ce64),
	.w6(32'h3c23d8c1),
	.w7(32'hbbc33320),
	.w8(32'hbb314df3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ee947),
	.w1(32'hba9c28a4),
	.w2(32'hbb56ec54),
	.w3(32'h3ba15880),
	.w4(32'hbb06f1a1),
	.w5(32'hbb1b3887),
	.w6(32'h3ba1930a),
	.w7(32'hbaf3ab40),
	.w8(32'hba806380),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d8694d),
	.w1(32'hb80977cb),
	.w2(32'h382a6d56),
	.w3(32'hb898c2db),
	.w4(32'hb95cd4d1),
	.w5(32'hb9177cf9),
	.w6(32'h38866219),
	.w7(32'h38b9bc23),
	.w8(32'h393ef2fc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f1c606),
	.w1(32'h38cddf77),
	.w2(32'h39718de7),
	.w3(32'h3924ce31),
	.w4(32'h394346fd),
	.w5(32'h391b71a3),
	.w6(32'h38b2c958),
	.w7(32'h375e28eb),
	.w8(32'hb93515c8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d39d6),
	.w1(32'hbb16efa2),
	.w2(32'h39bd7c78),
	.w3(32'hbb6c02f3),
	.w4(32'hbaa75127),
	.w5(32'h3ac750bc),
	.w6(32'hbb29ba9d),
	.w7(32'hb9d648d8),
	.w8(32'h3b1d7c4d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c517827),
	.w1(32'h3b2ed7e2),
	.w2(32'hbb968cc4),
	.w3(32'h3c4aaf5d),
	.w4(32'h39eeeff4),
	.w5(32'h3b4191e5),
	.w6(32'h3ca76cb5),
	.w7(32'h3b153f59),
	.w8(32'h3c2daf00),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a922b70),
	.w1(32'hbb7a9050),
	.w2(32'hba58b66b),
	.w3(32'h3b4ce0de),
	.w4(32'hbb4dba96),
	.w5(32'hb81c734d),
	.w6(32'h3bb85eab),
	.w7(32'h3a7affa3),
	.w8(32'h3b36d9cf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1651b1),
	.w1(32'hbc2b0eab),
	.w2(32'hbb5625c5),
	.w3(32'h39f7828c),
	.w4(32'hbb56b1c1),
	.w5(32'h3b49c89a),
	.w6(32'h3b0da139),
	.w7(32'h3b608dc0),
	.w8(32'h3c3fb076),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398273ca),
	.w1(32'hb834953f),
	.w2(32'hb850affa),
	.w3(32'h3916116d),
	.w4(32'hb9815568),
	.w5(32'hb9b91601),
	.w6(32'h3950dea6),
	.w7(32'hb9909f95),
	.w8(32'hb9d08d86),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e9134),
	.w1(32'hb7c1d445),
	.w2(32'hb8b75c8b),
	.w3(32'hb903fcce),
	.w4(32'hb7dc9142),
	.w5(32'hb8ac415a),
	.w6(32'hb945d309),
	.w7(32'hb8c8240a),
	.w8(32'hb909e7ee),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6319df),
	.w1(32'h3b23ec0d),
	.w2(32'h3c041106),
	.w3(32'hbbdd9e53),
	.w4(32'h3bc728fd),
	.w5(32'h3bb937ed),
	.w6(32'hbc633661),
	.w7(32'hba1d393e),
	.w8(32'h3bc89952),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c0b2a),
	.w1(32'hba195f50),
	.w2(32'h3a7fe24b),
	.w3(32'hba8a6d3c),
	.w4(32'hbad913bf),
	.w5(32'h392ef75d),
	.w6(32'hb9f37d1a),
	.w7(32'hbacaf2e7),
	.w8(32'h38ea0e57),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9434e5),
	.w1(32'hbc088e23),
	.w2(32'hba1d4512),
	.w3(32'hbbafa97d),
	.w4(32'h3ae81677),
	.w5(32'h3c274942),
	.w6(32'hbbf45b34),
	.w7(32'h3ac1ee2e),
	.w8(32'h3c34cd94),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8741180),
	.w1(32'hb7fbdd92),
	.w2(32'hb7c05cc8),
	.w3(32'hb892ad34),
	.w4(32'hb85ea5d3),
	.w5(32'hb869969c),
	.w6(32'hb8a573e2),
	.w7(32'hb8876dda),
	.w8(32'hb892016d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d3e97d),
	.w1(32'hb8b813cd),
	.w2(32'hb8a391c8),
	.w3(32'hb8d63a30),
	.w4(32'hb9500a3f),
	.w5(32'hb94b89a8),
	.w6(32'hb93cd09b),
	.w7(32'hb9536d6e),
	.w8(32'hb93625c2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e4b3f),
	.w1(32'hba3d6599),
	.w2(32'hba171997),
	.w3(32'h3aea0e85),
	.w4(32'hbad6663e),
	.w5(32'hbab23df4),
	.w6(32'h3b71fd1a),
	.w7(32'h39fc55c1),
	.w8(32'h3a8d6dfe),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e6868),
	.w1(32'hbabc25df),
	.w2(32'h3a0f4c70),
	.w3(32'h3aa8f103),
	.w4(32'hb8eb207f),
	.w5(32'h3ae69ab1),
	.w6(32'h3ab08a99),
	.w7(32'h3b048246),
	.w8(32'h3b84d36f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2a7ea),
	.w1(32'h3700c564),
	.w2(32'hb9cf5a71),
	.w3(32'hb9981b08),
	.w4(32'hb9af17df),
	.w5(32'hba4e9ee9),
	.w6(32'h399fad0c),
	.w7(32'h39527304),
	.w8(32'hb9b4ead9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b1cf3),
	.w1(32'h3b536c76),
	.w2(32'h3a4d6d95),
	.w3(32'h3ba2df9e),
	.w4(32'h3b9c6e5e),
	.w5(32'h3b0c481a),
	.w6(32'h3b8218bd),
	.w7(32'h39d4b272),
	.w8(32'hbaa54480),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c413d75),
	.w1(32'h3bfeef3a),
	.w2(32'h3c56bc30),
	.w3(32'h3afad202),
	.w4(32'hbbaed63e),
	.w5(32'hbb2f9642),
	.w6(32'h387e0606),
	.w7(32'hbb94d6f7),
	.w8(32'h3a40a03c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca36406),
	.w1(32'hbbf0b9f2),
	.w2(32'h3c062054),
	.w3(32'hbc357361),
	.w4(32'h3a74d89e),
	.w5(32'h3c5d3f54),
	.w6(32'hbb6c501f),
	.w7(32'h3c34b2ad),
	.w8(32'h3caf7290),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4eec2),
	.w1(32'hbbef5a2c),
	.w2(32'h3c56f363),
	.w3(32'hbc7fa037),
	.w4(32'h3abd666b),
	.w5(32'h3cbc4cc9),
	.w6(32'hbc478027),
	.w7(32'h3b5d8d96),
	.w8(32'h3cb47cf9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc695),
	.w1(32'hbaa60632),
	.w2(32'h393b83b0),
	.w3(32'h37c5e960),
	.w4(32'h3a0e93bb),
	.w5(32'h3a62bd41),
	.w6(32'h3a8110e5),
	.w7(32'h3af6ba45),
	.w8(32'h3b35f5b5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903a62e),
	.w1(32'h397e48e0),
	.w2(32'hb8cf9f59),
	.w3(32'h38b2da23),
	.w4(32'h3954897a),
	.w5(32'hb8ba8615),
	.w6(32'h389b3563),
	.w7(32'h39059ec9),
	.w8(32'hb8fc5bb4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920bdb7),
	.w1(32'h394d6bd3),
	.w2(32'h38cf5353),
	.w3(32'hb96811ca),
	.w4(32'h3941e463),
	.w5(32'h391cfe89),
	.w6(32'hb969df5c),
	.w7(32'h37e822c9),
	.w8(32'hb8161234),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a334320),
	.w1(32'hbaa7e4a5),
	.w2(32'h3a482e3a),
	.w3(32'h3ab2c687),
	.w4(32'hba289cb0),
	.w5(32'h3aa09a0e),
	.w6(32'h398ba335),
	.w7(32'hbaf07327),
	.w8(32'h3a4adc9c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1faf92),
	.w1(32'hbb7a9bd4),
	.w2(32'hba28dedb),
	.w3(32'h3c29ebab),
	.w4(32'hbbc951c7),
	.w5(32'hbb41a848),
	.w6(32'h3c0c65df),
	.w7(32'hbbf46200),
	.w8(32'hbb4e8306),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3373eb),
	.w1(32'hbbd52592),
	.w2(32'hbb1978d0),
	.w3(32'h3a8b574e),
	.w4(32'hbb3f6d82),
	.w5(32'h39112680),
	.w6(32'h3b0a5c8d),
	.w7(32'h3ac507e2),
	.w8(32'h3bd5b50c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e92d1c),
	.w1(32'hbbdf0f59),
	.w2(32'hbbcaacf8),
	.w3(32'h3bb74664),
	.w4(32'hbb39dfcc),
	.w5(32'hbb2858b0),
	.w6(32'h3bf16092),
	.w7(32'h3acb1086),
	.w8(32'h3b76d1af),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a257503),
	.w1(32'hbb5fd17a),
	.w2(32'hbaf8b9f2),
	.w3(32'h3b143296),
	.w4(32'hb972ac01),
	.w5(32'h3b14e859),
	.w6(32'h3b8a614c),
	.w7(32'h3b19f54d),
	.w8(32'h3b94c500),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25c6cb),
	.w1(32'h3b317aa8),
	.w2(32'hbb4095b9),
	.w3(32'h3c40a0f4),
	.w4(32'h3b272717),
	.w5(32'h3a1cbb99),
	.w6(32'h3c404237),
	.w7(32'hbb006508),
	.w8(32'h3a231996),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca78fa),
	.w1(32'h38853b7d),
	.w2(32'hb996d052),
	.w3(32'hb9bf75d4),
	.w4(32'h396f0476),
	.w5(32'h37c9d0a2),
	.w6(32'hb96878fc),
	.w7(32'h39617726),
	.w8(32'h3846867c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e689e1),
	.w1(32'hb93bad64),
	.w2(32'hb991f67c),
	.w3(32'h39a88c4d),
	.w4(32'h3a09ca28),
	.w5(32'h39c7279f),
	.w6(32'h39503ca4),
	.w7(32'h3a382848),
	.w8(32'h3a5c4748),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971ca24),
	.w1(32'h39f34dd0),
	.w2(32'h39bc66c4),
	.w3(32'h396f05c5),
	.w4(32'h39bdcf79),
	.w5(32'h39930de0),
	.w6(32'h390f1be5),
	.w7(32'h39e5fa9d),
	.w8(32'h39c86c9f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f034f),
	.w1(32'hb93c285d),
	.w2(32'hba95fd7a),
	.w3(32'h3b10792d),
	.w4(32'h385ca74c),
	.w5(32'h3a591dbd),
	.w6(32'h3aa809c9),
	.w7(32'hba4ff05b),
	.w8(32'h3ac1a355),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c3f35),
	.w1(32'hb7ce4fdc),
	.w2(32'hba8d7051),
	.w3(32'h3ae753b6),
	.w4(32'h388eafc6),
	.w5(32'h39e252d6),
	.w6(32'h3ac98013),
	.w7(32'hb898e04c),
	.w8(32'h399a2a0b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c527c4b),
	.w1(32'h3aa74e16),
	.w2(32'hbb37b40f),
	.w3(32'h3c1cb553),
	.w4(32'hbb6d081e),
	.w5(32'hbba46534),
	.w6(32'h3c2dd943),
	.w7(32'hbb90d9ea),
	.w8(32'hbb4e0100),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39866f48),
	.w1(32'hbac585ed),
	.w2(32'hba5c62e3),
	.w3(32'h3b0752a1),
	.w4(32'hba6305c9),
	.w5(32'h3a2c0fda),
	.w6(32'hb9d069b1),
	.w7(32'hbb2d3b3d),
	.w8(32'hb9c28a75),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eca6e6),
	.w1(32'hb9536b3b),
	.w2(32'h39502d6a),
	.w3(32'hb8fff283),
	.w4(32'hb9a0fb19),
	.w5(32'h37490c09),
	.w6(32'hb837fec2),
	.w7(32'h35f0c9b0),
	.w8(32'h39a62b5d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811144f),
	.w1(32'h351567c8),
	.w2(32'hb758c209),
	.w3(32'hb7d5f008),
	.w4(32'hb7c3a113),
	.w5(32'hb6f15767),
	.w6(32'hb88bb1e6),
	.w7(32'hb7ca4b13),
	.w8(32'hb6fdc8e3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3d09),
	.w1(32'hb9e592cd),
	.w2(32'h39d5f857),
	.w3(32'hb9dfe60e),
	.w4(32'h39cfbe01),
	.w5(32'h3a8522d6),
	.w6(32'hb999de62),
	.w7(32'h39488b0e),
	.w8(32'h3a320f51),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e5c4d),
	.w1(32'hba1674d6),
	.w2(32'h39f07a2b),
	.w3(32'hb9a7489d),
	.w4(32'hb8c99207),
	.w5(32'h3a58e752),
	.w6(32'hb94a8150),
	.w7(32'h38c519c4),
	.w8(32'h3a5ea237),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20e6f0),
	.w1(32'hba19dc41),
	.w2(32'hb9b731db),
	.w3(32'hba470c6c),
	.w4(32'hb9ec64f7),
	.w5(32'hb9382dab),
	.w6(32'hba3b8d33),
	.w7(32'hba5c2d34),
	.w8(32'hb9bfc2fc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b796dbb),
	.w1(32'hba5afd4d),
	.w2(32'hbb368bcd),
	.w3(32'h3b6780b0),
	.w4(32'hbad95c0b),
	.w5(32'hbac7936c),
	.w6(32'h3b2055ae),
	.w7(32'hbb1b08cd),
	.w8(32'hb9d8fb6b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815863),
	.w1(32'hbae654fe),
	.w2(32'hbb7cd559),
	.w3(32'h3b2461c6),
	.w4(32'hbb481acd),
	.w5(32'hb993aa95),
	.w6(32'hbae87c5f),
	.w7(32'hbc112a95),
	.w8(32'hbb16fdc6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380dd63a),
	.w1(32'h3780d02a),
	.w2(32'hb8a36f34),
	.w3(32'h37becb1d),
	.w4(32'h37c69d81),
	.w5(32'hb869861b),
	.w6(32'hb77f7819),
	.w7(32'h369095b7),
	.w8(32'hb84d0c32),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7efb9b9),
	.w1(32'hb6107b60),
	.w2(32'hb8621d6f),
	.w3(32'hb75a51e1),
	.w4(32'h3785db3d),
	.w5(32'hb809628b),
	.w6(32'hb8209333),
	.w7(32'h35c4ae92),
	.w8(32'hb801bfb8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79104b5),
	.w1(32'hb873b096),
	.w2(32'hb8b984ab),
	.w3(32'hb8f6cf1f),
	.w4(32'hb93f2e58),
	.w5(32'hb937e971),
	.w6(32'hb91a8906),
	.w7(32'hb9490652),
	.w8(32'hb92b193f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aefd99),
	.w1(32'hb7870ab9),
	.w2(32'hb8b06bc3),
	.w3(32'hb88a2a07),
	.w4(32'hb70d0ca7),
	.w5(32'hb8b2fd93),
	.w6(32'hb8dbc030),
	.w7(32'hb8175c45),
	.w8(32'hb8ea2a57),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c9a99),
	.w1(32'h3c02be52),
	.w2(32'hb8f474de),
	.w3(32'h3baa1233),
	.w4(32'hbbf79d69),
	.w5(32'hbc3a732f),
	.w6(32'h3c2eb964),
	.w7(32'hbb2cd415),
	.w8(32'hbbb26fd3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2d19),
	.w1(32'hbc12b197),
	.w2(32'hbc1a469b),
	.w3(32'h3c472c27),
	.w4(32'h3b13a1fd),
	.w5(32'h3b7c3c58),
	.w6(32'h3c314d03),
	.w7(32'hba0b7411),
	.w8(32'h3a8e8c0f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8647),
	.w1(32'hbbc6526e),
	.w2(32'hbb0e6ee2),
	.w3(32'h3bf8d673),
	.w4(32'hbb3a85c6),
	.w5(32'h3b765e5e),
	.w6(32'h3bcebd46),
	.w7(32'hbbc5a7a0),
	.w8(32'h3b071630),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34c42d),
	.w1(32'hbc350e2e),
	.w2(32'hbb239f48),
	.w3(32'h3ad96faa),
	.w4(32'hb9b48ffb),
	.w5(32'h3bbbc540),
	.w6(32'h3baeaf31),
	.w7(32'h3c12e1f8),
	.w8(32'h3c9accfc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376d128c),
	.w1(32'h3854df45),
	.w2(32'hb85cb9e3),
	.w3(32'h372d3010),
	.w4(32'h381d0476),
	.w5(32'hb8c54b96),
	.w6(32'hb8187d55),
	.w7(32'h369830f6),
	.w8(32'hb8f598e1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80670a3),
	.w1(32'h38519ca8),
	.w2(32'hb8ed07ff),
	.w3(32'hb85550ad),
	.w4(32'h37a87075),
	.w5(32'hb9292d2c),
	.w6(32'hb8e6acb9),
	.w7(32'hb7f615c5),
	.w8(32'hb9380cae),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f01792),
	.w1(32'h38a5d642),
	.w2(32'hb8ee1ba7),
	.w3(32'hb8c14991),
	.w4(32'h383aa918),
	.w5(32'hb936f2cb),
	.w6(32'hb8fc6691),
	.w7(32'hb84b4044),
	.w8(32'hb95d05ec),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af788fe),
	.w1(32'hba401d2e),
	.w2(32'hbabded45),
	.w3(32'h3af1710e),
	.w4(32'hba6bd634),
	.w5(32'hba750f29),
	.w6(32'h3ab858b8),
	.w7(32'hbaa91cea),
	.w8(32'hba4ddd55),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3838ff67),
	.w1(32'h3943246a),
	.w2(32'h37a66d4a),
	.w3(32'hb7f38e6e),
	.w4(32'h39257453),
	.w5(32'h3889bd1b),
	.w6(32'hb81d972e),
	.w7(32'h38c893ce),
	.w8(32'hb69cb207),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6601),
	.w1(32'h3b07c59e),
	.w2(32'hba4d47b1),
	.w3(32'h3b92aeff),
	.w4(32'h3b1f1b92),
	.w5(32'hbb414a66),
	.w6(32'h3bbd2e36),
	.w7(32'h3b04a12a),
	.w8(32'hb9da0b8d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec3ecd),
	.w1(32'h3b907345),
	.w2(32'hbaad6900),
	.w3(32'h3bdb17b0),
	.w4(32'h3b1360c0),
	.w5(32'hbb04a1ef),
	.w6(32'h3c22ba8b),
	.w7(32'h3a98a5dc),
	.w8(32'hba9ef310),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719cec),
	.w1(32'hbb678e8b),
	.w2(32'hbb0b1a55),
	.w3(32'h3a48e5ab),
	.w4(32'hbb30efcc),
	.w5(32'hbb2536f0),
	.w6(32'h3a88f424),
	.w7(32'h3b328161),
	.w8(32'h3bab3417),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93a4f2),
	.w1(32'h3a10860c),
	.w2(32'h391357f2),
	.w3(32'h3b83821e),
	.w4(32'hba8c89b8),
	.w5(32'h394dcd4e),
	.w6(32'h3b9b083a),
	.w7(32'hba1ce88c),
	.w8(32'h3a393195),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf842e),
	.w1(32'h3b8900ac),
	.w2(32'h3aaafb00),
	.w3(32'h3b34019e),
	.w4(32'h3a3b4ec1),
	.w5(32'hbb68439c),
	.w6(32'h3ba88c8e),
	.w7(32'h3b3b2f09),
	.w8(32'hbaf71e5d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad03c51),
	.w1(32'hbad5cea7),
	.w2(32'h3a76ab98),
	.w3(32'h3b235e88),
	.w4(32'hbacad600),
	.w5(32'hb8621149),
	.w6(32'h3abcfa76),
	.w7(32'hb98d4edc),
	.w8(32'h3aa05fa4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e84b),
	.w1(32'h3a128434),
	.w2(32'hba443b44),
	.w3(32'h3ba6fa0e),
	.w4(32'h3a474818),
	.w5(32'hb8d9fe04),
	.w6(32'h3b99eeb4),
	.w7(32'hb99ca286),
	.w8(32'h39beb55c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b323d5),
	.w1(32'hb73c0c36),
	.w2(32'hb7a48725),
	.w3(32'h37cdcb33),
	.w4(32'hb694e32c),
	.w5(32'hb7f69d7d),
	.w6(32'h3641a160),
	.w7(32'hb738390d),
	.w8(32'hb84b1890),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387547df),
	.w1(32'h382d2f49),
	.w2(32'h37a02aad),
	.w3(32'h369e0c97),
	.w4(32'hb7a56b6b),
	.w5(32'hb85b6c00),
	.w6(32'h38871039),
	.w7(32'h37ec63a8),
	.w8(32'hb78aad0a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad128f),
	.w1(32'hb91ee3d2),
	.w2(32'hb95e6094),
	.w3(32'h38d1321f),
	.w4(32'hb8bd6fa4),
	.w5(32'hb90144af),
	.w6(32'h382b3d9b),
	.w7(32'hb7e1f4fc),
	.w8(32'hb9187761),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae55e5b),
	.w1(32'hba30f8c6),
	.w2(32'h39a0b5e4),
	.w3(32'hba22c805),
	.w4(32'h3a198a67),
	.w5(32'h3aab4ca4),
	.w6(32'hba419319),
	.w7(32'h3a1251ea),
	.w8(32'h3a9d436b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9ead3),
	.w1(32'hbb6394cd),
	.w2(32'h3a5fd986),
	.w3(32'h3a97fde0),
	.w4(32'hbabe4839),
	.w5(32'h3b2e511f),
	.w6(32'h3b0269b0),
	.w7(32'h3b6cabe3),
	.w8(32'h3bd06c92),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07c216),
	.w1(32'hba64387b),
	.w2(32'hb97de955),
	.w3(32'hb992d103),
	.w4(32'hba78a3be),
	.w5(32'hb9815e11),
	.w6(32'h399dbeb9),
	.w7(32'hb96e5497),
	.w8(32'h397e6f4b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a999e),
	.w1(32'hbb7dfc16),
	.w2(32'hbba68ed1),
	.w3(32'h3ba946f0),
	.w4(32'h39a075b2),
	.w5(32'hbad34a31),
	.w6(32'h3b99228c),
	.w7(32'h3a7acfa7),
	.w8(32'h3a157851),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a10aa),
	.w1(32'h3882a669),
	.w2(32'hba9547be),
	.w3(32'h3bdc1d1d),
	.w4(32'h3b10745f),
	.w5(32'h3b920302),
	.w6(32'h3c3722e2),
	.w7(32'h3b231709),
	.w8(32'h3bb773d0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cc76b),
	.w1(32'hbb7e2563),
	.w2(32'h3ba5cd9f),
	.w3(32'hbbbb5558),
	.w4(32'h3b0931d1),
	.w5(32'h3c2a8f82),
	.w6(32'hbbc476df),
	.w7(32'h3a91724b),
	.w8(32'h3c1f73c1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c664af4),
	.w1(32'h3c0eb348),
	.w2(32'h3a979e23),
	.w3(32'h3ba9a84a),
	.w4(32'hb8b6a2b6),
	.w5(32'hbc03b8bd),
	.w6(32'h3c4528c0),
	.w7(32'h3b817573),
	.w8(32'hba1adf7e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe324b2),
	.w1(32'hbb93072e),
	.w2(32'h39b84670),
	.w3(32'hba77f9ca),
	.w4(32'h3a8b109f),
	.w5(32'h3b6d9e7f),
	.w6(32'hb936826c),
	.w7(32'h3adc3839),
	.w8(32'h3b75ccd2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f4834),
	.w1(32'h3a9d49b8),
	.w2(32'hbb4ff60b),
	.w3(32'h3c000a41),
	.w4(32'hbb5f8466),
	.w5(32'hbc01304c),
	.w6(32'h3c4a7c9f),
	.w7(32'h3a84cb0e),
	.w8(32'hbb0125c5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8836d),
	.w1(32'hba1e0987),
	.w2(32'hb9f913ee),
	.w3(32'h389e2f0d),
	.w4(32'hbb2637ba),
	.w5(32'hbb0d6dd4),
	.w6(32'h3b193f64),
	.w7(32'h3b25c362),
	.w8(32'h3b4dfe9c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08699e),
	.w1(32'hbb923c3b),
	.w2(32'h3af9c478),
	.w3(32'hbb341f1e),
	.w4(32'h3acc9ee8),
	.w5(32'h3bde85d3),
	.w6(32'hbab3c221),
	.w7(32'h3ba603dd),
	.w8(32'h3c1ccc63),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c11de),
	.w1(32'h396e19a5),
	.w2(32'hb90d8dfd),
	.w3(32'h395530e9),
	.w4(32'h3a02196c),
	.w5(32'hb89459e4),
	.w6(32'h38ce602f),
	.w7(32'h3989ad29),
	.w8(32'hb98431f5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75866),
	.w1(32'hbaa0f12d),
	.w2(32'hbb4372e7),
	.w3(32'h3be5539e),
	.w4(32'hbaf50bbe),
	.w5(32'hbaff9a19),
	.w6(32'h3c19994a),
	.w7(32'hba0e23d1),
	.w8(32'h3a9fcdc9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c0f49),
	.w1(32'h3a3e4810),
	.w2(32'hbb17cb9e),
	.w3(32'h3ae9e09b),
	.w4(32'h38a931a9),
	.w5(32'hbb0cdcbc),
	.w6(32'h3ba71ad6),
	.w7(32'h3b2c631d),
	.w8(32'h3aee69b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b65a1),
	.w1(32'h3b8f8693),
	.w2(32'hb9035890),
	.w3(32'h3c3132d8),
	.w4(32'h3ba52213),
	.w5(32'hbb8f3982),
	.w6(32'h3c407ce7),
	.w7(32'h3b28dabe),
	.w8(32'hbb263003),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9a1a8),
	.w1(32'h3abacd10),
	.w2(32'h3c17aab8),
	.w3(32'hba5fafa1),
	.w4(32'h3bdd8a49),
	.w5(32'h3c575b72),
	.w6(32'h3ae71c29),
	.w7(32'h3c2aa880),
	.w8(32'h3c82b621),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb927547),
	.w1(32'hbbef9c8f),
	.w2(32'hbb5ced90),
	.w3(32'h3b6939e5),
	.w4(32'hbb3137f8),
	.w5(32'h3a48e7ec),
	.w6(32'h3b82f76a),
	.w7(32'h3ad0bd6c),
	.w8(32'h3bbf1273),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04cf35),
	.w1(32'h3bb8210b),
	.w2(32'h3a063487),
	.w3(32'h3b5446aa),
	.w4(32'hba8b1eec),
	.w5(32'hbbdc23d3),
	.w6(32'h3bd74f09),
	.w7(32'hbb1e5f76),
	.w8(32'hbbecf981),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82f07d),
	.w1(32'hba958ef6),
	.w2(32'hbad7c072),
	.w3(32'hbaf0ebff),
	.w4(32'hbaa0da5d),
	.w5(32'hba764d69),
	.w6(32'hba84fecb),
	.w7(32'hba9ec5b7),
	.w8(32'hbaa61a1f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8671db),
	.w1(32'h3ba3e5b8),
	.w2(32'h3bad6306),
	.w3(32'h3c34767a),
	.w4(32'h3b4bd541),
	.w5(32'hbb100ea9),
	.w6(32'h3c16d3d6),
	.w7(32'h3b107b7c),
	.w8(32'h3bf26d85),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeff0e),
	.w1(32'h3b11924f),
	.w2(32'h3b372c08),
	.w3(32'h3b924056),
	.w4(32'h3b12663c),
	.w5(32'h3b2c0002),
	.w6(32'h3b71064e),
	.w7(32'h3b6c1c6e),
	.w8(32'h3a31406b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba305213),
	.w1(32'h38ba0063),
	.w2(32'h39bd97f6),
	.w3(32'hba22dec3),
	.w4(32'h3796b2a7),
	.w5(32'h39a38635),
	.w6(32'hba35c7b9),
	.w7(32'h36f589a5),
	.w8(32'h3992554a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09674e),
	.w1(32'h3a01fad7),
	.w2(32'h38990981),
	.w3(32'h3b162ed8),
	.w4(32'h39aba25e),
	.w5(32'hbaa02db7),
	.w6(32'h3b045f3f),
	.w7(32'h3b0a7655),
	.w8(32'h3b159f8b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7028a),
	.w1(32'hbaa0f4ea),
	.w2(32'h38ec1ce3),
	.w3(32'h3b55e4fb),
	.w4(32'hb985a3de),
	.w5(32'h3a18bb0b),
	.w6(32'h3bafb2fe),
	.w7(32'hb9459752),
	.w8(32'h3abcb3c4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85e23b),
	.w1(32'hbb91200f),
	.w2(32'hba13512f),
	.w3(32'h39f0fea1),
	.w4(32'hba89131c),
	.w5(32'h3a8b496f),
	.w6(32'h3a5363ff),
	.w7(32'h3aabb9b4),
	.w8(32'h3b8e0e2d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987327),
	.w1(32'hbaea34c8),
	.w2(32'h3b49ba7b),
	.w3(32'hbbc784bf),
	.w4(32'hba5ed2a3),
	.w5(32'h3bb398c6),
	.w6(32'hbbb60141),
	.w7(32'h3a2674bc),
	.w8(32'h3be26ad5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aab05),
	.w1(32'hbb5cbab5),
	.w2(32'hbb134dd7),
	.w3(32'hbab38336),
	.w4(32'hbad24b27),
	.w5(32'h398bd26f),
	.w6(32'h38c07fc9),
	.w7(32'h3b074936),
	.w8(32'h3baf1420),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50baee),
	.w1(32'hbb8306c1),
	.w2(32'hbc27a3b5),
	.w3(32'h3bcba223),
	.w4(32'h3bc869ed),
	.w5(32'hbadfc23d),
	.w6(32'h3bd13270),
	.w7(32'h3b29faf5),
	.w8(32'hba8cbc11),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19a77c),
	.w1(32'h3b68017f),
	.w2(32'h390a7a19),
	.w3(32'h3b8a6ccb),
	.w4(32'hbb4e6c54),
	.w5(32'hbbb92f5b),
	.w6(32'h3bb0406c),
	.w7(32'hba4a9e88),
	.w8(32'hbb03be89),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc431),
	.w1(32'hbb3ea763),
	.w2(32'hba84372a),
	.w3(32'h3aaf8bc5),
	.w4(32'hba297900),
	.w5(32'h3a2f03be),
	.w6(32'h3aee94f3),
	.w7(32'h3a40652b),
	.w8(32'h3b167c5a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c11f8),
	.w1(32'h39062329),
	.w2(32'hb7aab640),
	.w3(32'h3907891c),
	.w4(32'h38f60297),
	.w5(32'hb7b18575),
	.w6(32'h3955a63a),
	.w7(32'h39190bcd),
	.w8(32'h375a688b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80abe6),
	.w1(32'hba05bd93),
	.w2(32'hba51b191),
	.w3(32'hb803b220),
	.w4(32'hba004012),
	.w5(32'hba18135b),
	.w6(32'h3a59b337),
	.w7(32'h39cff488),
	.w8(32'h3908f918),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb677ac37),
	.w1(32'hb7d952c9),
	.w2(32'hb872e288),
	.w3(32'h36cf0962),
	.w4(32'h34eb047c),
	.w5(32'hb7454cb9),
	.w6(32'hb70b8e0d),
	.w7(32'hb6bf001d),
	.w8(32'hb7e73d6d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b05a9c),
	.w1(32'hb9a4e86e),
	.w2(32'hb95ac16e),
	.w3(32'hb93d3465),
	.w4(32'hb980fcd5),
	.w5(32'hb8ff0b32),
	.w6(32'hb983640a),
	.w7(32'hb9fb3e3d),
	.w8(32'hb9cb2b3d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab4697),
	.w1(32'hbba2b961),
	.w2(32'hbb3b1406),
	.w3(32'h3ad47fb7),
	.w4(32'hbb3aaa94),
	.w5(32'hbad4d697),
	.w6(32'h3b145c25),
	.w7(32'hba3d0102),
	.w8(32'h3a665dc7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0898a4),
	.w1(32'h395fcad8),
	.w2(32'h3a5fc764),
	.w3(32'hb88a7c58),
	.w4(32'h39272fdd),
	.w5(32'h3a80718d),
	.w6(32'hb9793d5a),
	.w7(32'hb88f4656),
	.w8(32'h3a39bf99),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ada3f),
	.w1(32'h3b01c203),
	.w2(32'hba5fdb79),
	.w3(32'h3b7f8021),
	.w4(32'h3adc0354),
	.w5(32'hba6872b9),
	.w6(32'h3b982787),
	.w7(32'h39af4cf7),
	.w8(32'hbabef062),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f902d),
	.w1(32'hbb31202e),
	.w2(32'h3b153932),
	.w3(32'hbb89d2b9),
	.w4(32'h3af1fdce),
	.w5(32'h3bc0bdc4),
	.w6(32'hbad4013a),
	.w7(32'h3c03cf32),
	.w8(32'h3c679fd4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cba7f),
	.w1(32'hb8b2d592),
	.w2(32'hb8a61d81),
	.w3(32'hb9353981),
	.w4(32'hb8fe1958),
	.w5(32'hb90b2487),
	.w6(32'hb9396312),
	.w7(32'hb8ef9197),
	.w8(32'h3711f218),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a516e9),
	.w1(32'h389a3288),
	.w2(32'h39193e11),
	.w3(32'hb8feb0e6),
	.w4(32'hb8c7c28b),
	.w5(32'hb79be8df),
	.w6(32'hb4d60091),
	.w7(32'hb671e25b),
	.w8(32'h390849e0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70b4928),
	.w1(32'hb7a329d1),
	.w2(32'h36b41a8e),
	.w3(32'hb7cf5034),
	.w4(32'hb838e783),
	.w5(32'hb800fb5b),
	.w6(32'hb841be51),
	.w7(32'hb88097dd),
	.w8(32'hb84047a7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1682e1),
	.w1(32'hb923baea),
	.w2(32'h399c2901),
	.w3(32'hb9b10aee),
	.w4(32'hb7c9fc7b),
	.w5(32'h3a119a88),
	.w6(32'h39879acc),
	.w7(32'h39f682ed),
	.w8(32'h3a32ca71),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f1f43),
	.w1(32'h3a775cce),
	.w2(32'hbbd2ce47),
	.w3(32'h3bfecfda),
	.w4(32'h3c02402b),
	.w5(32'hba67794d),
	.w6(32'h3bfff7af),
	.w7(32'h3aed5725),
	.w8(32'h3a53d594),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb8004),
	.w1(32'h3a29cb4b),
	.w2(32'hbaf203bc),
	.w3(32'h3bbd216d),
	.w4(32'hbb683fe9),
	.w5(32'hbb82b0a4),
	.w6(32'h3be579b1),
	.w7(32'hbb11ec5a),
	.w8(32'hbb29957d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac3532),
	.w1(32'h3a47bb25),
	.w2(32'hb9957b22),
	.w3(32'h39fe8120),
	.w4(32'hb879db0a),
	.w5(32'hba6d3667),
	.w6(32'h3a8becf6),
	.w7(32'h38ac9f0b),
	.w8(32'hb979bfa1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a542382),
	.w1(32'hba73bd2b),
	.w2(32'hba95ec1c),
	.w3(32'h3b108dbb),
	.w4(32'hb9c495ba),
	.w5(32'h38a62fb9),
	.w6(32'h3b203838),
	.w7(32'hb892d7c7),
	.w8(32'h3a9d6ab8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab339eb),
	.w1(32'hbab0de07),
	.w2(32'h38bbd56b),
	.w3(32'hba61bb6a),
	.w4(32'hba9c516a),
	.w5(32'h39bf8ee8),
	.w6(32'hba0be1b9),
	.w7(32'hb9e23e88),
	.w8(32'h3ae427a4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce880),
	.w1(32'hba65151d),
	.w2(32'hba8bb256),
	.w3(32'h3aff8c67),
	.w4(32'hbb143709),
	.w5(32'hba97c98d),
	.w6(32'h3b3e2c8a),
	.w7(32'hbab586da),
	.w8(32'hba110141),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b683eab),
	.w1(32'hb9861d2e),
	.w2(32'h3ae0b21d),
	.w3(32'h3aa20a34),
	.w4(32'hbb1d5fae),
	.w5(32'hbb00a814),
	.w6(32'h3a65fcf5),
	.w7(32'h3a9d8fe6),
	.w8(32'h3b844725),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1131d6),
	.w1(32'h3b81aa9d),
	.w2(32'hbac973c8),
	.w3(32'h3beeebe5),
	.w4(32'hba539515),
	.w5(32'hbb2f0109),
	.w6(32'h3c109277),
	.w7(32'hb987913f),
	.w8(32'hbacf339d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40a520),
	.w1(32'hbb5f9853),
	.w2(32'h3a02fea6),
	.w3(32'h3a085d60),
	.w4(32'h39603f01),
	.w5(32'h3b551bc2),
	.w6(32'h3aace9ca),
	.w7(32'h3b84c088),
	.w8(32'h3be2c53a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ea7c),
	.w1(32'h3a823376),
	.w2(32'hbb07cd14),
	.w3(32'h3b45f836),
	.w4(32'hbaa83331),
	.w5(32'hbb4ce92d),
	.w6(32'h3b975287),
	.w7(32'h3a832dbd),
	.w8(32'hb9aed6df),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c164102),
	.w1(32'h3b26f655),
	.w2(32'hbb195e87),
	.w3(32'h3c00a96d),
	.w4(32'h3aa38804),
	.w5(32'hb961f5ae),
	.w6(32'h3c0e6fdc),
	.w7(32'hba9eafba),
	.w8(32'h3907dac5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75b7b),
	.w1(32'hbb743efa),
	.w2(32'hbb4aa49e),
	.w3(32'h3b199260),
	.w4(32'h3a0fb7ce),
	.w5(32'h38ef1ca2),
	.w6(32'h3b88c3a4),
	.w7(32'h3b204b7d),
	.w8(32'h3b2cdf8e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84fbe5),
	.w1(32'h3abfa0e0),
	.w2(32'hb9fd79b4),
	.w3(32'h3b1cc3c3),
	.w4(32'hb9a9fb74),
	.w5(32'hbb0212b6),
	.w6(32'h3bbb8d64),
	.w7(32'h3aa59764),
	.w8(32'hb9807080),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8c6f0),
	.w1(32'hba1446de),
	.w2(32'hb9db8265),
	.w3(32'h3a4c7673),
	.w4(32'hb913da23),
	.w5(32'hb9a837df),
	.w6(32'h3a88064a),
	.w7(32'h3a08a0df),
	.w8(32'h3a3c6f06),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb64970),
	.w1(32'hbbe87691),
	.w2(32'hbb7688b0),
	.w3(32'hbbe595be),
	.w4(32'h3bf33ce3),
	.w5(32'h3c40dc54),
	.w6(32'hbbb7d0d4),
	.w7(32'h3c35a352),
	.w8(32'h3c90a5e7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8451ba),
	.w1(32'hba60a2eb),
	.w2(32'hbaa01f58),
	.w3(32'h3b17b0a0),
	.w4(32'h38a1d6dd),
	.w5(32'h3a2578bd),
	.w6(32'h3b1d4516),
	.w7(32'h3abf5e5e),
	.w8(32'h3ae40ae2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395383fd),
	.w1(32'h38b9e839),
	.w2(32'hb85bdf87),
	.w3(32'h396b7a2b),
	.w4(32'h38efa298),
	.w5(32'hb7cdb61f),
	.w6(32'h397851f1),
	.w7(32'h3957995f),
	.w8(32'hb87cf6ed),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946668e),
	.w1(32'h392e7efa),
	.w2(32'hb841ab7c),
	.w3(32'hb937102a),
	.w4(32'h38d84f46),
	.w5(32'hb82a63da),
	.w6(32'hb96913d6),
	.w7(32'h390687a2),
	.w8(32'h3805a5cb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae049e8),
	.w1(32'h3ab68562),
	.w2(32'h3a93dcc7),
	.w3(32'h3aaf754f),
	.w4(32'h3a8076f4),
	.w5(32'h3a6ea01f),
	.w6(32'h3b155b10),
	.w7(32'h3a8f8d23),
	.w8(32'h3a16216e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0720ee),
	.w1(32'hbb8d3299),
	.w2(32'hbaf85225),
	.w3(32'h399f5727),
	.w4(32'hbabe1ddb),
	.w5(32'h3abb86df),
	.w6(32'h3b54b901),
	.w7(32'h3ba06527),
	.w8(32'h3c01c789),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b240a5f),
	.w1(32'hbb833065),
	.w2(32'hbb355534),
	.w3(32'h3b707b94),
	.w4(32'hbb387eaa),
	.w5(32'hbb068ebe),
	.w6(32'h3b99aa82),
	.w7(32'hb9c859e3),
	.w8(32'h3a911ccd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831a779),
	.w1(32'h389def0f),
	.w2(32'hb7e95b66),
	.w3(32'h37d578c2),
	.w4(32'h3723319a),
	.w5(32'hb8078fce),
	.w6(32'h38322c20),
	.w7(32'hb85d953d),
	.w8(32'hb88229a0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e04f),
	.w1(32'hba23d542),
	.w2(32'h394df601),
	.w3(32'h3b90a6a7),
	.w4(32'hbac8bb32),
	.w5(32'hba8310da),
	.w6(32'h3bd3560b),
	.w7(32'h3aa58371),
	.w8(32'h3aa42fc5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a4eff),
	.w1(32'hbb1615c0),
	.w2(32'hb9aeedfe),
	.w3(32'h3aac7924),
	.w4(32'hba6f11dc),
	.w5(32'h387e3505),
	.w6(32'h3b4ab540),
	.w7(32'h3a987df3),
	.w8(32'h3aae7aa1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ab272),
	.w1(32'h3bb591b9),
	.w2(32'h3993715b),
	.w3(32'h3bb97cab),
	.w4(32'h3a04cb9e),
	.w5(32'hbbc621e2),
	.w6(32'h3bfff48d),
	.w7(32'hba10592c),
	.w8(32'hbaff3043),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd9329),
	.w1(32'hbb705d95),
	.w2(32'h3a6fb990),
	.w3(32'hbbcbd02c),
	.w4(32'hbba5825c),
	.w5(32'h3b75835a),
	.w6(32'hbbd8bea9),
	.w7(32'h3ab91b73),
	.w8(32'h3bf90185),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11e8a),
	.w1(32'hba8b7713),
	.w2(32'h3abee63b),
	.w3(32'h39fc0096),
	.w4(32'hba2ef1ba),
	.w5(32'h3b268a70),
	.w6(32'h3a51a5eb),
	.w7(32'h3a7d72d5),
	.w8(32'h3b68fe90),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba978540),
	.w1(32'hbabf1e9f),
	.w2(32'hba8ed1cc),
	.w3(32'hb91c24e9),
	.w4(32'hb9fcca12),
	.w5(32'hba2b0493),
	.w6(32'hba1e84ce),
	.w7(32'hba5e3473),
	.w8(32'hb9c37edb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688afc),
	.w1(32'hbb838c17),
	.w2(32'hbaaf3169),
	.w3(32'h3987442b),
	.w4(32'h3a0bcb68),
	.w5(32'h3b25e8b8),
	.w6(32'h393be081),
	.w7(32'h3a6ba0fd),
	.w8(32'h3b9571e2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb201e6d),
	.w1(32'hbb3d3612),
	.w2(32'h3ac2f9d0),
	.w3(32'hb9d1aa83),
	.w4(32'hbaa0b8db),
	.w5(32'h3b3e1ca7),
	.w6(32'hba475f5c),
	.w7(32'hb730f764),
	.w8(32'h3baa1aa5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87fa32),
	.w1(32'hbb3a028c),
	.w2(32'h3a61de4b),
	.w3(32'hbb1d6331),
	.w4(32'hba8a39d6),
	.w5(32'h3b256acf),
	.w6(32'hbadb2eb6),
	.w7(32'h39af497d),
	.w8(32'h3b869e5a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009721),
	.w1(32'h3a74943c),
	.w2(32'hb9d961ff),
	.w3(32'h3ab67ac7),
	.w4(32'h39f46636),
	.w5(32'hba53ee4a),
	.w6(32'h3b14b3ab),
	.w7(32'h38e31add),
	.w8(32'hb993d3fb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f21834),
	.w1(32'h3941ed96),
	.w2(32'h36d5d14d),
	.w3(32'h3749b64b),
	.w4(32'hb91a19fa),
	.w5(32'h379ad423),
	.w6(32'h399ef360),
	.w7(32'h3983496c),
	.w8(32'h3a3c6e9f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd56c),
	.w1(32'h3ad63f67),
	.w2(32'hbafdabd7),
	.w3(32'h3b561d32),
	.w4(32'hbb011fbf),
	.w5(32'hbb86d491),
	.w6(32'h3bcc3071),
	.w7(32'hba102934),
	.w8(32'hba4db1fd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6aef6),
	.w1(32'h3a862df2),
	.w2(32'h3a195beb),
	.w3(32'h39ccc06b),
	.w4(32'h3920ef60),
	.w5(32'hb9bc2766),
	.w6(32'h39a2ca33),
	.w7(32'h3a493334),
	.w8(32'h3966bb92),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7734b6),
	.w1(32'hbb85b29c),
	.w2(32'hbb5fb4fa),
	.w3(32'h3afdd346),
	.w4(32'h3b032975),
	.w5(32'h3a37bf63),
	.w6(32'hb92ff7cd),
	.w7(32'h398b2729),
	.w8(32'h3b07770b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391606c1),
	.w1(32'h39ea4b71),
	.w2(32'h3a616f44),
	.w3(32'hb8291d4e),
	.w4(32'h38fec72c),
	.w5(32'h3a1881fb),
	.w6(32'hb976d9da),
	.w7(32'hb946a040),
	.w8(32'h394a8935),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b7f4),
	.w1(32'hbb12155a),
	.w2(32'hb8b1a2a1),
	.w3(32'h39515739),
	.w4(32'h3a485f13),
	.w5(32'h3b14529c),
	.w6(32'h3aba1489),
	.w7(32'h39c46642),
	.w8(32'h3b805ef9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981e8d9),
	.w1(32'hb8c9e8e5),
	.w2(32'hb8831ea5),
	.w3(32'hb9bcbb4d),
	.w4(32'hb946de3f),
	.w5(32'hb8c9e4bd),
	.w6(32'hb98d749d),
	.w7(32'hb947cd01),
	.w8(32'hb90d30bd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a5d80),
	.w1(32'h39e59735),
	.w2(32'hb7e68e58),
	.w3(32'h3a13e66c),
	.w4(32'h39a9f0f0),
	.w5(32'h398994b7),
	.w6(32'h3a09473a),
	.w7(32'h397d4abc),
	.w8(32'h39af37a3),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb046ba3),
	.w1(32'hbae297f2),
	.w2(32'h3ad695d7),
	.w3(32'hba00e2c4),
	.w4(32'hb8c382a1),
	.w5(32'h3aeac760),
	.w6(32'h38c10345),
	.w7(32'h3aa2b83e),
	.w8(32'h3b6c23b1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7752d8),
	.w1(32'hbb9baac6),
	.w2(32'hbb942ae2),
	.w3(32'h3bbd3c8c),
	.w4(32'h3b0496e3),
	.w5(32'h3b17e2a9),
	.w6(32'h3c12770a),
	.w7(32'hbabc28ed),
	.w8(32'hb9d50f6e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac41338),
	.w1(32'hba8b6efc),
	.w2(32'h3a59a3cd),
	.w3(32'hbabf6e56),
	.w4(32'hbac36264),
	.w5(32'h39ca8da3),
	.w6(32'hb94d05a5),
	.w7(32'hba8b4120),
	.w8(32'h3a4e9063),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cab72),
	.w1(32'hbb811228),
	.w2(32'hb85f487c),
	.w3(32'h3af5092c),
	.w4(32'hb89d076b),
	.w5(32'h3b3cbad5),
	.w6(32'h3a75ea64),
	.w7(32'h3b22b4e4),
	.w8(32'h3bbd829d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40217),
	.w1(32'hbac837ba),
	.w2(32'hb9052a67),
	.w3(32'hba860c61),
	.w4(32'hbabd4474),
	.w5(32'h39d4adcd),
	.w6(32'hbb35fdc9),
	.w7(32'hbada57a3),
	.w8(32'hb998d536),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcfce7),
	.w1(32'hbbdd6b6e),
	.w2(32'hbb247d52),
	.w3(32'h3bbd4f83),
	.w4(32'hbc15aadc),
	.w5(32'hbb0e76dc),
	.w6(32'h3b7fa2c7),
	.w7(32'hbc18809c),
	.w8(32'hbb5128da),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40427a),
	.w1(32'hb98347a2),
	.w2(32'h3b0e1364),
	.w3(32'h3b0caebc),
	.w4(32'hbb29b8a0),
	.w5(32'hbb08e660),
	.w6(32'h3b94b907),
	.w7(32'hb8b231f6),
	.w8(32'h39986d2f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9dda9),
	.w1(32'hbb05a925),
	.w2(32'hbb5d14f4),
	.w3(32'h3bc76b5d),
	.w4(32'hbb7b381e),
	.w5(32'hbb8a9d89),
	.w6(32'h3be071ea),
	.w7(32'hbb43d1fa),
	.w8(32'hba8c747d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d57834),
	.w1(32'hb90ae62e),
	.w2(32'hb8e40bb9),
	.w3(32'hba3e12eb),
	.w4(32'hb9e9ba2a),
	.w5(32'hb9eac8d3),
	.w6(32'hba53b020),
	.w7(32'hba0cc8cc),
	.w8(32'hb9e5feaf),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f8af),
	.w1(32'hb8b7231f),
	.w2(32'hbb278089),
	.w3(32'h3b1f233a),
	.w4(32'hbb0c9dd2),
	.w5(32'hbb840f4e),
	.w6(32'h3b2b137e),
	.w7(32'hbac86996),
	.w8(32'hbadd1da9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a55732),
	.w1(32'h3771f6a1),
	.w2(32'hb875b4e3),
	.w3(32'hb7a0e9e4),
	.w4(32'hb734a8b2),
	.w5(32'hb8986b02),
	.w6(32'hb8594d65),
	.w7(32'hb86f93ab),
	.w8(32'hb8f062ca),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d22b45),
	.w1(32'hba4c302e),
	.w2(32'hba5af5b3),
	.w3(32'hb953a206),
	.w4(32'hba2f7e90),
	.w5(32'hba08b681),
	.w6(32'h3a79c2b3),
	.w7(32'h3a33291b),
	.w8(32'h3a63822d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913b52c),
	.w1(32'hba7a1740),
	.w2(32'hba68a045),
	.w3(32'h3a48f86a),
	.w4(32'hb98df60b),
	.w5(32'h37934492),
	.w6(32'h380c9c24),
	.w7(32'h39bc9713),
	.w8(32'h3a1c5ee2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba41dfd),
	.w1(32'hb838a679),
	.w2(32'hbb0f9e30),
	.w3(32'h3b660444),
	.w4(32'hbae57590),
	.w5(32'hbb1d83aa),
	.w6(32'h3b82c41a),
	.w7(32'hba71aa5d),
	.w8(32'h3a56df37),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ce9b9),
	.w1(32'h372b0384),
	.w2(32'hb7a25b01),
	.w3(32'h37461a10),
	.w4(32'h3784c8ca),
	.w5(32'hb7669914),
	.w6(32'hb7841cb4),
	.w7(32'h34544940),
	.w8(32'hb78ffb53),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b7c183),
	.w1(32'h389a65ff),
	.w2(32'h38b5c12a),
	.w3(32'hb6ba9bf2),
	.w4(32'h38b2598f),
	.w5(32'h38b052da),
	.w6(32'hb8c71ffa),
	.w7(32'h384365eb),
	.w8(32'h38da86aa),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d315),
	.w1(32'hbac7a507),
	.w2(32'hba8e3d89),
	.w3(32'h3832616b),
	.w4(32'hb918b7a6),
	.w5(32'hbaa155e3),
	.w6(32'hb9941873),
	.w7(32'h39a133fa),
	.w8(32'h3888b6e6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c359b),
	.w1(32'hbafee37d),
	.w2(32'h3b195934),
	.w3(32'h3b71be7d),
	.w4(32'hbb54dbdf),
	.w5(32'h3b37e585),
	.w6(32'h3b1974ee),
	.w7(32'hbaf7fb03),
	.w8(32'hba7ba03a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd573),
	.w1(32'h3ba23489),
	.w2(32'h3afef71a),
	.w3(32'h3bd8921c),
	.w4(32'h3b0f86ff),
	.w5(32'hba51c10f),
	.w6(32'h3b17cff7),
	.w7(32'h3ac32ce9),
	.w8(32'h3b2a7a2e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eee21f),
	.w1(32'hb9bc91c2),
	.w2(32'h37bacb1e),
	.w3(32'h3a01c879),
	.w4(32'hb9958167),
	.w5(32'h39d74e47),
	.w6(32'h39f3e8e2),
	.w7(32'h39df8efc),
	.w8(32'h3a1ca775),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c582934),
	.w1(32'hbaed8715),
	.w2(32'hbbe2139e),
	.w3(32'h3c67086b),
	.w4(32'hbb1110f1),
	.w5(32'hbba1292b),
	.w6(32'h3c1653d1),
	.w7(32'hbb5059f6),
	.w8(32'hbb1771d3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c663),
	.w1(32'hbba5774d),
	.w2(32'h3b91d98f),
	.w3(32'hbb827a06),
	.w4(32'hbbab81e9),
	.w5(32'h3a8628c4),
	.w6(32'hbb47dfaa),
	.w7(32'h3b15b38b),
	.w8(32'h3c063f0a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84c11f),
	.w1(32'h3b098176),
	.w2(32'h3aa81834),
	.w3(32'h3a90fade),
	.w4(32'h3a8c46bd),
	.w5(32'hba2c8658),
	.w6(32'h3ac1f634),
	.w7(32'h3ac6c69b),
	.w8(32'h39216a88),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386777ff),
	.w1(32'h382f4707),
	.w2(32'hb8199d9a),
	.w3(32'h388cc345),
	.w4(32'h37aad189),
	.w5(32'hb709b127),
	.w6(32'h37f8d050),
	.w7(32'h37c4b7e7),
	.w8(32'h371cc4a4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890df41),
	.w1(32'hb895c8f3),
	.w2(32'h378eb739),
	.w3(32'hb6ab2d5a),
	.w4(32'h367ce34c),
	.w5(32'h38c24cb7),
	.w6(32'hb8a300aa),
	.w7(32'h3882d8f9),
	.w8(32'h39093faf),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb773c9af),
	.w1(32'h37a4a1a3),
	.w2(32'hb7a10e5c),
	.w3(32'hb7641f15),
	.w4(32'h36864f24),
	.w5(32'hb82ed5ca),
	.w6(32'hb816b46a),
	.w7(32'hb78aae68),
	.w8(32'hb867a4ab),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398154ce),
	.w1(32'h3b191309),
	.w2(32'h3b437056),
	.w3(32'h3ac51408),
	.w4(32'h3b1ee348),
	.w5(32'h3ae7e730),
	.w6(32'h3b46f1e9),
	.w7(32'h3ae6560a),
	.w8(32'h3ab54fbb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd403e),
	.w1(32'hba4e887a),
	.w2(32'hb9853190),
	.w3(32'h3acd9edb),
	.w4(32'hba38621f),
	.w5(32'h39c52995),
	.w6(32'h3b4f787c),
	.w7(32'h383e6e9e),
	.w8(32'h3ab9b800),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada550a),
	.w1(32'hbb9c85cf),
	.w2(32'h3a273ab8),
	.w3(32'h3a4e762b),
	.w4(32'hbb964266),
	.w5(32'h38177fec),
	.w6(32'h3ab7dc9c),
	.w7(32'h3a2cee28),
	.w8(32'h3ba8c17f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd01a9),
	.w1(32'hbacf4c60),
	.w2(32'hbabad615),
	.w3(32'hb9a56d91),
	.w4(32'hb98e6220),
	.w5(32'h39c81452),
	.w6(32'h382217f4),
	.w7(32'h3989242d),
	.w8(32'h3a23372f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ebe33),
	.w1(32'hba6de877),
	.w2(32'hba31b378),
	.w3(32'h3b71f112),
	.w4(32'hbaf2537b),
	.w5(32'hba09f9d1),
	.w6(32'h3bd83a8a),
	.w7(32'hb9f75fd9),
	.w8(32'h3b180e5b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5be658),
	.w1(32'h39348f65),
	.w2(32'h39283919),
	.w3(32'h3b04b600),
	.w4(32'h3af0eded),
	.w5(32'h3a001f1e),
	.w6(32'h3a008e7e),
	.w7(32'hb9a2fe50),
	.w8(32'hba7588d6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816376a),
	.w1(32'hb791478f),
	.w2(32'hb8aef0ca),
	.w3(32'hb85aa705),
	.w4(32'hb8143b3f),
	.w5(32'hb8c324e9),
	.w6(32'hb8b4cfd6),
	.w7(32'hb87b29c7),
	.w8(32'hb8e4854d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51b42a),
	.w1(32'hb98c2bf2),
	.w2(32'h3ae9fd05),
	.w3(32'h3a998aac),
	.w4(32'hbac5b946),
	.w5(32'hba8b7b1f),
	.w6(32'h398de553),
	.w7(32'hba7d89ea),
	.w8(32'hbaca8888),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883283a),
	.w1(32'h379fbd1f),
	.w2(32'hb9137b44),
	.w3(32'hb8cd0ad8),
	.w4(32'hb6124a9c),
	.w5(32'hb92054dc),
	.w6(32'hb93b1c01),
	.w7(32'hb8acd652),
	.w8(32'hb94ce931),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2589c),
	.w1(32'hb99884e7),
	.w2(32'h390ba968),
	.w3(32'h3a6d6823),
	.w4(32'h3a1d1eec),
	.w5(32'h38d481f2),
	.w6(32'h3afd1c0c),
	.w7(32'h395632d4),
	.w8(32'h3a985423),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f3cc2),
	.w1(32'hbb70da81),
	.w2(32'h3ad65db6),
	.w3(32'hbb012bf4),
	.w4(32'hbad1dda7),
	.w5(32'h3b6c2c82),
	.w6(32'h39e0572c),
	.w7(32'h3b1d7b56),
	.w8(32'h3c05309f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0177a1),
	.w1(32'hbb5b8206),
	.w2(32'h394cacc9),
	.w3(32'h39c6db27),
	.w4(32'hba82170e),
	.w5(32'h3b0e71a2),
	.w6(32'h3ae39382),
	.w7(32'h3ad52c51),
	.w8(32'h3ba8b523),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e5a48),
	.w1(32'h36163178),
	.w2(32'h3a8664fc),
	.w3(32'hb9b5669d),
	.w4(32'h3980bf55),
	.w5(32'h3abaa1e0),
	.w6(32'hb98e5841),
	.w7(32'h39075259),
	.w8(32'h3aa5bd25),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83635c),
	.w1(32'hbb9e3f87),
	.w2(32'h39b3fbe0),
	.w3(32'hbb06bc0b),
	.w4(32'hbb0f2220),
	.w5(32'h3b150215),
	.w6(32'hb9a89215),
	.w7(32'h3b2b1519),
	.w8(32'h3c0c67eb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67f407),
	.w1(32'h3a0b8138),
	.w2(32'hb9714b75),
	.w3(32'h3b36d99c),
	.w4(32'hbac97867),
	.w5(32'hbb21d04a),
	.w6(32'h3b983fa2),
	.w7(32'hba0ebbee),
	.w8(32'hbae91a3d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae98ea1),
	.w1(32'hbbb07bc8),
	.w2(32'hbb770cb2),
	.w3(32'h3b403c34),
	.w4(32'hbb956d2d),
	.w5(32'hbb146ea8),
	.w6(32'h3b8b6109),
	.w7(32'hb920c4ff),
	.w8(32'h3b196339),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd37bd),
	.w1(32'hb8f72822),
	.w2(32'hb929464b),
	.w3(32'hb8bf2b71),
	.w4(32'hb8c082fb),
	.w5(32'hb93918e7),
	.w6(32'hb8e0ef38),
	.w7(32'hb87236f5),
	.w8(32'hb8b60666),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f7a62),
	.w1(32'h382e8bde),
	.w2(32'hb7a593df),
	.w3(32'hb818956d),
	.w4(32'h39999153),
	.w5(32'h3a0999c9),
	.w6(32'hb90c533c),
	.w7(32'h38e13486),
	.w8(32'h39a3af5a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb131cc0),
	.w1(32'hbb356461),
	.w2(32'hbb2fb1c5),
	.w3(32'h3ba124a0),
	.w4(32'h39132cde),
	.w5(32'h3a185e47),
	.w6(32'h3bf59ec8),
	.w7(32'h39aea17b),
	.w8(32'h3aaf05f3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7321c),
	.w1(32'hbb79a464),
	.w2(32'hbb242f9c),
	.w3(32'h3bb5f76b),
	.w4(32'h393fe991),
	.w5(32'h3b321cdf),
	.w6(32'h3c054e06),
	.w7(32'hba77c050),
	.w8(32'hb9a91b3b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd6639),
	.w1(32'hbb7decc1),
	.w2(32'hbab35ef4),
	.w3(32'h3b473a07),
	.w4(32'hbb34b7c9),
	.w5(32'hba627fb8),
	.w6(32'h3b801333),
	.w7(32'hb6818d0c),
	.w8(32'h3b4a9abe),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbda922),
	.w1(32'h3ba84934),
	.w2(32'hbb5b1981),
	.w3(32'h3b4d9d4f),
	.w4(32'h3b7fbcc2),
	.w5(32'hbaeac57f),
	.w6(32'h3b9f59f9),
	.w7(32'h3b79b1f0),
	.w8(32'hbb127bd3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45359a),
	.w1(32'h3a419f98),
	.w2(32'h38993f5d),
	.w3(32'h3a42b3e1),
	.w4(32'h39e8ce78),
	.w5(32'h3988d14a),
	.w6(32'h3a84472b),
	.w7(32'h3a6d08fb),
	.w8(32'h39e2b5cd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71e40f),
	.w1(32'h39da24f6),
	.w2(32'hba3908f1),
	.w3(32'h3a067dfe),
	.w4(32'hb9cbb078),
	.w5(32'hbaee63fa),
	.w6(32'h3a1516d9),
	.w7(32'hba085cca),
	.w8(32'hbacf1af5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ea8b0),
	.w1(32'h3b1f9e59),
	.w2(32'h3b84e17d),
	.w3(32'h3c31d8b2),
	.w4(32'h3c00f74e),
	.w5(32'h3bc06701),
	.w6(32'h3c0ca2aa),
	.w7(32'hb9935857),
	.w8(32'hbb0c73e8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f53fa),
	.w1(32'h3952adf2),
	.w2(32'hbba21963),
	.w3(32'h3c1cff5d),
	.w4(32'hba84ec1c),
	.w5(32'hbb4abd98),
	.w6(32'h3c147743),
	.w7(32'hbb12b9c9),
	.w8(32'hb9ba3962),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba61a5),
	.w1(32'h3b8cdcba),
	.w2(32'hba4e3df4),
	.w3(32'h3baf7c11),
	.w4(32'h3b4e6224),
	.w5(32'hbb10d5d3),
	.w6(32'h3c0b3713),
	.w7(32'h3a24c186),
	.w8(32'hba98a0e0),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5724),
	.w1(32'hbbad17c0),
	.w2(32'hb99a09ab),
	.w3(32'hbb4b9928),
	.w4(32'h3a240d8b),
	.w5(32'h3bb6429b),
	.w6(32'hbb02f24e),
	.w7(32'h3b32e24e),
	.w8(32'h3bfc32c3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb66912),
	.w1(32'hbb7d694c),
	.w2(32'h3b2361b9),
	.w3(32'hbb40bb46),
	.w4(32'hbacca344),
	.w5(32'h3b704661),
	.w6(32'hb9c95475),
	.w7(32'h3b975258),
	.w8(32'h3c39a129),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81dd2d7),
	.w1(32'hb7bcf927),
	.w2(32'hb81e5751),
	.w3(32'hb80fea1c),
	.w4(32'hb7b233da),
	.w5(32'hb80eb43e),
	.w6(32'hb83121cf),
	.w7(32'hb7e05760),
	.w8(32'hb81049ae),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811da35),
	.w1(32'hb74dff33),
	.w2(32'hb83993d1),
	.w3(32'hb830697d),
	.w4(32'hb7d82563),
	.w5(32'hb86dc198),
	.w6(32'hb881ae01),
	.w7(32'hb837f727),
	.w8(32'hb89a3724),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb2c37),
	.w1(32'hbb057bdc),
	.w2(32'hbb43979a),
	.w3(32'hba785b96),
	.w4(32'hba363442),
	.w5(32'hbadae8b3),
	.w6(32'h3a006bab),
	.w7(32'hb8d2e67e),
	.w8(32'h3997b63d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb703e9d7),
	.w1(32'h37ca6fa6),
	.w2(32'hb8155f71),
	.w3(32'hb807e79f),
	.w4(32'h377d34c2),
	.w5(32'hb82b5a1a),
	.w6(32'hb85bcd18),
	.w7(32'hb744ab1c),
	.w8(32'hb888bd64),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf7c08),
	.w1(32'h3ad61e9a),
	.w2(32'h3b0569a1),
	.w3(32'h3ac5b6c6),
	.w4(32'h3afab7db),
	.w5(32'h3aa0bc64),
	.w6(32'h3af1af70),
	.w7(32'h3a844bf8),
	.w8(32'h3a1c1ec8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b705add),
	.w1(32'h3a9ffa80),
	.w2(32'hbb3097cc),
	.w3(32'h3bb8ff26),
	.w4(32'h3b3034fd),
	.w5(32'hb961e74d),
	.w6(32'h3bf645cc),
	.w7(32'h3b0c7824),
	.w8(32'h394683a8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95875a),
	.w1(32'hbb23be30),
	.w2(32'hba6f287d),
	.w3(32'h3b0a3c87),
	.w4(32'h3a3decbc),
	.w5(32'h3adcd0dd),
	.w6(32'h3b2ec888),
	.w7(32'h3aba612b),
	.w8(32'h3b11786f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e8a4bc),
	.w1(32'hb80e8a84),
	.w2(32'hb82fa2ce),
	.w3(32'hb86fb616),
	.w4(32'hb87edc64),
	.w5(32'hb8aa68b2),
	.w6(32'hb8b7b1ca),
	.w7(32'hb8652ba4),
	.w8(32'hb8156901),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fe444),
	.w1(32'h3bcec212),
	.w2(32'h3ae4b7da),
	.w3(32'h3c329396),
	.w4(32'h3b7dbe2f),
	.w5(32'hbb74cf41),
	.w6(32'h3c4f5b97),
	.w7(32'h3965fdfa),
	.w8(32'hbbf7bcb7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51d0d2),
	.w1(32'hb835fc78),
	.w2(32'hbac844dd),
	.w3(32'h3b391289),
	.w4(32'hba9d1317),
	.w5(32'hbaf3f4b8),
	.w6(32'h3b701b5e),
	.w7(32'hba12f6f7),
	.w8(32'hb9f2fbb3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39825414),
	.w1(32'h38a416f4),
	.w2(32'h352ba51f),
	.w3(32'h398eed31),
	.w4(32'hb8dac5af),
	.w5(32'hb99531ca),
	.w6(32'h38f6f06c),
	.w7(32'hb9d8f67d),
	.w8(32'hb9ec536e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801466),
	.w1(32'h3b281edd),
	.w2(32'hba3af623),
	.w3(32'h3b62f87c),
	.w4(32'h3a83f789),
	.w5(32'hba97b444),
	.w6(32'h3ba01620),
	.w7(32'h39c78906),
	.w8(32'hba62af0d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ef444),
	.w1(32'hb8c9cebb),
	.w2(32'h36c58b8b),
	.w3(32'hb92006e6),
	.w4(32'hb92341a2),
	.w5(32'hb88f803f),
	.w6(32'hb835abb5),
	.w7(32'hb8b2e673),
	.w8(32'hb80cc999),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9144421),
	.w1(32'hb934f91e),
	.w2(32'hb9bf7cec),
	.w3(32'hb932d99f),
	.w4(32'hb9bdd721),
	.w5(32'hba0a36c9),
	.w6(32'h39d91ad3),
	.w7(32'h3824963d),
	.w8(32'hb913cdfc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e7a31c),
	.w1(32'hb80f8dfd),
	.w2(32'hb8ab147d),
	.w3(32'hb6044d5a),
	.w4(32'hb87e5d3e),
	.w5(32'hb8bc5acc),
	.w6(32'h32bd92e8),
	.w7(32'hb846f263),
	.w8(32'hb89b740b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6fcb5),
	.w1(32'hb848b426),
	.w2(32'hb78d9528),
	.w3(32'hb8325ddc),
	.w4(32'hb888d186),
	.w5(32'hb8acbc86),
	.w6(32'hb84238cb),
	.w7(32'hb849d442),
	.w8(32'hb91444f3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0bb9),
	.w1(32'hbb2abed8),
	.w2(32'hba66df25),
	.w3(32'hb9651164),
	.w4(32'h3a88253e),
	.w5(32'h3b02b444),
	.w6(32'h39c39025),
	.w7(32'h3abf993c),
	.w8(32'h3b2bb4f8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14379b),
	.w1(32'h3a0b1d56),
	.w2(32'hb8b6c581),
	.w3(32'h3b94a1f6),
	.w4(32'hbbb91f29),
	.w5(32'hbb8af285),
	.w6(32'h3c00070a),
	.w7(32'hbb59ce88),
	.w8(32'hb89cf296),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be546a5),
	.w1(32'h3b303404),
	.w2(32'hba5cde05),
	.w3(32'h3bceb8bf),
	.w4(32'hba51dc6b),
	.w5(32'hbb4dfa63),
	.w6(32'h3bd3373a),
	.w7(32'hbabbb378),
	.w8(32'hbb16f336),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4aed),
	.w1(32'h386ba08d),
	.w2(32'hbab2d606),
	.w3(32'h3b8f9bbf),
	.w4(32'hbb8a3970),
	.w5(32'hbb9eed20),
	.w6(32'h3badb15d),
	.w7(32'hbb608b55),
	.w8(32'hbb520085),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9980195),
	.w1(32'hb97ec17f),
	.w2(32'h38a9b3d8),
	.w3(32'hb9615f8c),
	.w4(32'hb9728351),
	.w5(32'h38ade6d2),
	.w6(32'hb8fca681),
	.w7(32'hb929258f),
	.w8(32'h38fb8942),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ab7f6),
	.w1(32'h38c0f6b3),
	.w2(32'hba2215f8),
	.w3(32'h3914a9bd),
	.w4(32'hb9dc9b94),
	.w5(32'hba5f6075),
	.w6(32'h39bca5bc),
	.w7(32'hb800a856),
	.w8(32'hb8ec4a6e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f6a64),
	.w1(32'h37e2e081),
	.w2(32'hb7e022fb),
	.w3(32'h38e82993),
	.w4(32'h37f26b77),
	.w5(32'hb89d655c),
	.w6(32'h37fec98d),
	.w7(32'hb7c97339),
	.w8(32'hb88c3b4d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c17641),
	.w1(32'hb731c7fc),
	.w2(32'hb86a3317),
	.w3(32'hb7717573),
	.w4(32'h3604e0dc),
	.w5(32'hb822f1c5),
	.w6(32'hb8129ea4),
	.w7(32'hb70f748e),
	.w8(32'hb8138757),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9331d),
	.w1(32'hb7776c34),
	.w2(32'hbb5462ec),
	.w3(32'h3b5f6418),
	.w4(32'hbb9096d4),
	.w5(32'hbb8a5b26),
	.w6(32'h3b6d4438),
	.w7(32'hbb3a307e),
	.w8(32'hbaa3c2e4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394516ca),
	.w1(32'h37a30925),
	.w2(32'h38a97dbb),
	.w3(32'h39512512),
	.w4(32'h3928e7a9),
	.w5(32'h391060a2),
	.w6(32'h38332d47),
	.w7(32'h39654aba),
	.w8(32'h396ebff3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf6993),
	.w1(32'hb917f977),
	.w2(32'h3acb1a35),
	.w3(32'hb9a2bad4),
	.w4(32'hb9b71b3c),
	.w5(32'h3ada2ca8),
	.w6(32'h38933d17),
	.w7(32'hb9b9c930),
	.w8(32'h3ad70994),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b9b9a),
	.w1(32'h3a5bb169),
	.w2(32'h3a31fdab),
	.w3(32'h3b2009c9),
	.w4(32'h39b909cf),
	.w5(32'h39f21a0e),
	.w6(32'h396303c7),
	.w7(32'hba738826),
	.w8(32'hba952bf1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883416a),
	.w1(32'h37d071e2),
	.w2(32'h3817115d),
	.w3(32'hb8a87952),
	.w4(32'h389aa06c),
	.w5(32'h39060c65),
	.w6(32'hb8a70ae5),
	.w7(32'h388428de),
	.w8(32'h390d488a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cee9f),
	.w1(32'hba6b7405),
	.w2(32'hba97c353),
	.w3(32'h3a2a3669),
	.w4(32'hba7755ec),
	.w5(32'hba04b661),
	.w6(32'h3a9dc07d),
	.w7(32'hb8cea657),
	.w8(32'h39f1cf58),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e2567),
	.w1(32'h39bc6599),
	.w2(32'h39ebf404),
	.w3(32'hb6fbaf5e),
	.w4(32'h383352b4),
	.w5(32'h39762741),
	.w6(32'h39cc9480),
	.w7(32'h398da24a),
	.w8(32'h39d5d41a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56ae57),
	.w1(32'h3aed2c68),
	.w2(32'hb9ad8296),
	.w3(32'h3b8ebf47),
	.w4(32'hbc0bc714),
	.w5(32'hbc1efed1),
	.w6(32'h3ba30a2f),
	.w7(32'hbbe7e404),
	.w8(32'hbb90643a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9003d),
	.w1(32'h3b8fae70),
	.w2(32'h3a5d9752),
	.w3(32'h375fe0e8),
	.w4(32'h3adab55c),
	.w5(32'h3a58c06a),
	.w6(32'h3b72bf74),
	.w7(32'h3af59213),
	.w8(32'h3aeda502),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c552fe),
	.w1(32'hbb46828c),
	.w2(32'hbbeb2b8d),
	.w3(32'h3c0d7daf),
	.w4(32'h3b62cc81),
	.w5(32'h3b2ec0bf),
	.w6(32'h3bc9d6ec),
	.w7(32'h3a9c91f0),
	.w8(32'hb8c54017),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule