module layer_8_featuremap_108(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c272e47),
	.w1(32'h3affb18a),
	.w2(32'hbab4b95c),
	.w3(32'h3c596cdb),
	.w4(32'h3a93fd33),
	.w5(32'hbb8d96e2),
	.w6(32'h3c830141),
	.w7(32'h3bf7b749),
	.w8(32'h3c387b3b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb33c9e),
	.w1(32'h3b875948),
	.w2(32'hbb6bc240),
	.w3(32'h3bddd210),
	.w4(32'hbbb12489),
	.w5(32'hbc4ec733),
	.w6(32'hbb5318f1),
	.w7(32'h3b2bb27c),
	.w8(32'h3afde9b9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2db79),
	.w1(32'h3aa0b3a2),
	.w2(32'h3c06189f),
	.w3(32'h3b65d419),
	.w4(32'hbae8cb4e),
	.w5(32'hbcc44e8b),
	.w6(32'h3a929cc9),
	.w7(32'h3bb202ef),
	.w8(32'hbc6d9d7d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd0507),
	.w1(32'hbcceff54),
	.w2(32'h3b8a8d51),
	.w3(32'h3bdbb90a),
	.w4(32'hbb180afd),
	.w5(32'hbcb2f000),
	.w6(32'hbc12dfef),
	.w7(32'h3c1cb1c5),
	.w8(32'h3c5692b5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d208e01),
	.w1(32'h3b443f4e),
	.w2(32'hbbb47c37),
	.w3(32'hbc823abd),
	.w4(32'hbc615514),
	.w5(32'hbae807fd),
	.w6(32'hbc080bf7),
	.w7(32'hbc377d06),
	.w8(32'hbcd68a16),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3da0b3),
	.w1(32'hbc920de1),
	.w2(32'hbbe3f7c2),
	.w3(32'h3c4c2c36),
	.w4(32'h3c16a9cb),
	.w5(32'h3a96ef83),
	.w6(32'hbc01857c),
	.w7(32'h3b1a21f9),
	.w8(32'h3caf3736),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee31e),
	.w1(32'h3c15c19d),
	.w2(32'h3b98465f),
	.w3(32'hbc3430b9),
	.w4(32'h3ba7f023),
	.w5(32'hbb1628be),
	.w6(32'hbc066dd4),
	.w7(32'h3c3bf2b8),
	.w8(32'h3cb9b284),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f5593),
	.w1(32'hbc28d863),
	.w2(32'hbbe10123),
	.w3(32'hbc53a9fb),
	.w4(32'h3a90f914),
	.w5(32'hbae85c2b),
	.w6(32'hbcc637ad),
	.w7(32'hba49ed2a),
	.w8(32'hbb8bc2e5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ebf64),
	.w1(32'h3c339b14),
	.w2(32'hbb013ea6),
	.w3(32'h3c3db4c3),
	.w4(32'h3c0c80ca),
	.w5(32'hbc0c72d9),
	.w6(32'h3ac13f76),
	.w7(32'hbb3362a8),
	.w8(32'h3a788b4e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed6346),
	.w1(32'h3bfdc8cc),
	.w2(32'h3c51badb),
	.w3(32'hba0c23f0),
	.w4(32'h3c846a02),
	.w5(32'hbc4803fb),
	.w6(32'h3b0c99da),
	.w7(32'h3ce28ee7),
	.w8(32'h3d672007),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d247eb4),
	.w1(32'h3c48d964),
	.w2(32'h3b460ba1),
	.w3(32'hbd644bd1),
	.w4(32'hbc6de7db),
	.w5(32'h38316256),
	.w6(32'hbda3a1b6),
	.w7(32'hbc9ea7c0),
	.w8(32'hbd10f3e6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc807fdd),
	.w1(32'h3ad1da51),
	.w2(32'hbc19df64),
	.w3(32'h3b000e64),
	.w4(32'hbc56018d),
	.w5(32'hbc6a66d3),
	.w6(32'h3d628eaf),
	.w7(32'hbb12efbf),
	.w8(32'hbc38b6b3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc028be2),
	.w1(32'h39986fcd),
	.w2(32'h3b3e1fc7),
	.w3(32'hbb8cef79),
	.w4(32'hbac17c8e),
	.w5(32'h3a4740fa),
	.w6(32'h3b57c14d),
	.w7(32'hbb2600a6),
	.w8(32'hb941d88b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95e0b2),
	.w1(32'hbacad981),
	.w2(32'hba96c606),
	.w3(32'hbab68bd8),
	.w4(32'hbaae3d4d),
	.w5(32'hba29a436),
	.w6(32'hbaafcbd7),
	.w7(32'hba296fab),
	.w8(32'hba165710),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d5497),
	.w1(32'h37387c9d),
	.w2(32'hb90b3a66),
	.w3(32'hb9235764),
	.w4(32'hb94220b0),
	.w5(32'hb93ba742),
	.w6(32'hb994fd93),
	.w7(32'hb97f287e),
	.w8(32'hb968f425),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade3add),
	.w1(32'hbad6edde),
	.w2(32'hbb478c56),
	.w3(32'hbb202b69),
	.w4(32'hbaeb7611),
	.w5(32'hbb48b625),
	.w6(32'hbaa55a85),
	.w7(32'hba9bfbd7),
	.w8(32'hbb20531c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabd3b8),
	.w1(32'hbb11e2c9),
	.w2(32'hbb5d9dd1),
	.w3(32'hba7fb757),
	.w4(32'hbb27aae1),
	.w5(32'hbb8b0ad7),
	.w6(32'hba711433),
	.w7(32'hbb487465),
	.w8(32'hbb9719bd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1a768),
	.w1(32'h3b88bbf2),
	.w2(32'h3b3f0066),
	.w3(32'hba0bae58),
	.w4(32'h39c1c66e),
	.w5(32'h3b2d82c5),
	.w6(32'hb9ddaa18),
	.w7(32'h3b1a3c62),
	.w8(32'h3ba2e76e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb778268),
	.w1(32'hbc5ccdd3),
	.w2(32'hbb861687),
	.w3(32'hbba93c11),
	.w4(32'hbc28ea99),
	.w5(32'hbb146630),
	.w6(32'h3b10c4b6),
	.w7(32'h3b26cfc2),
	.w8(32'h3c0ee0b3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9886db),
	.w1(32'hbc4f02b2),
	.w2(32'hbc9366bc),
	.w3(32'hbb5b2ae9),
	.w4(32'hbbc06abe),
	.w5(32'hbc472476),
	.w6(32'hbb10ebb7),
	.w7(32'hbb29c2fe),
	.w8(32'hbc04993d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a23e4),
	.w1(32'hbb1ba853),
	.w2(32'hbba30699),
	.w3(32'hb994d326),
	.w4(32'h3a009eb7),
	.w5(32'hbb8f4cd0),
	.w6(32'h3b2ebf67),
	.w7(32'h3b63c209),
	.w8(32'hb9df6f07),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bf2a2),
	.w1(32'h3c167935),
	.w2(32'h3c03ebeb),
	.w3(32'h3bc364be),
	.w4(32'h3bb9ab85),
	.w5(32'h3bb06bf3),
	.w6(32'h3bd96316),
	.w7(32'h3bb8408a),
	.w8(32'h39c30fdd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c465e54),
	.w1(32'hbb203853),
	.w2(32'hbc5f1d30),
	.w3(32'h3c17ee0e),
	.w4(32'hbbb6d46c),
	.w5(32'hbc69ac94),
	.w6(32'h3bdc4a4a),
	.w7(32'hbb8df8fd),
	.w8(32'hbc272e91),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0de875),
	.w1(32'h3a54d811),
	.w2(32'hba170207),
	.w3(32'hbad2bf11),
	.w4(32'hbab62c12),
	.w5(32'hbaf8ba71),
	.w6(32'hbb2b2e27),
	.w7(32'hbb861cda),
	.w8(32'hbb7ae35b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd91fa),
	.w1(32'hbbeab936),
	.w2(32'hbc77555e),
	.w3(32'hba86100f),
	.w4(32'hb9183fc7),
	.w5(32'hbc417628),
	.w6(32'hbabf80d6),
	.w7(32'hb970cbfc),
	.w8(32'hbc43bc94),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beffab1),
	.w1(32'h3b8d8b4d),
	.w2(32'h399cf595),
	.w3(32'h3be7c0d4),
	.w4(32'h3b5a8238),
	.w5(32'hbb3dd9b3),
	.w6(32'h3bba7514),
	.w7(32'h3b15274e),
	.w8(32'hba1a1f7d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee8a8f),
	.w1(32'h3aa934e7),
	.w2(32'h3a11f7fc),
	.w3(32'h3b022b71),
	.w4(32'h39e62bd5),
	.w5(32'hb8af4754),
	.w6(32'h3ab7b1a1),
	.w7(32'h388be56b),
	.w8(32'hb9eb2869),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6a2f80),
	.w1(32'hbd73798b),
	.w2(32'hbd58bdfb),
	.w3(32'hbc55e719),
	.w4(32'hbb9d782f),
	.w5(32'hbc5f0c2a),
	.w6(32'hbd4056e8),
	.w7(32'hbd05fee4),
	.w8(32'hbc997c56),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b787610),
	.w1(32'h3ac38eab),
	.w2(32'h37155b9e),
	.w3(32'h3b1922c8),
	.w4(32'h3a3f26c7),
	.w5(32'hb9bfdace),
	.w6(32'h3b8a98aa),
	.w7(32'h3b382127),
	.w8(32'h3ae346df),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5c76a),
	.w1(32'h3a87572f),
	.w2(32'hbaa07055),
	.w3(32'hba49fb51),
	.w4(32'hba7ec0f1),
	.w5(32'hbb2c7325),
	.w6(32'hbaa2e7fc),
	.w7(32'hbaaec2b1),
	.w8(32'hbb90096f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7320b8),
	.w1(32'h3bb42a90),
	.w2(32'h3ba71116),
	.w3(32'h3bbe61e4),
	.w4(32'h3bc2eb43),
	.w5(32'h3bd1945b),
	.w6(32'h3bfc4fc2),
	.w7(32'h3be0f6de),
	.w8(32'h3bcde54d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a472588),
	.w1(32'hb8b1b98d),
	.w2(32'hbb1eaddf),
	.w3(32'h3b1b7fc4),
	.w4(32'h3a989aac),
	.w5(32'hbad6db33),
	.w6(32'h3b0a64ce),
	.w7(32'h3a3c0277),
	.w8(32'hb9f512b3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a97f8c),
	.w1(32'hb97a9405),
	.w2(32'hb8e1e6db),
	.w3(32'hb9659d02),
	.w4(32'hb90bd394),
	.w5(32'hb85e4a64),
	.w6(32'hb984cfeb),
	.w7(32'hb9454fdb),
	.w8(32'hb914c12c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c8f6bc),
	.w1(32'hb7a76c95),
	.w2(32'h3904409a),
	.w3(32'h37c70092),
	.w4(32'hb76ccffa),
	.w5(32'h3904a524),
	.w6(32'hb73bdca5),
	.w7(32'hb6578c12),
	.w8(32'h390fd29c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba447ea5),
	.w1(32'h3a283ba2),
	.w2(32'hba266105),
	.w3(32'hba5683bd),
	.w4(32'h3ac17465),
	.w5(32'hba56521e),
	.w6(32'h39488ce7),
	.w7(32'h3a8a1d5c),
	.w8(32'hba9f7984),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17bd65),
	.w1(32'hbba407f9),
	.w2(32'hbb80a27e),
	.w3(32'hbb0d458b),
	.w4(32'hbba3b57b),
	.w5(32'hbb7ada8d),
	.w6(32'hba2f323b),
	.w7(32'hba9fab59),
	.w8(32'hba24e5f7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994de4a),
	.w1(32'hba36b28d),
	.w2(32'hbad939a8),
	.w3(32'hba87660f),
	.w4(32'hbad42274),
	.w5(32'hbb2bb4a7),
	.w6(32'hba8f775f),
	.w7(32'hbaa221cc),
	.w8(32'hbb1ddeab),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd06e61),
	.w1(32'h3ba5a970),
	.w2(32'h3a30ea08),
	.w3(32'h3ba9d66c),
	.w4(32'h3b77b195),
	.w5(32'h3a22d652),
	.w6(32'h3bb6ade4),
	.w7(32'h3b755e83),
	.w8(32'h39ba07b1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c9192),
	.w1(32'hb967958b),
	.w2(32'hb981e3b4),
	.w3(32'h37f68d6d),
	.w4(32'hb8b1ddc2),
	.w5(32'hb9553d26),
	.w6(32'hb79bf14d),
	.w7(32'hb92b61db),
	.w8(32'h37bed06b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39215a57),
	.w1(32'h3a2a2d45),
	.w2(32'h3a1aa423),
	.w3(32'h3a829891),
	.w4(32'h3ab452b1),
	.w5(32'h3ab1e821),
	.w6(32'h39ce785b),
	.w7(32'h3a5a9f26),
	.w8(32'h3a342f24),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace7d1),
	.w1(32'h39fb9d74),
	.w2(32'hbbd5cbeb),
	.w3(32'hba95dabd),
	.w4(32'hbba48f32),
	.w5(32'hbc2e4f5e),
	.w6(32'h3af432db),
	.w7(32'h3aa18f82),
	.w8(32'hbbc02c64),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0444ee),
	.w1(32'hbb2c2469),
	.w2(32'hba865370),
	.w3(32'hbb010ca2),
	.w4(32'hbb11b6d8),
	.w5(32'hba8bb594),
	.w6(32'hba3f6f07),
	.w7(32'hba19b6b1),
	.w8(32'h3a85de8a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a3bca),
	.w1(32'hba248b80),
	.w2(32'hba799774),
	.w3(32'hba35242a),
	.w4(32'hba6607ed),
	.w5(32'hbaa680a4),
	.w6(32'hba062dcb),
	.w7(32'hba0a5c3b),
	.w8(32'hba3ef044),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10f16f),
	.w1(32'hbb4c1d24),
	.w2(32'hbb80c03d),
	.w3(32'hbb169076),
	.w4(32'hbb67b761),
	.w5(32'hbbaa7491),
	.w6(32'hbb1e25e5),
	.w7(32'hbb2e2750),
	.w8(32'hbb6312a4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842028),
	.w1(32'hb8bc8a19),
	.w2(32'hbac0b2f7),
	.w3(32'h38b3b388),
	.w4(32'hbad3a3bd),
	.w5(32'hbad37025),
	.w6(32'h3b0b6053),
	.w7(32'h3ae47adb),
	.w8(32'h39bd8454),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2d5a7),
	.w1(32'hba16e195),
	.w2(32'h3aa1ccd0),
	.w3(32'h3990154c),
	.w4(32'h3ae30e9a),
	.w5(32'h3b2aea58),
	.w6(32'h3b46875a),
	.w7(32'h3b6b5a89),
	.w8(32'h3b8bbb7e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a73dae),
	.w1(32'h35310873),
	.w2(32'h3865c76e),
	.w3(32'hb777ca39),
	.w4(32'hb74a4e8b),
	.w5(32'h38597839),
	.w6(32'hb7f8b38a),
	.w7(32'hb7b70db4),
	.w8(32'h382af856),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888b0a1),
	.w1(32'hbbf9294e),
	.w2(32'hbc54771f),
	.w3(32'hbbbcc977),
	.w4(32'hbc236db4),
	.w5(32'hbc62e70f),
	.w6(32'hbb7a4049),
	.w7(32'hbb9b2137),
	.w8(32'hbbf8c80b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29b669),
	.w1(32'hba4434b1),
	.w2(32'hb78e1d10),
	.w3(32'hba2180e9),
	.w4(32'hb9d7ab91),
	.w5(32'h39e733f0),
	.w6(32'h3a4af370),
	.w7(32'h3a9cbff4),
	.w8(32'h3b01dce7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdae944),
	.w1(32'h3b51b9b4),
	.w2(32'h39b9c800),
	.w3(32'h3a6a8ee8),
	.w4(32'hbaed05ce),
	.w5(32'hbb191982),
	.w6(32'hb89caf09),
	.w7(32'hbb110bdb),
	.w8(32'hba97e425),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26762b),
	.w1(32'h3c09d697),
	.w2(32'h3b5be360),
	.w3(32'h3c34f60d),
	.w4(32'h3c1727d7),
	.w5(32'h3b9b05c9),
	.w6(32'h3c5f73de),
	.w7(32'h3c3c5357),
	.w8(32'h3b981473),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9030c9),
	.w1(32'hbca2ccdf),
	.w2(32'hbc9771c4),
	.w3(32'hbc24f209),
	.w4(32'hbc88528d),
	.w5(32'hbc8f63c3),
	.w6(32'hbb8e1345),
	.w7(32'hbbac59b0),
	.w8(32'hbb834298),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e481c),
	.w1(32'hbb3111ff),
	.w2(32'hbbb180c3),
	.w3(32'h3ad71a6d),
	.w4(32'hbb5963bf),
	.w5(32'hbbf8e172),
	.w6(32'hb95653db),
	.w7(32'hbb37da03),
	.w8(32'hbbc5dbaa),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdc43b),
	.w1(32'hbafa02ba),
	.w2(32'hbb1ecf3a),
	.w3(32'hbaabf557),
	.w4(32'hbb32c86f),
	.w5(32'hba83e538),
	.w6(32'h3b2cf617),
	.w7(32'h3abec9da),
	.w8(32'h3b2935f1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d42cb7),
	.w1(32'hb8c3aadf),
	.w2(32'hb71c2dc6),
	.w3(32'hb82db644),
	.w4(32'hb8d03211),
	.w5(32'hb8342aaf),
	.w6(32'hb79300b1),
	.w7(32'hb8a5d879),
	.w8(32'hb7ae0e2e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbc834),
	.w1(32'hb7191679),
	.w2(32'hbbf216b4),
	.w3(32'h3b8ff129),
	.w4(32'hbaf9deb9),
	.w5(32'hbbb81735),
	.w6(32'h3b21b8ca),
	.w7(32'h3a675675),
	.w8(32'h3a4bb05a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e87f01),
	.w1(32'h3a903ab9),
	.w2(32'h3abd0094),
	.w3(32'h3a3b8c1f),
	.w4(32'h3a7207fc),
	.w5(32'h3a4c345a),
	.w6(32'h3ab3e6a0),
	.w7(32'h38ba0928),
	.w8(32'hb9c7d9c8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f1e2d),
	.w1(32'hbae55ddf),
	.w2(32'hbb38b252),
	.w3(32'hbb8d9185),
	.w4(32'hbbf8b966),
	.w5(32'hbc06d458),
	.w6(32'hbba5d2e7),
	.w7(32'hbb6d846d),
	.w8(32'hbb39e577),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c8246),
	.w1(32'hba8b2076),
	.w2(32'hbac70e93),
	.w3(32'h37adf783),
	.w4(32'hba8a7330),
	.w5(32'hba873dc6),
	.w6(32'hbac7d6dc),
	.w7(32'hba2986bd),
	.w8(32'hb917fe18),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba285f08),
	.w1(32'hbaa56677),
	.w2(32'hbb46a443),
	.w3(32'hbac79a8c),
	.w4(32'hbb035cae),
	.w5(32'hbb9279da),
	.w6(32'hbb66541e),
	.w7(32'hbb02b588),
	.w8(32'hbb6b81e6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae72852),
	.w1(32'hbb2e5b1a),
	.w2(32'hbb9d8ed8),
	.w3(32'hbb0a8f39),
	.w4(32'hbb6b46cb),
	.w5(32'hbbd3ba30),
	.w6(32'hbb7aefd6),
	.w7(32'hbb8d626d),
	.w8(32'hbbd34408),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14b89f),
	.w1(32'h3a1b9382),
	.w2(32'h39bfe7ed),
	.w3(32'h3971494d),
	.w4(32'h39f860da),
	.w5(32'h399ca5e6),
	.w6(32'h38bc0f8e),
	.w7(32'h39ae268a),
	.w8(32'h39893861),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39fad3),
	.w1(32'hbaf08ab7),
	.w2(32'hbb741da8),
	.w3(32'hbb0f1677),
	.w4(32'hbb917418),
	.w5(32'hbba70cf8),
	.w6(32'h3bab86dd),
	.w7(32'h3b69e360),
	.w8(32'h3ac15f45),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895e7d),
	.w1(32'hbb04fa77),
	.w2(32'hbaa91ffd),
	.w3(32'hb9f531d8),
	.w4(32'hbb278f94),
	.w5(32'hbacad22f),
	.w6(32'hb9ebf9fa),
	.w7(32'hbaca6330),
	.w8(32'h38ffd38d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d999),
	.w1(32'h3a642eec),
	.w2(32'h3801a55f),
	.w3(32'h3a9f5a76),
	.w4(32'hb943932a),
	.w5(32'hba99ace7),
	.w6(32'h3a1acffa),
	.w7(32'hba2722c0),
	.w8(32'hba436044),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be862d),
	.w1(32'hbb0c77b0),
	.w2(32'hbb3c2a08),
	.w3(32'hba2883f6),
	.w4(32'hbb86390e),
	.w5(32'hbbc35fa2),
	.w6(32'h390e86e9),
	.w7(32'hbb2e7fe2),
	.w8(32'hbb911325),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2c0ab),
	.w1(32'hb923223b),
	.w2(32'hbaf69f7d),
	.w3(32'h3a83e403),
	.w4(32'h39503843),
	.w5(32'hbad386e2),
	.w6(32'hbaf3e209),
	.w7(32'hba95471f),
	.w8(32'hb93b4ee8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7dd42),
	.w1(32'h38907118),
	.w2(32'hbba73d16),
	.w3(32'h3b315506),
	.w4(32'hba825a7b),
	.w5(32'hbbe65d9f),
	.w6(32'h3aa1905f),
	.w7(32'hb9d5a7c5),
	.w8(32'hbbba5046),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a031e5f),
	.w1(32'h38ae2d81),
	.w2(32'hbb3e908c),
	.w3(32'hb933627b),
	.w4(32'hba84f7c5),
	.w5(32'hbb731cc3),
	.w6(32'hba0770f5),
	.w7(32'hbaabf439),
	.w8(32'hbb1ef3e4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960d330),
	.w1(32'hbbb4ddb2),
	.w2(32'hbc22a9af),
	.w3(32'hb976dc01),
	.w4(32'hbbaab4b0),
	.w5(32'hbc427664),
	.w6(32'hbbe6332e),
	.w7(32'hbb9a826a),
	.w8(32'hbbe99730),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52811b),
	.w1(32'h3a8cfa68),
	.w2(32'h3aad7639),
	.w3(32'h3ae4d1ba),
	.w4(32'h3acd5b96),
	.w5(32'h3adbc3c0),
	.w6(32'h3aebeff7),
	.w7(32'h3ab1e695),
	.w8(32'h3ae92ba5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32e04c),
	.w1(32'h3ab65ac8),
	.w2(32'h3a2b7e9c),
	.w3(32'h3aa08dbb),
	.w4(32'hb99e7e17),
	.w5(32'hba688020),
	.w6(32'h3a50250c),
	.w7(32'hb83c8498),
	.w8(32'hba0f008b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c7af3),
	.w1(32'h3a913b1c),
	.w2(32'hba11dfdc),
	.w3(32'h39ad49e2),
	.w4(32'hba858ecc),
	.w5(32'hbaccedf2),
	.w6(32'hb99e059f),
	.w7(32'hba91a5ef),
	.w8(32'hba2694a3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b386458),
	.w1(32'hb9146a26),
	.w2(32'hbc001689),
	.w3(32'hba8a7c9a),
	.w4(32'hbb6f75e4),
	.w5(32'hbc4429bc),
	.w6(32'hbb0ab437),
	.w7(32'hbb63bb0f),
	.w8(32'hbc03bdd5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8031c20),
	.w1(32'hb8873193),
	.w2(32'hb8294bf8),
	.w3(32'hb8183785),
	.w4(32'hb88f715f),
	.w5(32'hb8212c1e),
	.w6(32'hb7796c7b),
	.w7(32'hb83beccd),
	.w8(32'h3703f26b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2401bb),
	.w1(32'hbb0f60fb),
	.w2(32'hbbf54d64),
	.w3(32'h3aef236d),
	.w4(32'hba8635ad),
	.w5(32'hbbe29855),
	.w6(32'h3a1226cb),
	.w7(32'hbad775fa),
	.w8(32'hbc011956),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998e65e),
	.w1(32'hb9a26565),
	.w2(32'h3a9d9aab),
	.w3(32'hb88d9726),
	.w4(32'hba969184),
	.w5(32'h3c36a12d),
	.w6(32'hb9145700),
	.w7(32'hbabb7b48),
	.w8(32'h3bc14acd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0527a2),
	.w1(32'hbaa85598),
	.w2(32'hbb9d9722),
	.w3(32'h3b0d2355),
	.w4(32'hbac8ca16),
	.w5(32'hbbd3afb0),
	.w6(32'hbbe6753e),
	.w7(32'h3758bd51),
	.w8(32'hbba18fd2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cb7c),
	.w1(32'hbb533071),
	.w2(32'hbaf6cb68),
	.w3(32'hbba4c6ea),
	.w4(32'hbb92531f),
	.w5(32'hbba4fc97),
	.w6(32'hbbe41925),
	.w7(32'hba1b9652),
	.w8(32'h3a853d38),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccfa88),
	.w1(32'hbbbc3e15),
	.w2(32'hbbb3f02d),
	.w3(32'hbbac9666),
	.w4(32'hbb52b223),
	.w5(32'h3b6a16f7),
	.w6(32'hbbb9f6aa),
	.w7(32'h390eaffc),
	.w8(32'h3b675bea),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb3c6d),
	.w1(32'hbb0ec8a8),
	.w2(32'hbbcc7e91),
	.w3(32'hbbb490d3),
	.w4(32'h38895d33),
	.w5(32'h3b55b8d3),
	.w6(32'hba9aecc8),
	.w7(32'hba34d16a),
	.w8(32'h3b466ed1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39390c8b),
	.w1(32'h3ac9eb2c),
	.w2(32'hbb61a123),
	.w3(32'h3a1f2dcd),
	.w4(32'hbb29a627),
	.w5(32'hbbf2c050),
	.w6(32'hbbf46702),
	.w7(32'hbb35f937),
	.w8(32'hba25dea3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d755e3),
	.w1(32'hbb625d0e),
	.w2(32'hbbeea5bc),
	.w3(32'hbb8f3b6b),
	.w4(32'hba08f3a9),
	.w5(32'hb9155301),
	.w6(32'hbb3a1f1f),
	.w7(32'h3b506240),
	.w8(32'h3bbd2cb3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba949f9b),
	.w1(32'hbb81b1ee),
	.w2(32'hbc61a311),
	.w3(32'hbb5d5692),
	.w4(32'hbbe82426),
	.w5(32'hbc493328),
	.w6(32'h3b750ae0),
	.w7(32'h39746b5e),
	.w8(32'hbc34efce),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9454d7),
	.w1(32'hbb09b7b6),
	.w2(32'hbca28551),
	.w3(32'hbb281289),
	.w4(32'hbc02a4ba),
	.w5(32'hbc28e290),
	.w6(32'hbb76b8a3),
	.w7(32'hbc5fefd5),
	.w8(32'hbb670c6c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5dbb55),
	.w1(32'h3ae51347),
	.w2(32'hbc05ee91),
	.w3(32'hbb2b392f),
	.w4(32'hbb24f0d1),
	.w5(32'hbb9fa806),
	.w6(32'hbbcafb99),
	.w7(32'hbb058ba9),
	.w8(32'hbb8490cb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb90d77),
	.w1(32'hbb3dccc4),
	.w2(32'hbb9a8253),
	.w3(32'hbaf7c932),
	.w4(32'hbb137308),
	.w5(32'h3be7bc29),
	.w6(32'hba90bbde),
	.w7(32'hbb8d1500),
	.w8(32'h3963d506),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed0e14),
	.w1(32'hbb22432d),
	.w2(32'h3c038a88),
	.w3(32'hba50c54b),
	.w4(32'h3b94d4e5),
	.w5(32'h3c344276),
	.w6(32'hbb8dfe02),
	.w7(32'h3ca37978),
	.w8(32'h3c70c432),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5aa4),
	.w1(32'h39b23f37),
	.w2(32'hbb046f4e),
	.w3(32'h3b2459d5),
	.w4(32'h3ac03897),
	.w5(32'h3b5c9c5d),
	.w6(32'hb911a0b1),
	.w7(32'h3a6a6242),
	.w8(32'h3c08f74a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d0a3c),
	.w1(32'h3b71f2e2),
	.w2(32'hbbeba553),
	.w3(32'h3c13f975),
	.w4(32'h3bfba547),
	.w5(32'hbaf63e41),
	.w6(32'h3c182d9c),
	.w7(32'h3bb81d54),
	.w8(32'hbaad0a12),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2468bf),
	.w1(32'hbb6ba74b),
	.w2(32'hbb4ba7c5),
	.w3(32'hbbb61bac),
	.w4(32'hbaf44eab),
	.w5(32'hba055326),
	.w6(32'hbbb44f91),
	.w7(32'h3b9d17cf),
	.w8(32'h3a385cad),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb6fb6),
	.w1(32'h3b55c0d8),
	.w2(32'h3b2d4db1),
	.w3(32'hbb5e950c),
	.w4(32'hba6452da),
	.w5(32'h3b45d4a2),
	.w6(32'hbb941407),
	.w7(32'h3c7cb616),
	.w8(32'h3c983815),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2092ff),
	.w1(32'hba30b209),
	.w2(32'hbb096e5a),
	.w3(32'hba8c844f),
	.w4(32'hba96feba),
	.w5(32'hba7eefa3),
	.w6(32'hbb8b8e8b),
	.w7(32'hbadad3be),
	.w8(32'hba94c9b3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2290b2),
	.w1(32'h3b31afcc),
	.w2(32'hbbff84d7),
	.w3(32'hb9eb8623),
	.w4(32'h3bbb217d),
	.w5(32'hbb988918),
	.w6(32'h3a893cf9),
	.w7(32'h3b3e6d72),
	.w8(32'hbbab3d08),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63a7dc),
	.w1(32'h3a6c670d),
	.w2(32'h3a343b24),
	.w3(32'hba1ab3e5),
	.w4(32'hba021976),
	.w5(32'hbb0e4cac),
	.w6(32'hbbe385ee),
	.w7(32'h391723d2),
	.w8(32'hbb0b9055),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc115d23),
	.w1(32'hbb874946),
	.w2(32'hbbc3328e),
	.w3(32'hbb987be3),
	.w4(32'hbb7fa93f),
	.w5(32'h3a862a56),
	.w6(32'hbb08fa4a),
	.w7(32'h3b03b9dd),
	.w8(32'h3b13e935),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b170290),
	.w1(32'hbbb036f7),
	.w2(32'hbc1101d2),
	.w3(32'hba07b315),
	.w4(32'hbc009296),
	.w5(32'hbc30cd67),
	.w6(32'h3b636fbb),
	.w7(32'h3bedcc81),
	.w8(32'h3a9864c5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6323d2),
	.w1(32'h38906d43),
	.w2(32'hbb0af9b2),
	.w3(32'hba234607),
	.w4(32'h3bb71082),
	.w5(32'h3b9f6411),
	.w6(32'hb8f29137),
	.w7(32'h3bb67fac),
	.w8(32'h3bd7dadd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d2e8d),
	.w1(32'h3b654de0),
	.w2(32'hbae2383a),
	.w3(32'hbb03203d),
	.w4(32'h3ba6b875),
	.w5(32'hba86d7aa),
	.w6(32'hbb964118),
	.w7(32'h3b1c6b15),
	.w8(32'hbb8703e7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47d4ad),
	.w1(32'hbaa11695),
	.w2(32'hbbc2d563),
	.w3(32'hbb029a22),
	.w4(32'h3b7f6611),
	.w5(32'h3be9cf1f),
	.w6(32'hbad72f23),
	.w7(32'hba7040bf),
	.w8(32'h3c3c9cee),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3ed7f),
	.w1(32'hbb476feb),
	.w2(32'hbb67f519),
	.w3(32'h3bb65c1c),
	.w4(32'h3b37e228),
	.w5(32'h3c137897),
	.w6(32'h3ba41639),
	.w7(32'hbb0f1aee),
	.w8(32'hbac450e8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9581f06),
	.w1(32'hbb182c26),
	.w2(32'hbbc325ca),
	.w3(32'hb91fe27f),
	.w4(32'h3bf26e72),
	.w5(32'h3ba8330a),
	.w6(32'hbb8512a5),
	.w7(32'h3bf097ed),
	.w8(32'h3c073e70),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbb6bc),
	.w1(32'hbb6752f6),
	.w2(32'hbc38f3da),
	.w3(32'h3ab7df05),
	.w4(32'h3bba6034),
	.w5(32'hbb143d60),
	.w6(32'h3a7f21d5),
	.w7(32'hbaf1a8c4),
	.w8(32'hbc1893f6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec387),
	.w1(32'hbc033873),
	.w2(32'h3bcd0b77),
	.w3(32'hbb2970e6),
	.w4(32'h3c410721),
	.w5(32'h3c115a70),
	.w6(32'hbc1107b0),
	.w7(32'h3ba83d68),
	.w8(32'hb98c1636),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c200205),
	.w1(32'h3b8e70a5),
	.w2(32'hbba38355),
	.w3(32'hbb561fea),
	.w4(32'hbb2173b5),
	.w5(32'h3be4ba3f),
	.w6(32'hbb9f2119),
	.w7(32'hbb5603e1),
	.w8(32'h3a84a4f2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4213),
	.w1(32'hbc07d006),
	.w2(32'hbc981985),
	.w3(32'hbc228d9c),
	.w4(32'hbc13d627),
	.w5(32'hbc662a67),
	.w6(32'hbc557a58),
	.w7(32'hbc4a95c4),
	.w8(32'hbc1aac2c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f2187),
	.w1(32'hbb7d43c8),
	.w2(32'hbc66d759),
	.w3(32'hbb5f8eeb),
	.w4(32'hbb28a05a),
	.w5(32'hbc5e26db),
	.w6(32'hbba0d6f5),
	.w7(32'h3b00357d),
	.w8(32'hbbe899b7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b9e5d),
	.w1(32'hbc5440e4),
	.w2(32'hbb44ea1f),
	.w3(32'hbc4f9774),
	.w4(32'hbb79bea4),
	.w5(32'h3c338e88),
	.w6(32'hbc6a3661),
	.w7(32'hba97d9e9),
	.w8(32'h3bf07f6b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56044),
	.w1(32'h3c1326af),
	.w2(32'hba4b3407),
	.w3(32'h3bcf78c7),
	.w4(32'h3b09c713),
	.w5(32'hba8c9df3),
	.w6(32'hbb3b035c),
	.w7(32'hbae83a65),
	.w8(32'h399af3fb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5b8eb),
	.w1(32'h39709319),
	.w2(32'hbba40873),
	.w3(32'h3b138f41),
	.w4(32'h39482380),
	.w5(32'h3be04096),
	.w6(32'h39546dc8),
	.w7(32'hbaae4d0c),
	.w8(32'hbacd323c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5ebbf),
	.w1(32'hbc360236),
	.w2(32'hbbbd8af3),
	.w3(32'hbc129a0d),
	.w4(32'hbb970ff1),
	.w5(32'hbbdeb18a),
	.w6(32'hbb980f8d),
	.w7(32'hbb80cc90),
	.w8(32'h3a440d90),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c36c2),
	.w1(32'hbba61a27),
	.w2(32'hbbb00637),
	.w3(32'hbb92da4c),
	.w4(32'h3bbdc1fc),
	.w5(32'hbc002cda),
	.w6(32'hbab393f0),
	.w7(32'h3bc52e5e),
	.w8(32'h3b40de06),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1446f6),
	.w1(32'hbaa4b970),
	.w2(32'h3bb6c77e),
	.w3(32'h3b8d5562),
	.w4(32'h3b8539ba),
	.w5(32'h3c06dae6),
	.w6(32'h3b38154a),
	.w7(32'h3c10474d),
	.w8(32'h3be09561),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c73ae4),
	.w1(32'hbaf9e137),
	.w2(32'hbb5884f8),
	.w3(32'hbab2ca1a),
	.w4(32'h3bbce523),
	.w5(32'h3bae167a),
	.w6(32'hbb2afd2b),
	.w7(32'h3bb68961),
	.w8(32'h3b668a2c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfee56),
	.w1(32'hbbf30a4e),
	.w2(32'hbc485f9d),
	.w3(32'hbb985e4e),
	.w4(32'hb9ed4ef9),
	.w5(32'hb9d1e335),
	.w6(32'hbbc7b2ed),
	.w7(32'h3bf06911),
	.w8(32'h3b5c9e9d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcc405),
	.w1(32'hbb8a1ce7),
	.w2(32'hbac9c2c8),
	.w3(32'hb8d8b1ab),
	.w4(32'hbb6726f2),
	.w5(32'h3b6e66ed),
	.w6(32'hbbdb0fb8),
	.w7(32'hbb1f8552),
	.w8(32'h3914d1b0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb431e96),
	.w1(32'hbb02509a),
	.w2(32'hbc279046),
	.w3(32'hbaac28e3),
	.w4(32'hbbd8ff2d),
	.w5(32'hbbc051c4),
	.w6(32'hbbdf0db2),
	.w7(32'hbbece2ea),
	.w8(32'hbbe61f92),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c634),
	.w1(32'hbbee1105),
	.w2(32'hbb433edc),
	.w3(32'hbb423545),
	.w4(32'hbb173e18),
	.w5(32'h3b0a13d6),
	.w6(32'hbb995756),
	.w7(32'hba0532fd),
	.w8(32'hbac38181),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4dfb),
	.w1(32'h39fb1efc),
	.w2(32'h3a239646),
	.w3(32'h3a4aeefd),
	.w4(32'h3b0309fd),
	.w5(32'hbbbc4ed3),
	.w6(32'hbbe59f13),
	.w7(32'hbb57f7d5),
	.w8(32'h3a0db405),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d66c4),
	.w1(32'h3b1ad2c6),
	.w2(32'hbb83ab79),
	.w3(32'hbb2f005f),
	.w4(32'h3b0d7aca),
	.w5(32'h3b9a38b5),
	.w6(32'hbbce4a1d),
	.w7(32'h3ba6e12b),
	.w8(32'h3be356e2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409542),
	.w1(32'hbabb52e7),
	.w2(32'h3c0eb3b9),
	.w3(32'h3a812862),
	.w4(32'h3bab399f),
	.w5(32'h3baa08fa),
	.w6(32'h39eb08d6),
	.w7(32'h3c1e3699),
	.w8(32'h3c0e031e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ceafd),
	.w1(32'hbbd22e76),
	.w2(32'hbbe95015),
	.w3(32'hbb18f397),
	.w4(32'h3bccda7b),
	.w5(32'h3bfa4613),
	.w6(32'hbb8b8422),
	.w7(32'h3c3006e4),
	.w8(32'h3c1361ef),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f681d),
	.w1(32'hbb5dd803),
	.w2(32'h3a05574e),
	.w3(32'h3b57f8d2),
	.w4(32'hbb0d8be5),
	.w5(32'h3c1cb43e),
	.w6(32'h3b44775c),
	.w7(32'hba644074),
	.w8(32'h3b9ae09d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c711e),
	.w1(32'h3aa34377),
	.w2(32'hb910086f),
	.w3(32'h3ac5bc09),
	.w4(32'h3b7fc2f6),
	.w5(32'h3be12cb9),
	.w6(32'hbbf465e2),
	.w7(32'h3a07909c),
	.w8(32'h3b26b4dd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10ee6d),
	.w1(32'hbb13afbf),
	.w2(32'hbc53bc92),
	.w3(32'hbbc975b7),
	.w4(32'hba4a98ab),
	.w5(32'h3a7a3b33),
	.w6(32'hbbcca28a),
	.w7(32'h3b492ea0),
	.w8(32'h3a7250ee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80f25c),
	.w1(32'hbbc07736),
	.w2(32'h3b49bc68),
	.w3(32'hba6ccb08),
	.w4(32'h3ae494ac),
	.w5(32'h3aeec46b),
	.w6(32'hbbdfd3f0),
	.w7(32'h3be4af6f),
	.w8(32'h3b436317),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c39b1),
	.w1(32'hbb72d041),
	.w2(32'hbc093f58),
	.w3(32'hbb5f41e7),
	.w4(32'h3b6dbcbe),
	.w5(32'hb9d9da97),
	.w6(32'hb7bff016),
	.w7(32'h3bc9b040),
	.w8(32'h3b25b66e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1a23),
	.w1(32'hbbc0096e),
	.w2(32'hbac8ee91),
	.w3(32'hbbc0031c),
	.w4(32'hba44e80d),
	.w5(32'h3c0f4bf2),
	.w6(32'hba267c89),
	.w7(32'h39c842d2),
	.w8(32'hba82877f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule