module layer_8_featuremap_72(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a680ef8),
	.w1(32'hbb787748),
	.w2(32'h3b389e01),
	.w3(32'hbaf167ca),
	.w4(32'h3b2c0445),
	.w5(32'h3a962e2e),
	.w6(32'h3aef5e33),
	.w7(32'h3ad04add),
	.w8(32'h3a320b12),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39449654),
	.w1(32'hba14307c),
	.w2(32'h3acfe000),
	.w3(32'hba67693b),
	.w4(32'h396cdf79),
	.w5(32'h39eea3e4),
	.w6(32'h3a84b3e1),
	.w7(32'h3b2eba99),
	.w8(32'h39570347),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17dd55),
	.w1(32'hba02b829),
	.w2(32'hb98d6022),
	.w3(32'hbabd4973),
	.w4(32'hb9cfc94e),
	.w5(32'hb938e6f1),
	.w6(32'hb93e3a84),
	.w7(32'h3a4dba69),
	.w8(32'hbc5ad298),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56f6f1),
	.w1(32'hbb472ed7),
	.w2(32'hbc58e61d),
	.w3(32'hbae2abc0),
	.w4(32'hbbb81218),
	.w5(32'hbc5fb35b),
	.w6(32'hbb836f0e),
	.w7(32'hbc056166),
	.w8(32'h3b37284c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a0419),
	.w1(32'hbc068411),
	.w2(32'hbab49448),
	.w3(32'hb9d065ac),
	.w4(32'hbb221173),
	.w5(32'hba01772e),
	.w6(32'hb6b473b3),
	.w7(32'hbb3253ec),
	.w8(32'h3bd8f1c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d7ebe),
	.w1(32'hbaa86a15),
	.w2(32'h3c22a08f),
	.w3(32'hbbbf377d),
	.w4(32'hbb07bb13),
	.w5(32'h3b8d19e7),
	.w6(32'h3c1ef2ea),
	.w7(32'h3c15b38a),
	.w8(32'h3b657cc0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c3c23),
	.w1(32'hbb1bc44f),
	.w2(32'h3b943147),
	.w3(32'h39a0b7c4),
	.w4(32'h39a5cf72),
	.w5(32'h3b0fa0dc),
	.w6(32'h3b816a14),
	.w7(32'h3b8ba83c),
	.w8(32'h3ad78e9d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1b39f),
	.w1(32'hbc42f79f),
	.w2(32'hbb5f6252),
	.w3(32'hba1ac508),
	.w4(32'hbb42dd53),
	.w5(32'hbaa46c05),
	.w6(32'hbaf585d5),
	.w7(32'hbb92495d),
	.w8(32'h3b86c510),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afe9aa),
	.w1(32'hba1a7faa),
	.w2(32'h3bb0cafd),
	.w3(32'hba0eda7b),
	.w4(32'hb8db286a),
	.w5(32'h3b4efd91),
	.w6(32'h3b6d1a94),
	.w7(32'h3b9c5cb9),
	.w8(32'h3c9a9691),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c942a9b),
	.w1(32'h3d1e66c6),
	.w2(32'h3bf04631),
	.w3(32'hbb9ef081),
	.w4(32'hba634400),
	.w5(32'h3cbcbab3),
	.w6(32'hbb8bbb96),
	.w7(32'hbc0e01be),
	.w8(32'hbaf32983),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d6b08),
	.w1(32'hba9b1d28),
	.w2(32'hbb726cbe),
	.w3(32'hbbd65248),
	.w4(32'hbb397d15),
	.w5(32'hbb0b89aa),
	.w6(32'hbb3d157d),
	.w7(32'hbc1010e3),
	.w8(32'h3b0a9293),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a5530),
	.w1(32'hbb5b2cf0),
	.w2(32'h3a47d345),
	.w3(32'hba000cf7),
	.w4(32'hb9f21b82),
	.w5(32'h3a94d017),
	.w6(32'h3b47117b),
	.w7(32'h3b6bcec1),
	.w8(32'hb995aae1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92137f7),
	.w1(32'hbbb797f7),
	.w2(32'hba988264),
	.w3(32'hbab7872e),
	.w4(32'hbb2f3177),
	.w5(32'hb9fe39c2),
	.w6(32'h3ac50258),
	.w7(32'hb9a485af),
	.w8(32'h3c1359d1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a808691),
	.w1(32'hbab00216),
	.w2(32'h3c3b93ad),
	.w3(32'hbb903ffd),
	.w4(32'hba650b11),
	.w5(32'h3bc389dd),
	.w6(32'h3c463e72),
	.w7(32'h3c402a1c),
	.w8(32'h3b977bdb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add0c12),
	.w1(32'hbb655b53),
	.w2(32'h3c2648e1),
	.w3(32'hbb056b5c),
	.w4(32'hbb568436),
	.w5(32'h3ba4e467),
	.w6(32'h3be6edd8),
	.w7(32'h3bea7811),
	.w8(32'h3a5b704d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ccdac),
	.w1(32'h3b2870a2),
	.w2(32'hba4ac098),
	.w3(32'hba9ffc3a),
	.w4(32'h3990248f),
	.w5(32'h3b399898),
	.w6(32'hba16b01d),
	.w7(32'hbb13394f),
	.w8(32'hbc0dea19),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0ff00),
	.w1(32'h3b0d1822),
	.w2(32'hbd0c2226),
	.w3(32'h3b7e1ff7),
	.w4(32'h3cd256b1),
	.w5(32'hbab65b9b),
	.w6(32'hbbab9831),
	.w7(32'hbc420ec8),
	.w8(32'hbad0976b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5540a8),
	.w1(32'hbb9814ed),
	.w2(32'hbbb56143),
	.w3(32'hbad19c7e),
	.w4(32'hba74d38d),
	.w5(32'hbb3daa04),
	.w6(32'hb8805989),
	.w7(32'hbb3a59d0),
	.w8(32'hbb3ea176),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ba75),
	.w1(32'hbc94154f),
	.w2(32'hbc159683),
	.w3(32'hbb5ecfdc),
	.w4(32'hbbbfdd07),
	.w5(32'hbbca01b3),
	.w6(32'hbb8ab608),
	.w7(32'hbc359474),
	.w8(32'h3c07d390),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21bbfe),
	.w1(32'h3bc46870),
	.w2(32'hbcde6e03),
	.w3(32'hbbf3949e),
	.w4(32'hbc95908c),
	.w5(32'hbcaaec07),
	.w6(32'hbbba3e6b),
	.w7(32'hbc97c410),
	.w8(32'h3b3f6989),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004b42),
	.w1(32'hbbbd707d),
	.w2(32'hbb9e6793),
	.w3(32'h3c12fd4f),
	.w4(32'h3afc82eb),
	.w5(32'h397ed891),
	.w6(32'hbb98d2ad),
	.w7(32'hbb86d019),
	.w8(32'h3b6b5c0e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7702f8),
	.w1(32'hbc244e9a),
	.w2(32'hba2b0c29),
	.w3(32'hb9ec2557),
	.w4(32'hbb0d1429),
	.w5(32'h3aa4c870),
	.w6(32'h39bb9670),
	.w7(32'hba844076),
	.w8(32'h3c063197),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04b77a),
	.w1(32'h3b0ea7b2),
	.w2(32'hbbc0c571),
	.w3(32'h3cc313b7),
	.w4(32'h3c7ba8e0),
	.w5(32'h3c0aff74),
	.w6(32'h3b3d6052),
	.w7(32'h3bbeda8b),
	.w8(32'h3b8d52e3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65b395),
	.w1(32'hbbbafa27),
	.w2(32'h3a1e1baa),
	.w3(32'h39e27a0f),
	.w4(32'h3b94d79f),
	.w5(32'h3a44c69a),
	.w6(32'h3b2d9434),
	.w7(32'hbb191461),
	.w8(32'hb9bac60a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f35b5),
	.w1(32'h3b4f0305),
	.w2(32'hbb8ca5a5),
	.w3(32'h3bc2d8bd),
	.w4(32'h3bf5ce6d),
	.w5(32'h3ba6517a),
	.w6(32'h3aa7b2b9),
	.w7(32'hbafe06d0),
	.w8(32'h3bf6eb61),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2f6cb),
	.w1(32'h3ad296fc),
	.w2(32'hbbc217f4),
	.w3(32'h3cb3590f),
	.w4(32'h3c615949),
	.w5(32'h3bf128dd),
	.w6(32'h3b18c9c1),
	.w7(32'h3ba3906c),
	.w8(32'h3bd2edcc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccbcf0),
	.w1(32'h3a90db72),
	.w2(32'hbbb09048),
	.w3(32'h3c9856ee),
	.w4(32'h3c3ec07f),
	.w5(32'h3bc503c0),
	.w6(32'h3b00a3c9),
	.w7(32'h3b8cad83),
	.w8(32'h3b1eee3b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9319aa0),
	.w1(32'hbbd5592f),
	.w2(32'hbb10009a),
	.w3(32'h3c66ae7f),
	.w4(32'h3a9b7afb),
	.w5(32'h3a3b4f4c),
	.w6(32'hbb89ef5c),
	.w7(32'hba9b92c0),
	.w8(32'h3c23acd8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc403a84),
	.w1(32'h3d058de5),
	.w2(32'hbb92bc37),
	.w3(32'h3ad5148d),
	.w4(32'h3c582a43),
	.w5(32'h3940ce9c),
	.w6(32'hbb045c72),
	.w7(32'hbcb47a39),
	.w8(32'hba03f0a2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ffd55),
	.w1(32'hba99ef47),
	.w2(32'hb9215ef5),
	.w3(32'hbb01939c),
	.w4(32'hba87d8a9),
	.w5(32'hb886fbf7),
	.w6(32'h3a121420),
	.w7(32'h39cd2e7d),
	.w8(32'h3c1c265a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca001b0),
	.w1(32'hbc928cd3),
	.w2(32'hbc4e6b43),
	.w3(32'h3c2cc8a2),
	.w4(32'h3c2db898),
	.w5(32'h3b45abb1),
	.w6(32'h3bb25fa0),
	.w7(32'h3bbe5f2c),
	.w8(32'h3bc0b4cc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f4f17),
	.w1(32'hbc257fe9),
	.w2(32'hbc41a883),
	.w3(32'h3cc32ee0),
	.w4(32'h3c2ff82b),
	.w5(32'h3b9e4faa),
	.w6(32'hbbe56f91),
	.w7(32'hbbf35f1a),
	.w8(32'hb9c5ecf9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf29a30),
	.w1(32'hbb2b6b37),
	.w2(32'h3c87478e),
	.w3(32'h3c488dff),
	.w4(32'h3c00b71b),
	.w5(32'h3beff9e9),
	.w6(32'h3b39da00),
	.w7(32'h3a168f3a),
	.w8(32'h3bb4b306),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f6aa1),
	.w1(32'h3a28ce2d),
	.w2(32'hbc8fe997),
	.w3(32'h3c10eb65),
	.w4(32'hbc1ec8fc),
	.w5(32'hbb842020),
	.w6(32'h3cd03fed),
	.w7(32'h3ca1f2ba),
	.w8(32'h3bffcf13),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c8b49),
	.w1(32'hba96b06e),
	.w2(32'h3c251e13),
	.w3(32'hbb810e6b),
	.w4(32'hba696567),
	.w5(32'h3ba87148),
	.w6(32'h3c2ddb23),
	.w7(32'h3c288417),
	.w8(32'h3b28f2f4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d5c0a),
	.w1(32'hbc11647e),
	.w2(32'hba96c0bc),
	.w3(32'h3a16bd2a),
	.w4(32'hb78e12ef),
	.w5(32'hbb05fb87),
	.w6(32'h3ad1ce94),
	.w7(32'hb9f13190),
	.w8(32'h3a9f4975),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b521853),
	.w1(32'hbc50f94a),
	.w2(32'hbc2f8fc1),
	.w3(32'h3c0dca81),
	.w4(32'h3c0b0f6c),
	.w5(32'hbc0a01cd),
	.w6(32'hbbb63990),
	.w7(32'hbc0e6a49),
	.w8(32'hba185ea6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840ca0),
	.w1(32'hba6297f2),
	.w2(32'hba98f9b2),
	.w3(32'hbb2f9338),
	.w4(32'hba37c582),
	.w5(32'h398672de),
	.w6(32'hba704804),
	.w7(32'hba1a9390),
	.w8(32'h3c224ed6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc89cd8),
	.w1(32'hbc150b1e),
	.w2(32'h3cc9e252),
	.w3(32'hb8ad8a30),
	.w4(32'hbb006718),
	.w5(32'h3c64fb47),
	.w6(32'h3c80f46f),
	.w7(32'h3c8d26ff),
	.w8(32'hbabd7c07),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4c85),
	.w1(32'hbc0f5d91),
	.w2(32'hbbba990e),
	.w3(32'h3bdaac70),
	.w4(32'h3ae29ea4),
	.w5(32'hbabb3003),
	.w6(32'hbbbe99eb),
	.w7(32'hbb1aa462),
	.w8(32'h3b3088d3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d2541),
	.w1(32'h3a8d4527),
	.w2(32'hbb0fc7fe),
	.w3(32'h3c164897),
	.w4(32'h3bb907af),
	.w5(32'h3b3d5f96),
	.w6(32'h3a86bb50),
	.w7(32'h3aeb4095),
	.w8(32'h3a6b2b2c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7709884),
	.w1(32'hb88854ea),
	.w2(32'h37a4ab31),
	.w3(32'h39e8c271),
	.w4(32'h398dcb6c),
	.w5(32'hb9e45013),
	.w6(32'hb92f90f7),
	.w7(32'hba7c2a88),
	.w8(32'hbb27b15d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860a69),
	.w1(32'h38afec29),
	.w2(32'hbb086dae),
	.w3(32'hb912a372),
	.w4(32'h39b615c7),
	.w5(32'hbae2d608),
	.w6(32'h3b0d00ce),
	.w7(32'h38b1d6c1),
	.w8(32'h39b2dd69),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b138c),
	.w1(32'hb97a1849),
	.w2(32'hba02af0f),
	.w3(32'hb5b62d94),
	.w4(32'h38c72149),
	.w5(32'h37da3cbf),
	.w6(32'hba6d9613),
	.w7(32'hbaa83808),
	.w8(32'h3a7abb91),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25688c),
	.w1(32'h3a58685e),
	.w2(32'hb955d701),
	.w3(32'h39997490),
	.w4(32'h3a2015a7),
	.w5(32'h398b5cb9),
	.w6(32'h39724440),
	.w7(32'hba2a4cf9),
	.w8(32'hba2b665e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04d4bf),
	.w1(32'hb8910471),
	.w2(32'h37912f6f),
	.w3(32'h393a1b69),
	.w4(32'h3ada7b8e),
	.w5(32'h3a896764),
	.w6(32'hba002773),
	.w7(32'hba754623),
	.w8(32'hb9e523a4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ff89),
	.w1(32'hbb78f813),
	.w2(32'h3b4f2b1f),
	.w3(32'hb9123771),
	.w4(32'hbbe1d2fa),
	.w5(32'h3a51fbb5),
	.w6(32'h3b90a3b1),
	.w7(32'h3bc807f6),
	.w8(32'hbabd723c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919908f),
	.w1(32'hbaa1d679),
	.w2(32'hbb1cb79f),
	.w3(32'h3a4cf1e8),
	.w4(32'h3a055b75),
	.w5(32'hbb39004a),
	.w6(32'hbb71499a),
	.w7(32'hbafd1726),
	.w8(32'hbad9bb4b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34059a),
	.w1(32'hb97f5bc5),
	.w2(32'h3a4eaaf3),
	.w3(32'hbb26cd24),
	.w4(32'hba92e7d8),
	.w5(32'h3a24e167),
	.w6(32'hba547c2f),
	.w7(32'hb965f2a3),
	.w8(32'h3a295a7c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe4be0),
	.w1(32'h3a0bc4f1),
	.w2(32'hb9666c06),
	.w3(32'h3a3f8be2),
	.w4(32'h3a8fb722),
	.w5(32'h39480418),
	.w6(32'h38b3eaab),
	.w7(32'hba2954c5),
	.w8(32'h39b4b597),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f584bd),
	.w1(32'hb8802539),
	.w2(32'hb838f456),
	.w3(32'h3a1d639d),
	.w4(32'h39d3b67f),
	.w5(32'h39940eba),
	.w6(32'hb991c3b2),
	.w7(32'hba219b7f),
	.w8(32'h3a9ab538),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9fce4),
	.w1(32'hb996b969),
	.w2(32'hba1c9bee),
	.w3(32'h3a3e93dc),
	.w4(32'h39f2e590),
	.w5(32'h3a713bc4),
	.w6(32'hba8264f4),
	.w7(32'hbaf1c5b1),
	.w8(32'h3a9cb76b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a0053),
	.w1(32'hbb8f1e39),
	.w2(32'hbbbd2b1b),
	.w3(32'h3a846184),
	.w4(32'hbb18b457),
	.w5(32'hbb63da2c),
	.w6(32'hbb09869b),
	.w7(32'h3a59dd03),
	.w8(32'h3ad0d8d6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af28fa7),
	.w1(32'h3a4a6906),
	.w2(32'h3aeade09),
	.w3(32'h3ab60f04),
	.w4(32'h3aea67c0),
	.w5(32'h3b346713),
	.w6(32'h3aa6edad),
	.w7(32'h39fe6703),
	.w8(32'hba43e60f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab74172),
	.w1(32'hbba57107),
	.w2(32'hbb849147),
	.w3(32'hbaab7615),
	.w4(32'hbbc1ef9e),
	.w5(32'hbb0fca7b),
	.w6(32'h3ad5f948),
	.w7(32'h3ac6c676),
	.w8(32'hbadfe094),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e9a32),
	.w1(32'hb9be7dd6),
	.w2(32'hbbbc9952),
	.w3(32'h3b976c12),
	.w4(32'h3b018516),
	.w5(32'hbb131555),
	.w6(32'hbbb88265),
	.w7(32'hbbd7d3c5),
	.w8(32'hbaf9bf9c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1300b),
	.w1(32'hba44dae1),
	.w2(32'h3aabb5a0),
	.w3(32'h39da4c05),
	.w4(32'h3b0fe621),
	.w5(32'hbaa361b1),
	.w6(32'h3aab7913),
	.w7(32'h3ac79c3b),
	.w8(32'hb88b276b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b611d),
	.w1(32'h3a29086a),
	.w2(32'hbc08e0bc),
	.w3(32'h3a1e0fc0),
	.w4(32'hbae19dd3),
	.w5(32'hbaf8dbde),
	.w6(32'hbbd58039),
	.w7(32'h3a20c38e),
	.w8(32'hba3a1d5d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa81a3),
	.w1(32'hb988793d),
	.w2(32'h3a63919e),
	.w3(32'hbab2e85f),
	.w4(32'hba326e1f),
	.w5(32'h3927fe58),
	.w6(32'hba5a2959),
	.w7(32'h38df7740),
	.w8(32'hbb16ae0d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3291fd),
	.w1(32'hbb2380bb),
	.w2(32'h3a094e76),
	.w3(32'hbb13ea1a),
	.w4(32'hbb9aa24e),
	.w5(32'hbaa26a68),
	.w6(32'hb9e097e0),
	.w7(32'h3885f39c),
	.w8(32'hbb77ffbe),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f2ca1),
	.w1(32'hbb121b7a),
	.w2(32'h3ab4569c),
	.w3(32'h3b15885d),
	.w4(32'h3b4fff80),
	.w5(32'hbafaa62e),
	.w6(32'h39877925),
	.w7(32'h3b024faf),
	.w8(32'hba26b2c7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05305f),
	.w1(32'hba2df1d0),
	.w2(32'hba910168),
	.w3(32'h3aa70417),
	.w4(32'h3b09fd12),
	.w5(32'hba007ef7),
	.w6(32'hba70c179),
	.w7(32'hba7d1d06),
	.w8(32'h39f1441a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86f646),
	.w1(32'hba337163),
	.w2(32'hbaa81dbb),
	.w3(32'hb7b59209),
	.w4(32'h39ebe85a),
	.w5(32'hb8f20315),
	.w6(32'hbacddf0d),
	.w7(32'hbb2b8b91),
	.w8(32'h3af3a072),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89354a),
	.w1(32'h3baeb1d2),
	.w2(32'hbb42664d),
	.w3(32'h3ba4fb4b),
	.w4(32'hb8cb2af3),
	.w5(32'hbae7f531),
	.w6(32'hbb971c3c),
	.w7(32'hbad653a0),
	.w8(32'hb69b3c05),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997c985),
	.w1(32'hba225f57),
	.w2(32'hba83d5e5),
	.w3(32'hb989fb3a),
	.w4(32'hb6bd4b1c),
	.w5(32'hba17663d),
	.w6(32'hba8e25e2),
	.w7(32'hbab3cc26),
	.w8(32'h39759c14),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3728f16c),
	.w1(32'h37c197a4),
	.w2(32'h364beafb),
	.w3(32'hb8896b50),
	.w4(32'hb81f6c71),
	.w5(32'h396458a7),
	.w6(32'hb8c0b366),
	.w7(32'hb9a537cd),
	.w8(32'h39e407f0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bc838),
	.w1(32'hb98438f7),
	.w2(32'hb99362ba),
	.w3(32'h390077be),
	.w4(32'hb9506fde),
	.w5(32'h37cc8fe2),
	.w6(32'hb9caf303),
	.w7(32'hba364d28),
	.w8(32'hbaeade3e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0b22d),
	.w1(32'hb9c79bbc),
	.w2(32'h39c07ce2),
	.w3(32'h3b503b23),
	.w4(32'h3acbe6d6),
	.w5(32'hb9360053),
	.w6(32'hb8efd2ff),
	.w7(32'h384795a5),
	.w8(32'h3a2ecbf1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a099702),
	.w1(32'h3a28465d),
	.w2(32'hb9070db3),
	.w3(32'h39c2498b),
	.w4(32'h3a3ac52c),
	.w5(32'hb7e03663),
	.w6(32'h391d5b8e),
	.w7(32'hb9e315a0),
	.w8(32'h38cfd944),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f81450),
	.w1(32'hb943b50d),
	.w2(32'h3a26b6b1),
	.w3(32'h3989a7d8),
	.w4(32'h38e88a20),
	.w5(32'h377d6e97),
	.w6(32'hb9c0b91b),
	.w7(32'h3a31d5d2),
	.w8(32'h3a60a90d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a61e5e),
	.w1(32'h39053ff2),
	.w2(32'hb9d6de3c),
	.w3(32'hb9891a2c),
	.w4(32'h392b123d),
	.w5(32'hb90ce881),
	.w6(32'hb9e8dfb9),
	.w7(32'hba9794e8),
	.w8(32'h3a28dcad),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e151b2),
	.w1(32'h3a2d6ea9),
	.w2(32'hb94f32c2),
	.w3(32'h3a34f246),
	.w4(32'h3a796f2f),
	.w5(32'h37ed6ae6),
	.w6(32'hb8f62463),
	.w7(32'hba24b40b),
	.w8(32'h3ad0c522),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fa305),
	.w1(32'h3a03b400),
	.w2(32'hb8e0a653),
	.w3(32'hb8faad0e),
	.w4(32'hb7e05140),
	.w5(32'h38ffdb40),
	.w6(32'h39661b5c),
	.w7(32'hba71bec2),
	.w8(32'hbb2c0a95),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d92de),
	.w1(32'hb988a898),
	.w2(32'hbbbcdf9d),
	.w3(32'h39e48ae3),
	.w4(32'h3b0831f2),
	.w5(32'hbb865b06),
	.w6(32'hbbaddc20),
	.w7(32'hbb2e260b),
	.w8(32'h39d2e4a7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1220df),
	.w1(32'h39a1e1a9),
	.w2(32'hba6c7f14),
	.w3(32'h3ac4ac47),
	.w4(32'h3ac8a7d6),
	.w5(32'h38a0b3e5),
	.w6(32'hba81e038),
	.w7(32'hba731b74),
	.w8(32'h39ce3639),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36efe485),
	.w1(32'hb8d8d8e1),
	.w2(32'hb9cb8139),
	.w3(32'hb97964c2),
	.w4(32'h3718189a),
	.w5(32'hb8945055),
	.w6(32'hba12a68a),
	.w7(32'hba8c389b),
	.w8(32'h3a6ec6bb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f375ec),
	.w1(32'h39bc2f44),
	.w2(32'hb9d981dc),
	.w3(32'h3a13793e),
	.w4(32'h3a2f0b6d),
	.w5(32'hb8cf9771),
	.w6(32'hba08982a),
	.w7(32'hba8cb0bb),
	.w8(32'hb902618d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a0b6b),
	.w1(32'h389568f2),
	.w2(32'h3a9804b0),
	.w3(32'h38f8e691),
	.w4(32'hb95ad85a),
	.w5(32'hb9db319e),
	.w6(32'hba1d6881),
	.w7(32'h3a35f370),
	.w8(32'h39583b3d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cdbfd),
	.w1(32'h399067a2),
	.w2(32'h3979bb95),
	.w3(32'h3a3f5846),
	.w4(32'h3a594af2),
	.w5(32'h38a0e26f),
	.w6(32'hb9b7b6d9),
	.w7(32'hb8f04f4b),
	.w8(32'hb8f1db1a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bec2db),
	.w1(32'h39e7e365),
	.w2(32'hba405fbe),
	.w3(32'hb9da1d8b),
	.w4(32'hb8eddfa8),
	.w5(32'hba7bf79d),
	.w6(32'hb9a2d593),
	.w7(32'hb92c49f1),
	.w8(32'hbb20b0dc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d100c),
	.w1(32'hbb6ec85c),
	.w2(32'hbaf3a3d1),
	.w3(32'hbb39ee77),
	.w4(32'hbb3b3187),
	.w5(32'hbb871e83),
	.w6(32'hbb8eeb8d),
	.w7(32'hbb55eb64),
	.w8(32'h3980ee7d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b0fdf),
	.w1(32'hb7b15e12),
	.w2(32'hb9d88a8d),
	.w3(32'h39d0d7a7),
	.w4(32'h39b2ffda),
	.w5(32'h386145af),
	.w6(32'hba85f560),
	.w7(32'hba913468),
	.w8(32'h3a8d8233),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0d6d3),
	.w1(32'h3aa2f637),
	.w2(32'h3a79a020),
	.w3(32'h3a8a4639),
	.w4(32'h3a197275),
	.w5(32'hb9cb6153),
	.w6(32'h3a38f50c),
	.w7(32'h3923b89e),
	.w8(32'hbbbf09b4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aced0),
	.w1(32'hbb73c126),
	.w2(32'hb9c45c98),
	.w3(32'hbaf5d1da),
	.w4(32'hbb652409),
	.w5(32'hbba0b135),
	.w6(32'hba1f99df),
	.w7(32'h3b16b4e6),
	.w8(32'h3a508ae5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0469a),
	.w1(32'h3aa47bc9),
	.w2(32'h3ab5eb4b),
	.w3(32'h3ab524a8),
	.w4(32'h3b1f91bf),
	.w5(32'h3b2890bd),
	.w6(32'h3968ce0d),
	.w7(32'hba0e14cc),
	.w8(32'h3996bfbf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a086eb9),
	.w1(32'h39e4c061),
	.w2(32'hba535e91),
	.w3(32'h392d53df),
	.w4(32'h3a20798f),
	.w5(32'hb826739f),
	.w6(32'hba2f4363),
	.w7(32'hbadb8eea),
	.w8(32'hbaeef62a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae61d),
	.w1(32'hb9b6bfa2),
	.w2(32'h3a82ff76),
	.w3(32'hbb625758),
	.w4(32'hbac6a80d),
	.w5(32'h3a4d8147),
	.w6(32'hba93e5a7),
	.w7(32'hb994268e),
	.w8(32'h38988ac5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380ada),
	.w1(32'hbaa01789),
	.w2(32'hb98ebe30),
	.w3(32'h3a05221a),
	.w4(32'hba5850db),
	.w5(32'hba93ab14),
	.w6(32'hba3a5329),
	.w7(32'hba51f52a),
	.w8(32'hbb079d44),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6280d4),
	.w1(32'hb98fb7e0),
	.w2(32'h3b11371b),
	.w3(32'hbb59ca78),
	.w4(32'hbb8f90cb),
	.w5(32'hbb0e60cb),
	.w6(32'hb9db2792),
	.w7(32'hb9d28674),
	.w8(32'hbaf9a0aa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e983e),
	.w1(32'hb98dd864),
	.w2(32'h3a828d3c),
	.w3(32'hbb4d6499),
	.w4(32'hbaabe2e7),
	.w5(32'h3a4f1b36),
	.w6(32'hba82e007),
	.w7(32'hb938e091),
	.w8(32'hbace85c5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35e90a),
	.w1(32'hb969c50f),
	.w2(32'h3a5b952a),
	.w3(32'hbb331409),
	.w4(32'hba9a6d2d),
	.w5(32'h3a1e4c4d),
	.w6(32'hba642c64),
	.w7(32'hb93b3384),
	.w8(32'h3a90e913),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a936949),
	.w1(32'h3a4e099c),
	.w2(32'h3aaa1a5f),
	.w3(32'h385daefd),
	.w4(32'h3a75274e),
	.w5(32'h3b002ef5),
	.w6(32'h3a04c1e6),
	.w7(32'hb9ace6be),
	.w8(32'hbb5df795),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e0acc),
	.w1(32'hb930a4ed),
	.w2(32'hbbd4f723),
	.w3(32'hba502145),
	.w4(32'h3ac410b7),
	.w5(32'hbbd1ef4f),
	.w6(32'hbab3c7ab),
	.w7(32'hb98aab25),
	.w8(32'h39517c35),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958b662),
	.w1(32'hb7d23652),
	.w2(32'hb91763ad),
	.w3(32'h39b98f63),
	.w4(32'h3967b824),
	.w5(32'h388d198a),
	.w6(32'hb99e26ab),
	.w7(32'hb9f5cfac),
	.w8(32'hb99a7c7e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bf722),
	.w1(32'hba9a7f1e),
	.w2(32'h3ab17430),
	.w3(32'h3b21f346),
	.w4(32'h3a89808a),
	.w5(32'hbaa15b6f),
	.w6(32'hbb0ab9b8),
	.w7(32'h3b34c18e),
	.w8(32'h3939787f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67801b),
	.w1(32'h3a602cd1),
	.w2(32'h3af61a74),
	.w3(32'hb9793275),
	.w4(32'h3ab73d20),
	.w5(32'h3b198ad0),
	.w6(32'hba937b23),
	.w7(32'hbb1f6315),
	.w8(32'hba99aebd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cbb7),
	.w1(32'hbbadcc70),
	.w2(32'hbb2104fe),
	.w3(32'h3a9923ac),
	.w4(32'hba71ba99),
	.w5(32'hbb561677),
	.w6(32'hbb266ffb),
	.w7(32'hbaa998e7),
	.w8(32'h3abea047),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4749e),
	.w1(32'h3bbae645),
	.w2(32'h3b21c306),
	.w3(32'h3a9a4173),
	.w4(32'hbb542366),
	.w5(32'hbb377b41),
	.w6(32'h3b1d6757),
	.w7(32'h3b7eb65e),
	.w8(32'hb8cc7f19),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e44b64),
	.w1(32'hb8f96f54),
	.w2(32'h3a598b93),
	.w3(32'hb83342eb),
	.w4(32'hb9b4da7b),
	.w5(32'hba313ca2),
	.w6(32'hba210bbd),
	.w7(32'h3a23ea45),
	.w8(32'h3a364cf8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a411213),
	.w1(32'h398ff5b1),
	.w2(32'h39fe4b74),
	.w3(32'h3984135e),
	.w4(32'h3718bf66),
	.w5(32'hb985bddc),
	.w6(32'h3a1eaebc),
	.w7(32'h3971a632),
	.w8(32'hba524aec),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba575a33),
	.w1(32'hbb0de86e),
	.w2(32'h3a52150a),
	.w3(32'hbac6e312),
	.w4(32'hbb6d7864),
	.w5(32'hba64882b),
	.w6(32'h39091e6d),
	.w7(32'h39e94caa),
	.w8(32'h399031ea),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c85146),
	.w1(32'hba3a0f3b),
	.w2(32'hba196799),
	.w3(32'h3977a2b2),
	.w4(32'hb6b31f9d),
	.w5(32'hb7f545c7),
	.w6(32'hba562db1),
	.w7(32'hba96ac6c),
	.w8(32'h398b6a81),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7333a14),
	.w1(32'h3763ec72),
	.w2(32'hb960c79b),
	.w3(32'h3a8da5e4),
	.w4(32'h3ac45d8f),
	.w5(32'hb7dab0eb),
	.w6(32'hbac10a77),
	.w7(32'hba7bfbba),
	.w8(32'h39091e14),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3840256b),
	.w1(32'h39dd1323),
	.w2(32'h3aab0ce0),
	.w3(32'hba8e31fe),
	.w4(32'hb9eb6a23),
	.w5(32'h3a465d0e),
	.w6(32'hb7ff5a13),
	.w7(32'hba1695c2),
	.w8(32'hba4819ea),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a98d6e),
	.w1(32'hb90a3b3d),
	.w2(32'h39a054b6),
	.w3(32'hbaa46a32),
	.w4(32'hba138464),
	.w5(32'h398987f1),
	.w6(32'hb9c8f49f),
	.w7(32'hb8fcf000),
	.w8(32'h3b7418d5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d441a),
	.w1(32'hbb9ee7d2),
	.w2(32'hb8859df5),
	.w3(32'hbb5619f1),
	.w4(32'hba5a7e80),
	.w5(32'h3bb62795),
	.w6(32'hb81fb705),
	.w7(32'hbb46069f),
	.w8(32'hbafe0dda),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fc7e6),
	.w1(32'h3d44b7cb),
	.w2(32'h3d470f1d),
	.w3(32'hbc7d5d12),
	.w4(32'h3c6e310d),
	.w5(32'h3b0bfef8),
	.w6(32'h3cabfc16),
	.w7(32'h3bbddd94),
	.w8(32'h3a72c12b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826ed1),
	.w1(32'hbbb8f0d1),
	.w2(32'hb8206e37),
	.w3(32'hbbc1e92b),
	.w4(32'hbbd8bc91),
	.w5(32'h38bf295d),
	.w6(32'hbb5d326f),
	.w7(32'hba69de83),
	.w8(32'h3b738acc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8286a9),
	.w1(32'hbc37406c),
	.w2(32'hba29211d),
	.w3(32'hba9b19d8),
	.w4(32'hbb679d67),
	.w5(32'hba39df9b),
	.w6(32'hbae183fd),
	.w7(32'hba06bea9),
	.w8(32'h3864569a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bceb8b8),
	.w1(32'h3bd781bb),
	.w2(32'h3afb495f),
	.w3(32'hbbf83efc),
	.w4(32'hbc2dd647),
	.w5(32'h3ae6e05d),
	.w6(32'hbc34ea5e),
	.w7(32'hbc5ee5c9),
	.w8(32'hbca1a3d9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd75735),
	.w1(32'h3d876a23),
	.w2(32'h3c1e5554),
	.w3(32'h3a47ed77),
	.w4(32'h3c6d66ee),
	.w5(32'hba88dbae),
	.w6(32'h3c8cf7e9),
	.w7(32'h3c824613),
	.w8(32'hbbc8bad7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b404ba5),
	.w1(32'h3bd351c2),
	.w2(32'h3b770d13),
	.w3(32'hbc1e2c7c),
	.w4(32'hbbe89bab),
	.w5(32'hbb360bf2),
	.w6(32'hbc16cd4a),
	.w7(32'hbc9c686e),
	.w8(32'h3c736833),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66c752),
	.w1(32'h3b59e88a),
	.w2(32'hbb013c5f),
	.w3(32'h3c70eaba),
	.w4(32'h3c044cfa),
	.w5(32'h3be8fab9),
	.w6(32'h3c0e5314),
	.w7(32'h38094c3a),
	.w8(32'h3b00310a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349d49),
	.w1(32'hbc19b16d),
	.w2(32'h3b2b028c),
	.w3(32'hbbabb03b),
	.w4(32'hbb24b132),
	.w5(32'hbb02b8e8),
	.w6(32'hbb8484e8),
	.w7(32'hbb9273f8),
	.w8(32'h387b6d2d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f71a90),
	.w1(32'hb9341788),
	.w2(32'h3b34b573),
	.w3(32'hbb0172c4),
	.w4(32'hba8c03db),
	.w5(32'h3a9ee834),
	.w6(32'hba9bc360),
	.w7(32'h39ee841c),
	.w8(32'h3aa8c3c5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8f7ea),
	.w1(32'hb8fbb38d),
	.w2(32'h3b5ec5b7),
	.w3(32'hbbbf5159),
	.w4(32'hbb1def42),
	.w5(32'h3a014d25),
	.w6(32'hbb78140a),
	.w7(32'h3a05e041),
	.w8(32'h3ba05d08),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38d52d),
	.w1(32'h3d1a9140),
	.w2(32'hbbd95ffa),
	.w3(32'h3c3781a9),
	.w4(32'h3c4b29f0),
	.w5(32'hbba73e55),
	.w6(32'hbaf1c594),
	.w7(32'h3b0e7e4f),
	.w8(32'h3bcc98f8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f6e7d),
	.w1(32'hbab0401f),
	.w2(32'h3a8e0176),
	.w3(32'h3ab684f7),
	.w4(32'h3bbdce33),
	.w5(32'h3abaf504),
	.w6(32'h3b517d05),
	.w7(32'hbb4f770c),
	.w8(32'h3bd5f920),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03d41a),
	.w1(32'h3d06f68a),
	.w2(32'hbb282efc),
	.w3(32'h3ca51aef),
	.w4(32'h3d05a284),
	.w5(32'hbc1e4ea2),
	.w6(32'h3cbcc1f2),
	.w7(32'h38e771f5),
	.w8(32'h3b9eb813),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e142e),
	.w1(32'h3d93e781),
	.w2(32'h3c1ce979),
	.w3(32'h3a572516),
	.w4(32'h3c6dd96b),
	.w5(32'h3c2a3d9e),
	.w6(32'h3ca596a6),
	.w7(32'h3b381012),
	.w8(32'h3b2c0b8f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbddb2a),
	.w1(32'h3d11301d),
	.w2(32'h3d1ff9b6),
	.w3(32'h3cc9f96b),
	.w4(32'h3ce48ea6),
	.w5(32'hbc71491c),
	.w6(32'h3cb5886d),
	.w7(32'h3cb2f9e9),
	.w8(32'h3bc09c8d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94270c),
	.w1(32'h3dbcb666),
	.w2(32'h3c2f43a4),
	.w3(32'hbc220c5f),
	.w4(32'h3d0b33f8),
	.w5(32'h3c1c5101),
	.w6(32'h3b8e57da),
	.w7(32'h3b09a245),
	.w8(32'h3c7d386a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1daf02),
	.w1(32'h3b25b2f5),
	.w2(32'h3b93b43c),
	.w3(32'h3c89f5f6),
	.w4(32'h3bbaaf18),
	.w5(32'h3c3bb40b),
	.w6(32'h3c130d37),
	.w7(32'h3c1f1aa8),
	.w8(32'h3c428e61),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c473),
	.w1(32'hbc4246cc),
	.w2(32'hbb6ee9a5),
	.w3(32'hbbc84983),
	.w4(32'hbc1cde8d),
	.w5(32'h3a15d81e),
	.w6(32'h3b355227),
	.w7(32'hbb2a7986),
	.w8(32'hbb177890),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb25316),
	.w1(32'h3d4a53cc),
	.w2(32'h3d084abd),
	.w3(32'h3be814af),
	.w4(32'h3cd2b917),
	.w5(32'hbb9084af),
	.w6(32'h3aab9c91),
	.w7(32'h3a91eb88),
	.w8(32'hbbc33706),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7616c0),
	.w1(32'h3ba6c40b),
	.w2(32'h3bcf71be),
	.w3(32'hbc8c62ec),
	.w4(32'hbc417e0b),
	.w5(32'hbb814ac1),
	.w6(32'hbc59fa09),
	.w7(32'hbc72c539),
	.w8(32'h3bce41f4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999ae2c),
	.w1(32'hbbbf4cbb),
	.w2(32'h3adbd4db),
	.w3(32'hbba8c373),
	.w4(32'hbb513cdb),
	.w5(32'h3bad203c),
	.w6(32'hbaf40878),
	.w7(32'hbb104d53),
	.w8(32'hbcabab95),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81184d),
	.w1(32'h3d506fec),
	.w2(32'h3c899c18),
	.w3(32'hba604724),
	.w4(32'hbb4aa86b),
	.w5(32'hbb8bfe87),
	.w6(32'hbc887ac9),
	.w7(32'hbc30dfc5),
	.w8(32'hba9a0909),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule