module layer_10_featuremap_459(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837415),
	.w1(32'h39bbb612),
	.w2(32'hb9766ee7),
	.w3(32'hbb73e3c3),
	.w4(32'hb9641bd6),
	.w5(32'hbb21a56a),
	.w6(32'hbadecdf3),
	.w7(32'h39b15f53),
	.w8(32'h3a9cc2be),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109864),
	.w1(32'hbad25959),
	.w2(32'hbbad7456),
	.w3(32'h3a80d70e),
	.w4(32'hbae52bd0),
	.w5(32'hbb7a4786),
	.w6(32'h3a4f00d9),
	.w7(32'hbb0d8dfb),
	.w8(32'hbbb9fe7d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6d988),
	.w1(32'h39e66d89),
	.w2(32'h3b2501d0),
	.w3(32'hbb79d2e0),
	.w4(32'h3a54011b),
	.w5(32'h3b036f24),
	.w6(32'hbb8978bf),
	.w7(32'h3ad1c9b1),
	.w8(32'h3b698c9f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147387),
	.w1(32'h3b0a8cec),
	.w2(32'hba29660d),
	.w3(32'hb98cfca3),
	.w4(32'hba8dd1c0),
	.w5(32'hba3668a1),
	.w6(32'h3b0619b4),
	.w7(32'hba744933),
	.w8(32'hb9c2524a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d32f5),
	.w1(32'h3a840e88),
	.w2(32'h3af36494),
	.w3(32'h3ac9a152),
	.w4(32'h39d7c348),
	.w5(32'h3a76cafa),
	.w6(32'h3b08f58c),
	.w7(32'h3aa43232),
	.w8(32'h3b05d7a9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aa6ff),
	.w1(32'h3a136299),
	.w2(32'hbaa29960),
	.w3(32'hba371f0d),
	.w4(32'h3b1a007c),
	.w5(32'h3a921607),
	.w6(32'h39e73774),
	.w7(32'h3b16afa3),
	.w8(32'hba16ef64),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398245b7),
	.w1(32'h3a288d68),
	.w2(32'h3a7d7fde),
	.w3(32'hbae246ad),
	.w4(32'h3a5f6174),
	.w5(32'hba0161a3),
	.w6(32'hbab34142),
	.w7(32'hba2ff528),
	.w8(32'hb8f4f401),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61ff4f),
	.w1(32'hb8684360),
	.w2(32'hbabe72a3),
	.w3(32'h3a628076),
	.w4(32'hb933737f),
	.w5(32'hbb668982),
	.w6(32'hba20b225),
	.w7(32'hb9883e6b),
	.w8(32'hbb68f8d3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c78aa),
	.w1(32'h3acbdf06),
	.w2(32'h3aff9ce1),
	.w3(32'hba56e25e),
	.w4(32'h3a59f1f3),
	.w5(32'hba75ce5a),
	.w6(32'hba0375e8),
	.w7(32'h3b0de8e5),
	.w8(32'hbac141d3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f39e8),
	.w1(32'h3a3cd931),
	.w2(32'hba0366e9),
	.w3(32'h39b31ecb),
	.w4(32'h3a89f2d2),
	.w5(32'hbb089ffa),
	.w6(32'h3a0ceaf9),
	.w7(32'hb9a5d1f2),
	.w8(32'hba5e9a12),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953fae6),
	.w1(32'hba48c94f),
	.w2(32'h390ea6e2),
	.w3(32'hba25486f),
	.w4(32'hba2d60ef),
	.w5(32'hba2934ce),
	.w6(32'hba444144),
	.w7(32'hbafb1027),
	.w8(32'hbadbbf27),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a402def),
	.w1(32'h3a92ae06),
	.w2(32'h3ae39fa8),
	.w3(32'h3abe1aeb),
	.w4(32'h3aa3fe79),
	.w5(32'hb99b21f7),
	.w6(32'h3a2fcad9),
	.w7(32'h3a4c2d09),
	.w8(32'hb883aef8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f253),
	.w1(32'hbb1a9f51),
	.w2(32'hbb8e133f),
	.w3(32'hba15b61f),
	.w4(32'hbba11b8c),
	.w5(32'hbb58f04a),
	.w6(32'h3a7269da),
	.w7(32'hbba96e95),
	.w8(32'hbbd5b4ff),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf097d),
	.w1(32'h39154d23),
	.w2(32'h3b8826ab),
	.w3(32'hbbae50f1),
	.w4(32'h3a58132d),
	.w5(32'h3b6cfa22),
	.w6(32'hbb9ea770),
	.w7(32'h3b74fcc1),
	.w8(32'h3bb30138),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399687f6),
	.w1(32'h399aadb1),
	.w2(32'h3a112115),
	.w3(32'h3a483747),
	.w4(32'hba3ba713),
	.w5(32'h3abb9184),
	.w6(32'h3b250029),
	.w7(32'hba76a871),
	.w8(32'hb81c7c14),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1886fe),
	.w1(32'hb9b3d0b2),
	.w2(32'hba307411),
	.w3(32'hbae1195f),
	.w4(32'hba027f72),
	.w5(32'h39b234d0),
	.w6(32'hba6df021),
	.w7(32'h3944b811),
	.w8(32'h3ad3c454),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ab00f),
	.w1(32'hba0d7453),
	.w2(32'hba1a7de8),
	.w3(32'hbb1f5648),
	.w4(32'hba83c378),
	.w5(32'hba493dc2),
	.w6(32'hb8e50b3e),
	.w7(32'hbad6621f),
	.w8(32'hbb238402),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf80a38),
	.w1(32'h3aaf658d),
	.w2(32'h3a358b88),
	.w3(32'h3a373652),
	.w4(32'h3a5f30c1),
	.w5(32'h3a8a85bb),
	.w6(32'hba314ffb),
	.w7(32'h3a668d74),
	.w8(32'h3b06277c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab06197),
	.w1(32'hbb0a0798),
	.w2(32'hb95bcc83),
	.w3(32'h3b09dbd6),
	.w4(32'hbaf3a460),
	.w5(32'hbacc907c),
	.w6(32'h3b2a87e7),
	.w7(32'hba406556),
	.w8(32'hbabee922),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9993831),
	.w1(32'h3afbc2b0),
	.w2(32'h3ba40123),
	.w3(32'hba8340e1),
	.w4(32'h3a2882e5),
	.w5(32'h3bd2f3a1),
	.w6(32'hb9e71835),
	.w7(32'hba107bca),
	.w8(32'hb8c7a50e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefbd48),
	.w1(32'h3b11ba86),
	.w2(32'h3b6e1fcc),
	.w3(32'hba33b526),
	.w4(32'h3b1e7d4a),
	.w5(32'h3a0f4d13),
	.w6(32'h3b22aea1),
	.w7(32'h3b78c0a9),
	.w8(32'h3a2f7754),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bc93f),
	.w1(32'hbba49911),
	.w2(32'h3b4381fb),
	.w3(32'hbb0281cc),
	.w4(32'hbb984162),
	.w5(32'h3bbeafc1),
	.w6(32'h395f53b4),
	.w7(32'hbb3b15c2),
	.w8(32'h3b69bc88),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f947b),
	.w1(32'hba1fe82e),
	.w2(32'h3a673530),
	.w3(32'hba70ed26),
	.w4(32'hba27f2c4),
	.w5(32'h3b196273),
	.w6(32'hbabcb83e),
	.w7(32'h3a022a0d),
	.w8(32'h39d381d7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a521eee),
	.w1(32'hbaac939e),
	.w2(32'hbb1408b6),
	.w3(32'h3b70e34a),
	.w4(32'hbc002519),
	.w5(32'hbbf7de71),
	.w6(32'h3afcd46a),
	.w7(32'hbaf587b6),
	.w8(32'hbb4a7c69),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248923),
	.w1(32'hbba26612),
	.w2(32'hbb193650),
	.w3(32'hbc0f292f),
	.w4(32'hbbb77b07),
	.w5(32'hbaad7b60),
	.w6(32'hbb088570),
	.w7(32'hbb138441),
	.w8(32'hb7a7099f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeb735),
	.w1(32'h3ae98dc3),
	.w2(32'hbab74da9),
	.w3(32'hbaa11021),
	.w4(32'h3abd46c3),
	.w5(32'hbbcf742d),
	.w6(32'h3ab8d36d),
	.w7(32'h3b1662ec),
	.w8(32'hb9d920bd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d0c52),
	.w1(32'hb7471e7f),
	.w2(32'h3a795d53),
	.w3(32'hb8018f72),
	.w4(32'h3b58ce97),
	.w5(32'h39ad2fba),
	.w6(32'h3aadfaca),
	.w7(32'h3ac39836),
	.w8(32'h3ac65cee),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6191b),
	.w1(32'hba825ff5),
	.w2(32'hbb706edc),
	.w3(32'h39bed122),
	.w4(32'hba5a09ce),
	.w5(32'hbb67f48b),
	.w6(32'hba0465e9),
	.w7(32'hbabf4698),
	.w8(32'hbb12912e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20791d),
	.w1(32'hbb2b293f),
	.w2(32'hbb31783f),
	.w3(32'h39ae36e8),
	.w4(32'hbb0293d6),
	.w5(32'hbb743702),
	.w6(32'h3ab4ee08),
	.w7(32'hb98d2cd6),
	.w8(32'hbb28711b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae13d77),
	.w1(32'h3b0157cf),
	.w2(32'h3b2c96e7),
	.w3(32'hb8d9391a),
	.w4(32'h3acb14da),
	.w5(32'h3b005003),
	.w6(32'h3aa2d331),
	.w7(32'h3a9ba3f7),
	.w8(32'h39ffa2f6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45c9ad),
	.w1(32'h3aea455b),
	.w2(32'h3b8fce58),
	.w3(32'hba182715),
	.w4(32'h3b66ce3e),
	.w5(32'h3b728b88),
	.w6(32'hb9ce09e0),
	.w7(32'h3af7939d),
	.w8(32'h3aea7204),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac879e5),
	.w1(32'hbab6ac8f),
	.w2(32'hba843a07),
	.w3(32'h3b899f55),
	.w4(32'hba3a0605),
	.w5(32'h3a30b00e),
	.w6(32'h3b4f12ef),
	.w7(32'hbabd7564),
	.w8(32'h39c41379),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53b58d),
	.w1(32'hbab2b102),
	.w2(32'h39f8a146),
	.w3(32'hb948cae9),
	.w4(32'h39cfdbb6),
	.w5(32'hba8f5e83),
	.w6(32'hb920a80c),
	.w7(32'h3aa36507),
	.w8(32'hb9fe593f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3baef),
	.w1(32'hba92ef4a),
	.w2(32'h39b205fc),
	.w3(32'hba5d2e04),
	.w4(32'h398ad5c0),
	.w5(32'hb8fed1d0),
	.w6(32'hbb4d5c95),
	.w7(32'h383fc8fe),
	.w8(32'hba8854ee),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab349f1),
	.w1(32'h3ac4c9d6),
	.w2(32'h3b8618d5),
	.w3(32'h3b219a18),
	.w4(32'h3a84dce3),
	.w5(32'h3b0e140e),
	.w6(32'h3a530207),
	.w7(32'h3b607ac4),
	.w8(32'h3ae95299),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed9dde),
	.w1(32'h3aa7319e),
	.w2(32'h3ac71e36),
	.w3(32'h3b8ee9b1),
	.w4(32'h39bfa42c),
	.w5(32'h3a907ddb),
	.w6(32'h3b8b707f),
	.w7(32'h3a52dd40),
	.w8(32'h3abe5bd1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6de8c),
	.w1(32'hbb89c2ef),
	.w2(32'hbb4be7a0),
	.w3(32'h38fa19d9),
	.w4(32'hba488a43),
	.w5(32'hbb29e70b),
	.w6(32'h3ac89fee),
	.w7(32'hbad76929),
	.w8(32'hbb7d2a33),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f4681),
	.w1(32'hba2de20a),
	.w2(32'hbb293f76),
	.w3(32'h398d6f61),
	.w4(32'hba0da296),
	.w5(32'hb997fc25),
	.w6(32'hba9ddeec),
	.w7(32'hba587c0b),
	.w8(32'hbb6e7937),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3139f),
	.w1(32'h3ade75d6),
	.w2(32'h39d4b961),
	.w3(32'hbb48c98b),
	.w4(32'hbad09257),
	.w5(32'hbb6f5f25),
	.w6(32'hbb911516),
	.w7(32'h3abe332e),
	.w8(32'hb9cde54f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90638cf),
	.w1(32'hb989e3d8),
	.w2(32'hb936b8fa),
	.w3(32'hba33a025),
	.w4(32'h3ac12dce),
	.w5(32'h37a9f3de),
	.w6(32'h3ab0e651),
	.w7(32'h3aeffc59),
	.w8(32'hb98ddf6c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974e497),
	.w1(32'h3b17f5f6),
	.w2(32'hbaf0a672),
	.w3(32'h3b74b8c0),
	.w4(32'hb95516e0),
	.w5(32'hbae4b277),
	.w6(32'h3b3b7a40),
	.w7(32'h3ad53278),
	.w8(32'h3adcbe9e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c4bd0),
	.w1(32'hb99fa968),
	.w2(32'hb9e5a3ea),
	.w3(32'h3b9423a1),
	.w4(32'h38ed7f30),
	.w5(32'h3a67cc4d),
	.w6(32'h3b950c3a),
	.w7(32'hba973a89),
	.w8(32'hbafaea34),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6ae73),
	.w1(32'hba9a40a3),
	.w2(32'hbb9453ed),
	.w3(32'h3a54dacd),
	.w4(32'hbb2e2587),
	.w5(32'hb9b48b03),
	.w6(32'h3a1bb22e),
	.w7(32'hbb59b408),
	.w8(32'hbb4906a2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0090be),
	.w1(32'h3a63a5dd),
	.w2(32'hbb61807f),
	.w3(32'hbb144ce8),
	.w4(32'hb8e1dff2),
	.w5(32'hbbcf1cf7),
	.w6(32'hbac4e185),
	.w7(32'h3aa2cd3a),
	.w8(32'hbb99960d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba974eff),
	.w1(32'hbb14bd2b),
	.w2(32'hba92c174),
	.w3(32'h3a15780b),
	.w4(32'hbab3c97e),
	.w5(32'hba4145c7),
	.w6(32'h39b0a9ff),
	.w7(32'hbafaf1ca),
	.w8(32'hbaad1591),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00c46a),
	.w1(32'hba1b5dca),
	.w2(32'hbb1d0d0f),
	.w3(32'hbae529d6),
	.w4(32'hbac0859f),
	.w5(32'hbaec3afc),
	.w6(32'hb949a69b),
	.w7(32'hba41d6f1),
	.w8(32'hb9c6d3ed),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ef9aa),
	.w1(32'h3ad39def),
	.w2(32'h39e1b148),
	.w3(32'hbba09d2c),
	.w4(32'h3a1d7869),
	.w5(32'hbaa0b7d4),
	.w6(32'hbae683c3),
	.w7(32'h3b094d3a),
	.w8(32'h3a6f857a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c30911),
	.w1(32'hba317edd),
	.w2(32'h3aba4d95),
	.w3(32'h38c294fd),
	.w4(32'hb91eaff9),
	.w5(32'h3aedb02a),
	.w6(32'h37897c78),
	.w7(32'h3908fb23),
	.w8(32'h39f4e9a3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93a93c),
	.w1(32'h3b5bcc96),
	.w2(32'h3c015e10),
	.w3(32'h3acef05e),
	.w4(32'h3abd06fd),
	.w5(32'h3b279711),
	.w6(32'h3ae7422d),
	.w7(32'h3b7e6858),
	.w8(32'h3bba7f4d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae807c),
	.w1(32'h3aeeb71e),
	.w2(32'h3b14b3be),
	.w3(32'h3932338a),
	.w4(32'h3af33425),
	.w5(32'h3a59263b),
	.w6(32'h3b1e3e15),
	.w7(32'h3b068306),
	.w8(32'h3b8958d3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846c8c),
	.w1(32'h3b000054),
	.w2(32'hba005ec0),
	.w3(32'h3b4b427a),
	.w4(32'hbaaa7909),
	.w5(32'hbb4f0f12),
	.w6(32'h3b7caf45),
	.w7(32'h3ac1ff19),
	.w8(32'hbb158068),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62195d),
	.w1(32'hb9e88d50),
	.w2(32'h3b120c10),
	.w3(32'hba1a3ff1),
	.w4(32'hba247b0c),
	.w5(32'h3b407a84),
	.w6(32'hba3407c9),
	.w7(32'h398a3705),
	.w8(32'h3b09213d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d90f8),
	.w1(32'h3a076af3),
	.w2(32'h3aaaef54),
	.w3(32'hbb0e8ea4),
	.w4(32'h3a83c0a2),
	.w5(32'h3ad66e54),
	.w6(32'hbb2b3dc9),
	.w7(32'h3a8498c3),
	.w8(32'h3a8af045),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9061e0),
	.w1(32'h39ec39af),
	.w2(32'h38d2b9cb),
	.w3(32'h3ad513ec),
	.w4(32'h3b01b15a),
	.w5(32'h3a434f82),
	.w6(32'h3af5ce58),
	.w7(32'h3aec3699),
	.w8(32'hba8a71a7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20aadf),
	.w1(32'hb9e7572b),
	.w2(32'hbab9d482),
	.w3(32'h3ac98b99),
	.w4(32'h3a5f2b36),
	.w5(32'h3af35593),
	.w6(32'h3a70b7f3),
	.w7(32'hb92ac4bf),
	.w8(32'hbb32605e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945d574),
	.w1(32'hbb191b50),
	.w2(32'hbb86e11c),
	.w3(32'h3aa142d5),
	.w4(32'hba2fb4e8),
	.w5(32'hba627fc1),
	.w6(32'hbafc7648),
	.w7(32'h3a955e96),
	.w8(32'hbb9d1c2c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ed8f7),
	.w1(32'h3a79b21e),
	.w2(32'hba905aff),
	.w3(32'hbbb4d177),
	.w4(32'hb9251e0a),
	.w5(32'hbb3ee082),
	.w6(32'hbba93c1c),
	.w7(32'h3a0e2ac6),
	.w8(32'hba5ca429),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3d06b),
	.w1(32'hb77287b1),
	.w2(32'hba87a04b),
	.w3(32'hbb03517d),
	.w4(32'hba4be8a6),
	.w5(32'h3a3a2215),
	.w6(32'hb9839d12),
	.w7(32'hba2d7cf1),
	.w8(32'hbac15e15),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4231a2),
	.w1(32'hb8987a59),
	.w2(32'hbc0c3c87),
	.w3(32'h39e30085),
	.w4(32'hbac7af04),
	.w5(32'hbbc5da8c),
	.w6(32'hb7acf1c1),
	.w7(32'hbb339e6d),
	.w8(32'hbbe16e4e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded680),
	.w1(32'hba6acfb5),
	.w2(32'hba08f036),
	.w3(32'hbbe66600),
	.w4(32'h39aff0e0),
	.w5(32'hb98bf0f0),
	.w6(32'hbbcb95ab),
	.w7(32'hb9e37386),
	.w8(32'hbb5efd98),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ce6ac),
	.w1(32'h3b2afab1),
	.w2(32'h394644b2),
	.w3(32'hb9059dd6),
	.w4(32'h3b0ae7f1),
	.w5(32'hbb1dbfd2),
	.w6(32'hba6a2dda),
	.w7(32'h3aef720f),
	.w8(32'hbb252a93),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6abd2),
	.w1(32'h38796f47),
	.w2(32'hb91ea9c9),
	.w3(32'h3a832b8e),
	.w4(32'h381a9f9a),
	.w5(32'hbaf884e7),
	.w6(32'hb9e70626),
	.w7(32'h39443534),
	.w8(32'hbaaf3bdb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a98044),
	.w1(32'hbb211f62),
	.w2(32'hbbd8116b),
	.w3(32'hb9a67cf4),
	.w4(32'hbb955d85),
	.w5(32'hbbad4b35),
	.w6(32'hb92d00e5),
	.w7(32'hbb3df28d),
	.w8(32'hbb874e20),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0930f8),
	.w1(32'h3a7616dd),
	.w2(32'hb9127cd3),
	.w3(32'hbb253baa),
	.w4(32'hb83fd8e8),
	.w5(32'hbb5b5fe2),
	.w6(32'hba251a5b),
	.w7(32'hba9f5ea1),
	.w8(32'hbaef3188),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d8344),
	.w1(32'h3bb14552),
	.w2(32'h3b82478c),
	.w3(32'hb9d681cb),
	.w4(32'h3b72df85),
	.w5(32'h39d335a9),
	.w6(32'h39a27f67),
	.w7(32'h3bd5f450),
	.w8(32'h3b8270a2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b9aba),
	.w1(32'h3b735284),
	.w2(32'h3b4905a4),
	.w3(32'h3b2b2135),
	.w4(32'h3b3ad733),
	.w5(32'h3ab01013),
	.w6(32'h3badcd4c),
	.w7(32'h3b9a9635),
	.w8(32'h3b906d1f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e152f0),
	.w1(32'h3b0df6e6),
	.w2(32'h3aa71d3e),
	.w3(32'h3a35f9de),
	.w4(32'h3b1c607f),
	.w5(32'h3ac71012),
	.w6(32'h3b9958d2),
	.w7(32'h3affe2b2),
	.w8(32'h3aa0360e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0743f1),
	.w1(32'h3b3ba398),
	.w2(32'h39de38ba),
	.w3(32'h373cbd7e),
	.w4(32'h3b7730f3),
	.w5(32'hbb3da934),
	.w6(32'hb9ceb0b8),
	.w7(32'h3b5c5d5c),
	.w8(32'hbacccede),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9101a6),
	.w1(32'hbac47a97),
	.w2(32'hbab5728c),
	.w3(32'hbb39c548),
	.w4(32'h3997979f),
	.w5(32'hb8ccff16),
	.w6(32'hbb11c33a),
	.w7(32'h3ab36c6a),
	.w8(32'hbaf66468),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acffbbd),
	.w1(32'h3b64777e),
	.w2(32'h3b659dfe),
	.w3(32'h3a83a125),
	.w4(32'hbaddbc7e),
	.w5(32'h3b50833b),
	.w6(32'h398e312e),
	.w7(32'hbb6f08d5),
	.w8(32'h3bfe065b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b207cc9),
	.w1(32'hbae84bee),
	.w2(32'h3b0936be),
	.w3(32'hbb278fa7),
	.w4(32'h3a0e7f58),
	.w5(32'hbc0c217a),
	.w6(32'hbacc5b09),
	.w7(32'h3a0524c2),
	.w8(32'hbab40a2f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a895afb),
	.w1(32'h3ab07dcb),
	.w2(32'h3b39dd1f),
	.w3(32'h3ab6afea),
	.w4(32'hbb51a84f),
	.w5(32'hbb944f43),
	.w6(32'h3ace9caa),
	.w7(32'hba99c2ea),
	.w8(32'h3bd195df),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38eee4),
	.w1(32'hbbc88304),
	.w2(32'hb939fb56),
	.w3(32'h3c0792d8),
	.w4(32'hbb844bb1),
	.w5(32'h3b5cb1c9),
	.w6(32'h3c25255d),
	.w7(32'hba9a2c38),
	.w8(32'h3b948ab4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6291d),
	.w1(32'h3b059be7),
	.w2(32'hba617037),
	.w3(32'h3c270a11),
	.w4(32'h39e2580c),
	.w5(32'hbb1a7d5a),
	.w6(32'hbad0a5d2),
	.w7(32'hbaf03357),
	.w8(32'h3b20de1f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76d078),
	.w1(32'hb8ba333f),
	.w2(32'hbace65c2),
	.w3(32'h3b0e3e24),
	.w4(32'hba4d169d),
	.w5(32'hbbab388e),
	.w6(32'h3aa28a91),
	.w7(32'hbabc99ab),
	.w8(32'hbbb8ab25),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5d93a),
	.w1(32'h3c005981),
	.w2(32'hbb027678),
	.w3(32'h3aee93fd),
	.w4(32'h3c20b8d9),
	.w5(32'hbaffc99c),
	.w6(32'hbb00dff1),
	.w7(32'h3c63be7d),
	.w8(32'h3c57ae19),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58a551),
	.w1(32'hbb6a5772),
	.w2(32'hbb1f9cab),
	.w3(32'h3cb41b9b),
	.w4(32'hb9cd7619),
	.w5(32'hbad41f0a),
	.w6(32'h3bb0a022),
	.w7(32'hbb2fc623),
	.w8(32'hbb4d4d4a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce6d2f),
	.w1(32'h3be07698),
	.w2(32'hba874a0f),
	.w3(32'hbc2d7397),
	.w4(32'h3b4172da),
	.w5(32'hbc4c9893),
	.w6(32'hbbdb6294),
	.w7(32'h3b6f8fd6),
	.w8(32'h3bc34dcf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfe062),
	.w1(32'h3bb84b62),
	.w2(32'h3b29f8dc),
	.w3(32'h3ae173e5),
	.w4(32'h3c14c5d5),
	.w5(32'h3ac935e8),
	.w6(32'h3c036608),
	.w7(32'h3ae7c73c),
	.w8(32'hbae65853),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d4fa5),
	.w1(32'h3a8c69ee),
	.w2(32'h3becb90e),
	.w3(32'hbb6032eb),
	.w4(32'hbbaf9b58),
	.w5(32'hba7d0355),
	.w6(32'hbb0b28e9),
	.w7(32'hbba326df),
	.w8(32'h3b5a3793),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964c9bf),
	.w1(32'hbc0b6af0),
	.w2(32'hbc0ab75a),
	.w3(32'h3aa8e026),
	.w4(32'hbbc82382),
	.w5(32'hbb83fcb8),
	.w6(32'h3bbd079c),
	.w7(32'hbbebd58a),
	.w8(32'hbc29423a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50fb2d),
	.w1(32'hbb0f8df8),
	.w2(32'hbb577dd8),
	.w3(32'hbc0ca62f),
	.w4(32'hbb5a7098),
	.w5(32'hbb91cfbf),
	.w6(32'hbba4b01f),
	.w7(32'hbaa63faf),
	.w8(32'hbb219f1d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947ebff),
	.w1(32'h3afb32a8),
	.w2(32'h3b825662),
	.w3(32'hbad6a8c4),
	.w4(32'h3ae3a745),
	.w5(32'hbba14c64),
	.w6(32'h3929ef16),
	.w7(32'h3b1e3f17),
	.w8(32'hbaf88f96),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3696d654),
	.w1(32'h3a8c0f28),
	.w2(32'hbad28d94),
	.w3(32'hba9eae15),
	.w4(32'hba17ad53),
	.w5(32'hbab22bfa),
	.w6(32'h3b86ee97),
	.w7(32'hba0d2c0e),
	.w8(32'h3acd8f56),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea0baa),
	.w1(32'hbb9425dc),
	.w2(32'hb9a226a2),
	.w3(32'h3b45e238),
	.w4(32'hbb5f9584),
	.w5(32'hba29a054),
	.w6(32'hbbab0843),
	.w7(32'hb9839697),
	.w8(32'h3c0e4239),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d86a),
	.w1(32'hbb9c8323),
	.w2(32'hbbba60f4),
	.w3(32'h3b2868a3),
	.w4(32'hbb1cf612),
	.w5(32'hbc299044),
	.w6(32'h3c139c5b),
	.w7(32'hbc0601eb),
	.w8(32'h3a541c6a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb57e2f),
	.w1(32'hba283a86),
	.w2(32'h3940cc61),
	.w3(32'h39f39c52),
	.w4(32'h3b92af3a),
	.w5(32'hbad0dd28),
	.w6(32'hbc46d0dc),
	.w7(32'h3a9a44fc),
	.w8(32'h3ba322d0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca79c1),
	.w1(32'hbb8efa4b),
	.w2(32'hbb6c9e38),
	.w3(32'h3c2aa3a0),
	.w4(32'hbafb0a00),
	.w5(32'hbc11c669),
	.w6(32'h3bfea355),
	.w7(32'hb99365c0),
	.w8(32'h3bb3b346),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b6350),
	.w1(32'h3bb776fc),
	.w2(32'h3bb39e68),
	.w3(32'h3c0368be),
	.w4(32'h3bcac76a),
	.w5(32'h3bd02d64),
	.w6(32'h3be02732),
	.w7(32'hbad72c7a),
	.w8(32'hbb113f57),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3ebf6),
	.w1(32'h3a3c5ff4),
	.w2(32'hbc32ad83),
	.w3(32'hbbe3bd0f),
	.w4(32'h3b21067b),
	.w5(32'hbba7acfd),
	.w6(32'hbb7d7ac4),
	.w7(32'hbb057801),
	.w8(32'hbbbf0242),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62e253),
	.w1(32'h3b47b289),
	.w2(32'hbb0d34c5),
	.w3(32'hbc5ac837),
	.w4(32'h3b7659b0),
	.w5(32'hbb4f0e19),
	.w6(32'h39bbcbca),
	.w7(32'hba8571e2),
	.w8(32'hbb3c19a0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76255a),
	.w1(32'h3bad9a73),
	.w2(32'h3be2175a),
	.w3(32'hbc50ff6b),
	.w4(32'h3c3cbb3a),
	.w5(32'h39e2ed56),
	.w6(32'hbbbf9bb4),
	.w7(32'h3a9d7dce),
	.w8(32'hbae73003),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42a800),
	.w1(32'h3b31e7b4),
	.w2(32'h3b909ab3),
	.w3(32'h3bc5dbb9),
	.w4(32'h3b464b3d),
	.w5(32'hbbbc3f56),
	.w6(32'hbb9a4f0b),
	.w7(32'h39c63124),
	.w8(32'hbb92eb7a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acacac2),
	.w1(32'h3bae5aa0),
	.w2(32'h3c85e9df),
	.w3(32'hbba8eb18),
	.w4(32'h3c26d308),
	.w5(32'h3c1536a3),
	.w6(32'hbba3c573),
	.w7(32'h3b82585c),
	.w8(32'h392cf09a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf51ecd),
	.w1(32'h3b05332f),
	.w2(32'h3b378191),
	.w3(32'hb9c06ffa),
	.w4(32'h3b7a8dea),
	.w5(32'hba9ac63a),
	.w6(32'hba92c6f4),
	.w7(32'hbabec4a6),
	.w8(32'hbb0efea7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc2e9),
	.w1(32'h3ba8ddca),
	.w2(32'h3aacb576),
	.w3(32'h3c06d713),
	.w4(32'h3b79f82c),
	.w5(32'h3b33507f),
	.w6(32'h3c0a2787),
	.w7(32'h3a8afb50),
	.w8(32'h3bade95d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb675c0e),
	.w1(32'hbb2d2ff7),
	.w2(32'hbbb5e72b),
	.w3(32'hbbf76536),
	.w4(32'h3a47a17d),
	.w5(32'hbb9df4bb),
	.w6(32'hbb4c0626),
	.w7(32'hbb593290),
	.w8(32'h3c0184de),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17db10),
	.w1(32'hbb1b3c20),
	.w2(32'hbba224a4),
	.w3(32'h3ca4a675),
	.w4(32'hbb779487),
	.w5(32'hbbf19422),
	.w6(32'h3c42c84a),
	.w7(32'hbba9bb58),
	.w8(32'h3b0b6684),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c7dfa),
	.w1(32'hbbe2f919),
	.w2(32'hbc070371),
	.w3(32'hbc0b3ee0),
	.w4(32'hbb69c909),
	.w5(32'hbaf73c32),
	.w6(32'hbb7481bd),
	.w7(32'hba99716e),
	.w8(32'hba39f556),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918daeb),
	.w1(32'h3bcd6d1a),
	.w2(32'h3bf380a3),
	.w3(32'h3a8dfba9),
	.w4(32'h3bad0714),
	.w5(32'h3bc2a1d5),
	.w6(32'hb901599c),
	.w7(32'hba9c9301),
	.w8(32'hb9332273),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba3ff1),
	.w1(32'hbad093cc),
	.w2(32'hbba9baca),
	.w3(32'hb9f19a2c),
	.w4(32'hbb3baf57),
	.w5(32'hbc1de04e),
	.w6(32'hba064115),
	.w7(32'hbb8e9c1f),
	.w8(32'hbb3fff4d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03ccfc),
	.w1(32'hba9fe769),
	.w2(32'hbaed428c),
	.w3(32'h3c157c5c),
	.w4(32'hba028caa),
	.w5(32'hbb03946c),
	.w6(32'h3b1ac12c),
	.w7(32'hba13afe5),
	.w8(32'hbb0b2b2c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd91cc),
	.w1(32'hbbb0cb1f),
	.w2(32'h3b19e081),
	.w3(32'hbbd65906),
	.w4(32'hbc120bab),
	.w5(32'hbc1229fe),
	.w6(32'hbb45e2dc),
	.w7(32'hbc4bff3f),
	.w8(32'h3aaf976a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a3f67),
	.w1(32'hbba3a52f),
	.w2(32'h3b6c6f4a),
	.w3(32'h3bb1d7d1),
	.w4(32'hbc61ff4a),
	.w5(32'h3c5567da),
	.w6(32'h3bc9d9f0),
	.w7(32'hbbbca813),
	.w8(32'hb980cba4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d89c),
	.w1(32'hbb4d1618),
	.w2(32'h38bfb55d),
	.w3(32'hbba2f7be),
	.w4(32'hb9f0f2c8),
	.w5(32'hbb335794),
	.w6(32'hbc39ddf4),
	.w7(32'h3bddcb35),
	.w8(32'hbb466cdb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d84b5),
	.w1(32'hbb4983ce),
	.w2(32'hbae7671f),
	.w3(32'h3a588e6a),
	.w4(32'hba963d94),
	.w5(32'hbb825a71),
	.w6(32'h3ba674f9),
	.w7(32'h3a2c7cff),
	.w8(32'hba1fd572),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b97ace),
	.w1(32'h3ba297d4),
	.w2(32'h3c132bdd),
	.w3(32'h3b3090d4),
	.w4(32'h3bc117df),
	.w5(32'h3b45042b),
	.w6(32'h3bac1ad4),
	.w7(32'h3ad0d8af),
	.w8(32'h3b4db572),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd2f58),
	.w1(32'h3958965e),
	.w2(32'hbad7b9b3),
	.w3(32'hbb8d39ee),
	.w4(32'hb9df8499),
	.w5(32'hbb8908cf),
	.w6(32'hb88dd4e4),
	.w7(32'h3bba4f27),
	.w8(32'h3b908682),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69be8c),
	.w1(32'hbc32b361),
	.w2(32'hbb940e2e),
	.w3(32'hb7cca8f2),
	.w4(32'hbc76324e),
	.w5(32'hbc0a3d52),
	.w6(32'h3ba62240),
	.w7(32'hbc1566c2),
	.w8(32'hbb0f1b2b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7e0ae),
	.w1(32'h3b1bd39f),
	.w2(32'hbb222fcf),
	.w3(32'h3bacdf7f),
	.w4(32'hbb132863),
	.w5(32'hbc025692),
	.w6(32'h3b2143fa),
	.w7(32'hba559569),
	.w8(32'hb9650c01),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2c0c),
	.w1(32'h3af47edf),
	.w2(32'hbc301ed7),
	.w3(32'h3b878a3f),
	.w4(32'hbc57646a),
	.w5(32'h3b23ab58),
	.w6(32'h3bc27401),
	.w7(32'hbbc86b31),
	.w8(32'h3b8b5ec7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56964b),
	.w1(32'hbaeef3e6),
	.w2(32'hbbd71af6),
	.w3(32'h3af1bbcb),
	.w4(32'hbba91f30),
	.w5(32'hbc0d1cfb),
	.w6(32'h3b146898),
	.w7(32'hb9a03857),
	.w8(32'h3acdc745),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c8eac),
	.w1(32'hbba32385),
	.w2(32'hbbda3de3),
	.w3(32'h3c268c87),
	.w4(32'hbaa3b62c),
	.w5(32'hbbb30225),
	.w6(32'h3bb362c8),
	.w7(32'hbbcb1619),
	.w8(32'hbb98a337),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21998a),
	.w1(32'hbbd98748),
	.w2(32'hbc8e032a),
	.w3(32'h3bd93386),
	.w4(32'hbb752695),
	.w5(32'hbd0635eb),
	.w6(32'h3ba3fc60),
	.w7(32'hbaf11b68),
	.w8(32'h3a5d76b6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39877ee4),
	.w1(32'hbbd77f93),
	.w2(32'hb9f881cf),
	.w3(32'h3bc6cff1),
	.w4(32'hbb8341d1),
	.w5(32'hbb4a0e77),
	.w6(32'hbbf4daa9),
	.w7(32'hbb388058),
	.w8(32'hbb11dd0f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06644c),
	.w1(32'hbc308a91),
	.w2(32'hbc05f147),
	.w3(32'hb7ed6c6c),
	.w4(32'hbc0de159),
	.w5(32'hbc4be1b1),
	.w6(32'h3b4cda30),
	.w7(32'hbb1f40e1),
	.w8(32'h39ee5fc6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48ac4c),
	.w1(32'hbb4268a3),
	.w2(32'hbb12d6a7),
	.w3(32'h3c7a674d),
	.w4(32'h39f44dcd),
	.w5(32'hbb896a04),
	.w6(32'h3c561cf7),
	.w7(32'h3b97723d),
	.w8(32'hba8aab95),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18d91c),
	.w1(32'h3bf2cd13),
	.w2(32'h3c414844),
	.w3(32'hbb76544f),
	.w4(32'h3bc8defe),
	.w5(32'h3a9efcde),
	.w6(32'h3c026a70),
	.w7(32'hbb677e06),
	.w8(32'hba9671e7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e0e1c),
	.w1(32'h3ac5f4e1),
	.w2(32'hbb9ae728),
	.w3(32'hbb2d09d9),
	.w4(32'hb8e27e6b),
	.w5(32'hbbe2a702),
	.w6(32'h3bbaffc3),
	.w7(32'hbb854d2f),
	.w8(32'hbb97cae9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1acdf2),
	.w1(32'h3b1e5fef),
	.w2(32'hbb15f6be),
	.w3(32'h3ae82cfd),
	.w4(32'h3924d78e),
	.w5(32'h3b319f4c),
	.w6(32'hbb824fe7),
	.w7(32'hbb9a2f49),
	.w8(32'hba3300f4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b209),
	.w1(32'h3b559f49),
	.w2(32'h396af6cb),
	.w3(32'h3c2a3347),
	.w4(32'h3b501cce),
	.w5(32'hbaaba2a7),
	.w6(32'h3bd2a485),
	.w7(32'hba8d8738),
	.w8(32'hbbadddf2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc34f),
	.w1(32'h3b0d00c6),
	.w2(32'hbb9b2433),
	.w3(32'hbbdd7743),
	.w4(32'hbb73fa18),
	.w5(32'hbaaee1ef),
	.w6(32'hbba92c59),
	.w7(32'hbaf90a94),
	.w8(32'h3bc216ba),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd03a99),
	.w1(32'h3b804de0),
	.w2(32'h3b6c57e7),
	.w3(32'h3bb39368),
	.w4(32'h3bf93981),
	.w5(32'hbb0eb1fb),
	.w6(32'hb9dd6a67),
	.w7(32'h3958080f),
	.w8(32'hb98f270e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d4b2),
	.w1(32'hbb60e03d),
	.w2(32'hbb26f297),
	.w3(32'h3b6481b0),
	.w4(32'h3b075057),
	.w5(32'h3aec8e6d),
	.w6(32'hba196039),
	.w7(32'hbbe66c43),
	.w8(32'hbbadbb0f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0049b),
	.w1(32'hbab19a31),
	.w2(32'hbaaa7e6e),
	.w3(32'hbade4808),
	.w4(32'hbb385253),
	.w5(32'hbc47bec8),
	.w6(32'h39be334b),
	.w7(32'hbb8572f2),
	.w8(32'h3b993818),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39f13),
	.w1(32'hbbbce3b1),
	.w2(32'hbb641fe9),
	.w3(32'h3bde5497),
	.w4(32'hbb90dabb),
	.w5(32'hbaa29e70),
	.w6(32'h3b98c5c3),
	.w7(32'hbb2cb49a),
	.w8(32'h3b779585),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67c59c),
	.w1(32'h3b90a591),
	.w2(32'h3c1db522),
	.w3(32'h3c09cc57),
	.w4(32'h3bab0aff),
	.w5(32'h3b669cdd),
	.w6(32'h3ba0f16d),
	.w7(32'h3b08cbf0),
	.w8(32'h3bd5d4fe),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3efc47),
	.w1(32'hb9c38d45),
	.w2(32'hbbfe5922),
	.w3(32'hba71ef99),
	.w4(32'h3aa28ca1),
	.w5(32'hbb50c93e),
	.w6(32'hbbc9ec64),
	.w7(32'h3b8fd5eb),
	.w8(32'hbbd65975),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ddbed),
	.w1(32'hbab872d8),
	.w2(32'hbbe8b651),
	.w3(32'h3a7e8b99),
	.w4(32'hbbe90f27),
	.w5(32'hbb163e93),
	.w6(32'hbc414702),
	.w7(32'hbbad5913),
	.w8(32'hbbdb52f8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb4f9),
	.w1(32'hb9b11330),
	.w2(32'h3b0f2ff7),
	.w3(32'hbb8e1639),
	.w4(32'hb8a47376),
	.w5(32'hba8b06a3),
	.w6(32'hba22824c),
	.w7(32'hb9b716cf),
	.w8(32'h3a96ee7f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768113),
	.w1(32'hbb6b5bc1),
	.w2(32'h3a57e70b),
	.w3(32'h3bf8009e),
	.w4(32'hbbd9161a),
	.w5(32'hbc444497),
	.w6(32'h3c092bdf),
	.w7(32'hba739f55),
	.w8(32'hbb8ccfd7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88847),
	.w1(32'h3c07ee2f),
	.w2(32'h3b7771ad),
	.w3(32'hbbc7d816),
	.w4(32'h3b957579),
	.w5(32'h3a1f6c65),
	.w6(32'hbc1baad1),
	.w7(32'hbae9d779),
	.w8(32'h3b1af3a8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b598706),
	.w1(32'hbb93ee3e),
	.w2(32'hbb6b6b9c),
	.w3(32'h3c6e5547),
	.w4(32'hbc23b7b7),
	.w5(32'h3af2830c),
	.w6(32'h3c6372cd),
	.w7(32'hbb8b3eb8),
	.w8(32'hbbcdfcf3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404c3c),
	.w1(32'hbbb9b80e),
	.w2(32'hbb57d374),
	.w3(32'hbbf8c396),
	.w4(32'h3b5255a5),
	.w5(32'hbb5d0f65),
	.w6(32'h39929e33),
	.w7(32'hbbeb2e11),
	.w8(32'hbc1460c0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb47a6c),
	.w1(32'hbbaea8a2),
	.w2(32'hbc661de3),
	.w3(32'hbc131aed),
	.w4(32'hbb5b4876),
	.w5(32'hbc26d4ce),
	.w6(32'hbc10d003),
	.w7(32'h3b1149d0),
	.w8(32'h3bff4cfc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43c052),
	.w1(32'hbafd0af7),
	.w2(32'h3c11d6fa),
	.w3(32'h3bd431c6),
	.w4(32'h3b5c95ce),
	.w5(32'h3abd30bd),
	.w6(32'hbb80e2c4),
	.w7(32'hbbafdd8f),
	.w8(32'hbb555af8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27259),
	.w1(32'h3999f477),
	.w2(32'h3bbf6f2a),
	.w3(32'hbaafe666),
	.w4(32'hbae9536f),
	.w5(32'h3c6eaaf3),
	.w6(32'hbb371a6e),
	.w7(32'h3b47fc72),
	.w8(32'h3c5901cc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1ed94),
	.w1(32'hbc2b78bf),
	.w2(32'hbb83644a),
	.w3(32'h3c54335f),
	.w4(32'hbc4384e5),
	.w5(32'hbc1e36ba),
	.w6(32'h3bced9c6),
	.w7(32'hbbd01ccb),
	.w8(32'hbc11d17b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7093e),
	.w1(32'hba889273),
	.w2(32'hbb119db2),
	.w3(32'hba9a2437),
	.w4(32'h3addc20d),
	.w5(32'h3a89e951),
	.w6(32'hbabda095),
	.w7(32'h3a599078),
	.w8(32'hbb95d695),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab66776),
	.w1(32'hbb840cf6),
	.w2(32'hbaa772b4),
	.w3(32'h3c157e61),
	.w4(32'h3a75c038),
	.w5(32'h3aac5241),
	.w6(32'h3bcf1353),
	.w7(32'hba301bef),
	.w8(32'hb9d7b1cb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c5fdd),
	.w1(32'hbb569b9f),
	.w2(32'h3b24902f),
	.w3(32'h3ba81c8d),
	.w4(32'hb980bf62),
	.w5(32'hbc11be37),
	.w6(32'hbb393b41),
	.w7(32'h3bab670d),
	.w8(32'hbba8a096),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ccf3e),
	.w1(32'hbb473a78),
	.w2(32'h3c69960d),
	.w3(32'h3b2e39ec),
	.w4(32'hbbd690d6),
	.w5(32'h3c868063),
	.w6(32'h3be850ec),
	.w7(32'h3a9521b1),
	.w8(32'h3b16845c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15e00a),
	.w1(32'h3ac2efdd),
	.w2(32'h3acf18c0),
	.w3(32'hbc1af286),
	.w4(32'h3bc88342),
	.w5(32'hbb357660),
	.w6(32'hba05eeb1),
	.w7(32'h3acbd412),
	.w8(32'h3ba84d5e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78429e),
	.w1(32'h3b190eb9),
	.w2(32'hb8f735ff),
	.w3(32'h3c168fdf),
	.w4(32'h3b18d545),
	.w5(32'hbbb2fe51),
	.w6(32'h3c0877cc),
	.w7(32'h3b6726dd),
	.w8(32'h3b3b19d3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ca711),
	.w1(32'h3996dfb9),
	.w2(32'hbabbe3fa),
	.w3(32'h3b748c95),
	.w4(32'hbb882af9),
	.w5(32'hbbce0f28),
	.w6(32'h3b7950d3),
	.w7(32'hbb6ee020),
	.w8(32'hbaffba6d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb213eaa),
	.w1(32'hbb96c56c),
	.w2(32'hbb755d71),
	.w3(32'h3a2a7c59),
	.w4(32'hbb8c31a6),
	.w5(32'h3bdef9b7),
	.w6(32'h3b80054e),
	.w7(32'hba588383),
	.w8(32'hbacb7c39),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba542fd),
	.w1(32'hbb17e0ac),
	.w2(32'hbabb754f),
	.w3(32'hbb8a466b),
	.w4(32'hb9e3717b),
	.w5(32'hbbe8c9f5),
	.w6(32'hbac150ac),
	.w7(32'hbb66e858),
	.w8(32'h3b9e972a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98baa9),
	.w1(32'h3a031fe9),
	.w2(32'hbbb9c9e9),
	.w3(32'h3cd458ad),
	.w4(32'hbb1fe33e),
	.w5(32'hbbf69f24),
	.w6(32'h3c6ef0f7),
	.w7(32'hbb3b584d),
	.w8(32'hbb6d5133),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef1cda),
	.w1(32'hba25a3db),
	.w2(32'h3be4211f),
	.w3(32'h3ac92b00),
	.w4(32'h3b842364),
	.w5(32'hb91d74ef),
	.w6(32'h3c2385a9),
	.w7(32'hbb330f67),
	.w8(32'hbbadd318),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1724e4),
	.w1(32'h39a7f636),
	.w2(32'h3a666b9e),
	.w3(32'hb8d4de7d),
	.w4(32'hba20e147),
	.w5(32'hbb187ff1),
	.w6(32'h3a2c9c9d),
	.w7(32'hbb3d0e21),
	.w8(32'h3aad3e10),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb182298),
	.w1(32'h3b4b85af),
	.w2(32'h3bd6630c),
	.w3(32'hbc5d2848),
	.w4(32'h3ab0ea8c),
	.w5(32'h3b0f9a36),
	.w6(32'hbc079958),
	.w7(32'h3ace1225),
	.w8(32'hbaec6cf4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ad613),
	.w1(32'hbbc7c723),
	.w2(32'hbc20e334),
	.w3(32'hbb2f51a8),
	.w4(32'hbac292c0),
	.w5(32'hbc04b807),
	.w6(32'hbbc5a73e),
	.w7(32'hbb2863c7),
	.w8(32'hbbe51402),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf297b5),
	.w1(32'h3b340830),
	.w2(32'h3c2d63af),
	.w3(32'hbaea5994),
	.w4(32'h3a74ef0f),
	.w5(32'h3ba12ee3),
	.w6(32'hbb85b7e8),
	.w7(32'h3ae9ef42),
	.w8(32'h3ba7fa70),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab72d11),
	.w1(32'h3ba63742),
	.w2(32'h3c280104),
	.w3(32'h390f09a7),
	.w4(32'h3ae3e2e1),
	.w5(32'h3bb0805c),
	.w6(32'hbaf4f894),
	.w7(32'hbae867d0),
	.w8(32'hbab6338c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06b435),
	.w1(32'hbc515281),
	.w2(32'hbc3fcc1a),
	.w3(32'hbbd4a12b),
	.w4(32'hbc6a3217),
	.w5(32'h3ab727ab),
	.w6(32'hbaae667b),
	.w7(32'h3bb7d26d),
	.w8(32'h3c900dd0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd2cd4),
	.w1(32'hbb742b30),
	.w2(32'hbc34e76b),
	.w3(32'h3ca4961f),
	.w4(32'hbbcb06ef),
	.w5(32'hbc1e1494),
	.w6(32'h3c62f9d8),
	.w7(32'hbaa3d3a5),
	.w8(32'hbb7cd1f5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba910f1),
	.w1(32'hbb76bf10),
	.w2(32'hbab69902),
	.w3(32'hbbc73ef8),
	.w4(32'hbb7f6d97),
	.w5(32'h3bb68879),
	.w6(32'hbc0154af),
	.w7(32'h3c017f98),
	.w8(32'h3c3f57dc),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c668a50),
	.w1(32'h39d9395b),
	.w2(32'h3b983a9f),
	.w3(32'h3c0d3e23),
	.w4(32'h3afcf00c),
	.w5(32'h3ba0fa43),
	.w6(32'h3ab9894b),
	.w7(32'hbb10be22),
	.w8(32'hbaa75a23),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f57605),
	.w1(32'h3bb90d67),
	.w2(32'h3bc5ee0b),
	.w3(32'hbb171387),
	.w4(32'h3bc8c9a1),
	.w5(32'h3bf0b621),
	.w6(32'hbbe77ca1),
	.w7(32'hbace7c54),
	.w8(32'hbb5105c1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd538f2),
	.w1(32'h3956ae71),
	.w2(32'hba60c17d),
	.w3(32'hb9a3282b),
	.w4(32'hbb4383d3),
	.w5(32'hba7f2d85),
	.w6(32'hbc5feff3),
	.w7(32'h3ab68d89),
	.w8(32'hbb2419df),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb8b36),
	.w1(32'h3ada534e),
	.w2(32'h3b61dd4a),
	.w3(32'h3b7fc1f1),
	.w4(32'hba073b09),
	.w5(32'h3b4d7930),
	.w6(32'h3b21ddc1),
	.w7(32'hbab57eb3),
	.w8(32'h3bac4774),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c405259),
	.w1(32'h3bcb24f3),
	.w2(32'hba368092),
	.w3(32'h3c883a6f),
	.w4(32'hbac36dbd),
	.w5(32'h3a08206f),
	.w6(32'h3c09401a),
	.w7(32'h3a247361),
	.w8(32'h3b8f2b02),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d4ad3),
	.w1(32'h3bba2616),
	.w2(32'h3bedcf1a),
	.w3(32'h3b0eab76),
	.w4(32'hbb628acb),
	.w5(32'hbc15cb4e),
	.w6(32'hba8ed08b),
	.w7(32'h3bda3641),
	.w8(32'hbad10be9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb390aaa),
	.w1(32'h3b0b4420),
	.w2(32'hbb870588),
	.w3(32'hbc1d0810),
	.w4(32'h3bb3666f),
	.w5(32'hbbbc6737),
	.w6(32'h3b355c83),
	.w7(32'h3b223041),
	.w8(32'hbaf00a51),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ec56b),
	.w1(32'h3b09fe2f),
	.w2(32'h3bbf9db4),
	.w3(32'h3ab8969b),
	.w4(32'hbbbf67fd),
	.w5(32'h3c15c0b7),
	.w6(32'h3b8bbc5b),
	.w7(32'h3b908fc6),
	.w8(32'h3c67a1cc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8b54),
	.w1(32'hbc089f7d),
	.w2(32'hbb6687ed),
	.w3(32'h3cafa4d0),
	.w4(32'hbb0c528b),
	.w5(32'hba159e36),
	.w6(32'h3c562c06),
	.w7(32'h3aaa98bb),
	.w8(32'hba9c9bff),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb979b22),
	.w1(32'hbac9e500),
	.w2(32'hbc23a070),
	.w3(32'hbb82c4a2),
	.w4(32'hbb7469ee),
	.w5(32'hbc5fa154),
	.w6(32'h3b5c8be7),
	.w7(32'hbbbbca15),
	.w8(32'hbb3c540b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2d28d),
	.w1(32'hba5f15a9),
	.w2(32'hbbb708d3),
	.w3(32'hbb10e48d),
	.w4(32'hbbc3e09f),
	.w5(32'hbb42006b),
	.w6(32'hbb1223aa),
	.w7(32'hbbdf1be1),
	.w8(32'h3ac8f4c5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4226a),
	.w1(32'hbb95f5eb),
	.w2(32'h3c8bef8f),
	.w3(32'h3ae86b6a),
	.w4(32'h3c3ad860),
	.w5(32'h3ceedd56),
	.w6(32'h3b9ef049),
	.w7(32'hbb4ede51),
	.w8(32'h3b6722c7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b73a7),
	.w1(32'h3b9ddeb7),
	.w2(32'h3be1525c),
	.w3(32'hba07ec8c),
	.w4(32'h3c450a9a),
	.w5(32'h3beba701),
	.w6(32'hbbea5ea7),
	.w7(32'h3b8f18bd),
	.w8(32'hba9d69ed),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4d284),
	.w1(32'hbbd89110),
	.w2(32'hbb870187),
	.w3(32'h3b4e44cd),
	.w4(32'hbba05b11),
	.w5(32'hbb181c4f),
	.w6(32'hbba745bd),
	.w7(32'hb98273a8),
	.w8(32'h3b23a0a5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a99e9),
	.w1(32'hbb66ac92),
	.w2(32'hbbff2119),
	.w3(32'h3c23c7e8),
	.w4(32'hbb8b6446),
	.w5(32'hbc2dabdb),
	.w6(32'h3c35d1c5),
	.w7(32'hbc2b478b),
	.w8(32'hbc675679),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba77d9),
	.w1(32'hbba75032),
	.w2(32'hbb833d84),
	.w3(32'hba503c0a),
	.w4(32'hbb9aa4e7),
	.w5(32'h3c07bca6),
	.w6(32'h3a5e96e8),
	.w7(32'hbafe9795),
	.w8(32'h3c6a7a80),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba31719),
	.w1(32'h35f7b6c1),
	.w2(32'hba62bf59),
	.w3(32'h3c1b40b1),
	.w4(32'h3b073714),
	.w5(32'hba8df312),
	.w6(32'hbb517759),
	.w7(32'h3bc1cfa3),
	.w8(32'h3b108103),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f660),
	.w1(32'h3a95b82d),
	.w2(32'h3ad8ecfb),
	.w3(32'hbb481012),
	.w4(32'h3a3b40d5),
	.w5(32'hbc284f0b),
	.w6(32'hbba0dceb),
	.w7(32'hb9db4ffb),
	.w8(32'hbb0aa203),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d2bdd),
	.w1(32'hbb142562),
	.w2(32'hbb77d7ac),
	.w3(32'h3bb1e64b),
	.w4(32'hbb10f002),
	.w5(32'hb84580b0),
	.w6(32'h3aabd2a6),
	.w7(32'h3a87bb2a),
	.w8(32'h3c3637c2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c320714),
	.w1(32'h3b0a0f62),
	.w2(32'h3c0aee86),
	.w3(32'h3c9475a0),
	.w4(32'h3bfdda64),
	.w5(32'h3ab9dff6),
	.w6(32'h3c08872a),
	.w7(32'hbac8c033),
	.w8(32'hbac28cf9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe468b9),
	.w1(32'h3b6bf21f),
	.w2(32'hbba9e63f),
	.w3(32'hbc417cfb),
	.w4(32'h3be13130),
	.w5(32'hbc78c794),
	.w6(32'hbb234746),
	.w7(32'hbbada60b),
	.w8(32'hbc7e5b0a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08b1fe),
	.w1(32'hbae6a189),
	.w2(32'hbb0859c1),
	.w3(32'h3a5338df),
	.w4(32'hbbb91af1),
	.w5(32'hbc253aa2),
	.w6(32'h3b0ba7c5),
	.w7(32'hbb29e9bf),
	.w8(32'hbbbe890d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c7d83),
	.w1(32'hb91c31dc),
	.w2(32'h3b9419ba),
	.w3(32'hbc187132),
	.w4(32'h38fd2c9c),
	.w5(32'hbb512aa0),
	.w6(32'h3a957423),
	.w7(32'hbb8430b5),
	.w8(32'h3bbdd591),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c642931),
	.w1(32'h3bdaebd0),
	.w2(32'h3b0b7fee),
	.w3(32'h3cbaded3),
	.w4(32'h3b8644f3),
	.w5(32'hbb51871b),
	.w6(32'h3c0b6256),
	.w7(32'h3b709124),
	.w8(32'hbc1e8415),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeab81),
	.w1(32'hbbc38928),
	.w2(32'h3a576e24),
	.w3(32'hbc0b129c),
	.w4(32'hbbfa64ba),
	.w5(32'hbbc0d507),
	.w6(32'hbc2159ba),
	.w7(32'hbb2acdf4),
	.w8(32'hbb238923),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389023e6),
	.w1(32'hbb6e19e1),
	.w2(32'hbbcded2b),
	.w3(32'hbb7a7349),
	.w4(32'hbc09b1c3),
	.w5(32'hbbdd01b0),
	.w6(32'hbade2061),
	.w7(32'hbb20ab9b),
	.w8(32'h3b88caeb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc820a0b),
	.w1(32'hbbbc36eb),
	.w2(32'h3909d306),
	.w3(32'hbc1de120),
	.w4(32'hba8a819b),
	.w5(32'hbb54988f),
	.w6(32'hb9863ce4),
	.w7(32'hbb9af7e5),
	.w8(32'h3ba82514),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77775a),
	.w1(32'hbb374c19),
	.w2(32'hbbca807f),
	.w3(32'hbaee260c),
	.w4(32'hbbb95b44),
	.w5(32'hbb2388c7),
	.w6(32'h3ace633f),
	.w7(32'hbb0bb926),
	.w8(32'hbbd8e7fb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47d561),
	.w1(32'hbb19cd23),
	.w2(32'h3b4c7d74),
	.w3(32'hbb5f9378),
	.w4(32'hbb284b45),
	.w5(32'hbbbd9d19),
	.w6(32'hb9f09353),
	.w7(32'hbb779917),
	.w8(32'hbba26ee0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc7d20),
	.w1(32'hbb7f6721),
	.w2(32'hbb80d083),
	.w3(32'hbc074f56),
	.w4(32'hbac4d757),
	.w5(32'hbbd1cd3f),
	.w6(32'hbb9a27cc),
	.w7(32'h3bb60ffe),
	.w8(32'hbadfdbaf),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db830),
	.w1(32'hbb407e57),
	.w2(32'hbacf845b),
	.w3(32'hbc353366),
	.w4(32'hbb23f939),
	.w5(32'hbc3c0ba2),
	.w6(32'hbc0387d2),
	.w7(32'h3a2800a1),
	.w8(32'hbb94e992),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb798efd),
	.w1(32'h397995e1),
	.w2(32'hbbbd90df),
	.w3(32'h3b083efc),
	.w4(32'hbad14623),
	.w5(32'hbc5b8a37),
	.w6(32'hba625e3e),
	.w7(32'hbae30595),
	.w8(32'h3b6db14b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26269b),
	.w1(32'hbb905625),
	.w2(32'hbbef801c),
	.w3(32'h3b2eb182),
	.w4(32'hbb97c17c),
	.w5(32'hbb258417),
	.w6(32'h3c1bc1d8),
	.w7(32'hbbce570e),
	.w8(32'h3a805453),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3104a),
	.w1(32'hba844340),
	.w2(32'hbbc7a201),
	.w3(32'h3b04bda7),
	.w4(32'hba472c07),
	.w5(32'hbb03a2e9),
	.w6(32'h3bc29011),
	.w7(32'hbb338b63),
	.w8(32'hbb71be9d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d293),
	.w1(32'hbc1e8122),
	.w2(32'hbbc8e3bb),
	.w3(32'hba88fce4),
	.w4(32'hbbf15b03),
	.w5(32'h3b1984dc),
	.w6(32'h3b300778),
	.w7(32'hbb2a1bda),
	.w8(32'h3aacdf58),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13356c),
	.w1(32'h399d3909),
	.w2(32'hb9a8f83b),
	.w3(32'h3b42312e),
	.w4(32'h3b533eca),
	.w5(32'h399667ba),
	.w6(32'hbb234f5a),
	.w7(32'hb93364d7),
	.w8(32'hbbbae79b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d4bdb),
	.w1(32'hbb1091aa),
	.w2(32'hbb3ba7d8),
	.w3(32'hba36206e),
	.w4(32'h3b479bcc),
	.w5(32'h3a40a0c1),
	.w6(32'h3a2b453a),
	.w7(32'h3b9a69c4),
	.w8(32'hb7840a46),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23bb77),
	.w1(32'hbc1b79bc),
	.w2(32'hbc53588a),
	.w3(32'hbb56451c),
	.w4(32'hbc4d883c),
	.w5(32'hbba6d160),
	.w6(32'h3b7dca51),
	.w7(32'hbb81e657),
	.w8(32'h3a349ea1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ad83),
	.w1(32'hba9193c9),
	.w2(32'hbbbe6134),
	.w3(32'hbb8d79fa),
	.w4(32'h3a181b4e),
	.w5(32'hbc6f0b1c),
	.w6(32'h3bdc6749),
	.w7(32'hb81b14e2),
	.w8(32'hbb6ebc99),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080d64),
	.w1(32'h3a8b6540),
	.w2(32'hbb2160ea),
	.w3(32'hbc0e9081),
	.w4(32'hbc133cee),
	.w5(32'hbb13e08c),
	.w6(32'h3a1bf913),
	.w7(32'h39da4097),
	.w8(32'h3b7f2d2c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f602),
	.w1(32'hbab1a00a),
	.w2(32'h3b5fe41f),
	.w3(32'hbade278e),
	.w4(32'hbbd7294a),
	.w5(32'hbaf724c3),
	.w6(32'hbadf590f),
	.w7(32'hbb9183de),
	.w8(32'hbb86d879),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ec395),
	.w1(32'h3b1894ce),
	.w2(32'hb9d5c4ee),
	.w3(32'h3afa194e),
	.w4(32'hbadc66cb),
	.w5(32'hbb892d59),
	.w6(32'h3acff757),
	.w7(32'hbb2bbaac),
	.w8(32'hbb8d1baa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5fddb),
	.w1(32'hbbbcb437),
	.w2(32'hbae0fff4),
	.w3(32'h3a8c4ea3),
	.w4(32'hbbc49080),
	.w5(32'hbc158f76),
	.w6(32'hbad59ae7),
	.w7(32'h3b038144),
	.w8(32'hbb5a343e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81248),
	.w1(32'h3b279d1f),
	.w2(32'h3bb14dde),
	.w3(32'h3a58676c),
	.w4(32'hbb188b27),
	.w5(32'h3c4edf61),
	.w6(32'h3bc3a9a5),
	.w7(32'hbb8e8f21),
	.w8(32'h3be92da7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b573428),
	.w1(32'hbb113606),
	.w2(32'h3b1310cf),
	.w3(32'h3b9b7331),
	.w4(32'hbb4a92e2),
	.w5(32'hbb489090),
	.w6(32'h3b3632bf),
	.w7(32'hbbe0adae),
	.w8(32'hb9096630),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba996fb2),
	.w1(32'hba31bc59),
	.w2(32'h39de43d2),
	.w3(32'hbbcaa0c1),
	.w4(32'hbb5b1936),
	.w5(32'hb9e5a3ab),
	.w6(32'hbb24da93),
	.w7(32'hbb5f515d),
	.w8(32'h3af8a211),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d931e),
	.w1(32'h3acb91bc),
	.w2(32'h3af03299),
	.w3(32'hba421d2a),
	.w4(32'h3b14275e),
	.w5(32'h3bb84e48),
	.w6(32'hbaf7b152),
	.w7(32'h3924ae9a),
	.w8(32'h3c029329),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8333bb),
	.w1(32'hbb261af0),
	.w2(32'hbbb8e4bf),
	.w3(32'hb9942699),
	.w4(32'h39b9938f),
	.w5(32'hbbad1180),
	.w6(32'h3b0988bd),
	.w7(32'h3ac8c984),
	.w8(32'hb9d5795c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8baa9b),
	.w1(32'h3b96f25c),
	.w2(32'hbc2ab233),
	.w3(32'h3b5d36af),
	.w4(32'hbc558ce6),
	.w5(32'h3c94c79c),
	.w6(32'hbaee49a5),
	.w7(32'hbc367015),
	.w8(32'h3c387514),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb471f42),
	.w1(32'h3bb23cee),
	.w2(32'hbbd12aa9),
	.w3(32'hbc5b947d),
	.w4(32'hb7d5202b),
	.w5(32'h3bc81ef1),
	.w6(32'hbbcb95ff),
	.w7(32'hb98ea441),
	.w8(32'h3bab3484),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffe80f),
	.w1(32'h3b4151af),
	.w2(32'hbc0bbb89),
	.w3(32'hbb006d98),
	.w4(32'hbad39bc8),
	.w5(32'hbc06b6a2),
	.w6(32'h395cd486),
	.w7(32'hbb3ae8e9),
	.w8(32'h3b85dc87),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf33db0),
	.w1(32'hbaeb900a),
	.w2(32'h3c36a7b7),
	.w3(32'hbb6a9016),
	.w4(32'h3a5bbaae),
	.w5(32'h3b1b7369),
	.w6(32'hba5f9cf2),
	.w7(32'h3b8cc5b5),
	.w8(32'hbb3412f7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bead648),
	.w1(32'h3a99c771),
	.w2(32'h3ae2f2cc),
	.w3(32'h3b57c2fd),
	.w4(32'hbb34b30d),
	.w5(32'h3b0097c6),
	.w6(32'h3bae5afb),
	.w7(32'hbb15a213),
	.w8(32'hbb0f016a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a822954),
	.w1(32'hbb3c0539),
	.w2(32'h3b371d41),
	.w3(32'h3b33be05),
	.w4(32'hba9972a7),
	.w5(32'hbb7f1a5e),
	.w6(32'h3aea367f),
	.w7(32'hb9822ec1),
	.w8(32'hbc09ff21),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956b591),
	.w1(32'hb9b9bbcd),
	.w2(32'h3bc17603),
	.w3(32'hb9cb3edc),
	.w4(32'h3b0a1ad3),
	.w5(32'h3bf34dd8),
	.w6(32'h3b7b4c7e),
	.w7(32'h3b88ec87),
	.w8(32'h3b620e52),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44655c),
	.w1(32'hbb1d8c74),
	.w2(32'h3a6712ce),
	.w3(32'hba53cae8),
	.w4(32'hbb204ab2),
	.w5(32'h3924119f),
	.w6(32'h3a375e6c),
	.w7(32'hba16021c),
	.w8(32'hb9c62c26),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63c7ee),
	.w1(32'hbb2aa103),
	.w2(32'h3b09909f),
	.w3(32'hbab64146),
	.w4(32'hba360449),
	.w5(32'hbad9adf5),
	.w6(32'hbb402a94),
	.w7(32'h3b4f02d3),
	.w8(32'h3b9cac0e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c5ccb),
	.w1(32'h3c0ca5ff),
	.w2(32'hbbd75a68),
	.w3(32'h3aaba6ea),
	.w4(32'h3a33ae01),
	.w5(32'h3c2f3cbb),
	.w6(32'hba3ce4f0),
	.w7(32'hbb9f4c0f),
	.w8(32'h3c69792b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9469b78),
	.w1(32'h3bc9e019),
	.w2(32'hbb7f6a67),
	.w3(32'hbc0c1bab),
	.w4(32'h3ab06f5a),
	.w5(32'h3bb19f91),
	.w6(32'hbafa1bb6),
	.w7(32'hbc104252),
	.w8(32'h3c48bb57),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69e60a),
	.w1(32'hbb9ee29c),
	.w2(32'h3b0a026c),
	.w3(32'hbc2a0079),
	.w4(32'hba9e3ad8),
	.w5(32'hba60ef92),
	.w6(32'hb8d606e4),
	.w7(32'h3babca3f),
	.w8(32'h39490998),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c30e),
	.w1(32'h3bdee599),
	.w2(32'hbbbc8ef8),
	.w3(32'h3ab9e18c),
	.w4(32'h3be7945b),
	.w5(32'h3c0361b8),
	.w6(32'h3b8c493b),
	.w7(32'hbb0f4632),
	.w8(32'h3c1cad2b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98c18a),
	.w1(32'hbb0ff01a),
	.w2(32'h3ae239b4),
	.w3(32'h386d8034),
	.w4(32'hbbad13ba),
	.w5(32'hba215767),
	.w6(32'hba9fa8b9),
	.w7(32'hbbb586fb),
	.w8(32'hbb47c938),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf347b),
	.w1(32'hbb4d654b),
	.w2(32'h3a922f8a),
	.w3(32'hbaecd59c),
	.w4(32'h3ba447f8),
	.w5(32'hbb258c2d),
	.w6(32'hbab323fe),
	.w7(32'h3b77c1ed),
	.w8(32'h3a9967b2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d16bc),
	.w1(32'hbb4a6ebc),
	.w2(32'h3c15308b),
	.w3(32'hbabe3467),
	.w4(32'h3b570f2b),
	.w5(32'h3a108120),
	.w6(32'hba6e381b),
	.w7(32'h3b898cce),
	.w8(32'hbba8f7c4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc52a),
	.w1(32'hbacf7c52),
	.w2(32'h3bcbb4cd),
	.w3(32'h3c02fef0),
	.w4(32'hb9617a6e),
	.w5(32'h3bab7af0),
	.w6(32'h3b675279),
	.w7(32'h3a95595e),
	.w8(32'h3b384c4c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab485f6),
	.w1(32'h3aa3dd01),
	.w2(32'hba9db53a),
	.w3(32'hba3ce7be),
	.w4(32'h3aa5f893),
	.w5(32'hba20471b),
	.w6(32'h3b3bfb8a),
	.w7(32'h39658f85),
	.w8(32'h3b31a9f2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17f1dd),
	.w1(32'hbba12410),
	.w2(32'hbbbe7419),
	.w3(32'hbb7145a6),
	.w4(32'hb8c3e604),
	.w5(32'hbb9f6062),
	.w6(32'hba9e7225),
	.w7(32'hbb941df4),
	.w8(32'hbab680cb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25e9fd),
	.w1(32'hbb0943d4),
	.w2(32'hbbc7fb5d),
	.w3(32'h3a59b9eb),
	.w4(32'hbbb99297),
	.w5(32'hbbb55c24),
	.w6(32'hbb4564f5),
	.w7(32'hbbabd082),
	.w8(32'hbad61b5f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc41e),
	.w1(32'h3baa53bf),
	.w2(32'hbbc63628),
	.w3(32'hbc16906d),
	.w4(32'h3bbb6b60),
	.w5(32'h3b83649e),
	.w6(32'hbb08b8f0),
	.w7(32'h3b2749fe),
	.w8(32'h3c2b91b1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb224079),
	.w1(32'hbb391b3e),
	.w2(32'hbb5fe646),
	.w3(32'hbb8ba77b),
	.w4(32'hbbaf4bf4),
	.w5(32'hbb7516f7),
	.w6(32'hbb908afb),
	.w7(32'hbb250ae3),
	.w8(32'hbb536455),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb3586),
	.w1(32'h3aa09148),
	.w2(32'hbc00cd72),
	.w3(32'hbab3e9ca),
	.w4(32'h390e8f0b),
	.w5(32'h3b0c4f87),
	.w6(32'hbade6097),
	.w7(32'hbacd4978),
	.w8(32'hba5b4d7f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde395f),
	.w1(32'h3b7b94ca),
	.w2(32'hbb010dd3),
	.w3(32'h3931ecb6),
	.w4(32'hba29abfb),
	.w5(32'hbbee1ee0),
	.w6(32'hbb81790b),
	.w7(32'hbb56153b),
	.w8(32'hbb464b7d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafac9b),
	.w1(32'hbbc6d3da),
	.w2(32'hbb263c27),
	.w3(32'hbbd0cbdc),
	.w4(32'hbaa27d6c),
	.w5(32'h3a240b12),
	.w6(32'hbbd1891f),
	.w7(32'h3ab5db61),
	.w8(32'hba927aec),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b65a11),
	.w1(32'hbb1fbf22),
	.w2(32'hbbcc35ad),
	.w3(32'hbaaf43d5),
	.w4(32'hbb0644a7),
	.w5(32'hbbaef6e9),
	.w6(32'hbb897998),
	.w7(32'hbb3dae8c),
	.w8(32'hba22ffed),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42aa8f),
	.w1(32'hb747539a),
	.w2(32'hbb0a2956),
	.w3(32'hbc0017f1),
	.w4(32'hba4eb744),
	.w5(32'h3badea66),
	.w6(32'hbb21273b),
	.w7(32'hbb20d459),
	.w8(32'h397a1f10),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d6907),
	.w1(32'hbaff7e6b),
	.w2(32'h3b9991c7),
	.w3(32'hba0c01d2),
	.w4(32'h3b855670),
	.w5(32'hbc06553c),
	.w6(32'hbb2bc6bf),
	.w7(32'h3bfdcf8f),
	.w8(32'hbb03d2d7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082465),
	.w1(32'hb96c1d9f),
	.w2(32'h3b35ccc9),
	.w3(32'h3bae2833),
	.w4(32'hbb4eafc6),
	.w5(32'h3b1335c3),
	.w6(32'h3b14b9d5),
	.w7(32'h38379d23),
	.w8(32'h3af15737),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c8389),
	.w1(32'h3c3a6e12),
	.w2(32'hbb92662e),
	.w3(32'h3bce66b9),
	.w4(32'h3c47245b),
	.w5(32'h3a9dfd58),
	.w6(32'h3b6dcba2),
	.w7(32'h3accbcb8),
	.w8(32'hb9974cd2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f4ab),
	.w1(32'hbbfcaa3c),
	.w2(32'hba48f83e),
	.w3(32'hb937507c),
	.w4(32'hbbe15791),
	.w5(32'hbbae7cdf),
	.w6(32'h3acc45e7),
	.w7(32'hba7385a6),
	.w8(32'hbc00cfdd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04d2fc),
	.w1(32'hbbc39050),
	.w2(32'h3bb4b32c),
	.w3(32'hbb1bffbf),
	.w4(32'h3bcce5ff),
	.w5(32'hbba96ee9),
	.w6(32'h3a473ac4),
	.w7(32'h3be076c1),
	.w8(32'hbb0a769b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cbc7a),
	.w1(32'hbc14437c),
	.w2(32'h3b7cb014),
	.w3(32'h3bbaff9b),
	.w4(32'h3b03b7e9),
	.w5(32'hbaa165ce),
	.w6(32'hbba27cc7),
	.w7(32'h3b8ea454),
	.w8(32'h3a11e0c6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14783d),
	.w1(32'hb9fec82f),
	.w2(32'h39fa66cd),
	.w3(32'h3b9d9857),
	.w4(32'hba4fea38),
	.w5(32'hbb7b4f96),
	.w6(32'h3931feb0),
	.w7(32'h3aca9f53),
	.w8(32'hbaf16d73),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227ca6),
	.w1(32'hbadb56ac),
	.w2(32'hbb0da101),
	.w3(32'h3b25acce),
	.w4(32'hbb93b0ee),
	.w5(32'hbb4079c1),
	.w6(32'h3b62fa5c),
	.w7(32'hbb0d1ddd),
	.w8(32'hbb0878f2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa42206),
	.w1(32'h3b03329c),
	.w2(32'h3b66588c),
	.w3(32'hbb816ac1),
	.w4(32'hb8aedb89),
	.w5(32'h3a62af5f),
	.w6(32'hba877669),
	.w7(32'hbbd4ac9c),
	.w8(32'h3b4ae853),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc5831),
	.w1(32'hbbc31e2c),
	.w2(32'h3c17b8cd),
	.w3(32'hbb9a4fb5),
	.w4(32'hbac0cecc),
	.w5(32'h3bec469d),
	.w6(32'hbb11a2b8),
	.w7(32'hba7c19f1),
	.w8(32'hbb5b39ed),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaedbaa),
	.w1(32'hba9a4d9f),
	.w2(32'h3a3d1f7b),
	.w3(32'hbac236be),
	.w4(32'h3a62b00d),
	.w5(32'h3b9bd246),
	.w6(32'hbb907193),
	.w7(32'hbb5a17fb),
	.w8(32'h3b749c6d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3529),
	.w1(32'hba33e630),
	.w2(32'h3b503558),
	.w3(32'h3acf9f0c),
	.w4(32'hbc0acfc3),
	.w5(32'h3b3aff25),
	.w6(32'h3b0efd86),
	.w7(32'hbbf66d85),
	.w8(32'hbb7e1793),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5922),
	.w1(32'hba912d71),
	.w2(32'h3af0cdcc),
	.w3(32'hb9c95e12),
	.w4(32'h3b5b8dd2),
	.w5(32'h3ba3b910),
	.w6(32'hba08982d),
	.w7(32'hbb1c56e4),
	.w8(32'h3b339b7b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a74ff),
	.w1(32'hbbaa0229),
	.w2(32'h3b62f046),
	.w3(32'h3afbcf96),
	.w4(32'hbb3985fb),
	.w5(32'hbb4fccd8),
	.w6(32'h3a90f0db),
	.w7(32'h3a947178),
	.w8(32'hbbc5e2db),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc11c9d),
	.w1(32'h3b94f247),
	.w2(32'hbb9b9f79),
	.w3(32'h3bbf3729),
	.w4(32'hba9f5353),
	.w5(32'hbb1dec70),
	.w6(32'h3b3bbf3f),
	.w7(32'hbc423868),
	.w8(32'h3bfc7db7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6ffcf),
	.w1(32'h3b8fbb6c),
	.w2(32'h3b890531),
	.w3(32'hbc25704f),
	.w4(32'hba1bb75d),
	.w5(32'h3c89473d),
	.w6(32'hbb1d9a54),
	.w7(32'hbb3aee05),
	.w8(32'h3c183297),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d9f1),
	.w1(32'hba4dd389),
	.w2(32'h3b442925),
	.w3(32'hbbe8ea91),
	.w4(32'h3b85b24f),
	.w5(32'h3a87c41d),
	.w6(32'h3b8e289c),
	.w7(32'h3b7e8277),
	.w8(32'hbbbaa962),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e33cb1),
	.w1(32'h3aba0a56),
	.w2(32'h3b1e9c12),
	.w3(32'hb923e170),
	.w4(32'h3aab8bea),
	.w5(32'hbb4b35ab),
	.w6(32'h3af2797e),
	.w7(32'h3b08a987),
	.w8(32'hba324eed),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b197f74),
	.w1(32'hb97ce0dd),
	.w2(32'hbb7f4c90),
	.w3(32'h3bb9b5f2),
	.w4(32'hba2e0dbf),
	.w5(32'hbbb0cfa2),
	.w6(32'hbb488d19),
	.w7(32'h3a0f360e),
	.w8(32'hbaa66568),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4031cf),
	.w1(32'hbbc12918),
	.w2(32'hbab58f06),
	.w3(32'hbbadd163),
	.w4(32'hba6d409b),
	.w5(32'hbc0107a4),
	.w6(32'hbb2f527e),
	.w7(32'h3b9379a1),
	.w8(32'hbb81033a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc27a8a),
	.w1(32'hbbb538f7),
	.w2(32'h3c1055a2),
	.w3(32'h3b9e4e8e),
	.w4(32'h39962ebe),
	.w5(32'hbb740382),
	.w6(32'hb8a743f3),
	.w7(32'h3c1162ec),
	.w8(32'hba4a2938),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb874),
	.w1(32'hbbc52516),
	.w2(32'hbaa019d6),
	.w3(32'h3b88b5ca),
	.w4(32'hbbf748de),
	.w5(32'hbc09f2f4),
	.w6(32'h3acc471c),
	.w7(32'hba595c8b),
	.w8(32'hbc03ed1a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce886a),
	.w1(32'h3a062c20),
	.w2(32'hb9594761),
	.w3(32'hbb4e63e6),
	.w4(32'hbbff7e4c),
	.w5(32'hbbb76775),
	.w6(32'hbac82923),
	.w7(32'hba506544),
	.w8(32'h3aa02e79),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02126f),
	.w1(32'hb9947df3),
	.w2(32'h3b929a77),
	.w3(32'hbaf9b488),
	.w4(32'h3b38a1e9),
	.w5(32'hba13e45b),
	.w6(32'hbbb30a90),
	.w7(32'h3ab2f0bf),
	.w8(32'h392967e4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule