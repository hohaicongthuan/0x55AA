module layer_8_featuremap_249(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec5613),
	.w1(32'h3b65fdbd),
	.w2(32'h3b3e9566),
	.w3(32'hbb8acee9),
	.w4(32'h3a133465),
	.w5(32'hbbb2eba8),
	.w6(32'hb96d242b),
	.w7(32'hba63b4ff),
	.w8(32'hba8b8c61),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb691d82),
	.w1(32'hbbb4d2bc),
	.w2(32'hbc2f21c3),
	.w3(32'hbbe96cc4),
	.w4(32'h3b47b862),
	.w5(32'hbafc8c37),
	.w6(32'h3b8f0e52),
	.w7(32'hba4c9e13),
	.w8(32'h3bfcd3ce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ac1c9),
	.w1(32'hb7965f30),
	.w2(32'h3b762d1e),
	.w3(32'h3c10c3f4),
	.w4(32'h3ba3a193),
	.w5(32'h3b934e2b),
	.w6(32'hbb4d756d),
	.w7(32'h3a230e21),
	.w8(32'h3bb1213b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4095c),
	.w1(32'hbbdf75e2),
	.w2(32'hbb26213b),
	.w3(32'h3c07c9dd),
	.w4(32'h3b8f05ee),
	.w5(32'h3a9d8ba4),
	.w6(32'hbb8ffc14),
	.w7(32'h3b477e1a),
	.w8(32'h3c0c74f1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c1fe3),
	.w1(32'hbc430313),
	.w2(32'hbd19b46a),
	.w3(32'h39a5f3c6),
	.w4(32'hbbac2ae9),
	.w5(32'hbcd5fdd6),
	.w6(32'h3bf89758),
	.w7(32'hbb22798a),
	.w8(32'h3c2e8110),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc861566),
	.w1(32'hba4c12c3),
	.w2(32'h3b2b6090),
	.w3(32'hbbb0f3c3),
	.w4(32'hba83d671),
	.w5(32'hbb766aaa),
	.w6(32'h3afbaf83),
	.w7(32'h3bfaee6f),
	.w8(32'h3a9b4a85),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b7b6d),
	.w1(32'h3ae957f3),
	.w2(32'hbbb58a84),
	.w3(32'hbc25efc8),
	.w4(32'hbb28bfcd),
	.w5(32'hbbcf140e),
	.w6(32'h380e5f94),
	.w7(32'hba8555b5),
	.w8(32'hbbb5229d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcecd82),
	.w1(32'h3babd627),
	.w2(32'hbbdd1f33),
	.w3(32'hbc36af79),
	.w4(32'hbb081879),
	.w5(32'hbc4a96e7),
	.w6(32'h3c105c12),
	.w7(32'h3c3c3f2e),
	.w8(32'h3c214264),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb7524),
	.w1(32'hbc72e084),
	.w2(32'hbd60e298),
	.w3(32'hbbf88b18),
	.w4(32'hbbc9a881),
	.w5(32'hbd35cb88),
	.w6(32'h3c9425dd),
	.w7(32'hbb8f59c8),
	.w8(32'h3c01aaa6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ce59c),
	.w1(32'h3c8a7f9c),
	.w2(32'h3b1b2c1f),
	.w3(32'hbcafb2b5),
	.w4(32'h3c09225a),
	.w5(32'h3b800eeb),
	.w6(32'h3bcfdd40),
	.w7(32'h3b9bd7fa),
	.w8(32'h3a56fdbc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba597775),
	.w1(32'hbb07fa95),
	.w2(32'hbc97e891),
	.w3(32'h3a9f9c8f),
	.w4(32'hba8ea7ba),
	.w5(32'hbc7f22b5),
	.w6(32'h3b8f4f32),
	.w7(32'h3a833e55),
	.w8(32'h3bffaaa4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e59ad),
	.w1(32'hbb8cc12e),
	.w2(32'hbc5b5a6e),
	.w3(32'hbc87753e),
	.w4(32'hbbe112fc),
	.w5(32'hbc16e5a6),
	.w6(32'hbb2f2bc9),
	.w7(32'hbbd42530),
	.w8(32'hbbb2c041),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d14f),
	.w1(32'h3b21017a),
	.w2(32'h3b8472ed),
	.w3(32'hbbef22ad),
	.w4(32'h3bbc652e),
	.w5(32'h3b326dda),
	.w6(32'h3bbf7cd9),
	.w7(32'h3b8f6908),
	.w8(32'h3a93a451),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedad5f),
	.w1(32'h3b096c85),
	.w2(32'h3be0a061),
	.w3(32'hba2b1273),
	.w4(32'h3baebbe6),
	.w5(32'h3c14d710),
	.w6(32'hbb05dcee),
	.w7(32'h3ae60442),
	.w8(32'h3aba977e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1881d9),
	.w1(32'h3cf18f03),
	.w2(32'h3d7c1a60),
	.w3(32'h3aa0df43),
	.w4(32'h3c92bea2),
	.w5(32'h3d3fd3b0),
	.w6(32'h3c5b84f2),
	.w7(32'h3cd7835b),
	.w8(32'h3c6b0931),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d23b7f2),
	.w1(32'h3b882e89),
	.w2(32'hbbb9ab8c),
	.w3(32'h3cc80eed),
	.w4(32'h3ab98e75),
	.w5(32'hbc1f54b0),
	.w6(32'h3b7122ed),
	.w7(32'hbbb2fa46),
	.w8(32'hbb887664),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54b16d),
	.w1(32'hbb604f9c),
	.w2(32'hbc10c46d),
	.w3(32'hbc0d2928),
	.w4(32'hbb7ce3f1),
	.w5(32'hbb68de48),
	.w6(32'hbb034fc6),
	.w7(32'h3b6cd7e2),
	.w8(32'h3960105b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc14ecc),
	.w1(32'h3b6e5934),
	.w2(32'h3c297d94),
	.w3(32'hbc51deb7),
	.w4(32'h3ad7a353),
	.w5(32'h3bd058bd),
	.w6(32'h3a21316e),
	.w7(32'h3b0d6f25),
	.w8(32'h3baa1742),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbbf87),
	.w1(32'h3c0a7270),
	.w2(32'hbc842e1c),
	.w3(32'h3bfb66c7),
	.w4(32'h3b2f38ac),
	.w5(32'hbca2b829),
	.w6(32'h3a52a409),
	.w7(32'hbb60faeb),
	.w8(32'hbb05ae3f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e984),
	.w1(32'h3c62bca5),
	.w2(32'h3c49b846),
	.w3(32'hbc4b5930),
	.w4(32'h3b344dda),
	.w5(32'h3b03948a),
	.w6(32'h3b805859),
	.w7(32'h3bf9f82d),
	.w8(32'hbb459623),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23bd66),
	.w1(32'h3b8da27e),
	.w2(32'h3ba1ab47),
	.w3(32'hbc328713),
	.w4(32'h3c350afb),
	.w5(32'h3ca5d4a5),
	.w6(32'h3b5e826a),
	.w7(32'h3b3541f1),
	.w8(32'h3a304a62),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad36ee),
	.w1(32'h3b6fa32c),
	.w2(32'h3b38638a),
	.w3(32'h3bff7dfe),
	.w4(32'h3a03d01d),
	.w5(32'hbb223c9b),
	.w6(32'h3bd2d348),
	.w7(32'h3a792a88),
	.w8(32'h3b09aa9d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b728dbd),
	.w1(32'h3ca8ba49),
	.w2(32'h3a904f54),
	.w3(32'h3bf8e428),
	.w4(32'h3bc839d6),
	.w5(32'hbb844461),
	.w6(32'h3c2e9bab),
	.w7(32'h3bce8324),
	.w8(32'h3c06dcac),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ba2bf),
	.w1(32'h3bd509ae),
	.w2(32'h3b4f5d94),
	.w3(32'h3b272891),
	.w4(32'h3b9da5ca),
	.w5(32'h3b930bb9),
	.w6(32'h3ba6467c),
	.w7(32'h3c0af583),
	.w8(32'h3c241830),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f9f3),
	.w1(32'h3c16b49a),
	.w2(32'h3c2d58ea),
	.w3(32'h3b3d7d1a),
	.w4(32'h3b3985e9),
	.w5(32'h3bd5aedc),
	.w6(32'h3c4630b4),
	.w7(32'h3cadc0a0),
	.w8(32'h3c861a7e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60b44e),
	.w1(32'h3c457a69),
	.w2(32'h3bb422da),
	.w3(32'h3c2953cd),
	.w4(32'hbb69c1af),
	.w5(32'h3a85bc61),
	.w6(32'h3c233896),
	.w7(32'h3b418872),
	.w8(32'hba97b97b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef7dae),
	.w1(32'hbb420ed3),
	.w2(32'hbba03069),
	.w3(32'h3b4ea5ca),
	.w4(32'hbb907077),
	.w5(32'hbc460cdc),
	.w6(32'h3be26a5f),
	.w7(32'h3c2126fc),
	.w8(32'h3bf641a7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc964726),
	.w1(32'h3c1a505a),
	.w2(32'h3a9d2c86),
	.w3(32'hbc65e126),
	.w4(32'h3c813eb9),
	.w5(32'h3ae07b66),
	.w6(32'hbba3d7e0),
	.w7(32'hbbdd2b24),
	.w8(32'hbae89210),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16d0cc),
	.w1(32'hbb3ec33f),
	.w2(32'h3a4e6c97),
	.w3(32'hbc0a1ac2),
	.w4(32'hbba45d27),
	.w5(32'hba3fb3d6),
	.w6(32'hbaa2ff2d),
	.w7(32'h3baf24e2),
	.w8(32'h3c203514),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c329a),
	.w1(32'hbbb87af0),
	.w2(32'hbc1340b5),
	.w3(32'h3c124ca7),
	.w4(32'hbb6ac737),
	.w5(32'hbba0c467),
	.w6(32'hbb585274),
	.w7(32'hbbc65f4e),
	.w8(32'hbc202291),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc062d4b),
	.w1(32'h3c41d44e),
	.w2(32'h3bcfa9e2),
	.w3(32'hbbe691c6),
	.w4(32'h3c44deca),
	.w5(32'h3c3a40d3),
	.w6(32'h3b9e0318),
	.w7(32'h3b9b83b0),
	.w8(32'h3bc10ca5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47ae43),
	.w1(32'h3c59ba62),
	.w2(32'h3b8aeed2),
	.w3(32'h3c658924),
	.w4(32'h3bec45a1),
	.w5(32'hb9012623),
	.w6(32'h3c78f61f),
	.w7(32'h3c1341d7),
	.w8(32'h3c0fb0da),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3650d7ed),
	.w1(32'h3b62f935),
	.w2(32'h3a6ec6a5),
	.w3(32'h3b63664b),
	.w4(32'h3b8797e1),
	.w5(32'h3a3cb378),
	.w6(32'hbaeeebe1),
	.w7(32'h3b86358f),
	.w8(32'h3b19e613),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ef960),
	.w1(32'hbbb0d290),
	.w2(32'hbbcae468),
	.w3(32'hba88c79f),
	.w4(32'hbbf7c955),
	.w5(32'hbbf1a8b2),
	.w6(32'hbc0c8c82),
	.w7(32'hbbb86641),
	.w8(32'hbbe0f2a3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52b36c),
	.w1(32'hbbae83f0),
	.w2(32'hbc20d6db),
	.w3(32'hbc24fce7),
	.w4(32'h39e16242),
	.w5(32'hbab76566),
	.w6(32'h3a33b5d6),
	.w7(32'hbb4fd6fd),
	.w8(32'hba38d271),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ce06),
	.w1(32'h3b4215a1),
	.w2(32'h3a55e9f6),
	.w3(32'h3b3f28b7),
	.w4(32'h3a166046),
	.w5(32'h393037d6),
	.w6(32'hbac62669),
	.w7(32'hba6292d9),
	.w8(32'hbab0e1e0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0bffb),
	.w1(32'h3b286b1b),
	.w2(32'hbb37f005),
	.w3(32'h3b2a5124),
	.w4(32'h3ae93982),
	.w5(32'hbb86b326),
	.w6(32'h3b19275e),
	.w7(32'h3a289225),
	.w8(32'h38326993),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a308),
	.w1(32'h3cf2de1f),
	.w2(32'h3d860078),
	.w3(32'hbb46d982),
	.w4(32'h3cdc6241),
	.w5(32'h3d71d349),
	.w6(32'h3caca369),
	.w7(32'h3d0d3269),
	.w8(32'h3d01a4a8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5b48c6),
	.w1(32'h3be829b1),
	.w2(32'h3a43bddf),
	.w3(32'h3d2f9a30),
	.w4(32'h3be9a382),
	.w5(32'h3b009918),
	.w6(32'h3a82ff9a),
	.w7(32'hba520558),
	.w8(32'h3a2f13c6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840182),
	.w1(32'h3ad7bd67),
	.w2(32'hbbe4d95b),
	.w3(32'h3b2b2935),
	.w4(32'hbb9ea0fb),
	.w5(32'hbb36abfc),
	.w6(32'hba6e227c),
	.w7(32'hbbc5c06b),
	.w8(32'hba141f00),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f433c),
	.w1(32'hbb800847),
	.w2(32'hbc5ba134),
	.w3(32'h3b3537d3),
	.w4(32'h3b17c8ce),
	.w5(32'hbbc2c0ed),
	.w6(32'h398ccdb0),
	.w7(32'hbb435e77),
	.w8(32'h3aa53db4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79f735),
	.w1(32'h3cfce934),
	.w2(32'h3c32ef68),
	.w3(32'h3bd099ab),
	.w4(32'h3d01c47b),
	.w5(32'h3c1456d4),
	.w6(32'h3cba912b),
	.w7(32'h3c28c104),
	.w8(32'hba89a47f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911a14),
	.w1(32'hbb74f7f3),
	.w2(32'hbb8b30d0),
	.w3(32'hbb56f242),
	.w4(32'hbb88ecf3),
	.w5(32'hbaf60246),
	.w6(32'hba9b4e2f),
	.w7(32'h3b187fd8),
	.w8(32'h3b8f3f32),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02bb07),
	.w1(32'h3b33854a),
	.w2(32'h3a64050c),
	.w3(32'h3ba974f4),
	.w4(32'h3bfb34cb),
	.w5(32'hbb4f42bb),
	.w6(32'h3abc87b1),
	.w7(32'hba9f5105),
	.w8(32'hbac39b4f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a89b),
	.w1(32'h3c284e9a),
	.w2(32'hbb9fb951),
	.w3(32'h3b7adf81),
	.w4(32'h3aab61e0),
	.w5(32'hbc42552e),
	.w6(32'h3c4ac191),
	.w7(32'h3bc80990),
	.w8(32'h3c544bed),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b979e96),
	.w1(32'h3b9fe19b),
	.w2(32'hbb952bf2),
	.w3(32'hbaf52306),
	.w4(32'hb9dce7b2),
	.w5(32'hbc00bfa8),
	.w6(32'hbae97a9f),
	.w7(32'hbc28cca5),
	.w8(32'hbc7fec44),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc417d44),
	.w1(32'h3b852587),
	.w2(32'hbabd32a0),
	.w3(32'hbc8891ca),
	.w4(32'h3b299b13),
	.w5(32'h3b1fedea),
	.w6(32'h3ba86b2f),
	.w7(32'h3ba8afe9),
	.w8(32'h3b7f4b4b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21d05f),
	.w1(32'h3b7dc329),
	.w2(32'hbbbc9a84),
	.w3(32'h3b94d18f),
	.w4(32'h3b9bfb94),
	.w5(32'hba109b6a),
	.w6(32'hbb861a3c),
	.w7(32'h3a6b8834),
	.w8(32'h395ad464),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6fc2d),
	.w1(32'h3b042f53),
	.w2(32'h3b2ffd6e),
	.w3(32'h3bf51717),
	.w4(32'h3b9a4269),
	.w5(32'h3b5e361f),
	.w6(32'h3b161fd4),
	.w7(32'h3b239397),
	.w8(32'h3c093a18),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a7089),
	.w1(32'hbb28a098),
	.w2(32'hbbc6e954),
	.w3(32'h3c15023c),
	.w4(32'hbaa3d500),
	.w5(32'hbbc232ec),
	.w6(32'hbc4ad53d),
	.w7(32'hbae79fc5),
	.w8(32'hbb6cfda7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb513),
	.w1(32'hbc3ab98e),
	.w2(32'hbc9e51d7),
	.w3(32'hbb81fc09),
	.w4(32'hb81cd305),
	.w5(32'hbab6f14f),
	.w6(32'hbb448d63),
	.w7(32'hbc1f1608),
	.w8(32'hba38b9c7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941098d),
	.w1(32'h3bfc78d7),
	.w2(32'h39ef0cb4),
	.w3(32'h3c78fc1a),
	.w4(32'h3c1771a0),
	.w5(32'hbbeb510a),
	.w6(32'h3bf8b6c2),
	.w7(32'h3b6f4901),
	.w8(32'h3ba4bda2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa220bb),
	.w1(32'hbb8e3947),
	.w2(32'h3ca5a3b3),
	.w3(32'hb97ddfae),
	.w4(32'h3b8fca4f),
	.w5(32'h3cf90cbc),
	.w6(32'hbbc07843),
	.w7(32'hb9a524bc),
	.w8(32'h3c15f49f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc17ce),
	.w1(32'h3b95cd94),
	.w2(32'hbbd23c1a),
	.w3(32'h3cf9ad51),
	.w4(32'h39bbd6a5),
	.w5(32'hbbdda248),
	.w6(32'hbbb51a83),
	.w7(32'hbbe97254),
	.w8(32'hbbc00493),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62a8da),
	.w1(32'h39ba968e),
	.w2(32'hbb4a6a9f),
	.w3(32'hbb888f5a),
	.w4(32'h3ab1bd44),
	.w5(32'hbbb82926),
	.w6(32'h3ab46488),
	.w7(32'hbad3e046),
	.w8(32'h3b5763d4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8440c8),
	.w1(32'h3be5f8c0),
	.w2(32'hbb2345be),
	.w3(32'h3aea9a27),
	.w4(32'hba00e812),
	.w5(32'hba0bc85c),
	.w6(32'hbc015277),
	.w7(32'hbbd21ea4),
	.w8(32'hbc01f121),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b058dd3),
	.w1(32'h3a07d71f),
	.w2(32'h3ac23dc0),
	.w3(32'h3bc227da),
	.w4(32'hbbbe755c),
	.w5(32'hbbe1e77f),
	.w6(32'h3a9239ba),
	.w7(32'h3c0c2bd4),
	.w8(32'h3a9e33e1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cbe49),
	.w1(32'hbb1e2dd7),
	.w2(32'hbc21672f),
	.w3(32'hbbef59c9),
	.w4(32'hbb76fe8a),
	.w5(32'hbc4e626d),
	.w6(32'hbb866a06),
	.w7(32'hbbb6324d),
	.w8(32'hba8d5d9f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a296b8),
	.w1(32'h3c866f27),
	.w2(32'h3cdc350f),
	.w3(32'h39daf768),
	.w4(32'h3c3c7040),
	.w5(32'h3cc9e6c4),
	.w6(32'h3bd543a6),
	.w7(32'h3c4b0d64),
	.w8(32'h3be5b02e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85caf9),
	.w1(32'h3be33e9c),
	.w2(32'hbbba5867),
	.w3(32'h3c43ae12),
	.w4(32'h39bc600f),
	.w5(32'hb989c546),
	.w6(32'h3bb1a0b3),
	.w7(32'h3bfc159d),
	.w8(32'h3bf3070d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24fe5a),
	.w1(32'h3c390471),
	.w2(32'h3c213341),
	.w3(32'h3ba0e8b8),
	.w4(32'h3bf8c6b4),
	.w5(32'hba8148e4),
	.w6(32'h3c3d0490),
	.w7(32'h3c8a5366),
	.w8(32'h3c5c53d5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2c25c),
	.w1(32'h3bcf6433),
	.w2(32'h39aaec4f),
	.w3(32'h3b350823),
	.w4(32'h3c31ccb1),
	.w5(32'h3bf504eb),
	.w6(32'h3ba3aa5f),
	.w7(32'h3b33b4a3),
	.w8(32'h3b281fcc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd93b),
	.w1(32'hba8fcd3d),
	.w2(32'hbccd32cb),
	.w3(32'h3b96f459),
	.w4(32'hbb7e0d61),
	.w5(32'hbca4eba3),
	.w6(32'h3a3a0c76),
	.w7(32'hbbbb31e7),
	.w8(32'hbb927444),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40ace0),
	.w1(32'h3b275e89),
	.w2(32'h3ac3f90a),
	.w3(32'hbba6cadf),
	.w4(32'h3b881100),
	.w5(32'h3b54fa40),
	.w6(32'h3be09872),
	.w7(32'h3bbbcc3b),
	.w8(32'h3b753041),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a179181),
	.w1(32'h3d12e4f0),
	.w2(32'h3d8b3574),
	.w3(32'h3aa80c04),
	.w4(32'h3cfd3060),
	.w5(32'h3d762e09),
	.w6(32'h3ca312b3),
	.w7(32'h3d01e608),
	.w8(32'h3ca95a8e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d481d44),
	.w1(32'hbaed2fbc),
	.w2(32'hbc24eb53),
	.w3(32'h3d29150d),
	.w4(32'h38e698a7),
	.w5(32'hbbbe69f5),
	.w6(32'h3b28fb0f),
	.w7(32'hbbb198ef),
	.w8(32'hbb8375a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f001f),
	.w1(32'hbb6e0230),
	.w2(32'hb981e560),
	.w3(32'hbb6553ec),
	.w4(32'h3bc33796),
	.w5(32'h3b2adfe9),
	.w6(32'h3a4703ab),
	.w7(32'h394983c8),
	.w8(32'h3aa40508),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144ccc),
	.w1(32'h3c0d85df),
	.w2(32'hbb625fa7),
	.w3(32'hbb1d91f7),
	.w4(32'h3af4fac1),
	.w5(32'hbaa89327),
	.w6(32'h3b17f5f4),
	.w7(32'hb99ce332),
	.w8(32'hbaa8f07d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe39f1),
	.w1(32'hba13aa7a),
	.w2(32'h3c203dae),
	.w3(32'hbbc9c563),
	.w4(32'hbb985b92),
	.w5(32'hba85b214),
	.w6(32'hbb117bef),
	.w7(32'h38bffd7c),
	.w8(32'hba08eeda),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b09666),
	.w1(32'h3b3dfbf8),
	.w2(32'h3ae93a87),
	.w3(32'h3befde18),
	.w4(32'h3c197dad),
	.w5(32'h3bbfd9e7),
	.w6(32'h3c0ba34c),
	.w7(32'h3bcb4cea),
	.w8(32'h3c862f1f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14485d),
	.w1(32'hbb6d4f12),
	.w2(32'h3b929d4b),
	.w3(32'h3c776ba8),
	.w4(32'hba9f6b46),
	.w5(32'h3b3d7582),
	.w6(32'h3ba30572),
	.w7(32'h3c6e784f),
	.w8(32'h3ca52dc5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65ee10),
	.w1(32'h3917afdd),
	.w2(32'hb9f72ffa),
	.w3(32'h3c173660),
	.w4(32'h3bbe4493),
	.w5(32'h3b33d893),
	.w6(32'h3b126549),
	.w7(32'h3a2af186),
	.w8(32'h3b3a4406),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbb84b),
	.w1(32'h3b6d5d1b),
	.w2(32'h3bb4bbbb),
	.w3(32'h3b9786ab),
	.w4(32'hbb5c8bf0),
	.w5(32'h3af0bf71),
	.w6(32'hb88a8754),
	.w7(32'hba471c44),
	.w8(32'hbb336755),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c3b5a),
	.w1(32'hbb9349e9),
	.w2(32'hbc1f1d27),
	.w3(32'hbbb92710),
	.w4(32'hbc0db715),
	.w5(32'hbc2b5acb),
	.w6(32'hbbc2accb),
	.w7(32'hbbd20243),
	.w8(32'hbb7c7899),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e525a),
	.w1(32'h3c02a520),
	.w2(32'h3bd987fe),
	.w3(32'hba8e57b3),
	.w4(32'h32e460c3),
	.w5(32'h3b8971ec),
	.w6(32'hba06bb4a),
	.w7(32'h3b856be9),
	.w8(32'h3b4af8a2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c165869),
	.w1(32'hbad209da),
	.w2(32'hbbe8d747),
	.w3(32'h3bbb6767),
	.w4(32'hbbbee6e0),
	.w5(32'hbc2af8c9),
	.w6(32'hbb4f8eb9),
	.w7(32'hbc21e5be),
	.w8(32'hbb394143),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7958),
	.w1(32'hbb8c3d70),
	.w2(32'hbba3e7d3),
	.w3(32'hb96eac37),
	.w4(32'hbbc2ac8e),
	.w5(32'hbb63b696),
	.w6(32'hbb03d002),
	.w7(32'hbb05f89a),
	.w8(32'hbb1625ab),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4399c),
	.w1(32'h3c099baa),
	.w2(32'hb9d61d20),
	.w3(32'h3b9eb71b),
	.w4(32'h3bf3c8ec),
	.w5(32'hbada8fc8),
	.w6(32'h3bb653cb),
	.w7(32'h3ab9279d),
	.w8(32'hbb55ef37),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacf4d1),
	.w1(32'h3b9b7978),
	.w2(32'h3b73f43b),
	.w3(32'hbac3bfd2),
	.w4(32'h3c100a0f),
	.w5(32'hbb2d4943),
	.w6(32'h3917ad83),
	.w7(32'h3ba09ee4),
	.w8(32'h3c0788ab),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095976),
	.w1(32'h3b8e64c1),
	.w2(32'h3bacd348),
	.w3(32'h3b104584),
	.w4(32'h3b86b4e4),
	.w5(32'h3bb009ed),
	.w6(32'hbb76d287),
	.w7(32'hba4259a9),
	.w8(32'h39ddf212),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78ddee),
	.w1(32'hbbb2c26d),
	.w2(32'hbb2a1b63),
	.w3(32'h3b7278ac),
	.w4(32'h3ba575a6),
	.w5(32'h3b6515aa),
	.w6(32'hbb35a467),
	.w7(32'hba87b9c4),
	.w8(32'h3b8b276e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3f47b),
	.w1(32'hbb0ea133),
	.w2(32'h3a27fd5d),
	.w3(32'h3ba6b778),
	.w4(32'h3b70f081),
	.w5(32'h3ab3cbdb),
	.w6(32'hbb97c308),
	.w7(32'hbb166c6f),
	.w8(32'h3b5ed49b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17db45),
	.w1(32'h3b2c0efc),
	.w2(32'hbb3643f8),
	.w3(32'h38fc806b),
	.w4(32'h3c2930b3),
	.w5(32'hbaa8b1d8),
	.w6(32'h3bafb013),
	.w7(32'hb9dd7a53),
	.w8(32'hba12f625),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dfcb9),
	.w1(32'hbc11d1e9),
	.w2(32'hbc9931ca),
	.w3(32'hbb490afe),
	.w4(32'hbb9adcb4),
	.w5(32'hbcb7b4f5),
	.w6(32'h3a243f28),
	.w7(32'h3aa0d413),
	.w8(32'hbba29744),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb583f),
	.w1(32'h3bede2f3),
	.w2(32'h3b37e2bd),
	.w3(32'hbb7f197d),
	.w4(32'h3b7dc635),
	.w5(32'hbb3dc76c),
	.w6(32'hbaed7c4b),
	.w7(32'hba9b0be2),
	.w8(32'h3b6f661b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c087006),
	.w1(32'hbc122975),
	.w2(32'hbc35d2c4),
	.w3(32'h3bfe1469),
	.w4(32'h3b07ba98),
	.w5(32'hbc761aa4),
	.w6(32'h3a34d6da),
	.w7(32'hbadfa316),
	.w8(32'hba9ad0e9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ee9c3),
	.w1(32'h3af60558),
	.w2(32'hbacab86d),
	.w3(32'hbc1f22c9),
	.w4(32'h3b04cd32),
	.w5(32'hbaacd0e7),
	.w6(32'h3bdcc949),
	.w7(32'h3bec677f),
	.w8(32'h3c39d75f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ccd43d),
	.w1(32'h3c78b525),
	.w2(32'h3ba39144),
	.w3(32'hbada4680),
	.w4(32'h3baca5aa),
	.w5(32'hbb174693),
	.w6(32'h3cbaf064),
	.w7(32'h3cb92f0f),
	.w8(32'h3cc8459d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb442b),
	.w1(32'h3b1170f7),
	.w2(32'h3a9944e3),
	.w3(32'hb97d7fee),
	.w4(32'h3bac68c5),
	.w5(32'h3b613aae),
	.w6(32'h3baa479d),
	.w7(32'h3c054fc6),
	.w8(32'h3c02ce7f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f883e),
	.w1(32'h3b209c62),
	.w2(32'h3bb9284a),
	.w3(32'h3b8d1e93),
	.w4(32'h3bf3f960),
	.w5(32'h3c1f4212),
	.w6(32'h3b6aae36),
	.w7(32'h3c05203f),
	.w8(32'h3c20f886),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9dd3e),
	.w1(32'hba5aaedc),
	.w2(32'hbaf8885d),
	.w3(32'h3c331061),
	.w4(32'h3ba5d5c9),
	.w5(32'h3c102ccb),
	.w6(32'h3b41716d),
	.w7(32'h3bcf6b7a),
	.w8(32'h3b270f05),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b1320),
	.w1(32'hbb5de1be),
	.w2(32'hbc0d1e0c),
	.w3(32'h3bb971c4),
	.w4(32'hb9d490ad),
	.w5(32'hbb1981da),
	.w6(32'hbaf7c4cd),
	.w7(32'hbbce2ada),
	.w8(32'hbbb7c522),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d53ad),
	.w1(32'hbba238d9),
	.w2(32'hbc2855c1),
	.w3(32'hb956d5b6),
	.w4(32'hbb8f8ca9),
	.w5(32'hbc3f2e11),
	.w6(32'hba1175d7),
	.w7(32'hba6986c5),
	.w8(32'hb9819f2e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c88e),
	.w1(32'h3b1de57b),
	.w2(32'hbc21d38f),
	.w3(32'hbc1ea87f),
	.w4(32'h3bb4dc14),
	.w5(32'hbba8424a),
	.w6(32'h3baef69e),
	.w7(32'hbaaa6e8c),
	.w8(32'h3975925d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9570a2),
	.w1(32'h3a37c3e5),
	.w2(32'hbc40e525),
	.w3(32'hbb23c8f2),
	.w4(32'hbbe62f82),
	.w5(32'hbc649e77),
	.w6(32'hba407b97),
	.w7(32'h3accb0bb),
	.w8(32'h3b03100f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d88dfc),
	.w1(32'h3bad4237),
	.w2(32'hbb548186),
	.w3(32'h3bc13e12),
	.w4(32'hba04b954),
	.w5(32'hbbdc88dc),
	.w6(32'h3bbf10c8),
	.w7(32'hba44dad5),
	.w8(32'h3a9ac300),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48276e),
	.w1(32'h3af38a7e),
	.w2(32'h3b02fc74),
	.w3(32'hbb417483),
	.w4(32'hbb80d538),
	.w5(32'hbb4f8302),
	.w6(32'h3b4c9387),
	.w7(32'h3bd1d157),
	.w8(32'h3b92c825),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89dfec),
	.w1(32'h3b7e849f),
	.w2(32'h38bae850),
	.w3(32'h3bec72ea),
	.w4(32'h3b68c011),
	.w5(32'h3a4449bb),
	.w6(32'h39a2d576),
	.w7(32'h3a4d049e),
	.w8(32'h3b5076b1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d45d5),
	.w1(32'h3c0527ab),
	.w2(32'h3b5fea0c),
	.w3(32'h3a8b6f25),
	.w4(32'h3b04b256),
	.w5(32'h3b142d83),
	.w6(32'h3bb0a8f0),
	.w7(32'h394a329b),
	.w8(32'hba7ade59),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fde1a),
	.w1(32'hbb967352),
	.w2(32'hba2bc15b),
	.w3(32'hba854039),
	.w4(32'hbba4ca41),
	.w5(32'hbb4fd9aa),
	.w6(32'h3b72b54b),
	.w7(32'h3c35adcc),
	.w8(32'h3ba5d0ea),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57185),
	.w1(32'hbc146117),
	.w2(32'h3a0e5b2e),
	.w3(32'hbb78dcb2),
	.w4(32'h39be32b4),
	.w5(32'hbb08c005),
	.w6(32'hbb0fbf58),
	.w7(32'hb9f86649),
	.w8(32'hbb427423),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab03b5d),
	.w1(32'h3b2c80c0),
	.w2(32'hbac766cc),
	.w3(32'hbc0ab68f),
	.w4(32'h398b5a80),
	.w5(32'hbbdade56),
	.w6(32'h3c364490),
	.w7(32'h3c343bd6),
	.w8(32'h3be783e6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65b5a4),
	.w1(32'hba525b98),
	.w2(32'hbb045aba),
	.w3(32'hbc088a7a),
	.w4(32'hba4f4971),
	.w5(32'h3aa63ced),
	.w6(32'hbbb73fcd),
	.w7(32'h3883adfe),
	.w8(32'hbb76043b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d7bda),
	.w1(32'h3bf3d1c0),
	.w2(32'h3c61f33b),
	.w3(32'h3b80f446),
	.w4(32'h3aebdb18),
	.w5(32'h3bc82cfd),
	.w6(32'h3b6d0103),
	.w7(32'h3c41a51e),
	.w8(32'h3c7b9a0b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44ed1e),
	.w1(32'h3b8384f7),
	.w2(32'hbba1d1b1),
	.w3(32'h3b943b32),
	.w4(32'h3a394580),
	.w5(32'hbbe1b6ba),
	.w6(32'h3abeb6e2),
	.w7(32'h39ebab42),
	.w8(32'h3b3a5a4e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985e13),
	.w1(32'h3cad3ebc),
	.w2(32'h3d17d9bd),
	.w3(32'hbb980427),
	.w4(32'h3c8918d7),
	.w5(32'h3d05e35a),
	.w6(32'h3bbc532b),
	.w7(32'h3b5fc7ac),
	.w8(32'h3ad4e507),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce5248a),
	.w1(32'h3be26c39),
	.w2(32'h3c006560),
	.w3(32'h3ca99268),
	.w4(32'h3bc86368),
	.w5(32'h3b3732fb),
	.w6(32'h3c45a9ff),
	.w7(32'h3c899cd0),
	.w8(32'h3c5a1ded),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c108669),
	.w1(32'h3b3f404c),
	.w2(32'h3be139f1),
	.w3(32'h3bcde705),
	.w4(32'h3b97ebf6),
	.w5(32'hba49bea4),
	.w6(32'hbab966a5),
	.w7(32'h3b6b1d2b),
	.w8(32'h3bcee195),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d5f0),
	.w1(32'hb89a7e07),
	.w2(32'hbc0b68e6),
	.w3(32'h3b115793),
	.w4(32'hba62e60c),
	.w5(32'hbb5d157b),
	.w6(32'h3b0b16e8),
	.w7(32'h39f39523),
	.w8(32'h3965975d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3e014),
	.w1(32'hba3d19be),
	.w2(32'h3ad9e0bb),
	.w3(32'hbb937e65),
	.w4(32'h3b8eb785),
	.w5(32'h3be59b49),
	.w6(32'h3ac1c8ad),
	.w7(32'hba30035f),
	.w8(32'h3b97e371),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1eef1),
	.w1(32'h3b3a57a3),
	.w2(32'hbac7ee11),
	.w3(32'h3c241009),
	.w4(32'h3af80270),
	.w5(32'hbb2e4c5e),
	.w6(32'h3ad69020),
	.w7(32'h3aa89cbe),
	.w8(32'h3b231ab9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c8ab1),
	.w1(32'h3c1bab80),
	.w2(32'h3b81bf81),
	.w3(32'h3af1c044),
	.w4(32'h3c1c35ff),
	.w5(32'h3b0dc42c),
	.w6(32'h3c2087f2),
	.w7(32'h3bcdd3de),
	.w8(32'h3bcd9df3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14018b),
	.w1(32'hbc1164e7),
	.w2(32'hbcb561b5),
	.w3(32'hba0a3242),
	.w4(32'hbb5ad3fe),
	.w5(32'hbcb2cc6e),
	.w6(32'hbbdf840e),
	.w7(32'hbc5c0a3d),
	.w8(32'hbbdb49f6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc844fd0),
	.w1(32'h3b11721f),
	.w2(32'h3b16824e),
	.w3(32'hbc3565c6),
	.w4(32'hbbf6154f),
	.w5(32'hba009078),
	.w6(32'h3a5ec61f),
	.w7(32'h3b7565ed),
	.w8(32'h3c0f2298),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b262b00),
	.w1(32'h3bf863aa),
	.w2(32'h3b6c884e),
	.w3(32'h3b22312f),
	.w4(32'h3c3fd8ff),
	.w5(32'h3b9877c8),
	.w6(32'h3bae6f35),
	.w7(32'h3bcab872),
	.w8(32'h3b8b69f5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad45bcb),
	.w1(32'h3c21bfbe),
	.w2(32'h3cc4be88),
	.w3(32'h3b45acd6),
	.w4(32'h3c465223),
	.w5(32'h3cd0cfa8),
	.w6(32'h3ba287b3),
	.w7(32'h3c214f89),
	.w8(32'h3c2ab267),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb477b1),
	.w1(32'h3a8ca847),
	.w2(32'hbb981af4),
	.w3(32'h3caf55fe),
	.w4(32'hbb245c6a),
	.w5(32'hbbd101a1),
	.w6(32'h3b7b0b88),
	.w7(32'hba439e2e),
	.w8(32'hbadc961f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd09914),
	.w1(32'hbbb4c65c),
	.w2(32'hbc6ad514),
	.w3(32'hbbe39ab5),
	.w4(32'hbbbea207),
	.w5(32'hbc758b5c),
	.w6(32'hbae39fff),
	.w7(32'hbbf10270),
	.w8(32'hbbe03aa5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030b16),
	.w1(32'hb7c7c863),
	.w2(32'hbb6ba792),
	.w3(32'hbc068bc6),
	.w4(32'h3b670930),
	.w5(32'hbb5f2aaa),
	.w6(32'hba1fbbd1),
	.w7(32'h3bdd96e6),
	.w8(32'hbaa738cd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae574f3),
	.w1(32'h3b9396ca),
	.w2(32'h3b6208e4),
	.w3(32'hbb3c5f02),
	.w4(32'h3b1dddea),
	.w5(32'h39aad515),
	.w6(32'h3a1864e4),
	.w7(32'h3b066738),
	.w8(32'hb9ccba74),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8787a88),
	.w1(32'hbbcc3347),
	.w2(32'h39f0d9dd),
	.w3(32'h3a5a31c9),
	.w4(32'hba8e378f),
	.w5(32'hbb72f94a),
	.w6(32'hbc0ca672),
	.w7(32'hbb2863c7),
	.w8(32'hbbc70143),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc5486),
	.w1(32'h3c1c86f0),
	.w2(32'h3b86ca93),
	.w3(32'h3b793c4d),
	.w4(32'h3c0a9e33),
	.w5(32'hb94d377a),
	.w6(32'h3c24eb23),
	.w7(32'h3c0e5898),
	.w8(32'h3bda6424),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ae49),
	.w1(32'hbb9603e4),
	.w2(32'hbcd53c15),
	.w3(32'h3b9cbae6),
	.w4(32'h3ad8b7ee),
	.w5(32'hbc85dcec),
	.w6(32'h3b8e5de5),
	.w7(32'hbb8656f9),
	.w8(32'h3a515c99),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6547ea),
	.w1(32'hbae79799),
	.w2(32'hbc9ba104),
	.w3(32'hbbd7ddc0),
	.w4(32'hbb570f0b),
	.w5(32'hbc54bdce),
	.w6(32'h39d9e0b2),
	.w7(32'hbbd23e75),
	.w8(32'hbb23a9c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc869a6),
	.w1(32'h3bfb5bd2),
	.w2(32'h3ba132e3),
	.w3(32'hbb817b37),
	.w4(32'h3c07c95e),
	.w5(32'h3bbb5b27),
	.w6(32'h3bd1171a),
	.w7(32'h3c0101e2),
	.w8(32'h3c3cae3f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50ddfb),
	.w1(32'hbb059bb7),
	.w2(32'hbb35ad4c),
	.w3(32'h3c16d189),
	.w4(32'hbb1eebde),
	.w5(32'h3ad0eb90),
	.w6(32'hbb0f97b7),
	.w7(32'hbb6be836),
	.w8(32'hbb21ef36),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b984c53),
	.w1(32'hbb11b63f),
	.w2(32'hbb8decbf),
	.w3(32'hba4dbaa6),
	.w4(32'hbb1a89f8),
	.w5(32'hbba85316),
	.w6(32'hbb00c8de),
	.w7(32'hbbb1b9bb),
	.w8(32'hbabb7027),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9de957),
	.w1(32'h3bbdf23d),
	.w2(32'hbc12e2f1),
	.w3(32'h3b13aea0),
	.w4(32'h3bd4976d),
	.w5(32'hbc277770),
	.w6(32'h3a535739),
	.w7(32'hbbeec2aa),
	.w8(32'hbb3290ca),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule