module layer_10_featuremap_481(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1cff4),
	.w1(32'h3a1b314e),
	.w2(32'h3a9ef8db),
	.w3(32'hbc1af9b6),
	.w4(32'h3b121067),
	.w5(32'h3b2c2311),
	.w6(32'hbbeb8aee),
	.w7(32'hba8dec62),
	.w8(32'hbb5c4049),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f96e8),
	.w1(32'hbbde2ae3),
	.w2(32'h3aae7e8f),
	.w3(32'h3b8135ee),
	.w4(32'hbbf347a8),
	.w5(32'h3a1199e8),
	.w6(32'hbab0599f),
	.w7(32'hbbe19b73),
	.w8(32'h3c467db2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f5d47),
	.w1(32'hbb1eb431),
	.w2(32'h3a297ba7),
	.w3(32'h3c037d88),
	.w4(32'hbb398cd2),
	.w5(32'hbc396141),
	.w6(32'h3bb68b3c),
	.w7(32'hbb62c781),
	.w8(32'hbb1166ac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cf7cc),
	.w1(32'hbb98e88d),
	.w2(32'hbb8c5c4e),
	.w3(32'hbbdc3afd),
	.w4(32'h3a9fc4dc),
	.w5(32'h3cf90128),
	.w6(32'h39fb5861),
	.w7(32'h3b73bf37),
	.w8(32'h3c8406ff),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c88c4),
	.w1(32'h3b5005aa),
	.w2(32'hbaef2c26),
	.w3(32'h3c0669f3),
	.w4(32'h38ad2fc4),
	.w5(32'hbb926576),
	.w6(32'hbba5fa23),
	.w7(32'hbb361d37),
	.w8(32'hbaa92532),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0500d),
	.w1(32'h3a1cfaf8),
	.w2(32'h3c3b0a27),
	.w3(32'hbada5b84),
	.w4(32'h3b3ea85a),
	.w5(32'h3b9630b2),
	.w6(32'h3b2c1887),
	.w7(32'hbb84342f),
	.w8(32'hbb12f6c7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3c3ec),
	.w1(32'hbbd49072),
	.w2(32'hba7c2856),
	.w3(32'h3b7664b1),
	.w4(32'hbb7ac189),
	.w5(32'h3af99e8a),
	.w6(32'hba9c49a6),
	.w7(32'hb987ebb6),
	.w8(32'h3b961f67),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e1db5),
	.w1(32'h3bdaf7c3),
	.w2(32'hbb638a3a),
	.w3(32'h3c062907),
	.w4(32'hbaef41f2),
	.w5(32'hbc2976ae),
	.w6(32'h3c5aa2bb),
	.w7(32'h3c29cda9),
	.w8(32'h3bc1f9c2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ff2fb),
	.w1(32'hbb307870),
	.w2(32'h3abab862),
	.w3(32'hbbe02d1c),
	.w4(32'hba82c051),
	.w5(32'h3b1b4cff),
	.w6(32'h39e63746),
	.w7(32'h39b72f9e),
	.w8(32'h39ed7de4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d427a5),
	.w1(32'h3bd6c54f),
	.w2(32'h3c2028fe),
	.w3(32'h3ac4b467),
	.w4(32'h3b9a56c6),
	.w5(32'h3c7cf540),
	.w6(32'h3b6efbb8),
	.w7(32'h3b662b69),
	.w8(32'h3b449924),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a549972),
	.w1(32'hb897d330),
	.w2(32'h3b88f894),
	.w3(32'hba4414e9),
	.w4(32'h3bf14a4c),
	.w5(32'h3c143622),
	.w6(32'hbb25f879),
	.w7(32'h3bd0c3ce),
	.w8(32'h39b50240),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f86943),
	.w1(32'h3af31cb1),
	.w2(32'hba8fe8c2),
	.w3(32'h3b71f03f),
	.w4(32'h3903e51c),
	.w5(32'hbbbade65),
	.w6(32'h3a53ddb8),
	.w7(32'h3b1f3925),
	.w8(32'h3acebc64),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1033d8),
	.w1(32'h3baf2c6c),
	.w2(32'h3a574370),
	.w3(32'h3b999c5b),
	.w4(32'hbb095710),
	.w5(32'h3c8894bb),
	.w6(32'h3c301b28),
	.w7(32'h3b76703c),
	.w8(32'h3c79471b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae97802),
	.w1(32'hbb971a9d),
	.w2(32'hbbe24396),
	.w3(32'h3a373e50),
	.w4(32'hbba8b419),
	.w5(32'h3b7d9b7d),
	.w6(32'hba39e5fb),
	.w7(32'h3b87f043),
	.w8(32'h3bbdeadb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1d3d6),
	.w1(32'hba91bbe2),
	.w2(32'hbb962563),
	.w3(32'h3c0e8c2c),
	.w4(32'hbbcc8800),
	.w5(32'hbc2045fb),
	.w6(32'hbb26c665),
	.w7(32'hb963fe52),
	.w8(32'hbb9e5632),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2924),
	.w1(32'h3b5dcfa7),
	.w2(32'h3bf191bc),
	.w3(32'hbb68c77d),
	.w4(32'h3997bc39),
	.w5(32'hba96ef7e),
	.w6(32'h3bdf4027),
	.w7(32'h3beced91),
	.w8(32'h3a7ff221),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc62fd),
	.w1(32'hba932f42),
	.w2(32'hbb280e15),
	.w3(32'hbbc49d1c),
	.w4(32'h3abb33ba),
	.w5(32'h39ffe7c0),
	.w6(32'h3bcb50f0),
	.w7(32'h3a0e57ca),
	.w8(32'h3bd1acf9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e1b1d),
	.w1(32'h3bd0ed0e),
	.w2(32'h3c54577f),
	.w3(32'h3c17a7c1),
	.w4(32'h3b17f147),
	.w5(32'hb9e12f47),
	.w6(32'h3c9695f0),
	.w7(32'h3be1f9ef),
	.w8(32'hbc1ba44b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd933a),
	.w1(32'h3c006d16),
	.w2(32'h3b869f84),
	.w3(32'h3bf901d9),
	.w4(32'h3a25106f),
	.w5(32'hbb99e61f),
	.w6(32'h3bc205be),
	.w7(32'h3b168faf),
	.w8(32'hbbb56d62),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb320976),
	.w1(32'h3ac4fe81),
	.w2(32'h3b19a126),
	.w3(32'hbbb94fff),
	.w4(32'hbb4bfdf5),
	.w5(32'hbba1cf08),
	.w6(32'h3a1cbdcf),
	.w7(32'h3b8e7f61),
	.w8(32'h3b2782b0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82b69b),
	.w1(32'h3ad898a9),
	.w2(32'hbaacb1d8),
	.w3(32'hbb28b411),
	.w4(32'h3b8eb865),
	.w5(32'h3a001098),
	.w6(32'h3bce91e3),
	.w7(32'hb80131cd),
	.w8(32'h3a77979e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e25ee),
	.w1(32'hb97e5280),
	.w2(32'hbc02c732),
	.w3(32'hbb27d2de),
	.w4(32'hba447499),
	.w5(32'h391e11e8),
	.w6(32'hba9d204d),
	.w7(32'h3b38ead3),
	.w8(32'hb8ec61c1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969f5e),
	.w1(32'h3ba1642a),
	.w2(32'h3c8d7ec1),
	.w3(32'hb7cebecf),
	.w4(32'h3bff1f8a),
	.w5(32'h3bb1b18b),
	.w6(32'h3be9a2ee),
	.w7(32'h3c2d1817),
	.w8(32'h3aa079aa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3f11b),
	.w1(32'h3b16253c),
	.w2(32'h3b36cc32),
	.w3(32'h39744d64),
	.w4(32'hbb6a6863),
	.w5(32'h3acee5c1),
	.w6(32'hbb3b7a91),
	.w7(32'hbb62034a),
	.w8(32'hbadbff3f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb95238),
	.w1(32'h3aab0fb0),
	.w2(32'h3b1cc0c5),
	.w3(32'h3a59b6ac),
	.w4(32'h3baaa09f),
	.w5(32'hbb49ac8d),
	.w6(32'hbad626bd),
	.w7(32'h3b3c35f4),
	.w8(32'h3aab9998),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0769a4),
	.w1(32'h3badb37a),
	.w2(32'hbb0d9c44),
	.w3(32'hbc01a679),
	.w4(32'h398a41b3),
	.w5(32'hbbe35f86),
	.w6(32'hbc1fb258),
	.w7(32'h3a5380e3),
	.w8(32'hbbe22d9c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf18a1),
	.w1(32'h3bf4d67b),
	.w2(32'h3b97314c),
	.w3(32'hbc319a8a),
	.w4(32'h3bcbf8ce),
	.w5(32'h3a53f6ad),
	.w6(32'hbb23b313),
	.w7(32'h3a113cc4),
	.w8(32'h3a738aad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf8a4d),
	.w1(32'hbb8afe60),
	.w2(32'hb81b9b4f),
	.w3(32'hbb97eeff),
	.w4(32'hbb867002),
	.w5(32'hbabffbaf),
	.w6(32'h3bbff7d4),
	.w7(32'hbab871ed),
	.w8(32'hbaf8f88c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b9da6),
	.w1(32'h3b1bae10),
	.w2(32'h3bb2feab),
	.w3(32'hbb387e9e),
	.w4(32'h3c1354c8),
	.w5(32'hbbdc9ec0),
	.w6(32'hbafa7e27),
	.w7(32'hbbbf209d),
	.w8(32'hbc2e878b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa244f8),
	.w1(32'h3b92ca1f),
	.w2(32'h3b0c15c3),
	.w3(32'hbba06fae),
	.w4(32'h3b9e08f6),
	.w5(32'h3bbd74e9),
	.w6(32'h3b54bb6a),
	.w7(32'h3a61bf94),
	.w8(32'h3b0624fd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1de21b),
	.w1(32'h3b68de1c),
	.w2(32'h3ad77903),
	.w3(32'h38391103),
	.w4(32'hbb3f1abe),
	.w5(32'h3a1f71f9),
	.w6(32'hba6e47b7),
	.w7(32'hbb8afa2a),
	.w8(32'hbb725524),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af1e3d),
	.w1(32'hbb260084),
	.w2(32'hbb512bb3),
	.w3(32'h3b91ceb9),
	.w4(32'h3b4075a7),
	.w5(32'h3b596ac3),
	.w6(32'hb9d67c64),
	.w7(32'hba10657a),
	.w8(32'h3bc7d251),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c017912),
	.w1(32'hba6e482a),
	.w2(32'hbbcec037),
	.w3(32'h3ae55b88),
	.w4(32'hbab3aba2),
	.w5(32'hbc0c2d96),
	.w6(32'h3b5779f4),
	.w7(32'h3b04854b),
	.w8(32'h3b020cc2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3733f4),
	.w1(32'hbb80a19a),
	.w2(32'hbb4f1ba9),
	.w3(32'hbb4c8553),
	.w4(32'hbb34c097),
	.w5(32'hbacbc1c3),
	.w6(32'h3bd68220),
	.w7(32'h3babc6a2),
	.w8(32'h3b8b6731),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83ebc1),
	.w1(32'h3bb6d93c),
	.w2(32'h3b9017c0),
	.w3(32'h3b0b7e79),
	.w4(32'hba141217),
	.w5(32'h3c2ee007),
	.w6(32'h3bb55a87),
	.w7(32'h3c3c04f7),
	.w8(32'h3bed9509),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c000715),
	.w1(32'h3a7982da),
	.w2(32'h39f169dc),
	.w3(32'h3c866b0f),
	.w4(32'h3a885430),
	.w5(32'h3b184c2e),
	.w6(32'hbad503be),
	.w7(32'h3ae3a827),
	.w8(32'hba2444a8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f498c5),
	.w1(32'h3b12e78b),
	.w2(32'h3b906674),
	.w3(32'h3b2828f0),
	.w4(32'h3bac45d7),
	.w5(32'h3c0eb1f5),
	.w6(32'h3b150313),
	.w7(32'h3b532093),
	.w8(32'h3bbab414),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb659b4c),
	.w1(32'hbc1fff5c),
	.w2(32'hbbb7335e),
	.w3(32'hbbbd8a28),
	.w4(32'hbc7726e8),
	.w5(32'hbc08b50f),
	.w6(32'hbc1e91a2),
	.w7(32'hbc01c543),
	.w8(32'h3c36200d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad15a5b),
	.w1(32'hbc0182f4),
	.w2(32'h3b7d0d00),
	.w3(32'hbc2ea33f),
	.w4(32'hbc62d4e1),
	.w5(32'hbba3209c),
	.w6(32'hbc01b329),
	.w7(32'hbb9ccdeb),
	.w8(32'h3c0ee1e2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f86b34),
	.w1(32'hb8fd973f),
	.w2(32'hbb166658),
	.w3(32'hbb3e7f4f),
	.w4(32'hbaf18943),
	.w5(32'hba3227b4),
	.w6(32'hbb8f13c0),
	.w7(32'h3b496f15),
	.w8(32'h3a1464a3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9df876),
	.w1(32'h3b60f0f4),
	.w2(32'hbc34a583),
	.w3(32'hb93c071d),
	.w4(32'hbbc8c7d5),
	.w5(32'hbbf76f78),
	.w6(32'hbb960c52),
	.w7(32'h3bc6a406),
	.w8(32'h3c4543db),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf770f8),
	.w1(32'hbaf9f14b),
	.w2(32'hbbe75a92),
	.w3(32'h3c2c9df4),
	.w4(32'hbbc35202),
	.w5(32'hbb47b93f),
	.w6(32'hb955a787),
	.w7(32'hbafa9677),
	.w8(32'h3aa60c74),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6f0a9),
	.w1(32'hbb040e60),
	.w2(32'h3b059cb3),
	.w3(32'hbbdf638f),
	.w4(32'h39ea4bb5),
	.w5(32'h3cbd4376),
	.w6(32'hbbd9bf45),
	.w7(32'h3b2659f5),
	.w8(32'h3c52a1e8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053536),
	.w1(32'hbb374b23),
	.w2(32'h3b74b0a2),
	.w3(32'h3c6a9c58),
	.w4(32'hbaa43d8d),
	.w5(32'h3bf43aca),
	.w6(32'h3bea8e1a),
	.w7(32'h3c37f913),
	.w8(32'h3c8cc5ff),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ab2d0),
	.w1(32'hbaa2f279),
	.w2(32'h3b1a70f6),
	.w3(32'h3bd8a454),
	.w4(32'hbc006a88),
	.w5(32'hbac880ac),
	.w6(32'hb91b6dce),
	.w7(32'hbbd0c199),
	.w8(32'hbb65f6de),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4f5f2),
	.w1(32'h3b35e53f),
	.w2(32'h3ba7a094),
	.w3(32'hba916ba8),
	.w4(32'h39e159b7),
	.w5(32'h3b336c07),
	.w6(32'h3c049d64),
	.w7(32'h3b71e4c6),
	.w8(32'h3be6d02c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c24de),
	.w1(32'hbc446057),
	.w2(32'hbc0abbdc),
	.w3(32'h3a97e823),
	.w4(32'hbc5cf3b0),
	.w5(32'h3c881c6a),
	.w6(32'h3c62c66c),
	.w7(32'hbaf2d643),
	.w8(32'h3b97b02b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2037b),
	.w1(32'h3c44e5ef),
	.w2(32'h3bea4302),
	.w3(32'h3cd9bd4c),
	.w4(32'h3c6e2297),
	.w5(32'h3ba13da6),
	.w6(32'h3cc9b75c),
	.w7(32'h3cd2c3b4),
	.w8(32'h3c317747),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c93c2),
	.w1(32'hbbc5d4da),
	.w2(32'hbbdd8c1e),
	.w3(32'hbad27a0d),
	.w4(32'hbc09b8c8),
	.w5(32'hbbe8ff32),
	.w6(32'h3b11dceb),
	.w7(32'hb9c3df00),
	.w8(32'hbb3d2cb9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e475),
	.w1(32'h3b8b375a),
	.w2(32'h3a3b64c6),
	.w3(32'hbb5709e2),
	.w4(32'h3bdbd303),
	.w5(32'h3c3d3aee),
	.w6(32'h39b2fe57),
	.w7(32'h3b9b2f76),
	.w8(32'h3abc3e88),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd38e3),
	.w1(32'h3be04029),
	.w2(32'h3b06d32f),
	.w3(32'h3c486085),
	.w4(32'h3b9534a6),
	.w5(32'hbb3a2b3c),
	.w6(32'h3c515bbf),
	.w7(32'hbb01267d),
	.w8(32'hbb451bdf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f09fb),
	.w1(32'h3b221e91),
	.w2(32'hbbbc4d88),
	.w3(32'h3b937654),
	.w4(32'hba8e672b),
	.w5(32'hbbd37508),
	.w6(32'h3bea04b9),
	.w7(32'h39f0ddf2),
	.w8(32'h3b87d6d1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5120ba),
	.w1(32'h3b6dc282),
	.w2(32'h3bdf2343),
	.w3(32'hba7d078b),
	.w4(32'hbabb072e),
	.w5(32'h3ae37cce),
	.w6(32'h3a51e414),
	.w7(32'h3ae6ab0c),
	.w8(32'hbaea7fbe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04b283),
	.w1(32'hbaa7039f),
	.w2(32'hbb4feac2),
	.w3(32'h3c0251af),
	.w4(32'h3b800bc9),
	.w5(32'hbb867f09),
	.w6(32'h3c18d6bb),
	.w7(32'h3bfde4bf),
	.w8(32'hbc1c7954),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a67bb),
	.w1(32'h3b4ca37b),
	.w2(32'h39d8b517),
	.w3(32'h3ada29d2),
	.w4(32'hbb12241f),
	.w5(32'hbb811dea),
	.w6(32'hbbad18b2),
	.w7(32'h3b84d541),
	.w8(32'h3c13d79a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8751fc),
	.w1(32'hbb57b2bd),
	.w2(32'hbb9ced28),
	.w3(32'hbb8f6ad5),
	.w4(32'hbb3bae21),
	.w5(32'hbc3db4ca),
	.w6(32'hbab01766),
	.w7(32'hbb8044a9),
	.w8(32'hbbcbab04),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6890),
	.w1(32'h3bdc9daa),
	.w2(32'h398a3db2),
	.w3(32'hbb9d4694),
	.w4(32'hba426f99),
	.w5(32'hbad473c2),
	.w6(32'hbba84da3),
	.w7(32'hbbb0852b),
	.w8(32'hbba1752e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275b6d),
	.w1(32'h3ada8434),
	.w2(32'h3bb1dfac),
	.w3(32'h3a7d216e),
	.w4(32'h3b699381),
	.w5(32'hb8107c05),
	.w6(32'h3b8bdfe0),
	.w7(32'hbb6dfe4b),
	.w8(32'h3beddf71),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba236314),
	.w1(32'h3bb47ba5),
	.w2(32'h3ac3d4f3),
	.w3(32'h39d61736),
	.w4(32'h3b0bab99),
	.w5(32'h3ac8b8f3),
	.w6(32'hbae6d667),
	.w7(32'h3b221ec7),
	.w8(32'h3ba800ba),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b3e25),
	.w1(32'h3b4c5d86),
	.w2(32'h3b370f3a),
	.w3(32'hba245265),
	.w4(32'h3be6d51a),
	.w5(32'h3b8a9564),
	.w6(32'hb9015837),
	.w7(32'hba3d6360),
	.w8(32'h3b48173b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89309a),
	.w1(32'h3a8bf789),
	.w2(32'hbb043fc5),
	.w3(32'h3bf0589b),
	.w4(32'h3ab18a11),
	.w5(32'hbb8ca697),
	.w6(32'h3b8791e8),
	.w7(32'h3ab5957d),
	.w8(32'hbba427b6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b337d9d),
	.w1(32'hbb4c6106),
	.w2(32'hbba1c519),
	.w3(32'hbb214d0f),
	.w4(32'hbb42541f),
	.w5(32'hbbe707e9),
	.w6(32'hb9b0b7d2),
	.w7(32'h3b4cf82c),
	.w8(32'h3b76cec8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59a256),
	.w1(32'hbb5be053),
	.w2(32'hbc0ff79e),
	.w3(32'hbb5110da),
	.w4(32'h3b96cac3),
	.w5(32'h3b8f9f5b),
	.w6(32'hbb31ebc6),
	.w7(32'h3baac67a),
	.w8(32'hbbb16bf4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62005a),
	.w1(32'h3b55ec76),
	.w2(32'h3a9aa85b),
	.w3(32'hbaa1aef0),
	.w4(32'hba6b0598),
	.w5(32'h3b4e1bf1),
	.w6(32'hbc439b43),
	.w7(32'h3a8620aa),
	.w8(32'h3b898a60),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084a5d),
	.w1(32'h3ba2c2b5),
	.w2(32'h3a29e3f9),
	.w3(32'hbb753cd4),
	.w4(32'h39f396ec),
	.w5(32'h3a214b8d),
	.w6(32'h3b08ca4c),
	.w7(32'h3a0dc73a),
	.w8(32'hbb3189af),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0bd8),
	.w1(32'hbb3199da),
	.w2(32'hbb06344b),
	.w3(32'h3b50f4e4),
	.w4(32'hbc0ff260),
	.w5(32'hbc2537a8),
	.w6(32'h3a72c265),
	.w7(32'hbb75a6a9),
	.w8(32'h3aaa1edc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7831c),
	.w1(32'hbb51255d),
	.w2(32'hbba7bacd),
	.w3(32'hbbcc8169),
	.w4(32'h3ad6b76b),
	.w5(32'hbae8885b),
	.w6(32'h3a1a6858),
	.w7(32'h3bb79741),
	.w8(32'h3b66a272),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac70bc6),
	.w1(32'hbb78a893),
	.w2(32'hbb44750c),
	.w3(32'h3a6c2a2e),
	.w4(32'hbad35160),
	.w5(32'h3bb7a49d),
	.w6(32'h3ba621f3),
	.w7(32'h3b010607),
	.w8(32'h3c57735c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4475dc),
	.w1(32'hbb2add9e),
	.w2(32'hbb8b1285),
	.w3(32'hbb062855),
	.w4(32'hbab16bc8),
	.w5(32'hbb8a5714),
	.w6(32'h3bcadec9),
	.w7(32'hbb012490),
	.w8(32'h3b14675e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc206),
	.w1(32'hbb30ae50),
	.w2(32'hbb45c176),
	.w3(32'hbb8d1dd5),
	.w4(32'h39d46c11),
	.w5(32'hbb8b6592),
	.w6(32'hbba26013),
	.w7(32'hb89a1f9e),
	.w8(32'h3ac38f53),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefb5d0),
	.w1(32'hbb350c6a),
	.w2(32'hbb228f7f),
	.w3(32'hbb499a35),
	.w4(32'hbb83fccb),
	.w5(32'h3ab4a5b3),
	.w6(32'hbb7b8743),
	.w7(32'hbbce549c),
	.w8(32'hbb20602a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabd334),
	.w1(32'h3b2f5521),
	.w2(32'h3b961d4c),
	.w3(32'h39b77196),
	.w4(32'h3982f84a),
	.w5(32'h3b0a811f),
	.w6(32'h3a3691c2),
	.w7(32'hbb4ae72a),
	.w8(32'h3a5047b4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050ca3),
	.w1(32'hbabd3e29),
	.w2(32'hba536712),
	.w3(32'h3af7aab8),
	.w4(32'h3b810817),
	.w5(32'h3b04e6dc),
	.w6(32'hba001ed6),
	.w7(32'h38cd64c2),
	.w8(32'h3a947b71),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e249f),
	.w1(32'hbb98bf36),
	.w2(32'hbb56dd46),
	.w3(32'h3b0e88e8),
	.w4(32'h3b144a60),
	.w5(32'hbadc8914),
	.w6(32'h3ae73452),
	.w7(32'h3bc238bc),
	.w8(32'h39ed91a6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f150),
	.w1(32'h395ee50f),
	.w2(32'h3b9089b1),
	.w3(32'hbadaf782),
	.w4(32'hba7b77fc),
	.w5(32'h3b55b568),
	.w6(32'hb65c704b),
	.w7(32'hbb79adef),
	.w8(32'hbb0ab602),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb68b3c),
	.w1(32'h3b6ae83b),
	.w2(32'h3b7d2c49),
	.w3(32'h3b7ae28e),
	.w4(32'h3b2c4ce0),
	.w5(32'hbb51814f),
	.w6(32'h3b27d6d5),
	.w7(32'h3ae12eaf),
	.w8(32'hbbbe7a05),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ee8f),
	.w1(32'h3b1623a2),
	.w2(32'h3bb94d6c),
	.w3(32'h3b944579),
	.w4(32'h3c104a63),
	.w5(32'h3b415e51),
	.w6(32'h3c15a006),
	.w7(32'h3c12c467),
	.w8(32'h3b84d8c0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cb558),
	.w1(32'h3c0154e7),
	.w2(32'h3c231fa8),
	.w3(32'h3c7d033c),
	.w4(32'h3c1ad116),
	.w5(32'h3c71b0ef),
	.w6(32'h3c78db5c),
	.w7(32'h3be4b601),
	.w8(32'h3bacb2eb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eef5a),
	.w1(32'h3a9a9f5d),
	.w2(32'hbb2e4bb6),
	.w3(32'h3b46adef),
	.w4(32'hba61502e),
	.w5(32'hbb0bd506),
	.w6(32'h3b0a9d71),
	.w7(32'hbaa89956),
	.w8(32'hbb860788),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc280),
	.w1(32'hbacae65b),
	.w2(32'h3a24288f),
	.w3(32'hbbe40b8d),
	.w4(32'h3b26a728),
	.w5(32'h3c0c1e49),
	.w6(32'hbbf4875d),
	.w7(32'h3bb2e961),
	.w8(32'h3bda98ff),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c1ef),
	.w1(32'h3b06a8e0),
	.w2(32'h3b47b8c8),
	.w3(32'hb9e26b36),
	.w4(32'hbb4f2ba6),
	.w5(32'hbb4822ba),
	.w6(32'h39fa4c3a),
	.w7(32'hbbbde0ac),
	.w8(32'hbbb50928),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52a485),
	.w1(32'hbb6de1d9),
	.w2(32'hba954d36),
	.w3(32'h3a98d7ec),
	.w4(32'hbab69749),
	.w5(32'h3b209123),
	.w6(32'h38af739c),
	.w7(32'hba992709),
	.w8(32'hbae4cbc2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6436a),
	.w1(32'hbb503a49),
	.w2(32'hba8ebd7f),
	.w3(32'hbb85f850),
	.w4(32'hb966d801),
	.w5(32'h3a6a9b89),
	.w6(32'hbb7cc1ee),
	.w7(32'hbb0bb81d),
	.w8(32'hbb014712),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa2530),
	.w1(32'h3bcb4e10),
	.w2(32'h3b805583),
	.w3(32'hb95628e9),
	.w4(32'h3bd92a65),
	.w5(32'h3b0a8e8f),
	.w6(32'hbae5c447),
	.w7(32'h3ba943d4),
	.w8(32'hbae0d45e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadff360),
	.w1(32'h3b068d5c),
	.w2(32'h3b2d2464),
	.w3(32'hba8a5c7d),
	.w4(32'h3b2b3326),
	.w5(32'h3b651c81),
	.w6(32'hbb9f8d32),
	.w7(32'h3bc20ea7),
	.w8(32'h3b45a565),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144e25),
	.w1(32'h3b91c124),
	.w2(32'hbb3896c3),
	.w3(32'h3b39d6ea),
	.w4(32'h3b5b953d),
	.w5(32'hbb494719),
	.w6(32'hb9b0db17),
	.w7(32'h39481d9d),
	.w8(32'hbaddb515),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16348c),
	.w1(32'h3890aeac),
	.w2(32'hbbad7112),
	.w3(32'h3a3c4e44),
	.w4(32'hba332ad3),
	.w5(32'hbc00457d),
	.w6(32'h3a7bac55),
	.w7(32'hb757ccde),
	.w8(32'hbb1c6da9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ceac),
	.w1(32'hbb145d93),
	.w2(32'hbba4cf5c),
	.w3(32'hbbb2230a),
	.w4(32'hbbe422e8),
	.w5(32'hbc24f465),
	.w6(32'hbbf37a09),
	.w7(32'hbbdfc4f7),
	.w8(32'hbc29cb59),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6cdf7),
	.w1(32'hbaaf67ed),
	.w2(32'h3b0a2877),
	.w3(32'hbc0ae35a),
	.w4(32'hba74df5a),
	.w5(32'h3b7c69f6),
	.w6(32'hbbff6688),
	.w7(32'hbb7ac9c0),
	.w8(32'hba0e0573),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986e1b),
	.w1(32'h3b6da71e),
	.w2(32'h3c5a860b),
	.w3(32'h3bb5203b),
	.w4(32'h3918deeb),
	.w5(32'h3c79d85f),
	.w6(32'h3c6ade96),
	.w7(32'h3c27e188),
	.w8(32'h3b91d8ae),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c9ce4),
	.w1(32'hba9ef56c),
	.w2(32'h3aff33e8),
	.w3(32'h3c8a7d40),
	.w4(32'h3b08d2e8),
	.w5(32'h3bd0ba94),
	.w6(32'h3c63dda2),
	.w7(32'hb9caf1eb),
	.w8(32'h3b91f1ed),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea857),
	.w1(32'h3b6b77e8),
	.w2(32'h3b369bb8),
	.w3(32'hbb3b6281),
	.w4(32'hbb3e9f12),
	.w5(32'hbb43112b),
	.w6(32'h3a9fee9e),
	.w7(32'hbb2cc65d),
	.w8(32'hbb60e347),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9aad9),
	.w1(32'hbbe93a85),
	.w2(32'hbb332859),
	.w3(32'hbb9edd24),
	.w4(32'hbac61b60),
	.w5(32'h3b0a359a),
	.w6(32'hbb9b7ed1),
	.w7(32'hba520222),
	.w8(32'h3b0d7876),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10e46e),
	.w1(32'hbb89b7d8),
	.w2(32'hbb65087c),
	.w3(32'hbc32c07a),
	.w4(32'hbbfc369a),
	.w5(32'hbc05a992),
	.w6(32'hbbf958c2),
	.w7(32'hbc1c7ae5),
	.w8(32'hbbfb1366),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e0225),
	.w1(32'hbaa02550),
	.w2(32'hbb872777),
	.w3(32'hbb82d46c),
	.w4(32'hbb16f8bf),
	.w5(32'h3b8b1c36),
	.w6(32'hbbba6220),
	.w7(32'hbb87accd),
	.w8(32'h3b24014c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39bf3),
	.w1(32'hbbdef249),
	.w2(32'hbae3b188),
	.w3(32'hbad97d84),
	.w4(32'hbbfd08da),
	.w5(32'h3ade8a0b),
	.w6(32'hbb627a0b),
	.w7(32'hbba6d22b),
	.w8(32'hbb2cb1e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57887d),
	.w1(32'h3ab71bce),
	.w2(32'hbb22035f),
	.w3(32'hbbc18980),
	.w4(32'hbb1b95b9),
	.w5(32'hbb8adda1),
	.w6(32'hbb090996),
	.w7(32'hbb4f27e1),
	.w8(32'hbae5d5ce),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a280e33),
	.w1(32'h3b137528),
	.w2(32'h3c0c76c3),
	.w3(32'h3b962158),
	.w4(32'h3b13171f),
	.w5(32'h3c540a6b),
	.w6(32'h3b9f59fb),
	.w7(32'h3bd8017f),
	.w8(32'h3c1e69ef),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a119a3d),
	.w1(32'h3bce4909),
	.w2(32'h3c7f0152),
	.w3(32'h3bb2b219),
	.w4(32'h3c31f57a),
	.w5(32'h3d11b134),
	.w6(32'hb90d52b3),
	.w7(32'h3bff724e),
	.w8(32'h3cdf512a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0520d9),
	.w1(32'hba826d45),
	.w2(32'h3c156bad),
	.w3(32'h3ca5f352),
	.w4(32'h3b410424),
	.w5(32'h3a452b88),
	.w6(32'h3cded147),
	.w7(32'h3c96216d),
	.w8(32'h3b9bca5f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f14c),
	.w1(32'hbc02ebb2),
	.w2(32'hbb6fb460),
	.w3(32'hbc7ebeef),
	.w4(32'hbc10f0f0),
	.w5(32'hbaab5d1c),
	.w6(32'hbc8437d6),
	.w7(32'hbc5d87f0),
	.w8(32'h3b6d25ea),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f8f9),
	.w1(32'h398fda42),
	.w2(32'h3ab3583d),
	.w3(32'h3b8ccb35),
	.w4(32'h3ad7e5bc),
	.w5(32'h3bd84d83),
	.w6(32'h3bb07e9c),
	.w7(32'h3baa74df),
	.w8(32'h3bb5f87a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb561b5),
	.w1(32'hba3f0c81),
	.w2(32'h3b223cf9),
	.w3(32'hbb7b3992),
	.w4(32'hbb0974b7),
	.w5(32'h3aeee6bb),
	.w6(32'h39179a92),
	.w7(32'h39bd952c),
	.w8(32'hbbbc5685),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b20a2),
	.w1(32'h3b997504),
	.w2(32'h3bef381f),
	.w3(32'hbb65674e),
	.w4(32'hba887b2d),
	.w5(32'h3c1a5ce1),
	.w6(32'hbb5fb78d),
	.w7(32'hba633ef1),
	.w8(32'h3af8c95a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5220e0),
	.w1(32'h3c40a43b),
	.w2(32'h3c68b5df),
	.w3(32'h3cb52508),
	.w4(32'h3c53a70d),
	.w5(32'h3c346057),
	.w6(32'h3cc312d4),
	.w7(32'h3c83b281),
	.w8(32'h3c0cc61f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beed3d9),
	.w1(32'h3b12e5a1),
	.w2(32'h3b43d4dc),
	.w3(32'h3b6fe84c),
	.w4(32'h3b021782),
	.w5(32'h3b987953),
	.w6(32'h3a9389dc),
	.w7(32'hbad34079),
	.w8(32'h3a91e001),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb250210),
	.w1(32'h3a85efb8),
	.w2(32'hbad87b44),
	.w3(32'hbb699116),
	.w4(32'h3a5a8d08),
	.w5(32'h3ad7041f),
	.w6(32'hbba5c20e),
	.w7(32'hbabc13b2),
	.w8(32'hba8bca7a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ce421),
	.w1(32'h3b693e42),
	.w2(32'hbb286617),
	.w3(32'h3b698217),
	.w4(32'h3c1e1e8f),
	.w5(32'hbb08a099),
	.w6(32'h3ba1e19f),
	.w7(32'h3c805de8),
	.w8(32'h3bd2a109),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52ecd),
	.w1(32'h3c32df88),
	.w2(32'h3c34f876),
	.w3(32'h3b53fdd7),
	.w4(32'h3c3e1983),
	.w5(32'h3c43d8c7),
	.w6(32'h3bf020ed),
	.w7(32'h3c55685d),
	.w8(32'h3bdad597),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f49b),
	.w1(32'h3ada4dcd),
	.w2(32'h3a241146),
	.w3(32'h3bb89ab2),
	.w4(32'h38984f76),
	.w5(32'h3bd38bf1),
	.w6(32'h3b5f8cb4),
	.w7(32'hbb938532),
	.w8(32'h3c0b8ddf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff0fa9),
	.w1(32'h3ad29f4b),
	.w2(32'h3abdee94),
	.w3(32'h3abbc42c),
	.w4(32'hbbf869e1),
	.w5(32'hba114900),
	.w6(32'h3b933336),
	.w7(32'hbb0374a4),
	.w8(32'h3c134cfe),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9340a36),
	.w1(32'hbb3097dc),
	.w2(32'hba8d3be1),
	.w3(32'h3b559668),
	.w4(32'hbb9e355e),
	.w5(32'h3ad5eaa5),
	.w6(32'h3c1c899a),
	.w7(32'hbacc242a),
	.w8(32'h3b2fe4b7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adc602),
	.w1(32'hbac92e7f),
	.w2(32'hba81bbdd),
	.w3(32'h3b4381c8),
	.w4(32'h3a6ed741),
	.w5(32'hbb250a7b),
	.w6(32'h3b29c65d),
	.w7(32'h3b4deaa1),
	.w8(32'hbbaf5ca4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1079bb),
	.w1(32'hbb22b13a),
	.w2(32'hbacb4054),
	.w3(32'hbb2d56fb),
	.w4(32'hbae0a4fc),
	.w5(32'h3a56b4cf),
	.w6(32'hbbb00da5),
	.w7(32'h3b4cc706),
	.w8(32'h3be00aec),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb267ae0),
	.w1(32'h3b8fad9e),
	.w2(32'h3b9db8e4),
	.w3(32'h3b209ba5),
	.w4(32'h3bdeb87f),
	.w5(32'h3b899ba1),
	.w6(32'h3bda44c9),
	.w7(32'h3b3106fc),
	.w8(32'h3a958e9f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb026b66),
	.w1(32'hbb33d262),
	.w2(32'hbae0572c),
	.w3(32'hbb492935),
	.w4(32'hbb47d1aa),
	.w5(32'h39f1b17d),
	.w6(32'hbbf0fa3b),
	.w7(32'hbb3ba5ec),
	.w8(32'hb9b7f07d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964d1e),
	.w1(32'hbb9d2867),
	.w2(32'hba81d7d3),
	.w3(32'h3a9f243b),
	.w4(32'hbbc6b9a8),
	.w5(32'hbab0897f),
	.w6(32'h3a918e52),
	.w7(32'hbc2cf4a4),
	.w8(32'hbac5f63b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8711d2),
	.w1(32'h3b5da9a3),
	.w2(32'h3b95bfaa),
	.w3(32'h3b8bdd0b),
	.w4(32'h3acc225a),
	.w5(32'h3a644351),
	.w6(32'hba3341ff),
	.w7(32'hbb82f7bc),
	.w8(32'hbb62f25b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1de524),
	.w1(32'h3bbf4835),
	.w2(32'h3c245426),
	.w3(32'hba0afa83),
	.w4(32'h3b90b1fa),
	.w5(32'h3c1b6550),
	.w6(32'hbbae27c6),
	.w7(32'h3adc9862),
	.w8(32'h3b8fb8f6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48eb22),
	.w1(32'hbb0d0f11),
	.w2(32'hb9dd1150),
	.w3(32'h3bc9e8c9),
	.w4(32'h3afbfe5a),
	.w5(32'hb6852544),
	.w6(32'h3b7f5dde),
	.w7(32'h3b09d4a5),
	.w8(32'hba592817),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a4596),
	.w1(32'h3b1089f5),
	.w2(32'h3b69b288),
	.w3(32'hbb483518),
	.w4(32'h3bb167c4),
	.w5(32'h3bdbbfb5),
	.w6(32'hb9a5ff6e),
	.w7(32'h3af9bcc4),
	.w8(32'h3ba48693),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be26a8e),
	.w1(32'h3c12e8fd),
	.w2(32'h3c11e3ee),
	.w3(32'h3bdf6085),
	.w4(32'h3beea13f),
	.w5(32'h3a00373b),
	.w6(32'h3bc39562),
	.w7(32'h3b70c2c7),
	.w8(32'hbbd57067),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28e2a4),
	.w1(32'hbb7d2e6a),
	.w2(32'hbb90d9a9),
	.w3(32'hba78e410),
	.w4(32'hbb8431af),
	.w5(32'hbb346b2f),
	.w6(32'hbb6db7bf),
	.w7(32'hbabe24f4),
	.w8(32'h39b0f8b4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff8097),
	.w1(32'hbb85765a),
	.w2(32'hbbba7795),
	.w3(32'hbc0a515a),
	.w4(32'hbb130124),
	.w5(32'hbba87351),
	.w6(32'hbb9b3647),
	.w7(32'hbb2294f6),
	.w8(32'hbbd7ab51),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb37fa),
	.w1(32'h3b750bd2),
	.w2(32'h3c0713d2),
	.w3(32'hbc28541a),
	.w4(32'hbaa7b48f),
	.w5(32'hbacb1f55),
	.w6(32'hbc3a3e1d),
	.w7(32'hbab4e05b),
	.w8(32'hbb806928),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3ecaa),
	.w1(32'h3b77282a),
	.w2(32'h3ba63959),
	.w3(32'h3b9f2e20),
	.w4(32'h3b5def7d),
	.w5(32'h3c015035),
	.w6(32'hbb5a516c),
	.w7(32'hba4e2494),
	.w8(32'h3b686f62),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907cb74),
	.w1(32'h3bc4acbb),
	.w2(32'h3bee9404),
	.w3(32'h3b488e7c),
	.w4(32'h3bdc92f4),
	.w5(32'h3c0ef16a),
	.w6(32'h3a33f91a),
	.w7(32'h3b8a4f8a),
	.w8(32'h3c19056a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bd65a),
	.w1(32'hba079aac),
	.w2(32'hbb8571b1),
	.w3(32'h3b26efc1),
	.w4(32'hb95f1d2a),
	.w5(32'hb9cd4442),
	.w6(32'h3bf6f80e),
	.w7(32'hbb1c71b1),
	.w8(32'h3b9d26d9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b6659),
	.w1(32'h3b63a05f),
	.w2(32'h3b2f4d6f),
	.w3(32'h3b3a1f7e),
	.w4(32'h3aa6e01d),
	.w5(32'h3b835a69),
	.w6(32'h3c37f9cb),
	.w7(32'hba5c586b),
	.w8(32'hbaa67f7a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92b5ec),
	.w1(32'hbad7abe9),
	.w2(32'hbae17da6),
	.w3(32'h3b4ea085),
	.w4(32'h3b5aba00),
	.w5(32'h3b1c973b),
	.w6(32'h3acbae6f),
	.w7(32'h3bba2ce0),
	.w8(32'h3bc12e24),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c8ba9),
	.w1(32'h3ae31dab),
	.w2(32'h392366fc),
	.w3(32'h3b7edd4a),
	.w4(32'h3ac8ee3a),
	.w5(32'hb9466add),
	.w6(32'h3bbe140e),
	.w7(32'hbabbd497),
	.w8(32'h3adc4358),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5c5e),
	.w1(32'hb9b9e755),
	.w2(32'hba1ad822),
	.w3(32'h3b5b4fa2),
	.w4(32'h39bf1f89),
	.w5(32'hbbb18530),
	.w6(32'h3add7603),
	.w7(32'hba3e8ca9),
	.w8(32'hbbd1d77e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991390),
	.w1(32'hbb6c298d),
	.w2(32'hbb41a1e9),
	.w3(32'hbbaf44d9),
	.w4(32'hbbd3526f),
	.w5(32'hbbf91e1a),
	.w6(32'hbbdf3327),
	.w7(32'hbb93863f),
	.w8(32'hbbf9dcae),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ecf54),
	.w1(32'hbb98b6d8),
	.w2(32'hb8ee6cdb),
	.w3(32'hbbd0878d),
	.w4(32'hbadcab4a),
	.w5(32'h3b1a9f7c),
	.w6(32'hbbd13467),
	.w7(32'hbb4faa5e),
	.w8(32'h3b121625),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23577b),
	.w1(32'h3b607974),
	.w2(32'h3b9291cc),
	.w3(32'h3c3d9b1d),
	.w4(32'h3b8cfe7c),
	.w5(32'h3bb67044),
	.w6(32'h3c68907b),
	.w7(32'h3bad22bd),
	.w8(32'h3a0b379c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33cb08),
	.w1(32'hbc2964c1),
	.w2(32'hbb9625ee),
	.w3(32'hba36154a),
	.w4(32'hba19fc4a),
	.w5(32'h3b334411),
	.w6(32'hb9fe2e72),
	.w7(32'hbb82de76),
	.w8(32'h3a05f16e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750ebb),
	.w1(32'hbaedfd83),
	.w2(32'hba098086),
	.w3(32'h396d65b7),
	.w4(32'h3b189f3d),
	.w5(32'hb8ddda9e),
	.w6(32'h3b34fec2),
	.w7(32'h3b8b8033),
	.w8(32'hba2920d4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf15a5b),
	.w1(32'h3b858dbb),
	.w2(32'h3c1fd59e),
	.w3(32'hbb966cf3),
	.w4(32'hbb914307),
	.w5(32'hbbd26578),
	.w6(32'h3b02b07e),
	.w7(32'hbbb9922f),
	.w8(32'hbc288e12),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf93a7),
	.w1(32'hbbdc0726),
	.w2(32'hbbaf0378),
	.w3(32'hbbbdcf9b),
	.w4(32'hbbe56425),
	.w5(32'hbbb96b4a),
	.w6(32'hbc19f6e0),
	.w7(32'hbb3c35f7),
	.w8(32'hbb504fb4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fa534),
	.w1(32'h3b92a190),
	.w2(32'h3b810db6),
	.w3(32'hbbc1e619),
	.w4(32'h3b74d604),
	.w5(32'h3b4e10ce),
	.w6(32'hbb7de134),
	.w7(32'h3b2a0001),
	.w8(32'h3b5fe115),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b915e89),
	.w1(32'h3b62f9ba),
	.w2(32'h3b990aeb),
	.w3(32'h3b32a849),
	.w4(32'h3b64e51b),
	.w5(32'h3beaf80c),
	.w6(32'h3b87204d),
	.w7(32'h3b11842d),
	.w8(32'h39b8ec5d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb356941),
	.w1(32'h3a2d16fc),
	.w2(32'hba9072e4),
	.w3(32'hba9fba3c),
	.w4(32'hb92f3a28),
	.w5(32'h3ba1e5ad),
	.w6(32'hbc149d57),
	.w7(32'h3abeacf7),
	.w8(32'h3b7ca861),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ccbf),
	.w1(32'hbba57ec6),
	.w2(32'hbac7920b),
	.w3(32'hbb213672),
	.w4(32'hbbe63618),
	.w5(32'hbb07cf41),
	.w6(32'h39f867f3),
	.w7(32'hbbbbf9b3),
	.w8(32'hbb2f593e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c531),
	.w1(32'hba5704e2),
	.w2(32'hbb03dbe3),
	.w3(32'h3b625525),
	.w4(32'hbab9ca9d),
	.w5(32'h3a6a2446),
	.w6(32'hbb7e83e2),
	.w7(32'h3958c1d6),
	.w8(32'h3a944030),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3906a3),
	.w1(32'hba1c8cae),
	.w2(32'h3a294db5),
	.w3(32'h3a68d107),
	.w4(32'h3a544e78),
	.w5(32'h3acef7f3),
	.w6(32'hba3add37),
	.w7(32'h39c7314f),
	.w8(32'h3b385175),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2121e),
	.w1(32'hbb1d0e58),
	.w2(32'hbb272b28),
	.w3(32'h3b2b0ea4),
	.w4(32'hbb753da4),
	.w5(32'hb9dda47e),
	.w6(32'h3b53ad51),
	.w7(32'hba4fd1b6),
	.w8(32'h3ab9a946),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbed4dd),
	.w1(32'hba490745),
	.w2(32'hba01dbb8),
	.w3(32'hbbb44f79),
	.w4(32'hbb0b10c4),
	.w5(32'hbb47c87d),
	.w6(32'hbb784953),
	.w7(32'hbb37133b),
	.w8(32'hbb4694bc),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c647ce2),
	.w1(32'hb969217c),
	.w2(32'hbad72734),
	.w3(32'h3c3b613b),
	.w4(32'h3bff504f),
	.w5(32'hbb2d963c),
	.w6(32'h3c43e591),
	.w7(32'h3b95b477),
	.w8(32'h3a3a3b17),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3b37),
	.w1(32'h3ab0a824),
	.w2(32'hbac109f5),
	.w3(32'hbb2bb427),
	.w4(32'h3a2f444a),
	.w5(32'hbb186014),
	.w6(32'hbbb264fa),
	.w7(32'hba9c7bdc),
	.w8(32'hbb479185),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb39558),
	.w1(32'hba2603e4),
	.w2(32'hbb69040d),
	.w3(32'h3c506db6),
	.w4(32'hbaa38991),
	.w5(32'hbb8eec7f),
	.w6(32'h3c0d9f41),
	.w7(32'h3ad33929),
	.w8(32'hbac41ee8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba98a42),
	.w1(32'h3a5673df),
	.w2(32'hbb20ad4e),
	.w3(32'hb8a88f17),
	.w4(32'h39f15b96),
	.w5(32'h3a95e184),
	.w6(32'hbb85046e),
	.w7(32'h3a7f91e7),
	.w8(32'hb8f77f18),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84168c),
	.w1(32'h3be2b3cc),
	.w2(32'h3c3a27ee),
	.w3(32'hbaed5f3f),
	.w4(32'h3c42ea9d),
	.w5(32'h3bf82fad),
	.w6(32'h3ae4fec6),
	.w7(32'h3b5d4ee4),
	.w8(32'h3a9eccec),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961b6c1),
	.w1(32'hbad43333),
	.w2(32'h39eeeaba),
	.w3(32'hba066cc1),
	.w4(32'hbbf98cca),
	.w5(32'h3b045f3b),
	.w6(32'hbc075ba1),
	.w7(32'hbb684726),
	.w8(32'h3a53dc18),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7076d),
	.w1(32'hbbc06f8a),
	.w2(32'hbb7c7ad0),
	.w3(32'h3a4b9634),
	.w4(32'hbbd452fa),
	.w5(32'hbbb13955),
	.w6(32'h39f2ca61),
	.w7(32'hbb763dd3),
	.w8(32'hbb5d2b8d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8499),
	.w1(32'hba7926a4),
	.w2(32'hbc18eb32),
	.w3(32'hbabafa93),
	.w4(32'hbc065398),
	.w5(32'hbc2f6d92),
	.w6(32'hbb51d10f),
	.w7(32'hbc0e1cde),
	.w8(32'hbbf718cb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc16f0),
	.w1(32'h3c031687),
	.w2(32'h3bd5cd80),
	.w3(32'hbc10f87f),
	.w4(32'h3b9c5dea),
	.w5(32'h3a7a8945),
	.w6(32'hbbb4628f),
	.w7(32'hbac7bd0d),
	.w8(32'hbb86a14f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d816),
	.w1(32'hbb3b6687),
	.w2(32'hbb3d2599),
	.w3(32'hbc1c872a),
	.w4(32'hbbe91c0e),
	.w5(32'h3ae94d99),
	.w6(32'hbc23e6ed),
	.w7(32'hbc3999f2),
	.w8(32'hbb53456a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01f59f),
	.w1(32'hbb2e927b),
	.w2(32'hba8249a3),
	.w3(32'hb8dafe9e),
	.w4(32'hba6eee37),
	.w5(32'h3beeac21),
	.w6(32'hbb3f7463),
	.w7(32'hbb067989),
	.w8(32'h3b0eeb60),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8037ef),
	.w1(32'hbb0b90a1),
	.w2(32'hb999300f),
	.w3(32'h3b5e0739),
	.w4(32'h3b96a9cf),
	.w5(32'h3a42745f),
	.w6(32'h3bbd57ec),
	.w7(32'h3b1b89ed),
	.w8(32'h3b1dad65),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9195699),
	.w1(32'hbb273ae2),
	.w2(32'hb931b4ab),
	.w3(32'h3b47a36c),
	.w4(32'h3b4fccfc),
	.w5(32'h3b74591e),
	.w6(32'h3b12a704),
	.w7(32'hba09e350),
	.w8(32'h3988ec07),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e8c4b),
	.w1(32'h3a7a6cb0),
	.w2(32'h3b9096bc),
	.w3(32'h3abf3597),
	.w4(32'hbbabcb36),
	.w5(32'hbae8e639),
	.w6(32'h3b294acc),
	.w7(32'h39ce59a0),
	.w8(32'hbb1b303f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa21fb),
	.w1(32'h3bd75d27),
	.w2(32'h3c085442),
	.w3(32'hbaab902a),
	.w4(32'h3b9f50cb),
	.w5(32'h3c177335),
	.w6(32'h39eaf35f),
	.w7(32'hb8f86a87),
	.w8(32'hbb7759c8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b99af),
	.w1(32'hbac6f22c),
	.w2(32'h3afea5a7),
	.w3(32'hbaa7f242),
	.w4(32'hbad523f0),
	.w5(32'h3b55fcde),
	.w6(32'hbbdfbb4b),
	.w7(32'hbb27fcb3),
	.w8(32'hbbad2a93),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99743d),
	.w1(32'hbad0c68f),
	.w2(32'h3aabd138),
	.w3(32'hba6da03c),
	.w4(32'hbb122575),
	.w5(32'hbaab5b41),
	.w6(32'hbb793e14),
	.w7(32'hba7c85c7),
	.w8(32'hbb1a1ac5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7e104),
	.w1(32'h3b6519e8),
	.w2(32'hbb11c871),
	.w3(32'hbc480d54),
	.w4(32'h3a120b67),
	.w5(32'h3aca3e85),
	.w6(32'hbc0a2af6),
	.w7(32'h3ba940c3),
	.w8(32'h3b15cc64),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ff86),
	.w1(32'h3b0291fa),
	.w2(32'h3a689031),
	.w3(32'hbc3fc38b),
	.w4(32'h3bc9cc32),
	.w5(32'h3ba10760),
	.w6(32'hbc234159),
	.w7(32'h3b55b013),
	.w8(32'h3b777079),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa16bc7),
	.w1(32'hb992f7ee),
	.w2(32'hb9ff6b09),
	.w3(32'h39e7ae15),
	.w4(32'h3b8264dd),
	.w5(32'h3be6afd3),
	.w6(32'h393634a6),
	.w7(32'h3ba1a962),
	.w8(32'h3bf55da9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb0e0d),
	.w1(32'hbb9a128d),
	.w2(32'hbb2b98b9),
	.w3(32'hbbfc348d),
	.w4(32'hbbc780a0),
	.w5(32'hbc261677),
	.w6(32'hbbbaf3c1),
	.w7(32'hbc31a24e),
	.w8(32'hbc06ff53),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61815b),
	.w1(32'hbae103ac),
	.w2(32'h3ab96400),
	.w3(32'hbbc4c8be),
	.w4(32'hbaa14a39),
	.w5(32'h3ae0b6b8),
	.w6(32'hbb336128),
	.w7(32'hbbac3237),
	.w8(32'h3ac3da1c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8630d),
	.w1(32'hb6468902),
	.w2(32'hbb83181c),
	.w3(32'hbb70553c),
	.w4(32'hba24ec37),
	.w5(32'hbb8a356c),
	.w6(32'h39f1cafe),
	.w7(32'h3ab42233),
	.w8(32'hbabe6dd3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a68dc),
	.w1(32'h3b0d2b12),
	.w2(32'h3c3b11ab),
	.w3(32'hbb3f28e2),
	.w4(32'h3b87dc3d),
	.w5(32'h3c835c6f),
	.w6(32'hbb3fac7b),
	.w7(32'h3b11700c),
	.w8(32'h3c10818c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb88540),
	.w1(32'hbb9782d0),
	.w2(32'hba8955dc),
	.w3(32'h3c2f764f),
	.w4(32'hbb8dd299),
	.w5(32'hbb12226f),
	.w6(32'h3b98d4ce),
	.w7(32'hbbb3b11f),
	.w8(32'hba23d61e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be87735),
	.w1(32'h3bc2de99),
	.w2(32'h3a2282f6),
	.w3(32'h3ba918af),
	.w4(32'h3b07899a),
	.w5(32'hbb8aef36),
	.w6(32'h3c03cc9c),
	.w7(32'hb9e4e829),
	.w8(32'hbc20626e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba896ff8),
	.w1(32'h3ab933a9),
	.w2(32'h38ce122d),
	.w3(32'h39c82ebd),
	.w4(32'h3ac4448b),
	.w5(32'h3b9e9ced),
	.w6(32'h3b3c1eb5),
	.w7(32'h3b7079a9),
	.w8(32'h3b9bed65),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88138e),
	.w1(32'h3ba86a55),
	.w2(32'h3b6fca68),
	.w3(32'h3bad4ec7),
	.w4(32'h3b4d30a0),
	.w5(32'h3becac86),
	.w6(32'h3bfab5ef),
	.w7(32'h3b9eacc4),
	.w8(32'h3c54f190),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a4fb5),
	.w1(32'hbc04edc7),
	.w2(32'hbbc2192a),
	.w3(32'h3bacb1ac),
	.w4(32'hbb9a7aed),
	.w5(32'hba3f0098),
	.w6(32'h3c39b530),
	.w7(32'hbb85f8a9),
	.w8(32'h3a1d7a76),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09ccf5),
	.w1(32'hbbcd51ba),
	.w2(32'hbb432ef4),
	.w3(32'hbc04420b),
	.w4(32'hbc05c43e),
	.w5(32'hba90709f),
	.w6(32'hbbc0d99e),
	.w7(32'hbbd8edc4),
	.w8(32'h3ab9a13b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7257c),
	.w1(32'hbb710a7a),
	.w2(32'hbad90a85),
	.w3(32'h3b1a3e1a),
	.w4(32'h3be20509),
	.w5(32'h3b9a5f12),
	.w6(32'h3b577a55),
	.w7(32'h3b807df4),
	.w8(32'h3b4c68b8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fbdf2),
	.w1(32'hba93c9d0),
	.w2(32'h3b1dd5a1),
	.w3(32'hbb4b378c),
	.w4(32'h3a3d42a1),
	.w5(32'h3b3865b3),
	.w6(32'hbb9eb8bb),
	.w7(32'h3877c038),
	.w8(32'h3b434911),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03b1c4),
	.w1(32'h3a8583a8),
	.w2(32'h3a81ae6f),
	.w3(32'h3b38d318),
	.w4(32'h3bb5a90b),
	.w5(32'h3ab72710),
	.w6(32'hba96b90b),
	.w7(32'h3bb4deaa),
	.w8(32'h3b0941f0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d3e524),
	.w1(32'h3b3d91e9),
	.w2(32'h3b9a4202),
	.w3(32'h3bbe8b25),
	.w4(32'h3c0a12ac),
	.w5(32'h3bd8ddbf),
	.w6(32'h3bd529e5),
	.w7(32'h3bb12a0a),
	.w8(32'h3b21f2fe),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bec39d),
	.w1(32'h3b35562e),
	.w2(32'h3b90245e),
	.w3(32'hbb2d048c),
	.w4(32'h3b7c224b),
	.w5(32'h3bbc450f),
	.w6(32'hbb8f3d4c),
	.w7(32'hbb5b888a),
	.w8(32'hbb77d604),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a21c2),
	.w1(32'hbbbd90c3),
	.w2(32'hbbec86ea),
	.w3(32'h3b954b83),
	.w4(32'h3ad6aaed),
	.w5(32'hbb9ac00b),
	.w6(32'hba9a4162),
	.w7(32'h39f05800),
	.w8(32'hbb2cf773),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a30b),
	.w1(32'hba2c56ae),
	.w2(32'hbb34e625),
	.w3(32'hbc42cfd6),
	.w4(32'h39a6c0d5),
	.w5(32'h3a5b88ad),
	.w6(32'hbc1e145a),
	.w7(32'h3a452d7c),
	.w8(32'h3a8fed36),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fdf03),
	.w1(32'hbb4a4da7),
	.w2(32'h3a342862),
	.w3(32'hbac742fe),
	.w4(32'hbbe69f35),
	.w5(32'hbafd8cfd),
	.w6(32'hbb0ac9c2),
	.w7(32'hbbe9d6a0),
	.w8(32'hbbb5112a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814b1b),
	.w1(32'hba21fa38),
	.w2(32'h3a6dcffe),
	.w3(32'h3b2bb429),
	.w4(32'hba2cdbe2),
	.w5(32'hbb127f1a),
	.w6(32'h3b03679c),
	.w7(32'h3ac7386a),
	.w8(32'hbb888c4c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51b316),
	.w1(32'h3b5a89d4),
	.w2(32'h3b723837),
	.w3(32'h3b9c27b0),
	.w4(32'h3ba7cb0f),
	.w5(32'h3bb0cf28),
	.w6(32'h39e71723),
	.w7(32'hba111ab9),
	.w8(32'h3bbf2f1a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c834053),
	.w1(32'h3bb11613),
	.w2(32'hba997777),
	.w3(32'h3bc177f6),
	.w4(32'h3b394e31),
	.w5(32'hbc9e25c1),
	.w6(32'h3c00b1c5),
	.w7(32'hbb868a74),
	.w8(32'hbca3ca5d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a209d),
	.w1(32'hbc014f6a),
	.w2(32'hbbe45de3),
	.w3(32'hbc831429),
	.w4(32'hbb9ecaf4),
	.w5(32'h3b86b131),
	.w6(32'hbc9b2960),
	.w7(32'hba73ae20),
	.w8(32'h3cab5e9d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb811bc3),
	.w1(32'hb9066ef9),
	.w2(32'hb8366a1d),
	.w3(32'hbb015b8f),
	.w4(32'h3b693c56),
	.w5(32'hb964761d),
	.w6(32'h3bc7eb26),
	.w7(32'h3b8ce2c7),
	.w8(32'h3ae5642d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d231f9),
	.w1(32'h3b068186),
	.w2(32'h3b35aacd),
	.w3(32'hbad87792),
	.w4(32'h3ad7e932),
	.w5(32'hb96fab14),
	.w6(32'hbaf8fb6c),
	.w7(32'h3b42b6c1),
	.w8(32'h3a785398),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1203ec),
	.w1(32'h3ad2565c),
	.w2(32'h39c626c7),
	.w3(32'h3988a01b),
	.w4(32'h3aa4b24f),
	.w5(32'h389dd195),
	.w6(32'hb7121b87),
	.w7(32'hbb185168),
	.w8(32'hbb29dab5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b1152),
	.w1(32'hb8b002e2),
	.w2(32'h3a4d173e),
	.w3(32'hbb3a7d7e),
	.w4(32'hbad6d013),
	.w5(32'h391ed767),
	.w6(32'hbb3fcaec),
	.w7(32'hbb417cd8),
	.w8(32'hba594f88),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cedc5),
	.w1(32'h3b579411),
	.w2(32'h3ab9665a),
	.w3(32'hbb42351c),
	.w4(32'h3b8fd7e7),
	.w5(32'h3b64976b),
	.w6(32'hbbb911a0),
	.w7(32'h3bfd9a7e),
	.w8(32'h3b2945d5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3aea),
	.w1(32'hbbb1f255),
	.w2(32'hbb2719a2),
	.w3(32'hbafc9c89),
	.w4(32'hbbfa64d2),
	.w5(32'hb98f2c2a),
	.w6(32'h3b6c416a),
	.w7(32'h38d0263a),
	.w8(32'h3b506ca9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ff714),
	.w1(32'h3ba976ca),
	.w2(32'h3c098fcc),
	.w3(32'h3bda3c6c),
	.w4(32'h3bfb006f),
	.w5(32'h3d08b636),
	.w6(32'h3c30b0b4),
	.w7(32'h3c4cc463),
	.w8(32'h3cbea96b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8168fb),
	.w1(32'h3ba7c000),
	.w2(32'h3bca6292),
	.w3(32'h3c4d1887),
	.w4(32'h3c21f771),
	.w5(32'h3c3ac720),
	.w6(32'h3c8baff5),
	.w7(32'h3be8bb5b),
	.w8(32'h3c06d810),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45a2d6),
	.w1(32'h3b77ac6a),
	.w2(32'h3ac3b2c0),
	.w3(32'h3ad4c830),
	.w4(32'h3b2e3a9e),
	.w5(32'h3a815633),
	.w6(32'h39a1f03a),
	.w7(32'h3b63433d),
	.w8(32'hba048101),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4403b1),
	.w1(32'h3b2134af),
	.w2(32'h3a599a08),
	.w3(32'h3b31a505),
	.w4(32'h3af5a9aa),
	.w5(32'h3b24493b),
	.w6(32'h3b1d0ad6),
	.w7(32'h3afc4e73),
	.w8(32'h3973b457),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be8888),
	.w1(32'h39070b8c),
	.w2(32'h38239331),
	.w3(32'hba665cc4),
	.w4(32'h3a3a0531),
	.w5(32'h3b4b55f1),
	.w6(32'hbb01fbca),
	.w7(32'h3b0918ed),
	.w8(32'h3afd9eee),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2ba6d),
	.w1(32'h3b3cab5d),
	.w2(32'h3b0582c7),
	.w3(32'h3b0bd8fc),
	.w4(32'h3b1cbbcb),
	.w5(32'h3b0d9fe9),
	.w6(32'h3abf7bed),
	.w7(32'h3aa84ad0),
	.w8(32'h39d74bd0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21cc9f),
	.w1(32'hb9d447e7),
	.w2(32'hbaac949d),
	.w3(32'h39d60433),
	.w4(32'hba93165a),
	.w5(32'hba133a9e),
	.w6(32'hba328a73),
	.w7(32'h3871aa7a),
	.w8(32'h39f88a71),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853722),
	.w1(32'hbacf525f),
	.w2(32'hba09bb7a),
	.w3(32'h3aa8c1a5),
	.w4(32'hba525329),
	.w5(32'h3aa37762),
	.w6(32'h3b7c54cf),
	.w7(32'h3b453c7a),
	.w8(32'h3b8a0fb8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa3c4),
	.w1(32'hbbd494f7),
	.w2(32'hbb9e73c7),
	.w3(32'hbbedfda7),
	.w4(32'hbbea394e),
	.w5(32'hbb9fc5da),
	.w6(32'hbbe33bd9),
	.w7(32'hbbde5ab2),
	.w8(32'hbabbafc1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803fae),
	.w1(32'h3ab5f0a0),
	.w2(32'h3b53d51c),
	.w3(32'hbaba8d27),
	.w4(32'hba2ef6b2),
	.w5(32'h39c7cd01),
	.w6(32'hba079882),
	.w7(32'hba44a70a),
	.w8(32'h3ab54d66),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d20fd),
	.w1(32'hbaacec84),
	.w2(32'hba6b10cb),
	.w3(32'hba9047a8),
	.w4(32'hbafaca00),
	.w5(32'hbae176c6),
	.w6(32'h3936ef4b),
	.w7(32'hba9fda77),
	.w8(32'hbae340af),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361bc0),
	.w1(32'h3b35efc1),
	.w2(32'h3b993f49),
	.w3(32'hbb8b3370),
	.w4(32'h394462da),
	.w5(32'h3b876cc4),
	.w6(32'hbb31b572),
	.w7(32'h3ad0bcbd),
	.w8(32'h3b83654b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b4060),
	.w1(32'h3b058e42),
	.w2(32'h3aa1d3a1),
	.w3(32'h3b708152),
	.w4(32'h3acd482d),
	.w5(32'h39d51e0d),
	.w6(32'h3bab6048),
	.w7(32'h3aa24532),
	.w8(32'hbac7b46f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5f4d2),
	.w1(32'h3c3da4d0),
	.w2(32'h3c1f098f),
	.w3(32'h3c4a0189),
	.w4(32'h3c3f00fc),
	.w5(32'h3bdf3574),
	.w6(32'h3c5bf76b),
	.w7(32'h3c8273e2),
	.w8(32'h3bdcdb91),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b955565),
	.w1(32'hba10342f),
	.w2(32'h3a1a3e5d),
	.w3(32'h3b94357c),
	.w4(32'hb9d2b5f1),
	.w5(32'h3a821eca),
	.w6(32'h3ba09d9e),
	.w7(32'hba11b151),
	.w8(32'h3a13b416),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aabdf),
	.w1(32'h3a812a7f),
	.w2(32'h3a11cd00),
	.w3(32'h3aad397f),
	.w4(32'h3a575e53),
	.w5(32'h3a214bcd),
	.w6(32'h3a9d8551),
	.w7(32'h39d29d75),
	.w8(32'hba734e29),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25bd7a),
	.w1(32'hbac76c72),
	.w2(32'h3b085a01),
	.w3(32'hbaaad9d2),
	.w4(32'hb98a987a),
	.w5(32'h3b8a636b),
	.w6(32'h3af21e8b),
	.w7(32'h3b59d72d),
	.w8(32'h3b982eee),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b7b5),
	.w1(32'hb9c4268a),
	.w2(32'h3a418896),
	.w3(32'h3aa379e7),
	.w4(32'hbb363da8),
	.w5(32'hbabdde77),
	.w6(32'h3ba4b69b),
	.w7(32'hbaaba2c6),
	.w8(32'h396182e9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d68bbd),
	.w1(32'hba95950e),
	.w2(32'hbb02133a),
	.w3(32'hba2b6298),
	.w4(32'hba452380),
	.w5(32'h3aa2416b),
	.w6(32'hb9f9dfa6),
	.w7(32'hbaaff079),
	.w8(32'h3a9f0e38),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a4687),
	.w1(32'hbad4d370),
	.w2(32'hbb33aa87),
	.w3(32'hbae31f79),
	.w4(32'hbb055fe6),
	.w5(32'hbb909e53),
	.w6(32'hb8d542a4),
	.w7(32'hbad14c42),
	.w8(32'hbb67c1ee),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cd403),
	.w1(32'hba5a6b73),
	.w2(32'hba84a408),
	.w3(32'hbb160a3a),
	.w4(32'hbacfb008),
	.w5(32'h3b02023f),
	.w6(32'hbb186b83),
	.w7(32'hba2563ec),
	.w8(32'hb9ef494a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361e05),
	.w1(32'h3a505274),
	.w2(32'hb92607b6),
	.w3(32'h3a10f95a),
	.w4(32'h3a32b445),
	.w5(32'h39e1c069),
	.w6(32'hba91661b),
	.w7(32'h3a404f24),
	.w8(32'hb901286b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96996d6),
	.w1(32'hbb7a566f),
	.w2(32'h3a530818),
	.w3(32'h3a808f96),
	.w4(32'hba2c85d4),
	.w5(32'hba22d3a8),
	.w6(32'h3b634be9),
	.w7(32'h3a24738f),
	.w8(32'hba1805c9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fe694),
	.w1(32'h3bc8dbae),
	.w2(32'h3b35fb7f),
	.w3(32'h3be565a2),
	.w4(32'h3b332251),
	.w5(32'hbbbfd754),
	.w6(32'h3c2d6848),
	.w7(32'h3b1cee74),
	.w8(32'hbbde4c89),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26f0e2),
	.w1(32'h3b0cb974),
	.w2(32'h3b6d95c0),
	.w3(32'h3baab9ea),
	.w4(32'h3b9edb73),
	.w5(32'h3b846778),
	.w6(32'h3c15a4f9),
	.w7(32'h3bc9d3d6),
	.w8(32'h3b859ad2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fe46c9),
	.w1(32'hbac45783),
	.w2(32'hbaac211c),
	.w3(32'hba50c615),
	.w4(32'hbb151d57),
	.w5(32'h39346c93),
	.w6(32'hba9b44ea),
	.w7(32'hba792a42),
	.w8(32'h3a75e084),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09104f),
	.w1(32'hb908bd24),
	.w2(32'h39364710),
	.w3(32'hbb08f390),
	.w4(32'hbb3857f6),
	.w5(32'hba008fad),
	.w6(32'hbb2f0139),
	.w7(32'hbaa69f6d),
	.w8(32'h3adc0376),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fedcc),
	.w1(32'hba87a8e0),
	.w2(32'hbaf849c7),
	.w3(32'h39c5dc1e),
	.w4(32'hb9e8a0e7),
	.w5(32'hba6c6f5f),
	.w6(32'h3b0092e0),
	.w7(32'h3a5d0ee9),
	.w8(32'hba82f22b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e2efc),
	.w1(32'hb96c3135),
	.w2(32'hbad147b8),
	.w3(32'h3a160599),
	.w4(32'hba193e12),
	.w5(32'h3ab90707),
	.w6(32'hba646d39),
	.w7(32'hb9c69354),
	.w8(32'hba7b40fd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c9443),
	.w1(32'hbab2db4b),
	.w2(32'hbb24df20),
	.w3(32'h39ab296a),
	.w4(32'hbace784a),
	.w5(32'h3a362183),
	.w6(32'hbaad234d),
	.w7(32'h3a2d81dc),
	.w8(32'h3ae74db5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38bd96),
	.w1(32'hba717012),
	.w2(32'h3aab8f13),
	.w3(32'h3a831e1c),
	.w4(32'hba88659c),
	.w5(32'h3ac574c0),
	.w6(32'h3a152710),
	.w7(32'hbadb7b44),
	.w8(32'h37e1191d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1855fc),
	.w1(32'hbaaf5859),
	.w2(32'hba0d3a29),
	.w3(32'h3a60c702),
	.w4(32'hba41b69c),
	.w5(32'hb9f2efb8),
	.w6(32'h3a5dda83),
	.w7(32'hbae09d45),
	.w8(32'hbac4c6d5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba871b9d),
	.w1(32'h3a0a5d06),
	.w2(32'h3b63df20),
	.w3(32'hbab3f3c4),
	.w4(32'hba28b27b),
	.w5(32'h38af2ca2),
	.w6(32'hb8aafb45),
	.w7(32'h39b32973),
	.w8(32'h3b8b5b6f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa777ee),
	.w1(32'h3a95db30),
	.w2(32'h3af85913),
	.w3(32'hbaf3d22b),
	.w4(32'hba372c83),
	.w5(32'h3a84c1e5),
	.w6(32'h3a8a2914),
	.w7(32'h3ab85fec),
	.w8(32'h3b5ba920),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5507b0),
	.w1(32'h3a0521a1),
	.w2(32'hb9a9c498),
	.w3(32'hb96d0475),
	.w4(32'hba2dfdac),
	.w5(32'hba521858),
	.w6(32'hb8a79683),
	.w7(32'hba42a9e4),
	.w8(32'hbad6604e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9141d0),
	.w1(32'h39f9625b),
	.w2(32'h3b85d177),
	.w3(32'h3bff2750),
	.w4(32'h3b0f6249),
	.w5(32'h3b76bfa1),
	.w6(32'h3c2d6bbf),
	.w7(32'h3bab6c72),
	.w8(32'h39de8093),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ea86),
	.w1(32'hbb040184),
	.w2(32'hba107043),
	.w3(32'h3b2a04c0),
	.w4(32'hbb0331a4),
	.w5(32'hba907e53),
	.w6(32'h3ace7d26),
	.w7(32'h391bb56c),
	.w8(32'hba1f9f4c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02e726),
	.w1(32'h3b079d80),
	.w2(32'h3acfc2aa),
	.w3(32'hb9e9cd86),
	.w4(32'h3ade1997),
	.w5(32'h3b293949),
	.w6(32'hba6b60b5),
	.w7(32'h39e377aa),
	.w8(32'h3a1c00f9),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b263f15),
	.w1(32'h3b4caf56),
	.w2(32'h3b01c18c),
	.w3(32'h3b7b05e0),
	.w4(32'h3b4d04a8),
	.w5(32'h3a4ba127),
	.w6(32'h3b97dc0e),
	.w7(32'h3b6b04b7),
	.w8(32'h3ace3e33),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81d9c8),
	.w1(32'h38ede92b),
	.w2(32'hb8bb7fec),
	.w3(32'h3aa52859),
	.w4(32'h398f6620),
	.w5(32'hb6542b6c),
	.w6(32'h3a962abe),
	.w7(32'hb9ecba2d),
	.w8(32'hb9e67011),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ca41a),
	.w1(32'h3a47954a),
	.w2(32'hba865a77),
	.w3(32'hba1419f6),
	.w4(32'h38c28f3e),
	.w5(32'hbaa7bc62),
	.w6(32'h39e104ea),
	.w7(32'hb9f604f3),
	.w8(32'hbb1c2a7b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9425ff),
	.w1(32'hba081d96),
	.w2(32'hbab463e9),
	.w3(32'hbad08168),
	.w4(32'hba59b7e8),
	.w5(32'hba6359ec),
	.w6(32'hbad3c750),
	.w7(32'hbaa9d083),
	.w8(32'hba9c9f63),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba067735),
	.w1(32'hba7b412f),
	.w2(32'hb9a382d6),
	.w3(32'hba3ccc91),
	.w4(32'hba5839a3),
	.w5(32'hbac32716),
	.w6(32'hba2e201d),
	.w7(32'hb9d2f3cf),
	.w8(32'hba43cd89),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39683e89),
	.w1(32'hb7887ebd),
	.w2(32'hb90d9094),
	.w3(32'hba66d64b),
	.w4(32'hba999b03),
	.w5(32'h3918d3b2),
	.w6(32'hb8e64ebb),
	.w7(32'hba2f2df7),
	.w8(32'h388b875b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a6247),
	.w1(32'h3afd9468),
	.w2(32'h3b4503be),
	.w3(32'hb9478102),
	.w4(32'hbaca1eb1),
	.w5(32'h3a75def7),
	.w6(32'h3b6a8fa6),
	.w7(32'hba7ec577),
	.w8(32'h3a2ce2ad),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a332ba9),
	.w1(32'h3a68f761),
	.w2(32'h3a70bb9d),
	.w3(32'hba4b671f),
	.w4(32'hbb1f0394),
	.w5(32'hba04728c),
	.w6(32'hba8cc2eb),
	.w7(32'hbb0735c4),
	.w8(32'hba627af9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3970b),
	.w1(32'hb95c68bc),
	.w2(32'hbb064d12),
	.w3(32'h3bd9ad07),
	.w4(32'h3a619591),
	.w5(32'hbb867f96),
	.w6(32'h3b8720f9),
	.w7(32'h3a9dbb61),
	.w8(32'hbb879e5b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27da90),
	.w1(32'h39831580),
	.w2(32'h3adf8d98),
	.w3(32'hbb48b130),
	.w4(32'h3938b0a7),
	.w5(32'hb905844b),
	.w6(32'hb9e21cef),
	.w7(32'h3a5d1f34),
	.w8(32'h39b4395e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39931b3d),
	.w1(32'h3ab940f4),
	.w2(32'h3a9c672f),
	.w3(32'hba038140),
	.w4(32'h3ab68164),
	.w5(32'h3ab06a98),
	.w6(32'h37e98956),
	.w7(32'h3a73bbe7),
	.w8(32'h3a2fa7c2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49af45),
	.w1(32'hb9615d3c),
	.w2(32'h3883b478),
	.w3(32'h39ae922f),
	.w4(32'h3a0028de),
	.w5(32'hbaa51526),
	.w6(32'h3a06a5f3),
	.w7(32'hb8a0e485),
	.w8(32'hba54d7b6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd47ab),
	.w1(32'hb8c0c3a5),
	.w2(32'hb9c7e2d4),
	.w3(32'hba344656),
	.w4(32'h39fae2a7),
	.w5(32'hba4fae33),
	.w6(32'hb9297db5),
	.w7(32'hb8448054),
	.w8(32'hb86a982a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4109d8),
	.w1(32'hbb190b78),
	.w2(32'hbb20cca6),
	.w3(32'hbac2026a),
	.w4(32'hbb89c633),
	.w5(32'hbabdb406),
	.w6(32'hb91b4ef4),
	.w7(32'hbb65d160),
	.w8(32'hbb0ef290),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf29a59),
	.w1(32'hbacfcba7),
	.w2(32'hb9e20e7c),
	.w3(32'hbb1f457b),
	.w4(32'hbacd816b),
	.w5(32'h3a1784c1),
	.w6(32'hbb46db86),
	.w7(32'hba0e6e1c),
	.w8(32'hba6f772c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3218c5),
	.w1(32'h3a68c56e),
	.w2(32'h3ac7e9d7),
	.w3(32'h3a0a07ab),
	.w4(32'h3a9277af),
	.w5(32'h3ab21421),
	.w6(32'hb729644f),
	.w7(32'h3b0b4095),
	.w8(32'h3b56b526),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a519d0e),
	.w1(32'h39feb833),
	.w2(32'hbb1af707),
	.w3(32'h39e9b077),
	.w4(32'hb9d25a48),
	.w5(32'hba2eb63b),
	.w6(32'h3a2a7ed8),
	.w7(32'hba76e96b),
	.w8(32'hbaf374a3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9207c7),
	.w1(32'hb89006ba),
	.w2(32'h396f047f),
	.w3(32'hbacbd5b0),
	.w4(32'hb9c0abb5),
	.w5(32'h3b2d678a),
	.w6(32'hb8063eba),
	.w7(32'h3a589a6d),
	.w8(32'h3ab40237),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c0161),
	.w1(32'h3a14b4ba),
	.w2(32'h3afc7f22),
	.w3(32'h3b3fe046),
	.w4(32'h3adb00ea),
	.w5(32'h3af0a01b),
	.w6(32'h3b92d649),
	.w7(32'h3b589114),
	.w8(32'h3aaaae7a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add8ba0),
	.w1(32'hb9238e7c),
	.w2(32'hba9ee192),
	.w3(32'h3b0ec2de),
	.w4(32'h3a0f0f8e),
	.w5(32'h39c39276),
	.w6(32'h3b05813f),
	.w7(32'hba6b57f9),
	.w8(32'hb990c7e0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0080ba),
	.w1(32'hba3f45ae),
	.w2(32'hba47bbd8),
	.w3(32'h38d1c540),
	.w4(32'hbb0ad45b),
	.w5(32'hb9aa7443),
	.w6(32'h3b03e480),
	.w7(32'hba1954df),
	.w8(32'hb9b4a272),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6bf3a),
	.w1(32'hbb0c94d6),
	.w2(32'hba4ce96c),
	.w3(32'hb8f8e667),
	.w4(32'hbaddae11),
	.w5(32'hbb639670),
	.w6(32'h3af4b538),
	.w7(32'hbb3dc95d),
	.w8(32'hbb9e2912),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70700c),
	.w1(32'hbbadeb0f),
	.w2(32'hbbfead04),
	.w3(32'hbbdba04e),
	.w4(32'hbba404ad),
	.w5(32'hbb57e7ef),
	.w6(32'hbb756a0b),
	.w7(32'hbad29884),
	.w8(32'hba3c2d67),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule