module layer_10_featuremap_452(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0406a3),
	.w1(32'h3b9082c4),
	.w2(32'h3ba69676),
	.w3(32'hbbcfce61),
	.w4(32'h3c18aa91),
	.w5(32'hb8c4e5af),
	.w6(32'hbae9c963),
	.w7(32'hbb69ce55),
	.w8(32'hbc374d54),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26dc65),
	.w1(32'hbc31a756),
	.w2(32'hbc4c0233),
	.w3(32'hbb20dd79),
	.w4(32'hbb7b023b),
	.w5(32'h3b3acdc3),
	.w6(32'hbbb0de6e),
	.w7(32'h39b55a9a),
	.w8(32'h3b4903c4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a804c),
	.w1(32'h38ece1dd),
	.w2(32'h3ab5abd6),
	.w3(32'hbb488ce5),
	.w4(32'hbad4e2da),
	.w5(32'hbbfc78f9),
	.w6(32'h3a212cd8),
	.w7(32'hbb37d711),
	.w8(32'hbbf51a60),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8ca8f),
	.w1(32'hbbb58a21),
	.w2(32'hbc46d5d3),
	.w3(32'hbbeb3ee3),
	.w4(32'hbc064c24),
	.w5(32'h3c092632),
	.w6(32'hbb43d687),
	.w7(32'hbb6394c0),
	.w8(32'h3ba3bc4e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb44ea2),
	.w1(32'h3bc8edf2),
	.w2(32'h3b27761a),
	.w3(32'h3c38af6b),
	.w4(32'h3bac3c81),
	.w5(32'hbc01a24b),
	.w6(32'hbbd0a0ca),
	.w7(32'h3b74e339),
	.w8(32'hba506911),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6768f0),
	.w1(32'hbba26ac6),
	.w2(32'hbb864bb5),
	.w3(32'hb9e9a904),
	.w4(32'hbb5cd5e5),
	.w5(32'h3b90a27e),
	.w6(32'h3b406780),
	.w7(32'hbac4c8b0),
	.w8(32'hb9f0e4dc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad722aa),
	.w1(32'h3b881a8f),
	.w2(32'h3c42ee75),
	.w3(32'h3c0bd182),
	.w4(32'hbae438e1),
	.w5(32'h3ca284c0),
	.w6(32'hba1dec60),
	.w7(32'h3c8ea8cc),
	.w8(32'h3c3b9f37),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe33e8b),
	.w1(32'h3c9a2963),
	.w2(32'h3bf6c54d),
	.w3(32'h3c16930c),
	.w4(32'hbc2f8ff8),
	.w5(32'hbc320a3b),
	.w6(32'h3c87e720),
	.w7(32'h3b35ec6a),
	.w8(32'h3b812bed),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b040f81),
	.w1(32'hbaf4e19d),
	.w2(32'hbb958920),
	.w3(32'h3beabf06),
	.w4(32'hb9d0289a),
	.w5(32'h3b1df1b5),
	.w6(32'h3bf54a10),
	.w7(32'hb99fc77b),
	.w8(32'hbaf40565),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ebced),
	.w1(32'h3bf6b737),
	.w2(32'h3b49815c),
	.w3(32'hbbf95317),
	.w4(32'hbbd81626),
	.w5(32'h3b429d5b),
	.w6(32'hbc1f25b6),
	.w7(32'hbb7d833c),
	.w8(32'h3bbe8d48),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbd7a0),
	.w1(32'h3b20d464),
	.w2(32'hbbd67034),
	.w3(32'h3c0ca74d),
	.w4(32'h3bef9c67),
	.w5(32'h3bd0c5a4),
	.w6(32'h3ba91376),
	.w7(32'h3ba0472a),
	.w8(32'h3a88bc8c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb113bce),
	.w1(32'h3b64f585),
	.w2(32'h3cc0c54f),
	.w3(32'h3b3a8bde),
	.w4(32'h3c384e4b),
	.w5(32'h3ba1d19a),
	.w6(32'hba1d36d3),
	.w7(32'h3b92d316),
	.w8(32'h3bd957d0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc9dbb),
	.w1(32'h3c306758),
	.w2(32'h3be32734),
	.w3(32'hbc9aba2f),
	.w4(32'hbb17e55b),
	.w5(32'h3bbcedf7),
	.w6(32'hba9a6b5f),
	.w7(32'h3bc21ea8),
	.w8(32'h3b881344),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e426),
	.w1(32'h3c60c6c7),
	.w2(32'h3baebe5e),
	.w3(32'hbaab4059),
	.w4(32'h3a289497),
	.w5(32'hbbec962d),
	.w6(32'h3bac9719),
	.w7(32'h3c23185c),
	.w8(32'hbc07b3e1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa07374),
	.w1(32'hbc000bb4),
	.w2(32'hbbc0ef95),
	.w3(32'hbb63433d),
	.w4(32'h3b521739),
	.w5(32'hbbc7bf7a),
	.w6(32'hbb42dd85),
	.w7(32'hbaa73b76),
	.w8(32'hbbc424e2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15aaa8),
	.w1(32'h3c3d4bf4),
	.w2(32'h3bfdc9db),
	.w3(32'hbc13d4de),
	.w4(32'h3b1bb124),
	.w5(32'hbc0419fb),
	.w6(32'hbbbcc223),
	.w7(32'hbb470654),
	.w8(32'hbc99f7cf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1834e5),
	.w1(32'hbbbf9ab3),
	.w2(32'hbbd066ec),
	.w3(32'hbc46d6ec),
	.w4(32'hbb8fa2cf),
	.w5(32'hbba12193),
	.w6(32'hbbc89d58),
	.w7(32'hbba341cb),
	.w8(32'hbaeb64d9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4752),
	.w1(32'h3c6b3577),
	.w2(32'h3c472c05),
	.w3(32'hbc9478e9),
	.w4(32'h3c5a609e),
	.w5(32'h3cb77c1f),
	.w6(32'hbc1f0db7),
	.w7(32'h3a921664),
	.w8(32'hbc2a5041),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ed129),
	.w1(32'h3c050298),
	.w2(32'h3a4d5942),
	.w3(32'hb960d105),
	.w4(32'h3a4686af),
	.w5(32'hbba7049b),
	.w6(32'hbc8c0862),
	.w7(32'hbb9e264a),
	.w8(32'hbb3336ee),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81badd),
	.w1(32'hb9faf533),
	.w2(32'h3c027185),
	.w3(32'hbc63e383),
	.w4(32'h3c2ceec7),
	.w5(32'h3c8f58c4),
	.w6(32'hbb64373a),
	.w7(32'hbb23ac0a),
	.w8(32'hba267a90),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873ac9),
	.w1(32'h3b82f54c),
	.w2(32'hbb354bb4),
	.w3(32'h3b263f2e),
	.w4(32'hbb4c6f9d),
	.w5(32'hbc282c77),
	.w6(32'hbbe3ff70),
	.w7(32'hbade4c0d),
	.w8(32'h3af50715),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d1e04),
	.w1(32'hbbc12ac1),
	.w2(32'h3b149891),
	.w3(32'h39f444b5),
	.w4(32'hbbcf86c7),
	.w5(32'h3b658f21),
	.w6(32'h3c933f2a),
	.w7(32'h3ae1c720),
	.w8(32'h3c3b4f43),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c838732),
	.w1(32'hbb69003b),
	.w2(32'hb910cf34),
	.w3(32'hba0baf86),
	.w4(32'hbb778db4),
	.w5(32'h3d1255a9),
	.w6(32'hbb8258a0),
	.w7(32'h3be03f93),
	.w8(32'h3c2124c6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b352576),
	.w1(32'hb9fea8de),
	.w2(32'hbb34ace1),
	.w3(32'h3be01f30),
	.w4(32'h3b9a7f2e),
	.w5(32'h39a05461),
	.w6(32'hbabb6222),
	.w7(32'hb9455305),
	.w8(32'hbb1302e6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e237),
	.w1(32'hbc97e5e0),
	.w2(32'hbcfd3dab),
	.w3(32'h3c150baa),
	.w4(32'hbc22a637),
	.w5(32'h3c586d9e),
	.w6(32'h3c0bbac5),
	.w7(32'hbbe46b1f),
	.w8(32'h3a1ad2eb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97345c),
	.w1(32'hbbc51d78),
	.w2(32'hbbeaf86a),
	.w3(32'h3b165345),
	.w4(32'hbb3e4714),
	.w5(32'hbb9b2d2a),
	.w6(32'hbbcc4da6),
	.w7(32'h3b93ed78),
	.w8(32'h3cc54f63),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1580d4),
	.w1(32'hb8acf857),
	.w2(32'h3afd03ea),
	.w3(32'h3ca97c9e),
	.w4(32'hbbac36eb),
	.w5(32'h3bc2565b),
	.w6(32'h3c940b14),
	.w7(32'hbbabdc4a),
	.w8(32'hbb2a61a2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39bf8d),
	.w1(32'h3bfca2ec),
	.w2(32'hbaaa321b),
	.w3(32'hbbd9dc86),
	.w4(32'h3c2f9288),
	.w5(32'h3c8ad6e8),
	.w6(32'hbb8563d9),
	.w7(32'hbb802987),
	.w8(32'h3c260905),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc716),
	.w1(32'hbb34ebda),
	.w2(32'h3c417f00),
	.w3(32'h3c212897),
	.w4(32'h3c4d0790),
	.w5(32'h3d1fcd29),
	.w6(32'hba3ab468),
	.w7(32'h3b277135),
	.w8(32'hbbba2e8f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe2b28),
	.w1(32'hbc1c9b3e),
	.w2(32'hbc5a826f),
	.w3(32'hbb6b56a6),
	.w4(32'h3c4a525d),
	.w5(32'hbc3056d8),
	.w6(32'hbb02c40e),
	.w7(32'h3bde3951),
	.w8(32'h3baea6d6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37ec2),
	.w1(32'hbb69141f),
	.w2(32'hbaae3d18),
	.w3(32'hb9daafbd),
	.w4(32'h3c76d131),
	.w5(32'h3c632e0b),
	.w6(32'h3c0b495b),
	.w7(32'h3b297533),
	.w8(32'hba8adfb1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c248337),
	.w1(32'hbb88666f),
	.w2(32'hb81fd426),
	.w3(32'hbc694280),
	.w4(32'hbb883dc5),
	.w5(32'hbba61add),
	.w6(32'hbb8f42ef),
	.w7(32'hba9ed96f),
	.w8(32'hba8a4653),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb761e7e),
	.w1(32'hbb2270a7),
	.w2(32'hbb3c6b18),
	.w3(32'hbb9d073b),
	.w4(32'hbb4ec537),
	.w5(32'hbbfddf84),
	.w6(32'hbbba4e24),
	.w7(32'h3c073470),
	.w8(32'h3c20f543),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acba9),
	.w1(32'hbc2ac4ab),
	.w2(32'hbbb9997a),
	.w3(32'h3b094f03),
	.w4(32'hbad06bf3),
	.w5(32'h3bba1a81),
	.w6(32'h3c44d392),
	.w7(32'h3b1bafa1),
	.w8(32'h3b1cb0d5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b7cd),
	.w1(32'h3b9e19cc),
	.w2(32'h3b31866a),
	.w3(32'h3bd68976),
	.w4(32'hbad300fd),
	.w5(32'hbbad84f5),
	.w6(32'hb96560ba),
	.w7(32'h3b2eef9e),
	.w8(32'h3c2134e3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060745),
	.w1(32'hba1fbbca),
	.w2(32'h3bf8db6f),
	.w3(32'h3c0f3da1),
	.w4(32'h3a604c53),
	.w5(32'h3c647e9b),
	.w6(32'h3b49f891),
	.w7(32'h3bd83e8d),
	.w8(32'h3beea8e9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df699b),
	.w1(32'hbc8e5717),
	.w2(32'h3c6b0c63),
	.w3(32'h3c290922),
	.w4(32'hbcb8664f),
	.w5(32'h3a7e77cb),
	.w6(32'hbca3847c),
	.w7(32'hbc59f82c),
	.w8(32'h3c942d38),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc802b4c),
	.w1(32'hbc8ebbd2),
	.w2(32'hbcc59e29),
	.w3(32'h3c7a5156),
	.w4(32'h3c3b629b),
	.w5(32'hbc19dfc9),
	.w6(32'h3c928e1b),
	.w7(32'h3c0f9f9e),
	.w8(32'h3a945df7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167a71),
	.w1(32'h3b9d85ce),
	.w2(32'hbc6fe27e),
	.w3(32'h3bdaf0c9),
	.w4(32'h3ca265d0),
	.w5(32'h3c087ff0),
	.w6(32'h3ba90921),
	.w7(32'h3c42ffb0),
	.w8(32'h3ae87d26),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9f604),
	.w1(32'hbb9d1675),
	.w2(32'hbc2c20b1),
	.w3(32'hbc154c15),
	.w4(32'hbb941c4d),
	.w5(32'hbc3d9292),
	.w6(32'hbb5bfe80),
	.w7(32'hbb3db7db),
	.w8(32'h3ae199d0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb21b95),
	.w1(32'hbbb4919b),
	.w2(32'h3b021251),
	.w3(32'h3b95d9e7),
	.w4(32'hb8f46145),
	.w5(32'hbc47582c),
	.w6(32'hbb155d2e),
	.w7(32'h3b52e0ce),
	.w8(32'h3a36abcc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93823a),
	.w1(32'h3ade79d1),
	.w2(32'h3969179a),
	.w3(32'h3bdf2c2c),
	.w4(32'h3b7b8130),
	.w5(32'hbbc7fb85),
	.w6(32'h3b777bd5),
	.w7(32'hb8bc31df),
	.w8(32'hb9dbf643),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ab6a),
	.w1(32'hbb237126),
	.w2(32'hbbac29fd),
	.w3(32'hbb800cb1),
	.w4(32'h3b22c949),
	.w5(32'h3b97dcc4),
	.w6(32'h3ab75313),
	.w7(32'h3abf7c5e),
	.w8(32'h3c4f4a0f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab11a5),
	.w1(32'h3c77b00a),
	.w2(32'hba83a895),
	.w3(32'h3a9a385f),
	.w4(32'h3b7e6aec),
	.w5(32'hbc474f89),
	.w6(32'h3a4bdf35),
	.w7(32'hbc1942a0),
	.w8(32'hbc903722),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61cc17),
	.w1(32'hbc68b02c),
	.w2(32'hbc4c9fdb),
	.w3(32'hbbd54bc7),
	.w4(32'hbbca38a3),
	.w5(32'h3bb078c0),
	.w6(32'hbbc4b450),
	.w7(32'hba3fb7ae),
	.w8(32'h3ba18c94),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff9bae),
	.w1(32'hbc4eb8a7),
	.w2(32'hbbb3b366),
	.w3(32'hba3ccc72),
	.w4(32'h3ae47790),
	.w5(32'h3ae28688),
	.w6(32'h3a4b9310),
	.w7(32'hbc32ad01),
	.w8(32'hbc666743),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe709e2),
	.w1(32'h3b293aee),
	.w2(32'hbbed557e),
	.w3(32'hbc87a01b),
	.w4(32'hbbb3264c),
	.w5(32'hbbe5b33a),
	.w6(32'hbc268f2e),
	.w7(32'hba0f5d40),
	.w8(32'hbba70b4b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7499d1),
	.w1(32'h3c544f15),
	.w2(32'h3c76d5c7),
	.w3(32'hbbeb7981),
	.w4(32'hb9b78ad5),
	.w5(32'h3cb02b12),
	.w6(32'h36f0b9b0),
	.w7(32'h3bfadc28),
	.w8(32'h3b9467d5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1754b8),
	.w1(32'h3b983a78),
	.w2(32'h39ec3bbe),
	.w3(32'hbb597ef3),
	.w4(32'hbbca03d0),
	.w5(32'hbc1f8430),
	.w6(32'hbbc564fd),
	.w7(32'hba971c79),
	.w8(32'h3c1566f2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7272d0d),
	.w1(32'h3ba57e07),
	.w2(32'hb9390ea9),
	.w3(32'h3bb9014b),
	.w4(32'h3badfcbe),
	.w5(32'hbbc00e72),
	.w6(32'h3bea6d8e),
	.w7(32'h3c18a1f6),
	.w8(32'h3c3ad3ae),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428705),
	.w1(32'h3a94333e),
	.w2(32'h3b2a4323),
	.w3(32'h3bb6e24e),
	.w4(32'h3b352754),
	.w5(32'h3c15acba),
	.w6(32'hbb5752ea),
	.w7(32'h3c025f0c),
	.w8(32'h3b2fa8cc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6774e0),
	.w1(32'hbae86f88),
	.w2(32'hbc17efce),
	.w3(32'hbb2592f6),
	.w4(32'hba81e771),
	.w5(32'hbbd23ac4),
	.w6(32'h3b972551),
	.w7(32'hba6cf57d),
	.w8(32'hbb1e18b0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ccbc2),
	.w1(32'hbb4e2d3d),
	.w2(32'hba5f2ed2),
	.w3(32'h391eedc3),
	.w4(32'h3ab1d9a8),
	.w5(32'h3bc27c15),
	.w6(32'hbb763db9),
	.w7(32'h393e67ec),
	.w8(32'h3a7ef516),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a313d),
	.w1(32'h3ca63ecb),
	.w2(32'h3c4bc64a),
	.w3(32'h3b2ae621),
	.w4(32'h3bc23267),
	.w5(32'hbbe836fb),
	.w6(32'hbbd0d71b),
	.w7(32'h3ad983e2),
	.w8(32'h3bacab52),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cde574),
	.w1(32'h3b3203ca),
	.w2(32'h39be6f24),
	.w3(32'h3c1115b6),
	.w4(32'hbab0f126),
	.w5(32'hbbc8a4ff),
	.w6(32'h3c30952b),
	.w7(32'hbb4bcbe1),
	.w8(32'h3afca31a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba167c0b),
	.w1(32'h3a909732),
	.w2(32'hb73d42b6),
	.w3(32'hbb1de3b6),
	.w4(32'h3be4f075),
	.w5(32'hba596911),
	.w6(32'h39d5fa75),
	.w7(32'h3a5b8358),
	.w8(32'h39e90e70),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d3ee),
	.w1(32'h3a6b28ac),
	.w2(32'h3a577be6),
	.w3(32'hbb990628),
	.w4(32'h3ad753f2),
	.w5(32'hbc0c752e),
	.w6(32'hbb765c7f),
	.w7(32'h3834d073),
	.w8(32'hbb8907b6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07cda3),
	.w1(32'hb9b36cd4),
	.w2(32'hbab196ac),
	.w3(32'hbbbd9194),
	.w4(32'h3c40d397),
	.w5(32'h3a1b8882),
	.w6(32'h39dac558),
	.w7(32'h3bd25f9c),
	.w8(32'h39714af0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f097a1),
	.w1(32'h3b39d2b8),
	.w2(32'hbbd8efe3),
	.w3(32'h3c3e8a77),
	.w4(32'h3b0d2aec),
	.w5(32'hbc1d4126),
	.w6(32'h3c0fc0c1),
	.w7(32'hbb9b531c),
	.w8(32'hbbfd3323),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90329b),
	.w1(32'h3b661b20),
	.w2(32'h3bc392ef),
	.w3(32'hbbc34041),
	.w4(32'hbbbc69d7),
	.w5(32'h3acd83a1),
	.w6(32'h3acac87b),
	.w7(32'hb946481f),
	.w8(32'h3c5c3f78),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b507f69),
	.w1(32'h3a7aaa20),
	.w2(32'hbb0fc15e),
	.w3(32'hbb35830c),
	.w4(32'h399413a5),
	.w5(32'hba08c736),
	.w6(32'h3bbb3eec),
	.w7(32'h3aedd6a6),
	.w8(32'hbb17f6ea),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f9d7c),
	.w1(32'h39fcb7a8),
	.w2(32'hbb51f7f7),
	.w3(32'hbbf5665f),
	.w4(32'h3bebbe94),
	.w5(32'hbc17cb85),
	.w6(32'h3bfab343),
	.w7(32'h3bcca3cb),
	.w8(32'hbb17bcf9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b729d57),
	.w1(32'hbb800bf6),
	.w2(32'hbb820fbf),
	.w3(32'h3b438396),
	.w4(32'h3b8e2322),
	.w5(32'h3c8a59c5),
	.w6(32'h3b7f73de),
	.w7(32'h3a29fecf),
	.w8(32'h3b090503),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ff6c),
	.w1(32'h3b4d07f1),
	.w2(32'h3b5f03b0),
	.w3(32'h3c2c1f1d),
	.w4(32'h3ba2c9ae),
	.w5(32'hbbcabd7b),
	.w6(32'hbbc2a173),
	.w7(32'h3b2e5339),
	.w8(32'h3b6ceb30),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97c566),
	.w1(32'h3b9fa799),
	.w2(32'h3acf785d),
	.w3(32'hbb3d9ab6),
	.w4(32'hb95ecb89),
	.w5(32'hbc2324b7),
	.w6(32'h3b66b950),
	.w7(32'hbb7cbf8b),
	.w8(32'hba50c6c6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf650d),
	.w1(32'h37051d7f),
	.w2(32'hba105b36),
	.w3(32'h3b25b1b5),
	.w4(32'h3abea7a2),
	.w5(32'h3c0d1e7c),
	.w6(32'hbb4a34d5),
	.w7(32'h3b0ff3b5),
	.w8(32'h3c2518ee),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda8f01),
	.w1(32'h3cbd85f1),
	.w2(32'h3c8f2a74),
	.w3(32'hbb5380bb),
	.w4(32'hba877bd3),
	.w5(32'hbbd09a5b),
	.w6(32'h3b9a3b4a),
	.w7(32'hb9dda815),
	.w8(32'hbbe86350),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc678acb),
	.w1(32'hbb846fc2),
	.w2(32'h38fad9c4),
	.w3(32'h3b880ded),
	.w4(32'hba8cbe0d),
	.w5(32'hba2409c5),
	.w6(32'h3c4880c9),
	.w7(32'h3bc57c66),
	.w8(32'hbc10bc9a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16319d),
	.w1(32'hba1563b8),
	.w2(32'hbc13b56d),
	.w3(32'h3b63238a),
	.w4(32'hbb417193),
	.w5(32'h3bf2c168),
	.w6(32'h3bd71739),
	.w7(32'h3a75e239),
	.w8(32'hbc7b020f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93cd97),
	.w1(32'hbccfa65d),
	.w2(32'hbcc91ede),
	.w3(32'hbc050f54),
	.w4(32'h3bba07c6),
	.w5(32'hbb296421),
	.w6(32'hbb712f1c),
	.w7(32'h3ba2fb23),
	.w8(32'hbb35b523),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f40c1),
	.w1(32'hba42d0b5),
	.w2(32'hba01d962),
	.w3(32'h3a8d66a6),
	.w4(32'hb8d7ff48),
	.w5(32'hba0f5e98),
	.w6(32'hba373bba),
	.w7(32'hb93f2c21),
	.w8(32'h39136edf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39388eef),
	.w1(32'h35c83f10),
	.w2(32'hba0a7617),
	.w3(32'hb924e7ac),
	.w4(32'hba05ebfb),
	.w5(32'hba5bef7d),
	.w6(32'h3974700d),
	.w7(32'hb9dd5f67),
	.w8(32'hbaa7d3ec),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933aa74),
	.w1(32'hba3f82dc),
	.w2(32'hbab5869f),
	.w3(32'hb9ceca7f),
	.w4(32'hba9f4678),
	.w5(32'hbaf22a27),
	.w6(32'hb903350b),
	.w7(32'hba1f2caa),
	.w8(32'hbb0b969b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d0aa7),
	.w1(32'h3b78d577),
	.w2(32'h3b12fd6e),
	.w3(32'hbb2c2d18),
	.w4(32'h3b11120c),
	.w5(32'h3a866596),
	.w6(32'hb9b09d92),
	.w7(32'h3a59091f),
	.w8(32'hba8b4f10),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952d1e3),
	.w1(32'hba43e307),
	.w2(32'hba304471),
	.w3(32'h39d9fa50),
	.w4(32'hbaf2f440),
	.w5(32'hb9b7cd1f),
	.w6(32'h39f84438),
	.w7(32'hba3de807),
	.w8(32'hb9a3a0b8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac383f9),
	.w1(32'h3c1c4bf6),
	.w2(32'h3c3da0ba),
	.w3(32'h3aa4431c),
	.w4(32'hbab439bf),
	.w5(32'h3bb3e797),
	.w6(32'hbace0ab3),
	.w7(32'h3b3bb89e),
	.w8(32'h3b83b3cf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc079d82),
	.w1(32'h3bcd2c76),
	.w2(32'h3c353cd1),
	.w3(32'hbb1a2f5d),
	.w4(32'hb9974a34),
	.w5(32'h3bf1c5b8),
	.w6(32'hbae0e441),
	.w7(32'hba8ee8c0),
	.w8(32'h3909fea2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04074b),
	.w1(32'hbbff34c0),
	.w2(32'hbbc6254d),
	.w3(32'h391cf3b7),
	.w4(32'hbaeaf0b9),
	.w5(32'hbb342823),
	.w6(32'hbafec546),
	.w7(32'hbb06f1e2),
	.w8(32'hbb0cf2e0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a269400),
	.w1(32'h3b051ff4),
	.w2(32'hbb38d286),
	.w3(32'hbb506604),
	.w4(32'hb9965b0f),
	.w5(32'hbb8a3ef7),
	.w6(32'hb9bc9be6),
	.w7(32'hbaec04be),
	.w8(32'hbb981910),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba424409),
	.w1(32'h3c05db34),
	.w2(32'h3c0d1d15),
	.w3(32'hbb9e0aa0),
	.w4(32'hba5ba64b),
	.w5(32'h3b260d75),
	.w6(32'hbad45081),
	.w7(32'hba494896),
	.w8(32'hb7de9bc4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a0468),
	.w1(32'h3b92e635),
	.w2(32'h39af7c7d),
	.w3(32'hb99b9310),
	.w4(32'h3b58dbef),
	.w5(32'h3b0254c5),
	.w6(32'hba68522f),
	.w7(32'h3ad15de8),
	.w8(32'h3a64fcde),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69a5a1),
	.w1(32'h3bd0a563),
	.w2(32'h3bb1d140),
	.w3(32'h3764558e),
	.w4(32'h3b0629cb),
	.w5(32'h3b0b4db6),
	.w6(32'hbaa32e73),
	.w7(32'h3addf21b),
	.w8(32'h3ad44986),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914fb8d),
	.w1(32'h36e61977),
	.w2(32'h3a10fcc5),
	.w3(32'hb919d964),
	.w4(32'h39f7e56b),
	.w5(32'hb8691bf8),
	.w6(32'hb92e5c9c),
	.w7(32'h35855ff1),
	.w8(32'hb86e3c86),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e72bc),
	.w1(32'hbaa68b13),
	.w2(32'hba738eaf),
	.w3(32'h381cdc98),
	.w4(32'hbad50475),
	.w5(32'hbaa980a8),
	.w6(32'h397524b9),
	.w7(32'hbaf18c93),
	.w8(32'hb9f80ece),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9825f2e),
	.w1(32'h398aee96),
	.w2(32'hba3cf7ad),
	.w3(32'h395a7e16),
	.w4(32'h380ab9c4),
	.w5(32'hbacaf07c),
	.w6(32'hb9da81c6),
	.w7(32'h3927ab4a),
	.w8(32'hb983f527),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8430ba2),
	.w1(32'hba4f3cb9),
	.w2(32'hbaecd023),
	.w3(32'h3b060a9e),
	.w4(32'h3abc27bd),
	.w5(32'h3934d746),
	.w6(32'h3a3cdf3d),
	.w7(32'h3ad86a9b),
	.w8(32'h3941367f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf703a0),
	.w1(32'hbc1f301d),
	.w2(32'hbbc76bb2),
	.w3(32'h3b2f9065),
	.w4(32'h3a0be9d1),
	.w5(32'hba37af20),
	.w6(32'h3b2925b4),
	.w7(32'hb9f746a3),
	.w8(32'h3a98d8a3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9889858),
	.w1(32'hb8c2b1c0),
	.w2(32'h3a1888c2),
	.w3(32'h39c0b390),
	.w4(32'h392a8edc),
	.w5(32'h3ada3e45),
	.w6(32'hb9912f5e),
	.w7(32'h3975b269),
	.w8(32'hb92d2949),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e972a),
	.w1(32'hbc603363),
	.w2(32'hbc10fdf1),
	.w3(32'hb9ccd133),
	.w4(32'hbc060ae4),
	.w5(32'hbb136126),
	.w6(32'hbb1466ca),
	.w7(32'hbba86139),
	.w8(32'hbb861ebb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf81b0),
	.w1(32'h3be4d473),
	.w2(32'h3bf1272c),
	.w3(32'hbbcd085e),
	.w4(32'h3aeeca54),
	.w5(32'h3b3056d2),
	.w6(32'hbbbd1e23),
	.w7(32'h3adf9f56),
	.w8(32'hb9cdde2f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b695246),
	.w1(32'h39aba5e9),
	.w2(32'hbb29bb1a),
	.w3(32'h3beaf325),
	.w4(32'h3bcc81fd),
	.w5(32'h3b013cae),
	.w6(32'hba319db4),
	.w7(32'h3af49f62),
	.w8(32'h3a982864),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ea3d6),
	.w1(32'h3c19fd07),
	.w2(32'h3c3780b2),
	.w3(32'hbc0e2a6e),
	.w4(32'hbc064cf8),
	.w5(32'h3a92a12a),
	.w6(32'hbc07861e),
	.w7(32'h3c18a13c),
	.w8(32'h3ad8e720),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03c80e),
	.w1(32'h3af9c1c5),
	.w2(32'hbb1c72ce),
	.w3(32'h3bbc1e7e),
	.w4(32'h3c0040df),
	.w5(32'h3b95c7ca),
	.w6(32'h3ba0a479),
	.w7(32'h3be23313),
	.w8(32'h3b471224),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61e0bb),
	.w1(32'h3bc13e54),
	.w2(32'h3a537470),
	.w3(32'hbc53599c),
	.w4(32'h3a86387d),
	.w5(32'hbbbd9371),
	.w6(32'hbb88c0c6),
	.w7(32'hba89541c),
	.w8(32'hbc151506),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b8666),
	.w1(32'h3ade56c9),
	.w2(32'h39aef0bf),
	.w3(32'hbacff96a),
	.w4(32'hbb23d532),
	.w5(32'hbb0ea849),
	.w6(32'h39ba7645),
	.w7(32'hb952e678),
	.w8(32'hbbb5a5f3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b27c5),
	.w1(32'hbbc6a352),
	.w2(32'hbc141911),
	.w3(32'h3b4b0683),
	.w4(32'h3bd1c39d),
	.w5(32'h3a1d76de),
	.w6(32'hb9300585),
	.w7(32'h3b2c5bd4),
	.w8(32'hbac216e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6bd99),
	.w1(32'h39cc46fa),
	.w2(32'hb97f8170),
	.w3(32'h3a747b05),
	.w4(32'h3a8bf15f),
	.w5(32'hba1779fd),
	.w6(32'h3aaadc77),
	.w7(32'h3aac326f),
	.w8(32'hb94e5b41),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e6a53),
	.w1(32'h3bafa3cc),
	.w2(32'h3b6d9c1e),
	.w3(32'hbb8b609d),
	.w4(32'h3b882984),
	.w5(32'h3b430c9d),
	.w6(32'hbb32c40e),
	.w7(32'h3b17f2a4),
	.w8(32'h3a265c89),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1809f7),
	.w1(32'h3c46f8e8),
	.w2(32'h3c806f65),
	.w3(32'hbb75d973),
	.w4(32'hbb13197e),
	.w5(32'h3bc00c81),
	.w6(32'hbbdea0d2),
	.w7(32'h3a0492b0),
	.w8(32'hbab69bd7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4262e0),
	.w1(32'hbcaa301e),
	.w2(32'h3bbfd916),
	.w3(32'h3b859b28),
	.w4(32'hbcbf6ec9),
	.w5(32'hba906e52),
	.w6(32'hbaf1edaf),
	.w7(32'hbbee2c77),
	.w8(32'h3b0d94d3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82070c),
	.w1(32'hbca0708d),
	.w2(32'hbc8b9ee1),
	.w3(32'h3b96c25b),
	.w4(32'hb9c8f365),
	.w5(32'hbbf358a1),
	.w6(32'hb89ed20f),
	.w7(32'h3bc7a215),
	.w8(32'hba0f64b4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb5966),
	.w1(32'hbc508ef9),
	.w2(32'hbc1b2d7d),
	.w3(32'h3a230e9e),
	.w4(32'h3a800f5f),
	.w5(32'hbae2a77e),
	.w6(32'hb92a528c),
	.w7(32'h3ac3e624),
	.w8(32'h39f7926f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2d2bf),
	.w1(32'h3be93614),
	.w2(32'h3c216ff0),
	.w3(32'hbaf77863),
	.w4(32'hbc5bde49),
	.w5(32'h391201e6),
	.w6(32'hbc095f02),
	.w7(32'hbaf3e6e3),
	.w8(32'h3bdfb6bf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ea222),
	.w1(32'hb9417a76),
	.w2(32'h3a47d5b1),
	.w3(32'hbac88bb3),
	.w4(32'h397d18ea),
	.w5(32'h3a5652ed),
	.w6(32'h3ad959b5),
	.w7(32'h3b29d930),
	.w8(32'h3b6e8ce0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c271411),
	.w1(32'hbc3f8298),
	.w2(32'h3bf75a0b),
	.w3(32'h3c6497ec),
	.w4(32'hbcc768fb),
	.w5(32'hba9372a4),
	.w6(32'hbc286f1c),
	.w7(32'hbc95a6c8),
	.w8(32'hba17a996),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdf6e6),
	.w1(32'h3b9a4c40),
	.w2(32'h3bfa2068),
	.w3(32'h3b2e918f),
	.w4(32'hba0b54f5),
	.w5(32'h3bcf64fa),
	.w6(32'hbaf47e5b),
	.w7(32'h3a950aff),
	.w8(32'h3c0aa97e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39163e06),
	.w1(32'hba256bd3),
	.w2(32'hb94fcc2d),
	.w3(32'h39cd02da),
	.w4(32'h396d2494),
	.w5(32'hb9bdbfa4),
	.w6(32'h39c05e3c),
	.w7(32'h394ff80d),
	.w8(32'hb7c5c93c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc649),
	.w1(32'hb9c4cbf4),
	.w2(32'hba7a6393),
	.w3(32'h3b13ad4c),
	.w4(32'h3ac90d7d),
	.w5(32'hbad9db6f),
	.w6(32'h3b83669c),
	.w7(32'h3b1a2dd8),
	.w8(32'h39b57301),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8ab91),
	.w1(32'h3c01d977),
	.w2(32'h3bd3ba1d),
	.w3(32'hbb34684b),
	.w4(32'h3b60cb0e),
	.w5(32'h3b985273),
	.w6(32'hbb3c4c1a),
	.w7(32'h3b735912),
	.w8(32'h3b4a1b32),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a2ec),
	.w1(32'hbbad9c9a),
	.w2(32'hbbb19681),
	.w3(32'h3af18a58),
	.w4(32'h3b52104e),
	.w5(32'h3a81c0a3),
	.w6(32'hba5986ec),
	.w7(32'h3b041b80),
	.w8(32'h3968f17e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b916),
	.w1(32'h3ba69528),
	.w2(32'hbaa5c9f7),
	.w3(32'h3ac54c44),
	.w4(32'h3c2154e0),
	.w5(32'h3b6fa336),
	.w6(32'hbb8aa504),
	.w7(32'h3bda9c7b),
	.w8(32'h3b9ceb54),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08c94a),
	.w1(32'hbc125843),
	.w2(32'hbc1b568c),
	.w3(32'hbb8ef792),
	.w4(32'hbb71d588),
	.w5(32'hbba8bacb),
	.w6(32'hbb83677b),
	.w7(32'hbb3ef373),
	.w8(32'hbacd77d1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09d0ae),
	.w1(32'hbc2d4ac8),
	.w2(32'hbb996256),
	.w3(32'h3bd1d12a),
	.w4(32'hbc160a71),
	.w5(32'hba9bb400),
	.w6(32'h3b61932c),
	.w7(32'hb98bf07a),
	.w8(32'hbb823452),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f2c66),
	.w1(32'h3c174b6d),
	.w2(32'h3b094455),
	.w3(32'hb9af95b8),
	.w4(32'h3ab0ce31),
	.w5(32'hbbc53ac9),
	.w6(32'hba7ee46e),
	.w7(32'hba4e986d),
	.w8(32'hbc0ae6a2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749eed),
	.w1(32'hbb34ec3a),
	.w2(32'hbb3c59f9),
	.w3(32'hbb6205a7),
	.w4(32'h3902e63d),
	.w5(32'hba9f31b6),
	.w6(32'hbb432530),
	.w7(32'hba68f8d0),
	.w8(32'hbaca8677),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39155691),
	.w1(32'hba521260),
	.w2(32'hbaa6afd4),
	.w3(32'hb9b50ee1),
	.w4(32'hba243e53),
	.w5(32'hba418eae),
	.w6(32'h38841398),
	.w7(32'hba1ac05d),
	.w8(32'hba4fe406),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8a97b),
	.w1(32'hb9bf5304),
	.w2(32'hb9802d3e),
	.w3(32'hba9fcc90),
	.w4(32'hbaa3aae4),
	.w5(32'hbaed64f0),
	.w6(32'h3a89362b),
	.w7(32'h3a4d2cf8),
	.w8(32'hba350a81),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c99ab0),
	.w1(32'h3aafe33d),
	.w2(32'h39e77f12),
	.w3(32'hb944f09c),
	.w4(32'h3a45adf5),
	.w5(32'h3a4e8fcc),
	.w6(32'h3803bb0f),
	.w7(32'hba2e461e),
	.w8(32'h394d8d96),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57a1c3),
	.w1(32'h3b02e2db),
	.w2(32'h3af8a4c1),
	.w3(32'h3aa3481a),
	.w4(32'h3b04bd92),
	.w5(32'h3b2c888d),
	.w6(32'h39fb37f3),
	.w7(32'h3b1f64bc),
	.w8(32'h3b1434ed),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a531),
	.w1(32'hbbb37ea0),
	.w2(32'hbba745ce),
	.w3(32'hb983774e),
	.w4(32'h39a8a8e7),
	.w5(32'hba38b6a7),
	.w6(32'hb9cc47e0),
	.w7(32'hb97b6016),
	.w8(32'hb9936e97),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac4b0f),
	.w1(32'hb9c9af38),
	.w2(32'hbaf3439e),
	.w3(32'hb9dde9df),
	.w4(32'hba0d93c3),
	.w5(32'hba66dd15),
	.w6(32'hb9b8134c),
	.w7(32'h3a503dec),
	.w8(32'hba44a763),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d8809),
	.w1(32'h3bc09923),
	.w2(32'h3bfd609b),
	.w3(32'hbab52fd7),
	.w4(32'hbaeaf96e),
	.w5(32'h3b3bf6ad),
	.w6(32'hbb06fa4f),
	.w7(32'h3adb7f3b),
	.w8(32'h3ab765bb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18eb78),
	.w1(32'hbc7fe7ad),
	.w2(32'hbc94fc3a),
	.w3(32'hbaa4d4a5),
	.w4(32'h3a032efa),
	.w5(32'hbc02a7ae),
	.w6(32'h3b0dd098),
	.w7(32'h3a9d0321),
	.w8(32'hbba1706a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2a0c3),
	.w1(32'hba6e6f2d),
	.w2(32'hb99ed7f1),
	.w3(32'h394490bd),
	.w4(32'hba6b3304),
	.w5(32'hba40795f),
	.w6(32'h39fd8728),
	.w7(32'hba5cc0f6),
	.w8(32'hb9b02b4f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bfddc),
	.w1(32'h392fe2ef),
	.w2(32'hb96c7b6d),
	.w3(32'h3933e2b0),
	.w4(32'hba442e46),
	.w5(32'h39e314f3),
	.w6(32'hb993d0cc),
	.w7(32'hb9c1a2af),
	.w8(32'h3776ae4c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25eb9f),
	.w1(32'hba57b7f0),
	.w2(32'hba07b2b9),
	.w3(32'h38ad7b24),
	.w4(32'hba87b735),
	.w5(32'hba51eb5d),
	.w6(32'hb9bf667c),
	.w7(32'hb9adff99),
	.w8(32'hb927a707),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab11a4),
	.w1(32'h39215d60),
	.w2(32'h390590b2),
	.w3(32'hbaa245e4),
	.w4(32'h3adb1294),
	.w5(32'h3b394563),
	.w6(32'hba8ab7f3),
	.w7(32'h3a5b8a37),
	.w8(32'h3b08e7c0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc947197),
	.w1(32'hbb87c984),
	.w2(32'h3c1cddf5),
	.w3(32'h3bbb6e99),
	.w4(32'h3b6938f7),
	.w5(32'h3c35345a),
	.w6(32'h3c0a5cbd),
	.w7(32'h3c48755b),
	.w8(32'h3bc42628),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2cce3),
	.w1(32'h3c492158),
	.w2(32'h3bd0032f),
	.w3(32'hbb821b20),
	.w4(32'h3ba47fea),
	.w5(32'h3b220a03),
	.w6(32'hbafde9d1),
	.w7(32'h3b5348c7),
	.w8(32'hb9fce992),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f52b5),
	.w1(32'h3af9a196),
	.w2(32'h3b1008a0),
	.w3(32'h38f7a059),
	.w4(32'hba1f4b6e),
	.w5(32'h3a984803),
	.w6(32'hba19a833),
	.w7(32'hba5c9a63),
	.w8(32'h3a8002ce),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f32d1),
	.w1(32'hbac77882),
	.w2(32'hbb0a3bd2),
	.w3(32'h3b64df04),
	.w4(32'h3a1a553f),
	.w5(32'hb8a8231f),
	.w6(32'h3b2ae583),
	.w7(32'h3b34d1db),
	.w8(32'hba9114b1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e18fdb),
	.w1(32'h38aef1d9),
	.w2(32'h39281554),
	.w3(32'h3a691e96),
	.w4(32'h3aaddd81),
	.w5(32'hba827998),
	.w6(32'hba607e9c),
	.w7(32'h38f985c0),
	.w8(32'h38aa5bc8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a363bca),
	.w1(32'h3a8d1a1c),
	.w2(32'hb979b39b),
	.w3(32'hbb72598a),
	.w4(32'hb9654ab1),
	.w5(32'hbaf9e87f),
	.w6(32'hbaf5d7a7),
	.w7(32'hba37d5ab),
	.w8(32'hbb3fed44),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0e0ed),
	.w1(32'h3a72fd2a),
	.w2(32'hbab75ef2),
	.w3(32'h3ac51b4a),
	.w4(32'h3b0a40ba),
	.w5(32'hbb17dfe7),
	.w6(32'h3a95edef),
	.w7(32'hbacc713d),
	.w8(32'hbb83ac73),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c317b50),
	.w1(32'h3c9301eb),
	.w2(32'h3c82e83f),
	.w3(32'hbb30e491),
	.w4(32'h3b15dc71),
	.w5(32'h3bf03c6b),
	.w6(32'hbaee10df),
	.w7(32'h3b880cde),
	.w8(32'h3b4bbd34),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09258),
	.w1(32'hbbbe6b28),
	.w2(32'hbb9bb09d),
	.w3(32'hb8c59982),
	.w4(32'h3ad1ce30),
	.w5(32'h3a1283d5),
	.w6(32'hba882dca),
	.w7(32'hb9057593),
	.w8(32'hb8be0ddc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71ed0f),
	.w1(32'h3ac0be7c),
	.w2(32'h3b77dcb0),
	.w3(32'hb9872b1b),
	.w4(32'hbb0651fd),
	.w5(32'hb977224e),
	.w6(32'hbadcd6ce),
	.w7(32'hba9fdbb3),
	.w8(32'hbacc433c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52830),
	.w1(32'h3c064f6a),
	.w2(32'h3c173932),
	.w3(32'hbb40f259),
	.w4(32'h3a486486),
	.w5(32'h3bec8a64),
	.w6(32'hbbf5bdf3),
	.w7(32'hb6778978),
	.w8(32'h398af0cd),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc36b),
	.w1(32'hbc2b0d82),
	.w2(32'hbb921da0),
	.w3(32'hbab9cb55),
	.w4(32'hbbb3c931),
	.w5(32'h38e1a8af),
	.w6(32'hb98d2678),
	.w7(32'hbb5fcbdb),
	.w8(32'hbb2a8829),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f27d2),
	.w1(32'h3b93d529),
	.w2(32'h3bc2a11b),
	.w3(32'hbb4d29be),
	.w4(32'hba8507ef),
	.w5(32'h3acabd20),
	.w6(32'hbb624ad5),
	.w7(32'h3a91589a),
	.w8(32'h3b043051),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3656),
	.w1(32'hbad07a99),
	.w2(32'h39ca0e53),
	.w3(32'h39b62e36),
	.w4(32'hba1a68cd),
	.w5(32'hb99df00b),
	.w6(32'h389e47f4),
	.w7(32'h390eafaa),
	.w8(32'h3aea9181),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e6ce),
	.w1(32'hbae1882e),
	.w2(32'hbc8b71ca),
	.w3(32'h3b440cf8),
	.w4(32'h3b93ecff),
	.w5(32'hbb4fd374),
	.w6(32'h39d309a9),
	.w7(32'h3b730582),
	.w8(32'hbb4e6962),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae80952),
	.w1(32'hba8dfe3b),
	.w2(32'hbb03c46d),
	.w3(32'hba5eaf89),
	.w4(32'h3b1449c0),
	.w5(32'hba874bae),
	.w6(32'h3a2b8f69),
	.w7(32'h3b09fc04),
	.w8(32'hbaaf6d03),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e914f),
	.w1(32'hb90c73f3),
	.w2(32'hb941b686),
	.w3(32'hba2ec269),
	.w4(32'h3959fcde),
	.w5(32'h39b652e0),
	.w6(32'hba1755ca),
	.w7(32'h370b6261),
	.w8(32'h3882291b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388026e6),
	.w1(32'hb92f8c75),
	.w2(32'hba630580),
	.w3(32'h3999093e),
	.w4(32'hba486326),
	.w5(32'hba0b430b),
	.w6(32'h3a7bbcf6),
	.w7(32'hb9706372),
	.w8(32'hb8712a62),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4dbff),
	.w1(32'h3aeaa2e7),
	.w2(32'h3b1685f9),
	.w3(32'hbb008adb),
	.w4(32'hbaaad712),
	.w5(32'h39082f9c),
	.w6(32'hbadaa91f),
	.w7(32'hbaf4a8da),
	.w8(32'hba9d18cb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd31e6d),
	.w1(32'hbbe6988d),
	.w2(32'hbb02214f),
	.w3(32'h3ad55186),
	.w4(32'h3926d51a),
	.w5(32'h3b13af2b),
	.w6(32'h3ac1b5f3),
	.w7(32'h39ed01ef),
	.w8(32'h3b8652cb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5cd29),
	.w1(32'h3a3ad89b),
	.w2(32'hb84507f9),
	.w3(32'hbafccfa2),
	.w4(32'hbb0eaff5),
	.w5(32'hba2f1f10),
	.w6(32'hba60ef43),
	.w7(32'hbaef3cba),
	.w8(32'hbade7061),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39140607),
	.w1(32'hb8d6fa12),
	.w2(32'h39604305),
	.w3(32'hb7c35585),
	.w4(32'h3936ff88),
	.w5(32'h390c96c5),
	.w6(32'hba7137fb),
	.w7(32'h39456200),
	.w8(32'h3a4571ff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a1a5),
	.w1(32'h3bf63e19),
	.w2(32'h3b9f4d80),
	.w3(32'hbab32ca5),
	.w4(32'h3af3eb09),
	.w5(32'h3afadf73),
	.w6(32'h3977a9a9),
	.w7(32'h3aeca17e),
	.w8(32'h3b00a558),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89fa67e),
	.w1(32'h393dc067),
	.w2(32'hb94df564),
	.w3(32'h3ab3b093),
	.w4(32'hba16b528),
	.w5(32'hbabab1f6),
	.w6(32'h38b9df78),
	.w7(32'h39d341ac),
	.w8(32'hbaf416f4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b049ea0),
	.w1(32'h3c3b2865),
	.w2(32'h3c6c2d6b),
	.w3(32'hbc35a220),
	.w4(32'hbbb570b3),
	.w5(32'h39873bae),
	.w6(32'hbc0b9445),
	.w7(32'h3a81ca8f),
	.w8(32'h3b0e6b86),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07cbae),
	.w1(32'h3b65edc3),
	.w2(32'hbb8adb3b),
	.w3(32'hbb0e1b15),
	.w4(32'h3c6fd9ae),
	.w5(32'h3c4924ce),
	.w6(32'h3b98eefb),
	.w7(32'h3c1595b2),
	.w8(32'h3b995637),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ee337),
	.w1(32'hbb97e1ed),
	.w2(32'hbb337f5d),
	.w3(32'h3af73943),
	.w4(32'h3a4079b7),
	.w5(32'h39b01b48),
	.w6(32'h3b7b7931),
	.w7(32'h3aa47ccd),
	.w8(32'hb9791a5e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a3690),
	.w1(32'hba966a7b),
	.w2(32'h3a076c37),
	.w3(32'h3965fdd6),
	.w4(32'hb89f8da7),
	.w5(32'h3a2031ca),
	.w6(32'hb97dff68),
	.w7(32'h3ad18a87),
	.w8(32'h3b2a71f3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55dca),
	.w1(32'hbbbec58a),
	.w2(32'hbbb8ad7b),
	.w3(32'hbad54e5e),
	.w4(32'hba942477),
	.w5(32'hbaa746f4),
	.w6(32'hbab5a750),
	.w7(32'hbaa5d16a),
	.w8(32'hbac6cc62),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae67c5e),
	.w1(32'hbb92fd05),
	.w2(32'hbb4c16f6),
	.w3(32'hb8c09942),
	.w4(32'hbb18b602),
	.w5(32'hbaf379e2),
	.w6(32'hbb38e21d),
	.w7(32'hbbb9e7a4),
	.w8(32'hbb60c3b1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7badbe),
	.w1(32'hbb8e1a60),
	.w2(32'hbb8e4a1f),
	.w3(32'h39d91aed),
	.w4(32'h3a9307b9),
	.w5(32'hba0c8925),
	.w6(32'h38dca3fa),
	.w7(32'h3a44d1d0),
	.w8(32'hb966bc28),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06de4e),
	.w1(32'h3b477502),
	.w2(32'h3b59ef50),
	.w3(32'h3a259e66),
	.w4(32'hba819559),
	.w5(32'h3aa341c6),
	.w6(32'h365c9c78),
	.w7(32'hb8f9c430),
	.w8(32'h3aff0c56),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64229),
	.w1(32'hba875703),
	.w2(32'hbaa5474c),
	.w3(32'h3a0c389d),
	.w4(32'h37247bc7),
	.w5(32'hba2689ff),
	.w6(32'h39fc8111),
	.w7(32'h39e85801),
	.w8(32'hb98c9e0d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a3fbb),
	.w1(32'h3b35954b),
	.w2(32'h3b2c07f2),
	.w3(32'hbbaacdd2),
	.w4(32'h3a5caacf),
	.w5(32'h3a257a45),
	.w6(32'hbbb53032),
	.w7(32'hbab9fd7a),
	.w8(32'h3b1bf126),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ad089),
	.w1(32'h3b6ccf02),
	.w2(32'h3b8175d0),
	.w3(32'hba88854f),
	.w4(32'h3aaf3487),
	.w5(32'h3ac5edd5),
	.w6(32'hbb42627a),
	.w7(32'h3abaa0fc),
	.w8(32'hba3d1f8a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9aff02),
	.w1(32'hbb5ef875),
	.w2(32'hbbb87942),
	.w3(32'h3b034f95),
	.w4(32'h3b806da3),
	.w5(32'hb761bccd),
	.w6(32'h3aa6937e),
	.w7(32'h3a1603e8),
	.w8(32'hba2f0ab9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e3387),
	.w1(32'hb9f3d382),
	.w2(32'hbaada2c9),
	.w3(32'h3b04d50e),
	.w4(32'h39ae19d1),
	.w5(32'hba9b9ab8),
	.w6(32'h3a93535a),
	.w7(32'hb964f4b6),
	.w8(32'hba8ad82c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7b9cf),
	.w1(32'hba5ce0fc),
	.w2(32'h3b431ecf),
	.w3(32'h3b98d6dd),
	.w4(32'h3bbc374e),
	.w5(32'h3b94b698),
	.w6(32'h3bebf54d),
	.w7(32'h3bee5888),
	.w8(32'h3b00b41f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e909f5),
	.w1(32'h38d648ff),
	.w2(32'h3a48c9d6),
	.w3(32'hb9a32993),
	.w4(32'hb736c2ac),
	.w5(32'hb98aa87c),
	.w6(32'hb9b3f170),
	.w7(32'h39ecba89),
	.w8(32'h3a87b503),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe9133),
	.w1(32'h3a5cdbf9),
	.w2(32'h3a30359a),
	.w3(32'h3ab5fc6a),
	.w4(32'h3a0b4345),
	.w5(32'h3a3c96c5),
	.w6(32'h3abf3c03),
	.w7(32'h3a09e183),
	.w8(32'h39d93bf6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3da2c0),
	.w1(32'hbb952b45),
	.w2(32'hbbbb7f2c),
	.w3(32'hba8a42b5),
	.w4(32'h3acd1a5d),
	.w5(32'hba2eba5d),
	.w6(32'hbb2f5ef6),
	.w7(32'h3ab445a8),
	.w8(32'h3af6d6be),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a26df),
	.w1(32'h391581ad),
	.w2(32'h3c3123ce),
	.w3(32'hbbe69552),
	.w4(32'h3a8cc069),
	.w5(32'h3c22d56e),
	.w6(32'hbc42c734),
	.w7(32'h3b3d4718),
	.w8(32'h3b92044e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7432ec6),
	.w1(32'h39badd23),
	.w2(32'h3a2585ee),
	.w3(32'h382cf785),
	.w4(32'h3a27e107),
	.w5(32'hba06d862),
	.w6(32'h39b7dab8),
	.w7(32'h3a7a51a9),
	.w8(32'h39210a64),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826220),
	.w1(32'hbc018adb),
	.w2(32'hbc01b96f),
	.w3(32'hba5cbea3),
	.w4(32'hba3fdb03),
	.w5(32'hbb7d3e9f),
	.w6(32'hb97801b6),
	.w7(32'hba3c77ff),
	.w8(32'hbb2fcd55),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b4acd),
	.w1(32'h3bcf7115),
	.w2(32'h3bdfd7a8),
	.w3(32'hbac32e84),
	.w4(32'h3bd7c114),
	.w5(32'h3bf27944),
	.w6(32'hba2fe6c4),
	.w7(32'h3a232aeb),
	.w8(32'h39e32dc3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5068b),
	.w1(32'h3c792c7c),
	.w2(32'h3ad7a906),
	.w3(32'hb8f23e15),
	.w4(32'h3c05aa6f),
	.w5(32'h3af479bb),
	.w6(32'h3b2623bc),
	.w7(32'h3b942fb3),
	.w8(32'hbb989abc),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28d22a),
	.w1(32'h3c0649eb),
	.w2(32'h3b6267d8),
	.w3(32'hbb30668d),
	.w4(32'hb9a3b7ea),
	.w5(32'hb9eb4cbc),
	.w6(32'hbb757f52),
	.w7(32'hbb29fb38),
	.w8(32'hbb1b6c78),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fddc0),
	.w1(32'h3be65673),
	.w2(32'h3baacfb8),
	.w3(32'hbb89374e),
	.w4(32'h3b226a26),
	.w5(32'h3b73c788),
	.w6(32'hbb9cd8f5),
	.w7(32'h3b2ea49e),
	.w8(32'h3b0a4b21),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982155),
	.w1(32'hb975fa43),
	.w2(32'hbaaaf749),
	.w3(32'h39eecc31),
	.w4(32'hb960121b),
	.w5(32'h38b52f8d),
	.w6(32'hba017ad1),
	.w7(32'h381793ff),
	.w8(32'hb8f47e48),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a52de),
	.w1(32'h3b8a4cdf),
	.w2(32'hb91eb859),
	.w3(32'hbb8b4a45),
	.w4(32'h3b1512c7),
	.w5(32'hbb1bfa76),
	.w6(32'hbb6090cc),
	.w7(32'hba2ff676),
	.w8(32'hbb2c789c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398596e8),
	.w1(32'h3a0eb076),
	.w2(32'h39f15c59),
	.w3(32'h3a2f47aa),
	.w4(32'h3a4f483a),
	.w5(32'h39a3f250),
	.w6(32'h3a2f36e9),
	.w7(32'h3a29b018),
	.w8(32'hba12ef88),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b189d37),
	.w1(32'h3a2b7201),
	.w2(32'h3a9d0d22),
	.w3(32'h3ac64d07),
	.w4(32'h399487a0),
	.w5(32'h3a239293),
	.w6(32'h3a431041),
	.w7(32'h38fddaec),
	.w8(32'h3a112173),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8244c5),
	.w1(32'hbb476906),
	.w2(32'hbb1de54e),
	.w3(32'h39728ab0),
	.w4(32'hbae508ab),
	.w5(32'hba74db05),
	.w6(32'h3adeeb5a),
	.w7(32'hba494205),
	.w8(32'h39146fc8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be47d45),
	.w1(32'h3c0a104d),
	.w2(32'h3a57eec9),
	.w3(32'hbbb8dae2),
	.w4(32'h3ae49bab),
	.w5(32'hbb6f2451),
	.w6(32'h3a0c8183),
	.w7(32'h3ae214ec),
	.w8(32'hbbf42fb3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391723cc),
	.w1(32'hba16ac66),
	.w2(32'hba159a16),
	.w3(32'h3a810867),
	.w4(32'h3a190a75),
	.w5(32'h39b5e848),
	.w6(32'h3a50ff47),
	.w7(32'h3a1c6bc9),
	.w8(32'hb9d9c7ee),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b74ef),
	.w1(32'hb8c64e7c),
	.w2(32'hba795810),
	.w3(32'h3a317e47),
	.w4(32'h397f89d0),
	.w5(32'hba80ebea),
	.w6(32'h3a273799),
	.w7(32'h3a84ab0b),
	.w8(32'h3960ff01),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc388),
	.w1(32'hbbb6263e),
	.w2(32'hbbb5e6c8),
	.w3(32'hb9ff4489),
	.w4(32'h3a9abdfa),
	.w5(32'hbb1932d6),
	.w6(32'h3b29a645),
	.w7(32'hb9c68773),
	.w8(32'hbafa4bf9),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d2ab5),
	.w1(32'h3c0a61dd),
	.w2(32'h3bebf3ce),
	.w3(32'h3be23451),
	.w4(32'hb9ac773d),
	.w5(32'h3be3b394),
	.w6(32'h3b9e00f1),
	.w7(32'h3a9130e2),
	.w8(32'h3c1198fd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc03d3b),
	.w1(32'hbbc18fb1),
	.w2(32'h3c47014d),
	.w3(32'h3c6053e8),
	.w4(32'hbbad61e4),
	.w5(32'h3b65c637),
	.w6(32'h3bca5b7f),
	.w7(32'hbb7060d9),
	.w8(32'h3ba39f0e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ae666),
	.w1(32'hba2499f1),
	.w2(32'hba0a5876),
	.w3(32'h3a2b32cb),
	.w4(32'hba65d644),
	.w5(32'hb9d28f0f),
	.w6(32'h3a2da649),
	.w7(32'h3857f355),
	.w8(32'hb8926c90),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d534),
	.w1(32'h3c3398d8),
	.w2(32'h3a1884ac),
	.w3(32'hbba50399),
	.w4(32'h3ba98b74),
	.w5(32'h3b24d9b6),
	.w6(32'hbb0a9201),
	.w7(32'h3c328a08),
	.w8(32'hb7b4e2cc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ef51f),
	.w1(32'h3bdc6a90),
	.w2(32'hbbbf510e),
	.w3(32'hbbee7508),
	.w4(32'h3b81bd34),
	.w5(32'h3b20fd41),
	.w6(32'hb9692ef0),
	.w7(32'hbb48741f),
	.w8(32'hbc10a68d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cfa79),
	.w1(32'h3b84d69d),
	.w2(32'h3c0f7a05),
	.w3(32'hbb0058bd),
	.w4(32'hba1cd194),
	.w5(32'h3b5143b9),
	.w6(32'hbab973a9),
	.w7(32'h3b76e195),
	.w8(32'h3b74742a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadb324),
	.w1(32'hba02939a),
	.w2(32'h390c8ea3),
	.w3(32'hba12ed6a),
	.w4(32'h38b40c48),
	.w5(32'hba7b0e4e),
	.w6(32'hba2f3f72),
	.w7(32'hb950fd61),
	.w8(32'hba0347bc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8574fd3),
	.w1(32'h385b37ce),
	.w2(32'h3a2df6ea),
	.w3(32'h38b05f82),
	.w4(32'h3a03dd26),
	.w5(32'h3abdba6e),
	.w6(32'h39c53376),
	.w7(32'h3a001541),
	.w8(32'h3a00e82b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1171ac),
	.w1(32'h3a805d83),
	.w2(32'h3a85fd50),
	.w3(32'h3a2225a8),
	.w4(32'h3a1c6da1),
	.w5(32'h3a4f1ff8),
	.w6(32'h3a27d506),
	.w7(32'h3a4e9cd3),
	.w8(32'h3a56b6df),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b2b78),
	.w1(32'h3b637347),
	.w2(32'h3c4457eb),
	.w3(32'h3b04d9b9),
	.w4(32'h3924655c),
	.w5(32'h3c00c72d),
	.w6(32'hba04e693),
	.w7(32'h3b9b5e79),
	.w8(32'h3c03c32b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c4590),
	.w1(32'hbb09a0f1),
	.w2(32'h397fa302),
	.w3(32'hbaff123d),
	.w4(32'hbab73895),
	.w5(32'h3ab4aeea),
	.w6(32'hbb1aa782),
	.w7(32'hbadcd286),
	.w8(32'hba22dc96),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb7378),
	.w1(32'hbc27d8d0),
	.w2(32'hbbe03f8e),
	.w3(32'h3a98ede1),
	.w4(32'hbb138867),
	.w5(32'hbb37cdcc),
	.w6(32'h3adc5b86),
	.w7(32'hbb06601a),
	.w8(32'h3a7a6989),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf988c5),
	.w1(32'hbad7cde2),
	.w2(32'hbb4e97ec),
	.w3(32'h395437b3),
	.w4(32'hb9180ea8),
	.w5(32'hbb1e2049),
	.w6(32'hba07c7ad),
	.w7(32'h37a49daf),
	.w8(32'hbaf61bd9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad41c3a),
	.w1(32'h3bc36564),
	.w2(32'h3b9d6817),
	.w3(32'hbb2fcb39),
	.w4(32'h3b472af5),
	.w5(32'h3b53df4f),
	.w6(32'hbb256bad),
	.w7(32'h3b79cba2),
	.w8(32'h3b3b6538),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a11e8e),
	.w1(32'hbb3de1cb),
	.w2(32'h3acf9019),
	.w3(32'h3b90e8be),
	.w4(32'hba5710f0),
	.w5(32'h3b4265bb),
	.w6(32'h3b2a99ed),
	.w7(32'hba7a46a2),
	.w8(32'h3b4e62e0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82f5c2f),
	.w1(32'h3979fcbf),
	.w2(32'h39415e67),
	.w3(32'h36e2e8bf),
	.w4(32'h399a65de),
	.w5(32'h39f0905e),
	.w6(32'hb849cfd4),
	.w7(32'h39af7746),
	.w8(32'h39f60881),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c435fc5),
	.w1(32'h3b8d91c0),
	.w2(32'h3ac69244),
	.w3(32'h3bf4dadb),
	.w4(32'hb8d73813),
	.w5(32'hbb631c02),
	.w6(32'h3b3923d7),
	.w7(32'hb9d76425),
	.w8(32'hbb8d1c7a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b6efd),
	.w1(32'hb93ee4c2),
	.w2(32'hb72f332a),
	.w3(32'hb9e1dfdf),
	.w4(32'hb955ecf4),
	.w5(32'hb9157a55),
	.w6(32'hb943198b),
	.w7(32'hb9314609),
	.w8(32'hb8fca7e7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d750e),
	.w1(32'h3aad8eb5),
	.w2(32'h3a4b3e1c),
	.w3(32'hbad4e1ec),
	.w4(32'h3aa2084f),
	.w5(32'h3a957c25),
	.w6(32'hbb04560b),
	.w7(32'h3a8af71b),
	.w8(32'h3a9fb00a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1a072),
	.w1(32'hbc1a9722),
	.w2(32'hbc237be4),
	.w3(32'h3abe87eb),
	.w4(32'h3b70775a),
	.w5(32'hbab113aa),
	.w6(32'h3b6c34cb),
	.w7(32'h3b56e723),
	.w8(32'hb8f1f0bf),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2cfdf),
	.w1(32'hbb95d463),
	.w2(32'hbb7a2394),
	.w3(32'h3a28dc95),
	.w4(32'hba1bf186),
	.w5(32'hbae1e803),
	.w6(32'hb964b29e),
	.w7(32'hbab1e20b),
	.w8(32'hbaac3381),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d20e91),
	.w1(32'hba5266d9),
	.w2(32'hbacefc73),
	.w3(32'h38f9ce71),
	.w4(32'hba23a97c),
	.w5(32'hba6f6c73),
	.w6(32'h3a105de0),
	.w7(32'hba0ae14d),
	.w8(32'hba933d5e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a74a9),
	.w1(32'hbbc0327b),
	.w2(32'hbc0b6970),
	.w3(32'h39e634f9),
	.w4(32'h3a107400),
	.w5(32'hbb34f28c),
	.w6(32'hba7b0a82),
	.w7(32'hbb252922),
	.w8(32'hbb665b29),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b159c0a),
	.w1(32'h3b958c01),
	.w2(32'h3b2bc05a),
	.w3(32'hbb2d539c),
	.w4(32'h3a9702d8),
	.w5(32'hba696626),
	.w6(32'hbb450001),
	.w7(32'hb90df343),
	.w8(32'hba03aeaf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56a8e7),
	.w1(32'h3b214b35),
	.w2(32'h3ac8c2ea),
	.w3(32'hbb683092),
	.w4(32'h3a1855c8),
	.w5(32'h3a5e1668),
	.w6(32'hbb70139b),
	.w7(32'h3a2d2d26),
	.w8(32'h3835bc1d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b62dc),
	.w1(32'h396441e2),
	.w2(32'h395960a1),
	.w3(32'h39fba854),
	.w4(32'h38228d37),
	.w5(32'h38c72f54),
	.w6(32'h3a0e6e4d),
	.w7(32'hb83588de),
	.w8(32'h37887f25),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9b047),
	.w1(32'h39026138),
	.w2(32'h38840756),
	.w3(32'h38b78334),
	.w4(32'h396cabbf),
	.w5(32'h39a8d5e4),
	.w6(32'hb8f58dd9),
	.w7(32'hb907533b),
	.w8(32'h390fe89e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc781438),
	.w1(32'hbbcccb14),
	.w2(32'h3b48fd6c),
	.w3(32'h3a589ac5),
	.w4(32'h3b8ed781),
	.w5(32'h3c203392),
	.w6(32'hbba0e6e1),
	.w7(32'h3a771683),
	.w8(32'h3b176908),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4cafa),
	.w1(32'hbb4670c4),
	.w2(32'h39f19790),
	.w3(32'hbac175f4),
	.w4(32'h3b023eff),
	.w5(32'h3b825d74),
	.w6(32'hbb9dd2d8),
	.w7(32'h3b74b5a8),
	.w8(32'h3aaf49b8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6d3b),
	.w1(32'hbc0310ce),
	.w2(32'hbbd4dcba),
	.w3(32'hbb707bc2),
	.w4(32'hbb07ccdb),
	.w5(32'hb995c261),
	.w6(32'hbae98ff5),
	.w7(32'hbb23a1c0),
	.w8(32'hbae09f8b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a3946),
	.w1(32'h3c0ff80e),
	.w2(32'h3c6fce2c),
	.w3(32'hbbe84e4f),
	.w4(32'hbb1b9fcb),
	.w5(32'h3ba3b10a),
	.w6(32'hbb8c0e24),
	.w7(32'h3bbbe6e6),
	.w8(32'h3b1dbc3a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4ec9a),
	.w1(32'hb950242f),
	.w2(32'hba0088bb),
	.w3(32'h3a22bdf2),
	.w4(32'h39f27a86),
	.w5(32'h3a0497a9),
	.w6(32'h3abe091c),
	.w7(32'h3a96d3e3),
	.w8(32'hba39bcf5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198672),
	.w1(32'h3aea693d),
	.w2(32'h3a2017be),
	.w3(32'hba1b831d),
	.w4(32'hb99928ee),
	.w5(32'hba4336e5),
	.w6(32'hb93e814f),
	.w7(32'h3a54e208),
	.w8(32'hbac7fe17),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba092e0),
	.w1(32'hbbb6a385),
	.w2(32'h3cd9b641),
	.w3(32'h3c31c545),
	.w4(32'h395f41ce),
	.w5(32'h3cc26717),
	.w6(32'hbb13abbd),
	.w7(32'h3bdb1478),
	.w8(32'h3c8cd0fe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d83d8),
	.w1(32'h3be46fb1),
	.w2(32'h3b7ef464),
	.w3(32'hbbc25138),
	.w4(32'h3ac211fa),
	.w5(32'h3b533b30),
	.w6(32'hbb6a155d),
	.w7(32'h3b3bae43),
	.w8(32'h39e217f8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecbc0),
	.w1(32'h3b85f3a0),
	.w2(32'h3bf5749d),
	.w3(32'hbb77f9e7),
	.w4(32'hbb98ec91),
	.w5(32'h3ba8238a),
	.w6(32'hbbbd2e2e),
	.w7(32'hb9b5d96d),
	.w8(32'h3b4562c5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e5494),
	.w1(32'hbbf5eac2),
	.w2(32'hbc2a8c14),
	.w3(32'h3b5470d0),
	.w4(32'h3b42ed92),
	.w5(32'hbad8290f),
	.w6(32'h3b628c21),
	.w7(32'h3b3caaa8),
	.w8(32'hb981f301),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab71a06),
	.w1(32'hbbd551c6),
	.w2(32'hbc307b43),
	.w3(32'h3b717add),
	.w4(32'h3b99a6df),
	.w5(32'hba43c1c7),
	.w6(32'h3af30b46),
	.w7(32'h3af960df),
	.w8(32'hba7149df),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940f857),
	.w1(32'hb73a14c0),
	.w2(32'h38d5e11d),
	.w3(32'h387e55d2),
	.w4(32'h392abfa5),
	.w5(32'h39866d07),
	.w6(32'h39476f25),
	.w7(32'h39bebed6),
	.w8(32'h39906732),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396925d3),
	.w1(32'hb8d5195c),
	.w2(32'h390f8c0e),
	.w3(32'h399b1f62),
	.w4(32'hb98ce3ab),
	.w5(32'hb92f1d77),
	.w6(32'h39dfdd19),
	.w7(32'hb8bdebc1),
	.w8(32'h391b9086),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9b187),
	.w1(32'hbaa05055),
	.w2(32'hb920a270),
	.w3(32'hba3f783a),
	.w4(32'h3a55dff2),
	.w5(32'h3a224161),
	.w6(32'h39b2a8c3),
	.w7(32'h3ac1c6f4),
	.w8(32'hba9fadfe),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998ab88),
	.w1(32'hb86e4d62),
	.w2(32'h39efcc6c),
	.w3(32'hb9aea508),
	.w4(32'hb99a3560),
	.w5(32'h3903ad3b),
	.w6(32'hb9a32d56),
	.w7(32'hb9a591df),
	.w8(32'hb86f7fc8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac17e35),
	.w1(32'h3ba88610),
	.w2(32'h3bcf73a1),
	.w3(32'h3b4107b6),
	.w4(32'h3b660029),
	.w5(32'h3bb3dcac),
	.w6(32'hb8ce0100),
	.w7(32'h3b952306),
	.w8(32'h3ba4038d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d18c9),
	.w1(32'hbb27ab59),
	.w2(32'hba70a7d8),
	.w3(32'hbb731494),
	.w4(32'hbb1d5d58),
	.w5(32'h3b5b6775),
	.w6(32'hbb091ae1),
	.w7(32'h3b4c2006),
	.w8(32'hba0a143f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bda8),
	.w1(32'hbaa27aac),
	.w2(32'hba84ef16),
	.w3(32'hb9e976e5),
	.w4(32'hba2f383f),
	.w5(32'h3a0f1efe),
	.w6(32'hbacc591d),
	.w7(32'hb9217e85),
	.w8(32'h396cfa98),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5ecf9),
	.w1(32'hb8b35202),
	.w2(32'hb7c781d0),
	.w3(32'hb9997608),
	.w4(32'hb97651fa),
	.w5(32'hb812670a),
	.w6(32'hb86616b4),
	.w7(32'hb91baa12),
	.w8(32'h3858efcb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad722a),
	.w1(32'h3c672254),
	.w2(32'h3c7a861b),
	.w3(32'h3a082b8d),
	.w4(32'hbb04b1eb),
	.w5(32'h3bb94c55),
	.w6(32'hbbd88632),
	.w7(32'h3aba4f66),
	.w8(32'h3b7b19cc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03f547),
	.w1(32'h3b2f2af4),
	.w2(32'h3b2aa318),
	.w3(32'hbafef49c),
	.w4(32'h3ab95c2e),
	.w5(32'h3addabc4),
	.w6(32'hba5e449e),
	.w7(32'h3b41cb26),
	.w8(32'h3aed05a9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9567e02),
	.w1(32'hb7a07ea8),
	.w2(32'hb8bd6e12),
	.w3(32'hb99d3ede),
	.w4(32'hb9b357e5),
	.w5(32'hb908ea72),
	.w6(32'hb9a2f05e),
	.w7(32'h34e83c24),
	.w8(32'hb92f398a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b3086),
	.w1(32'h3c1536a6),
	.w2(32'h3be46b57),
	.w3(32'hbb39cc88),
	.w4(32'h3b02858e),
	.w5(32'h3b8e11ff),
	.w6(32'hbb4e183a),
	.w7(32'h3b0bb12f),
	.w8(32'h3b2084c9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940db78),
	.w1(32'h3a11c91f),
	.w2(32'h3a2bca91),
	.w3(32'h38b59d3c),
	.w4(32'h39d1dc44),
	.w5(32'h39ff1352),
	.w6(32'hb702223d),
	.w7(32'h39a64380),
	.w8(32'h39ef3a53),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c9bee),
	.w1(32'h3a04e69d),
	.w2(32'h3a226207),
	.w3(32'h39c0313d),
	.w4(32'hb8a1a798),
	.w5(32'h39ee77b4),
	.w6(32'h3a4fcf5d),
	.w7(32'h3a3b23fb),
	.w8(32'h39e6a0a1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92be84c),
	.w1(32'h393ac30c),
	.w2(32'h3969b234),
	.w3(32'h3916c713),
	.w4(32'hb837e4ce),
	.w5(32'h39c138ee),
	.w6(32'hb70565c5),
	.w7(32'h394cb2dd),
	.w8(32'h394bfed6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f26a7),
	.w1(32'hb988747d),
	.w2(32'hb9d446ed),
	.w3(32'h3999ee73),
	.w4(32'hb9e8f062),
	.w5(32'hb9a65dcc),
	.w6(32'h395f7cbf),
	.w7(32'h384c1aac),
	.w8(32'h36329adc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1b2be),
	.w1(32'hbb3fa1ac),
	.w2(32'hbafed941),
	.w3(32'h3a898e87),
	.w4(32'h3a946a4c),
	.w5(32'h3a4447e4),
	.w6(32'h3a17f4d6),
	.w7(32'h3aba8f68),
	.w8(32'h3767f1be),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f2a8b),
	.w1(32'h3c92614b),
	.w2(32'h3c045d0b),
	.w3(32'hbb8a0b78),
	.w4(32'h3b8b39c1),
	.w5(32'h3ba1526e),
	.w6(32'hbb3ffc55),
	.w7(32'h3b810e30),
	.w8(32'hbb069c1b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc9acd),
	.w1(32'h3bc1c91c),
	.w2(32'h3b426a10),
	.w3(32'hbbc065f1),
	.w4(32'h37a7929c),
	.w5(32'h3a1103c8),
	.w6(32'hbbc35204),
	.w7(32'hba9a723d),
	.w8(32'h39243a3e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39c38d),
	.w1(32'h3c767aad),
	.w2(32'h3c405783),
	.w3(32'hbb549ae6),
	.w4(32'h3b9abda7),
	.w5(32'h3bdbf16d),
	.w6(32'hbbab0d42),
	.w7(32'h3b05bc27),
	.w8(32'h3a28aa87),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53d821),
	.w1(32'h39dcfe8f),
	.w2(32'hb8b84597),
	.w3(32'h3a89f41c),
	.w4(32'h3a0c2a49),
	.w5(32'h38b23ca7),
	.w6(32'h3a9d37b4),
	.w7(32'h3a161fab),
	.w8(32'hb847d8f1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a701e6),
	.w1(32'h39d72832),
	.w2(32'h3a13a46c),
	.w3(32'hb95254c3),
	.w4(32'h396bcc44),
	.w5(32'hb87add88),
	.w6(32'h3a3e7ae4),
	.w7(32'h394bbaaa),
	.w8(32'hb738fe1b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdbca2),
	.w1(32'hb8c0231b),
	.w2(32'hb7f96578),
	.w3(32'hb97ba0de),
	.w4(32'hb88df187),
	.w5(32'h390c1fdf),
	.w6(32'hb9116cee),
	.w7(32'hb94a6005),
	.w8(32'hb85ce329),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f9f3e9),
	.w1(32'h39249045),
	.w2(32'h399ad8aa),
	.w3(32'h394b1b58),
	.w4(32'h39154cc1),
	.w5(32'h3958627e),
	.w6(32'hb70fc173),
	.w7(32'h3a0c8516),
	.w8(32'h39b86197),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2b5cd),
	.w1(32'h3b40333d),
	.w2(32'hba838f84),
	.w3(32'hbb388939),
	.w4(32'h3b30642f),
	.w5(32'hbb60d05b),
	.w6(32'h39ad8c7d),
	.w7(32'h39c7e2f2),
	.w8(32'hbbe3c4fb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62c3c0),
	.w1(32'hb75f75a9),
	.w2(32'hba039599),
	.w3(32'hba7725cd),
	.w4(32'hba028183),
	.w5(32'hba87bd77),
	.w6(32'hba348f91),
	.w7(32'hb9a98c7d),
	.w8(32'hba271b7e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab86c7f),
	.w1(32'h3a084d1c),
	.w2(32'h39ba0232),
	.w3(32'h3b0ba53e),
	.w4(32'h3a24566e),
	.w5(32'h3989df27),
	.w6(32'h3b00498d),
	.w7(32'h3a2da5df),
	.w8(32'hb922c924),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7fc5b),
	.w1(32'h3b2bd9a1),
	.w2(32'hba520b23),
	.w3(32'h3bbb5306),
	.w4(32'h3a85f0ec),
	.w5(32'hba760c13),
	.w6(32'h3b53b2e5),
	.w7(32'hba49a028),
	.w8(32'h38bc511e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a40b65),
	.w1(32'h38bf395e),
	.w2(32'h3871964c),
	.w3(32'h39cc4fe1),
	.w4(32'h38322c95),
	.w5(32'hb8bdde6f),
	.w6(32'h398ff0df),
	.w7(32'hb914392b),
	.w8(32'hb975e3d1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a364eb7),
	.w1(32'h3b06e591),
	.w2(32'h3ad96eee),
	.w3(32'hba735d30),
	.w4(32'h3a4f4462),
	.w5(32'h3a848285),
	.w6(32'hba42992a),
	.w7(32'h3a7cbf5e),
	.w8(32'h3a4e16ef),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398de940),
	.w1(32'h38542b39),
	.w2(32'h38b0e0dd),
	.w3(32'h3a5c5de6),
	.w4(32'h340abd76),
	.w5(32'h385285c7),
	.w6(32'h3a7768e0),
	.w7(32'h3a8f778e),
	.w8(32'h3a70e8e7),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a4100),
	.w1(32'h3c999be4),
	.w2(32'h3b1ab61f),
	.w3(32'hbc05305a),
	.w4(32'h3bb07f4d),
	.w5(32'hbbf9c4e6),
	.w6(32'hbb2b49b2),
	.w7(32'h3aad76aa),
	.w8(32'hbc514d59),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853151b),
	.w1(32'h39cfab20),
	.w2(32'h39c8d6f4),
	.w3(32'h38be95b0),
	.w4(32'h39fb79f9),
	.w5(32'h3a29da92),
	.w6(32'h398e5c4a),
	.w7(32'h3a054b67),
	.w8(32'h399359e2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32f374),
	.w1(32'hbc61ae05),
	.w2(32'hbbf69775),
	.w3(32'h3b0ca676),
	.w4(32'hbb30b40f),
	.w5(32'hba1153e6),
	.w6(32'h3a4c4eff),
	.w7(32'hbb113af0),
	.w8(32'hbb43a3ea),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule