module layer_6_featuremap_114(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b659),
	.w1(32'hbabf27cf),
	.w2(32'h3ac0d8a6),
	.w3(32'hbaa2c4dd),
	.w4(32'hbaaae6d9),
	.w5(32'h3a219df4),
	.w6(32'hba34fccd),
	.w7(32'h3b9f8480),
	.w8(32'h3b5ac6a0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21cef5),
	.w1(32'h3b22803a),
	.w2(32'h3bf7ccaf),
	.w3(32'h3a5ff357),
	.w4(32'h3ba66eed),
	.w5(32'h3c48d5e6),
	.w6(32'hbbada9fd),
	.w7(32'h3bc08e89),
	.w8(32'h3c6d3356),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31a3ff),
	.w1(32'h3c833f4e),
	.w2(32'h3d1b6845),
	.w3(32'hbca2b52c),
	.w4(32'hba9db74c),
	.w5(32'h3cb45cd5),
	.w6(32'hbca906e9),
	.w7(32'h3d34f54d),
	.w8(32'hba21ab41),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd11fb5c),
	.w1(32'hbb93f8d0),
	.w2(32'hbbd1e79b),
	.w3(32'hbad1dad0),
	.w4(32'hbbfaab2b),
	.w5(32'h3a02cc93),
	.w6(32'hbb5f5b2b),
	.w7(32'hbbcda353),
	.w8(32'h3b335a70),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45839e),
	.w1(32'h3b7a4274),
	.w2(32'h3bf5d1ca),
	.w3(32'hbc22e63d),
	.w4(32'hbc18c638),
	.w5(32'h3cb3c23e),
	.w6(32'h3b0da341),
	.w7(32'h3c2d4f6c),
	.w8(32'h3ca6948e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06b0d8),
	.w1(32'h3a3621ee),
	.w2(32'h3a6d1700),
	.w3(32'h3bb1c122),
	.w4(32'h3b6977fa),
	.w5(32'hbb2cbc00),
	.w6(32'h3b8b9b61),
	.w7(32'h3b443c3d),
	.w8(32'hbae81675),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980e761),
	.w1(32'h3be56fba),
	.w2(32'hba0f3366),
	.w3(32'h3b6fc77b),
	.w4(32'hbad13cb6),
	.w5(32'h3bb45919),
	.w6(32'h3b6d7782),
	.w7(32'h3aaffbab),
	.w8(32'h3bc16961),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3ec52),
	.w1(32'hbc688e52),
	.w2(32'hbc451536),
	.w3(32'h3c88f110),
	.w4(32'hbcd40a80),
	.w5(32'hbc222ec4),
	.w6(32'hbb98825a),
	.w7(32'hbcd01151),
	.w8(32'hbb9e2825),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b0d1f),
	.w1(32'h3a5863c9),
	.w2(32'h3c5aeffb),
	.w3(32'hbc9d4055),
	.w4(32'hbbf19d56),
	.w5(32'h3bfd592e),
	.w6(32'hbc8c1b72),
	.w7(32'h3c85a260),
	.w8(32'h3b58d658),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b143836),
	.w1(32'h3bc5e503),
	.w2(32'hbba6fab3),
	.w3(32'h3c44d1d3),
	.w4(32'hbb08d25b),
	.w5(32'hbbd70a8a),
	.w6(32'h3c265466),
	.w7(32'hbb6c2b6b),
	.w8(32'hbbca6465),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b210c),
	.w1(32'h3c8b9e21),
	.w2(32'h3c02fc2f),
	.w3(32'hbc820464),
	.w4(32'h3cc6faff),
	.w5(32'h3b4a2e13),
	.w6(32'h3c1b60a7),
	.w7(32'h3d52b77a),
	.w8(32'hbc6968bb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf1b9d5),
	.w1(32'hbb6dc8c0),
	.w2(32'h3a06f5ba),
	.w3(32'h3c488faa),
	.w4(32'h3c18f692),
	.w5(32'h3adad616),
	.w6(32'h3b96759e),
	.w7(32'h3baa5ca4),
	.w8(32'hb99236a6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5a723),
	.w1(32'hba48a81f),
	.w2(32'hbb9ad126),
	.w3(32'hbad02fa3),
	.w4(32'hbc1eb019),
	.w5(32'h3b1daddf),
	.w6(32'hbb67c76b),
	.w7(32'hbb34791a),
	.w8(32'h3b0d74f3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16cb5d),
	.w1(32'hb9be5884),
	.w2(32'h3b697581),
	.w3(32'hbc0f0e5a),
	.w4(32'hba15c5d6),
	.w5(32'h3ba98adf),
	.w6(32'hbc45356c),
	.w7(32'h3c3fe1cb),
	.w8(32'h3c7148e7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6d4cc),
	.w1(32'hbc52a84e),
	.w2(32'h3bb0b6c4),
	.w3(32'hbbe14fae),
	.w4(32'h3ad8f50d),
	.w5(32'h3c2e5727),
	.w6(32'hbc80c17d),
	.w7(32'h3c022292),
	.w8(32'h3c8087c3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c233f),
	.w1(32'hba6eac6b),
	.w2(32'h3b83685c),
	.w3(32'hbb86a7dc),
	.w4(32'hbb5395ad),
	.w5(32'h3a819614),
	.w6(32'hbbb60ea1),
	.w7(32'h3aaa92c4),
	.w8(32'h3b8e3420),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eae1b),
	.w1(32'hbc84f470),
	.w2(32'h3b893439),
	.w3(32'hbc97215d),
	.w4(32'h3c8104d1),
	.w5(32'hbba94606),
	.w6(32'hbc8387ce),
	.w7(32'h3c8b573b),
	.w8(32'hbc707d8c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca909d3),
	.w1(32'h3b5245cc),
	.w2(32'hbae1679c),
	.w3(32'h3c1bc8a3),
	.w4(32'h3b9e8e91),
	.w5(32'hbad1e159),
	.w6(32'h3be76c60),
	.w7(32'h39c0f684),
	.w8(32'hbb25ae05),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc1a6d),
	.w1(32'hba1d9de4),
	.w2(32'hbb06e296),
	.w3(32'h3b8750a0),
	.w4(32'hbb0c3ebf),
	.w5(32'hbb90e369),
	.w6(32'h3b30a514),
	.w7(32'hbb26746d),
	.w8(32'hbb14c6fb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac50558),
	.w1(32'h3b950f65),
	.w2(32'h3c896ebb),
	.w3(32'hbc2f661f),
	.w4(32'h3ce6a6a6),
	.w5(32'hbc9b06b4),
	.w6(32'h3bedc8a6),
	.w7(32'h3d0b2c33),
	.w8(32'hbcd092cf),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b8bfe),
	.w1(32'h3a3fbd86),
	.w2(32'h3b6bd52a),
	.w3(32'hbb162fb0),
	.w4(32'h3b18d000),
	.w5(32'h3af86e52),
	.w6(32'hbad9b1ca),
	.w7(32'h3bb81974),
	.w8(32'h3b051e0e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae85de0),
	.w1(32'hbbbb59c0),
	.w2(32'hbc82131f),
	.w3(32'hbc186616),
	.w4(32'h3b70d902),
	.w5(32'h3abd9e62),
	.w6(32'hbc086079),
	.w7(32'hbaca70bc),
	.w8(32'hba62f17b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0b27),
	.w1(32'hbb8b5585),
	.w2(32'h3b56c784),
	.w3(32'h3abfc69d),
	.w4(32'h3cb3d0ec),
	.w5(32'h3c0620f0),
	.w6(32'h3a12a9ea),
	.w7(32'h3b631140),
	.w8(32'h3ba3f40b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8c342),
	.w1(32'hbc76e474),
	.w2(32'hbc86996d),
	.w3(32'hbc918339),
	.w4(32'hbcdcf06e),
	.w5(32'h3cadfcd8),
	.w6(32'hbd194d49),
	.w7(32'hbcd47f4c),
	.w8(32'h3d075421),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c314db0),
	.w1(32'hbc176b72),
	.w2(32'hbcc3f8ea),
	.w3(32'hbc6c04ef),
	.w4(32'hbc46c1a5),
	.w5(32'h3c24c8d9),
	.w6(32'hbcbce962),
	.w7(32'hbc680a55),
	.w8(32'h3bbea098),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3073),
	.w1(32'hbc59430d),
	.w2(32'h3bfffd74),
	.w3(32'hbc01adb5),
	.w4(32'hbbc633d7),
	.w5(32'hbcbbbba9),
	.w6(32'hbc4e2af4),
	.w7(32'h3bf13d38),
	.w8(32'hbc928483),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63fdfd),
	.w1(32'h38487e5e),
	.w2(32'hbc42c3e2),
	.w3(32'hbb8ed33f),
	.w4(32'hbacbdcd3),
	.w5(32'h3c5af73b),
	.w6(32'hbbcb114e),
	.w7(32'hbba098fa),
	.w8(32'h3b672bef),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc61c16),
	.w1(32'hba541359),
	.w2(32'hbb57177b),
	.w3(32'hbb493fd0),
	.w4(32'hbb89c25b),
	.w5(32'hbb93394c),
	.w6(32'hbb6b4826),
	.w7(32'hbb13b9ec),
	.w8(32'hbb13e808),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb632384),
	.w1(32'hbb076e3c),
	.w2(32'h3ba64271),
	.w3(32'hbb8bf42e),
	.w4(32'h3acd8f3d),
	.w5(32'h3b69df11),
	.w6(32'hbb92f6bc),
	.w7(32'h3b3e439b),
	.w8(32'h3b9cd71f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb132b3),
	.w1(32'h3c666fa8),
	.w2(32'h3cf65c93),
	.w3(32'h3be9983d),
	.w4(32'h3b9d2bd3),
	.w5(32'h3bd01602),
	.w6(32'h3c29017b),
	.w7(32'hb905b248),
	.w8(32'hbbff0a7f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfde092),
	.w1(32'hba4a1fb1),
	.w2(32'hbb900bfd),
	.w3(32'hbc623f93),
	.w4(32'h3b4b584d),
	.w5(32'h3c7d6680),
	.w6(32'hba24899a),
	.w7(32'h3cca0078),
	.w8(32'h3c28aa9c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ea393),
	.w1(32'h3c151622),
	.w2(32'hbd0bd0d0),
	.w3(32'h3ce40fba),
	.w4(32'hbc820eb4),
	.w5(32'hbbcc4d2b),
	.w6(32'h3cb115bd),
	.w7(32'hbd15c69a),
	.w8(32'hbc71e308),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea94da),
	.w1(32'hbc15bf11),
	.w2(32'h3c63218f),
	.w3(32'hbcf5e6fd),
	.w4(32'h3c507b33),
	.w5(32'hbc1d5361),
	.w6(32'hbd238c3c),
	.w7(32'h3cd7269c),
	.w8(32'hbc83020b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd3f53),
	.w1(32'hbc4150b3),
	.w2(32'h3c4fb53a),
	.w3(32'hbc9c26a4),
	.w4(32'h3bd814c0),
	.w5(32'h3c0fa59f),
	.w6(32'hbc6ce633),
	.w7(32'h3c1f698e),
	.w8(32'hbbde41ea),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa0ef),
	.w1(32'h3aca7d67),
	.w2(32'hbbbf2190),
	.w3(32'h3bd58d89),
	.w4(32'h3a4a9a77),
	.w5(32'hbae3dadb),
	.w6(32'h3b987bfe),
	.w7(32'hbb643af4),
	.w8(32'hbba10fb3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc081f3e),
	.w1(32'hbbd12ef6),
	.w2(32'hbbe71c98),
	.w3(32'hb6e5a968),
	.w4(32'hbc5aa327),
	.w5(32'hbbd16131),
	.w6(32'hbc1220c1),
	.w7(32'hbc90017e),
	.w8(32'hbb869a22),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbc2c1),
	.w1(32'h3ae2ea2b),
	.w2(32'h3ae2e2d8),
	.w3(32'hb922cc6b),
	.w4(32'h3b92998b),
	.w5(32'h3a873c1d),
	.w6(32'h3b864e8a),
	.w7(32'h3b2cb2e3),
	.w8(32'hbaa14fc6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb814613),
	.w1(32'hbb1029f6),
	.w2(32'h3b78ff58),
	.w3(32'hb9f890da),
	.w4(32'h39cbb4a7),
	.w5(32'hbba05830),
	.w6(32'hba67c043),
	.w7(32'h3b5382b4),
	.w8(32'hbb4fb5bc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc82d6),
	.w1(32'h3c3ee48c),
	.w2(32'h3bb3948c),
	.w3(32'hbbaabb2d),
	.w4(32'hbb4ba452),
	.w5(32'h3c69a4af),
	.w6(32'h3b70411a),
	.w7(32'h3cc87997),
	.w8(32'h3c8e8159),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a972160),
	.w1(32'hbb8bae18),
	.w2(32'hb71c935e),
	.w3(32'hbcee619f),
	.w4(32'h3c412096),
	.w5(32'hbb592785),
	.w6(32'hbceeefc7),
	.w7(32'h3b2a2d8b),
	.w8(32'hbbe20ec5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37f84a),
	.w1(32'h3c71bc0d),
	.w2(32'hbd101700),
	.w3(32'h3c5950c4),
	.w4(32'h3c98a9b6),
	.w5(32'hbc93796b),
	.w6(32'h3d18fead),
	.w7(32'hb8ece9ac),
	.w8(32'hbcb98671),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133ecb),
	.w1(32'hbaf6f68e),
	.w2(32'hbb88eded),
	.w3(32'hbac8e806),
	.w4(32'hbbf94dd5),
	.w5(32'hb9498169),
	.w6(32'hbadcd9c2),
	.w7(32'hbb93e733),
	.w8(32'h3b21f8d2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b437004),
	.w1(32'h3be008b5),
	.w2(32'hbb57bdb9),
	.w3(32'h3bc840d7),
	.w4(32'h3bf4f072),
	.w5(32'h3b839e6a),
	.w6(32'h3c54cdab),
	.w7(32'h3bdd1bee),
	.w8(32'hb9fb0615),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf453af),
	.w1(32'h39cc4ad0),
	.w2(32'h3c59b7d3),
	.w3(32'h3bef3836),
	.w4(32'h3b8da594),
	.w5(32'h3aba5c35),
	.w6(32'h3c854fd1),
	.w7(32'hbc08ce8c),
	.w8(32'hbc14a3fa),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd156),
	.w1(32'hbbafbf49),
	.w2(32'hbb9a75a6),
	.w3(32'hbc3f2a75),
	.w4(32'h39d0ac08),
	.w5(32'h3be319a4),
	.w6(32'hbc0c1200),
	.w7(32'hba0064dd),
	.w8(32'h3bc4f4ba),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0bca5),
	.w1(32'h3c2d2d5c),
	.w2(32'hbd20dcc8),
	.w3(32'hbc337500),
	.w4(32'h3cffbaa9),
	.w5(32'h3bfefb15),
	.w6(32'h3c756ca4),
	.w7(32'h3d079d4a),
	.w8(32'hbd27e26d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd59f627),
	.w1(32'hbc471661),
	.w2(32'hbbedbe67),
	.w3(32'h3c24a1d7),
	.w4(32'hbb0be470),
	.w5(32'hbbac455e),
	.w6(32'hbc16be22),
	.w7(32'hbbe01c18),
	.w8(32'hbc08351a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72c25f),
	.w1(32'h3bf347f1),
	.w2(32'h3bb99271),
	.w3(32'hbc194cfc),
	.w4(32'h3b831b97),
	.w5(32'hb9c84fce),
	.w6(32'h3b59abed),
	.w7(32'h3d1300ce),
	.w8(32'hbc57cb8d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee8d12),
	.w1(32'hbc26b3ac),
	.w2(32'hba77c60a),
	.w3(32'hbb86c426),
	.w4(32'hbba6f72a),
	.w5(32'hbae57628),
	.w6(32'hbbc60b9d),
	.w7(32'hbb58cccf),
	.w8(32'h3b861b80),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53465a),
	.w1(32'h3badd03c),
	.w2(32'h3c46eb60),
	.w3(32'hba98b36c),
	.w4(32'hbb96e3f2),
	.w5(32'h3a98b868),
	.w6(32'hbbb3ffbc),
	.w7(32'h3c572951),
	.w8(32'h3ae0d8c7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a813f),
	.w1(32'hbb12b522),
	.w2(32'h3915662a),
	.w3(32'hba884cf5),
	.w4(32'hbb63127f),
	.w5(32'h3ab43468),
	.w6(32'hbb43001b),
	.w7(32'h3b058ece),
	.w8(32'h3bb97225),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f73c6),
	.w1(32'hbbde10fd),
	.w2(32'hbba7616c),
	.w3(32'hbb191d63),
	.w4(32'hbbd00b13),
	.w5(32'hbc2efeaa),
	.w6(32'hbb85bb45),
	.w7(32'hbb82aa2b),
	.w8(32'hbbe1c53c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf98bdc),
	.w1(32'hbc18cddf),
	.w2(32'hbb7b2579),
	.w3(32'hbc1b79ee),
	.w4(32'hbbc30e0c),
	.w5(32'h3bac2a7a),
	.w6(32'hbc49d915),
	.w7(32'hbae6b530),
	.w8(32'h3c274bdd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6469),
	.w1(32'h3a99108d),
	.w2(32'h3c704e07),
	.w3(32'hb9cecdd6),
	.w4(32'h3aeae55c),
	.w5(32'h3c17d4de),
	.w6(32'hbba10a6c),
	.w7(32'h3c27d092),
	.w8(32'h3c862425),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e9c80),
	.w1(32'h3ab892f1),
	.w2(32'hb99e0b56),
	.w3(32'h3a909378),
	.w4(32'hbb6dc0ca),
	.w5(32'h3b4af0fb),
	.w6(32'hbae64911),
	.w7(32'hbafb82b3),
	.w8(32'h3c1c2079),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad65e5c),
	.w1(32'hbb2c0b19),
	.w2(32'h3b574d89),
	.w3(32'h3c090e4b),
	.w4(32'hbafbc76e),
	.w5(32'hbc9cc488),
	.w6(32'h3c6208fb),
	.w7(32'h3c7fea09),
	.w8(32'h3ba7ffc5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c707d20),
	.w1(32'h3b1966a3),
	.w2(32'h3b93075b),
	.w3(32'hbb9ff0d4),
	.w4(32'hbb7b06a3),
	.w5(32'hbb1082fa),
	.w6(32'h3a31bd82),
	.w7(32'hbb54cc18),
	.w8(32'hbbc9d0dc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0489e),
	.w1(32'hbc243a8f),
	.w2(32'hbc61c65f),
	.w3(32'h3bd547e4),
	.w4(32'h3c3d3d55),
	.w5(32'h3b0c4a97),
	.w6(32'h3b80aef6),
	.w7(32'h3c6e7c14),
	.w8(32'h3b4ffedf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c624f3d),
	.w1(32'hbb659ba2),
	.w2(32'hbbcc946d),
	.w3(32'hba80911a),
	.w4(32'hbadb6bc8),
	.w5(32'hbaf0e9bb),
	.w6(32'hbb770ca2),
	.w7(32'hbb82a264),
	.w8(32'hbb0286f8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42dde1),
	.w1(32'hbcf6dbb3),
	.w2(32'hbcfda173),
	.w3(32'h3c887cc9),
	.w4(32'h3caf2c62),
	.w5(32'h3c8f8437),
	.w6(32'hbc3ddf3f),
	.w7(32'h3a225b2b),
	.w8(32'h3c32a6ab),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e7d9),
	.w1(32'hbbb136f0),
	.w2(32'hbc48c285),
	.w3(32'hbafedf2b),
	.w4(32'hbac91f33),
	.w5(32'hbba08808),
	.w6(32'hbbef4149),
	.w7(32'hbc377a57),
	.w8(32'hbc03f4be),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe70e72),
	.w1(32'hbc6f9ad7),
	.w2(32'hbcacb982),
	.w3(32'hbc92d5bb),
	.w4(32'hbcab33d0),
	.w5(32'hbc52c2ba),
	.w6(32'hbca70908),
	.w7(32'hbcf19c8d),
	.w8(32'hbcd07dde),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf921bd),
	.w1(32'hbc05d35c),
	.w2(32'h3cf81d4f),
	.w3(32'h3b8e4a04),
	.w4(32'h3b19e41f),
	.w5(32'h3c0e6d7a),
	.w6(32'h3c05a61a),
	.w7(32'h3ba5fe9a),
	.w8(32'hbce665c7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8e3e2),
	.w1(32'hbc889e65),
	.w2(32'hbc7d57b1),
	.w3(32'h3bf575df),
	.w4(32'h3c5abb2e),
	.w5(32'h3bcdd74e),
	.w6(32'hbc033642),
	.w7(32'h3bd95610),
	.w8(32'h3c4634e4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule