module layer_10_featuremap_139(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352306f7),
	.w1(32'h371c757b),
	.w2(32'h36cdc294),
	.w3(32'hb61063eb),
	.w4(32'h358ea317),
	.w5(32'h3717c561),
	.w6(32'h371259d2),
	.w7(32'h3672b234),
	.w8(32'hb56fee97),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3718ede1),
	.w1(32'hb7c39c04),
	.w2(32'h37a3c5bd),
	.w3(32'hb6388920),
	.w4(32'hb6f57a6c),
	.w5(32'h383d1c47),
	.w6(32'hb72f9a5d),
	.w7(32'h36a06e2c),
	.w8(32'h375debea),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5bdf2f5),
	.w1(32'h3676ec7d),
	.w2(32'h3594ae9f),
	.w3(32'hb59172f5),
	.w4(32'h357763fb),
	.w5(32'h35ed21de),
	.w6(32'h36adf281),
	.w7(32'h3520f1cc),
	.w8(32'h355122d7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363c02ad),
	.w1(32'hb78ae504),
	.w2(32'h369c1d1b),
	.w3(32'hb6fecc44),
	.w4(32'h3651a874),
	.w5(32'hb6acac49),
	.w6(32'h3661a0cb),
	.w7(32'hb786344d),
	.w8(32'hb674083e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65be1ce),
	.w1(32'hb6739d74),
	.w2(32'h374fa4da),
	.w3(32'hb6ad896c),
	.w4(32'hb6afbb1f),
	.w5(32'h36cae839),
	.w6(32'hb782feba),
	.w7(32'hb7a4622e),
	.w8(32'h34c487dd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361088aa),
	.w1(32'hb5b85ca5),
	.w2(32'hb67c23e6),
	.w3(32'hb2b5af90),
	.w4(32'hb393c58f),
	.w5(32'hb6c0e40a),
	.w6(32'h366bc7be),
	.w7(32'h36697637),
	.w8(32'h366ba94e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846d9e8),
	.w1(32'h38e861f7),
	.w2(32'h38787e08),
	.w3(32'h382d9318),
	.w4(32'h392517e0),
	.w5(32'h38f68e43),
	.w6(32'h39259ab9),
	.w7(32'h39394579),
	.w8(32'h38b2b290),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdafbe),
	.w1(32'h38eaacb1),
	.w2(32'hb8c704fe),
	.w3(32'hb96117e8),
	.w4(32'hb9339853),
	.w5(32'hb7d71db0),
	.w6(32'h39bb78ab),
	.w7(32'hb89e1e87),
	.w8(32'hb937215b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d064d4),
	.w1(32'h38296964),
	.w2(32'h36995f23),
	.w3(32'hb80b1565),
	.w4(32'hb822a148),
	.w5(32'hb708fbf2),
	.w6(32'hb858022d),
	.w7(32'hb7f920d5),
	.w8(32'hb638ff58),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385e148b),
	.w1(32'h38d14ced),
	.w2(32'h380baa82),
	.w3(32'hb8556406),
	.w4(32'hb7d8be73),
	.w5(32'hb82f7d93),
	.w6(32'hb8d95617),
	.w7(32'hb93c540b),
	.w8(32'hb7c9e940),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b55421),
	.w1(32'h373f2f61),
	.w2(32'h3764507c),
	.w3(32'h37ef1f24),
	.w4(32'h3762cd01),
	.w5(32'h3593d63a),
	.w6(32'hb7bacba5),
	.w7(32'hb86e55f5),
	.w8(32'h36c0b88f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902866a),
	.w1(32'h3877f58b),
	.w2(32'h38296c05),
	.w3(32'hb897d84b),
	.w4(32'h3924c3a9),
	.w5(32'h386209d3),
	.w6(32'h3927dcac),
	.w7(32'h392af781),
	.w8(32'h3878e4aa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824a012),
	.w1(32'h37f0d0a3),
	.w2(32'hb83935f3),
	.w3(32'hb89bc5f5),
	.w4(32'hb8cf3945),
	.w5(32'hb91edc24),
	.w6(32'hb885676d),
	.w7(32'hb915d460),
	.w8(32'hb87e6ca9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d50f44),
	.w1(32'h37f1256a),
	.w2(32'h38915758),
	.w3(32'hb69a09ba),
	.w4(32'h358c1a31),
	.w5(32'h38926ca7),
	.w6(32'hb81357c4),
	.w7(32'hb86a32b0),
	.w8(32'hb804d449),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4e570),
	.w1(32'hb73b6c70),
	.w2(32'hb7aef2a4),
	.w3(32'hb886fd01),
	.w4(32'hb8b0e494),
	.w5(32'hb7d8ef09),
	.w6(32'hb8c9ab46),
	.w7(32'hb8ac463d),
	.w8(32'hb8082cc2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aa5e33),
	.w1(32'hb899ac7f),
	.w2(32'hb93347ad),
	.w3(32'hb78a85fc),
	.w4(32'hb85e8440),
	.w5(32'hb9583dc8),
	.w6(32'hb8ca76f3),
	.w7(32'hb8d7c1f3),
	.w8(32'hb926ec41),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3646713e),
	.w1(32'hb6cb6cac),
	.w2(32'hb58ec81d),
	.w3(32'h3666ca42),
	.w4(32'hb61e100f),
	.w5(32'hb66351c2),
	.w6(32'h37135227),
	.w7(32'hb784086e),
	.w8(32'hb7969438),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ad5b2),
	.w1(32'h38b10aa5),
	.w2(32'hb9846c4d),
	.w3(32'h37836d8a),
	.w4(32'hb9187fba),
	.w5(32'hb9977b97),
	.w6(32'h39459bc9),
	.w7(32'h36b372f2),
	.w8(32'hb95b977d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5914b03),
	.w1(32'hb593aabf),
	.w2(32'hb8ffc366),
	.w3(32'hb898429f),
	.w4(32'hb8e4aa6a),
	.w5(32'hb918f19d),
	.w6(32'h38947a3c),
	.w7(32'hb7ae0671),
	.w8(32'hb8758010),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6507fac),
	.w1(32'hb69756e7),
	.w2(32'h3619345d),
	.w3(32'hb60aed73),
	.w4(32'h360e8aa9),
	.w5(32'h36f31760),
	.w6(32'h35e7ae29),
	.w7(32'h362d1a15),
	.w8(32'h36a4a8e4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb642b536),
	.w1(32'h354cb896),
	.w2(32'h34e1c0eb),
	.w3(32'h3592d1ee),
	.w4(32'hb45e464e),
	.w5(32'hb6108f16),
	.w6(32'h36a8a654),
	.w7(32'h3623586c),
	.w8(32'hb62b6c41),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79eaafa),
	.w1(32'hb6057dca),
	.w2(32'h375754f3),
	.w3(32'hb5982489),
	.w4(32'h353ed44d),
	.w5(32'h36ce118b),
	.w6(32'h37735e9d),
	.w7(32'h3733952d),
	.w8(32'h36761e33),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb9d8f),
	.w1(32'h38859809),
	.w2(32'hb89342a0),
	.w3(32'h39077837),
	.w4(32'h3848db37),
	.w5(32'hb9b7b7e2),
	.w6(32'h39054c6e),
	.w7(32'hb84491f8),
	.w8(32'hb8bd413a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379cfa60),
	.w1(32'hb6f18304),
	.w2(32'hb7f0728d),
	.w3(32'hb833a232),
	.w4(32'hb8977588),
	.w5(32'hb7f32dd0),
	.w6(32'hb86c1a8a),
	.w7(32'hb85e4296),
	.w8(32'h380b0c70),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90025f7),
	.w1(32'hb7d812dd),
	.w2(32'h37b3818d),
	.w3(32'hb893c7cc),
	.w4(32'hb6bcf51d),
	.w5(32'h38d52371),
	.w6(32'hb8cecfc6),
	.w7(32'h385bedc4),
	.w8(32'h38e9e979),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f05457),
	.w1(32'hb704919e),
	.w2(32'hb78c7b7c),
	.w3(32'hb7eeae01),
	.w4(32'hb8885e96),
	.w5(32'hb81d90ab),
	.w6(32'hb854c5fb),
	.w7(32'hb8a0fe4f),
	.w8(32'hb8098394),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb682735f),
	.w1(32'hb65f4eb0),
	.w2(32'hb6522792),
	.w3(32'hb6064c49),
	.w4(32'hb5f243f8),
	.w5(32'hb65bdfe3),
	.w6(32'hb5422440),
	.w7(32'hb57d3794),
	.w8(32'hb620602c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c0be0),
	.w1(32'hb7e5d52f),
	.w2(32'h362a9008),
	.w3(32'hb9622472),
	.w4(32'h38faf251),
	.w5(32'hb7940a66),
	.w6(32'hb981b538),
	.w7(32'hb92b6aa8),
	.w8(32'hb9015f87),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb2882),
	.w1(32'hb7ea58e1),
	.w2(32'hb775f805),
	.w3(32'hb6db35d1),
	.w4(32'hb73c8f52),
	.w5(32'hb60bca09),
	.w6(32'h365f6d80),
	.w7(32'hb7d05035),
	.w8(32'hb7e323ca),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916b735),
	.w1(32'hb89a306c),
	.w2(32'hb8ada572),
	.w3(32'hb92ba455),
	.w4(32'hb8c388de),
	.w5(32'hb7c325a7),
	.w6(32'hb9c93218),
	.w7(32'hb98fba46),
	.w8(32'hb8d72708),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73e4130),
	.w1(32'hb6160d18),
	.w2(32'hb68b5642),
	.w3(32'hb756a030),
	.w4(32'hb63c1fad),
	.w5(32'hb6925495),
	.w6(32'h3527a300),
	.w7(32'hb644499b),
	.w8(32'hb661d262),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ef75c4),
	.w1(32'hb693d297),
	.w2(32'hb3d5cc4e),
	.w3(32'hb6e85e37),
	.w4(32'hb6d9c834),
	.w5(32'hb618d78f),
	.w6(32'hb6906407),
	.w7(32'hb70586bc),
	.w8(32'h34708d24),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379c56eb),
	.w1(32'hb6be685d),
	.w2(32'hb81821bd),
	.w3(32'hb81fe023),
	.w4(32'hb889f0eb),
	.w5(32'hb81c3c5d),
	.w6(32'h37594fc6),
	.w7(32'hb83b5a7c),
	.w8(32'hb780c8b8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37904d85),
	.w1(32'h3804b39a),
	.w2(32'h37725cf0),
	.w3(32'hb748ae32),
	.w4(32'hb56a7d4b),
	.w5(32'h376cce35),
	.w6(32'hb7f88c77),
	.w7(32'hb7621bb3),
	.w8(32'hb52d84a9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8121c00),
	.w1(32'hb75d17eb),
	.w2(32'hb69edb7b),
	.w3(32'hb80eafd8),
	.w4(32'hb77483f3),
	.w5(32'hb7a1e458),
	.w6(32'hb73f9674),
	.w7(32'hb7ed4763),
	.w8(32'hb79fce47),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f7c72),
	.w1(32'h368220ff),
	.w2(32'h382235e0),
	.w3(32'h379cd3d8),
	.w4(32'h36863cd0),
	.w5(32'hb675a5db),
	.w6(32'h38b02b37),
	.w7(32'h389fe0c9),
	.w8(32'hb7b3c71c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b248a),
	.w1(32'h3923f7c5),
	.w2(32'h39d4afd7),
	.w3(32'hb80cdc8d),
	.w4(32'h3936a116),
	.w5(32'h39c23cff),
	.w6(32'h39d18041),
	.w7(32'h3994a979),
	.w8(32'h395a0c81),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937df0d),
	.w1(32'hb7ffe3e5),
	.w2(32'h3905590f),
	.w3(32'hb8c24bf7),
	.w4(32'h3854a93e),
	.w5(32'h392c314c),
	.w6(32'hb77f4660),
	.w7(32'h38c980da),
	.w8(32'h386c5356),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927a3cf),
	.w1(32'h3884ff8c),
	.w2(32'h39357f99),
	.w3(32'hb868ea71),
	.w4(32'h38de56a0),
	.w5(32'h39408a5f),
	.w6(32'hb88c9838),
	.w7(32'h3822d3d6),
	.w8(32'h38f0cbcf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a0592),
	.w1(32'hb8225dd4),
	.w2(32'hb7a7f14c),
	.w3(32'hb85929e6),
	.w4(32'hb82b4205),
	.w5(32'hb7cfd800),
	.w6(32'hb7b37404),
	.w7(32'hb7a17cee),
	.w8(32'hb7940d47),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368c81b6),
	.w1(32'h37a847b2),
	.w2(32'hb70f2140),
	.w3(32'hb6958bf0),
	.w4(32'h37955e44),
	.w5(32'hb7227ede),
	.w6(32'h376a9274),
	.w7(32'hb6f429f4),
	.w8(32'hb789499e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77eaef0),
	.w1(32'hb675ef32),
	.w2(32'hb6f29486),
	.w3(32'hb6f4a4a5),
	.w4(32'h3683e849),
	.w5(32'hb6f0609c),
	.w6(32'hb4404434),
	.w7(32'hb54a2e84),
	.w8(32'hb6d5fc09),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37158f8a),
	.w1(32'hb7cf2ce1),
	.w2(32'hb6f6a86a),
	.w3(32'h36a2d749),
	.w4(32'hb72a8e59),
	.w5(32'hb7817eb6),
	.w6(32'hb6adf095),
	.w7(32'hb8000a70),
	.w8(32'hb82ac0da),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36daf559),
	.w1(32'h37fbdc48),
	.w2(32'hb90284b8),
	.w3(32'hb95596f2),
	.w4(32'hb8fd320b),
	.w5(32'hb95f576c),
	.w6(32'hb960e504),
	.w7(32'hb939dade),
	.w8(32'hb8dc0a96),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6af11),
	.w1(32'hb8542c7d),
	.w2(32'hb789f375),
	.w3(32'hb8fa924b),
	.w4(32'hb90da4a5),
	.w5(32'hb6aeaf81),
	.w6(32'hb93219d8),
	.w7(32'hb8fc3682),
	.w8(32'h382a7298),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c39244),
	.w1(32'hb7e76bed),
	.w2(32'hb79e0ea9),
	.w3(32'hb86878b0),
	.w4(32'hb8ecf48e),
	.w5(32'hb7aed648),
	.w6(32'hb89f9e1d),
	.w7(32'hb7e1131c),
	.w8(32'h38c6cd78),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38573495),
	.w1(32'h38309336),
	.w2(32'hb7381f7c),
	.w3(32'hb4ac0eb7),
	.w4(32'h381ad3d3),
	.w5(32'hb799208a),
	.w6(32'hb782f8bb),
	.w7(32'h37dcfc07),
	.w8(32'h380a46ce),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a842a),
	.w1(32'hb7228af2),
	.w2(32'hb956db15),
	.w3(32'hb85f6d87),
	.w4(32'hb8e576ca),
	.w5(32'hb9523525),
	.w6(32'h3941000d),
	.w7(32'hb8593b62),
	.w8(32'hb918e47c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6880b05),
	.w1(32'h35e12cc0),
	.w2(32'hb6194929),
	.w3(32'hb700b20e),
	.w4(32'h36572d31),
	.w5(32'hb65d866d),
	.w6(32'hb5a6a153),
	.w7(32'h3695739c),
	.w8(32'h34f1c9f0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37799067),
	.w1(32'h37d2a691),
	.w2(32'hb785126c),
	.w3(32'h384fcfcc),
	.w4(32'h3856f8e0),
	.w5(32'hb778565c),
	.w6(32'h37d6449d),
	.w7(32'h3757f30d),
	.w8(32'hb73f45b3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3696249b),
	.w1(32'h36fdfb1d),
	.w2(32'hb742430f),
	.w3(32'hb65627c5),
	.w4(32'hb7675149),
	.w5(32'hb642d9e5),
	.w6(32'hb764290f),
	.w7(32'hb776ce22),
	.w8(32'hb68968db),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1639c),
	.w1(32'hb81bd130),
	.w2(32'hb7b4de69),
	.w3(32'hb7615f6b),
	.w4(32'hb881536c),
	.w5(32'hb7b961ff),
	.w6(32'hb7aaff13),
	.w7(32'hb84a0462),
	.w8(32'hb8151599),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb710acdd),
	.w1(32'h36a6f9ba),
	.w2(32'hb7c1089a),
	.w3(32'hb6f56f03),
	.w4(32'h371dac77),
	.w5(32'hb6583c38),
	.w6(32'h3790b4ea),
	.w7(32'h37cf66d6),
	.w8(32'h37697075),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb771172c),
	.w1(32'h38321613),
	.w2(32'hb917be52),
	.w3(32'hb908251d),
	.w4(32'hb8c40c60),
	.w5(32'hb9935a48),
	.w6(32'hb732cba2),
	.w7(32'hb939f763),
	.w8(32'hb946eb32),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ed32e4),
	.w1(32'h3784b157),
	.w2(32'hb7c16ad4),
	.w3(32'hb776fe9a),
	.w4(32'hb796a4fd),
	.w5(32'hb73e310f),
	.w6(32'h36f3d92b),
	.w7(32'h3738c2d3),
	.w8(32'h37f99f5f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7389ad5),
	.w1(32'h36f8bf5c),
	.w2(32'hb6efa586),
	.w3(32'hb790a22c),
	.w4(32'hb6d6df1b),
	.w5(32'hb785ed76),
	.w6(32'hb73a072e),
	.w7(32'hb7d3cf74),
	.w8(32'hb7fac783),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7028fd6),
	.w1(32'h35068dad),
	.w2(32'hb6da68cc),
	.w3(32'hb6d676b8),
	.w4(32'hb48fd3b5),
	.w5(32'hb6d7b522),
	.w6(32'h356c7a6d),
	.w7(32'hb6125632),
	.w8(32'hb6edcda8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d0e5b2),
	.w1(32'hb6c51f7b),
	.w2(32'h37268e9b),
	.w3(32'hb7762838),
	.w4(32'h36e20eea),
	.w5(32'h3649c6ca),
	.w6(32'hb75d5dcf),
	.w7(32'h3685e71b),
	.w8(32'h3683a3d3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66968f3),
	.w1(32'hb722c0dc),
	.w2(32'hb71bd634),
	.w3(32'h36f99d20),
	.w4(32'hb70a221d),
	.w5(32'hb7286100),
	.w6(32'hb615d907),
	.w7(32'hb7489490),
	.w8(32'hb7b5b6ea),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb734089f),
	.w1(32'h33ff1d76),
	.w2(32'h369815d1),
	.w3(32'hb7fdd5d8),
	.w4(32'hb7370348),
	.w5(32'hb7877600),
	.w6(32'hb833fca5),
	.w7(32'hb7a87d8b),
	.w8(32'hb6823595),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d88d4b),
	.w1(32'h37944af2),
	.w2(32'hb84a95e7),
	.w3(32'h36e9c879),
	.w4(32'h3733175e),
	.w5(32'hb8b3ffeb),
	.w6(32'h384f57b3),
	.w7(32'h37d78ed7),
	.w8(32'hb7f60014),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb862f655),
	.w1(32'h379609cb),
	.w2(32'hb8e13bc7),
	.w3(32'hb7eecc5b),
	.w4(32'hb7632cad),
	.w5(32'hb9199cf7),
	.w6(32'hb903991c),
	.w7(32'hb8e11ac3),
	.w8(32'hb8c2f414),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6101517),
	.w1(32'h37380beb),
	.w2(32'h35f4e4f8),
	.w3(32'hb6705b7a),
	.w4(32'h36fb9fd3),
	.w5(32'h361cad04),
	.w6(32'h3726bdb6),
	.w7(32'h361eae70),
	.w8(32'hb58bbd90),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b3ed37),
	.w1(32'h35ef94c2),
	.w2(32'hb569c489),
	.w3(32'hb5c78989),
	.w4(32'h353692bf),
	.w5(32'hb5047e2f),
	.w6(32'hb57c3d86),
	.w7(32'hb69300da),
	.w8(32'hb68090e7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c9f298),
	.w1(32'hb6fdd97d),
	.w2(32'hb722cc6a),
	.w3(32'hb6cb0a62),
	.w4(32'hb72098b3),
	.w5(32'hb71fe1eb),
	.w6(32'hb62f8e3b),
	.w7(32'hb66ddd61),
	.w8(32'hb65f987f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb586756a),
	.w1(32'hb5cf9be8),
	.w2(32'h369ab32c),
	.w3(32'hb5700b64),
	.w4(32'h355a73ae),
	.w5(32'h35abe34d),
	.w6(32'hb5897b76),
	.w7(32'h36dab6c8),
	.w8(32'hb5eb7dde),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7df17d6),
	.w1(32'hb8f63c60),
	.w2(32'hb9472ec1),
	.w3(32'hb967aa6f),
	.w4(32'hb890b59d),
	.w5(32'hb9a645e6),
	.w6(32'hb8a4de77),
	.w7(32'hb9ab8818),
	.w8(32'hb9a5eefe),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ffb378),
	.w1(32'hb63f043e),
	.w2(32'hb80c42ac),
	.w3(32'h38b1e0c9),
	.w4(32'hb8658626),
	.w5(32'hb80a7b20),
	.w6(32'h394937d3),
	.w7(32'h3904a865),
	.w8(32'h38dd6298),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88296fc),
	.w1(32'h377ba9e2),
	.w2(32'hb884af75),
	.w3(32'h3898cb54),
	.w4(32'hb87dea39),
	.w5(32'hb8a3b976),
	.w6(32'h389479e2),
	.w7(32'h385555e0),
	.w8(32'h389336d4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960a316),
	.w1(32'h35fa6840),
	.w2(32'h39832705),
	.w3(32'hb91867a7),
	.w4(32'hb5e89df7),
	.w5(32'h395bc33b),
	.w6(32'hb97b3381),
	.w7(32'hb8b49be1),
	.w8(32'h38f41f8b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b90f78),
	.w1(32'hb484c055),
	.w2(32'hb6c278f8),
	.w3(32'h36b097b4),
	.w4(32'hb67c50ac),
	.w5(32'hb6a7b52c),
	.w6(32'hb608270f),
	.w7(32'hb69a11e1),
	.w8(32'hb6c8d28a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6be96f3),
	.w1(32'hb4fbe92a),
	.w2(32'hb6cb99c1),
	.w3(32'hb69bbe91),
	.w4(32'hb4f6ec1f),
	.w5(32'hb6df0656),
	.w6(32'h3520e80a),
	.w7(32'hb598872c),
	.w8(32'hb5e730d3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64f870d),
	.w1(32'hb60fa6e1),
	.w2(32'hb65f3dec),
	.w3(32'hb556b024),
	.w4(32'h351adaf2),
	.w5(32'hb6918985),
	.w6(32'h351c9dee),
	.w7(32'h3623edbc),
	.w8(32'hb51257f4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36667bdc),
	.w1(32'hb7b390cd),
	.w2(32'hb89cd64c),
	.w3(32'hb8a2eabf),
	.w4(32'hb8943b58),
	.w5(32'hb8423ead),
	.w6(32'hb6645599),
	.w7(32'hb7777ced),
	.w8(32'hb81c99bd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4bff9ff),
	.w1(32'h36907c5f),
	.w2(32'hb5e9e9b4),
	.w3(32'h351e97a5),
	.w4(32'h36a2e1cf),
	.w5(32'hb60bacbf),
	.w6(32'h36db778d),
	.w7(32'h36467c6d),
	.w8(32'hb5275bd1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bcc91b),
	.w1(32'hb792f4e0),
	.w2(32'hb83236de),
	.w3(32'hb89391be),
	.w4(32'hb75917ee),
	.w5(32'hb8740840),
	.w6(32'h38d700a7),
	.w7(32'h36a826bb),
	.w8(32'hb8040519),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378aacaa),
	.w1(32'hb80cbbbd),
	.w2(32'hb8882b3d),
	.w3(32'hb8811203),
	.w4(32'hb8fbd13e),
	.w5(32'hb8c7f764),
	.w6(32'h397088c1),
	.w7(32'h391992d7),
	.w8(32'hb62e504a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902aded),
	.w1(32'hb8b48082),
	.w2(32'hb7e94553),
	.w3(32'hb9112811),
	.w4(32'hb90202e0),
	.w5(32'hb81e9bf7),
	.w6(32'hb91faea2),
	.w7(32'hb8d2a496),
	.w8(32'h3783f2ad),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3820ff13),
	.w1(32'h3891c246),
	.w2(32'hb7f213c2),
	.w3(32'hb8b8f908),
	.w4(32'hb890f301),
	.w5(32'hb8641a60),
	.w6(32'hb8a130f8),
	.w7(32'hb90a8793),
	.w8(32'hb8916b08),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f5ff6f),
	.w1(32'hb85126f0),
	.w2(32'h3667bc9b),
	.w3(32'hb8e975a9),
	.w4(32'hb7ed18c4),
	.w5(32'hb7964f03),
	.w6(32'hb8321f21),
	.w7(32'hb8d556b9),
	.w8(32'hb868744b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b2404f),
	.w1(32'h3800b7be),
	.w2(32'hb7062a60),
	.w3(32'hb8741251),
	.w4(32'hb7805537),
	.w5(32'hb750b9d9),
	.w6(32'hb88a4323),
	.w7(32'hb85cf454),
	.w8(32'h360d6d0d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a6148),
	.w1(32'h3737232a),
	.w2(32'hb7cc09c9),
	.w3(32'hb823437a),
	.w4(32'hb7b25dd3),
	.w5(32'hb857ee34),
	.w6(32'h38a41658),
	.w7(32'h37c1eba4),
	.w8(32'hb79b7d4e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a927f6),
	.w1(32'h35e351b0),
	.w2(32'hb62a5adf),
	.w3(32'hb63439cf),
	.w4(32'h368d2544),
	.w5(32'hb4f4c512),
	.w6(32'h362f0d81),
	.w7(32'hb5c63be7),
	.w8(32'hb676443f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ce5152),
	.w1(32'h36a8f012),
	.w2(32'h36019305),
	.w3(32'hb58e9b31),
	.w4(32'h36084d53),
	.w5(32'h361d8c62),
	.w6(32'h36b72367),
	.w7(32'h36afe91b),
	.w8(32'h36de8d67),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3610edde),
	.w1(32'h375e364b),
	.w2(32'hb54515ca),
	.w3(32'h35359661),
	.w4(32'h379ee7fe),
	.w5(32'h35a6378f),
	.w6(32'h373b617e),
	.w7(32'hb67e55b0),
	.w8(32'hb6db8b49),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71e55c6),
	.w1(32'h37738a7a),
	.w2(32'h37116be8),
	.w3(32'h3715bd64),
	.w4(32'h37acf76a),
	.w5(32'h374b8ed0),
	.w6(32'h36bcb145),
	.w7(32'h372fa9bf),
	.w8(32'h36b5c19d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e99567),
	.w1(32'hb85b90a3),
	.w2(32'h37fa1ac5),
	.w3(32'hb8e93acb),
	.w4(32'hb8a977b5),
	.w5(32'hb806f8c2),
	.w6(32'hb8e809e8),
	.w7(32'hb878b8f3),
	.w8(32'h380a57d4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7597b4d),
	.w1(32'hb7d400da),
	.w2(32'hb824322f),
	.w3(32'hb7db3843),
	.w4(32'hb76cb90d),
	.w5(32'hb72c78fb),
	.w6(32'hb575cbb3),
	.w7(32'hb79485d2),
	.w8(32'hb7b1360b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89923ac),
	.w1(32'h382fec16),
	.w2(32'h36f8b080),
	.w3(32'hb7ce3131),
	.w4(32'hb8b0dc68),
	.w5(32'hb8d39a1d),
	.w6(32'hb922a328),
	.w7(32'hb8ca6e70),
	.w8(32'hb7d29551),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ae754b),
	.w1(32'h37cb665d),
	.w2(32'hb887cd69),
	.w3(32'hb58c55b5),
	.w4(32'h38297173),
	.w5(32'hb8d2abca),
	.w6(32'h39388ba3),
	.w7(32'h3892f53e),
	.w8(32'hb8087e49),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a271ba),
	.w1(32'hb783e305),
	.w2(32'h38aadc97),
	.w3(32'hb9004bba),
	.w4(32'h377b984f),
	.w5(32'h38277489),
	.w6(32'hb8a5aec8),
	.w7(32'hb7ec051f),
	.w8(32'h38942ef5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9043dfe),
	.w1(32'h389b7bec),
	.w2(32'h38c60507),
	.w3(32'hb6c9745f),
	.w4(32'h37efabcd),
	.w5(32'hb92bd72a),
	.w6(32'hb91f9296),
	.w7(32'hb8d7e1e4),
	.w8(32'hb8932ac2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a4bfe0),
	.w1(32'hb7c61a55),
	.w2(32'h388d6acc),
	.w3(32'hb87f399c),
	.w4(32'hb786283d),
	.w5(32'h3847b93e),
	.w6(32'h3797a840),
	.w7(32'h38014862),
	.w8(32'h38cb9878),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39671cea),
	.w1(32'h39622fa2),
	.w2(32'hb8dd5eb0),
	.w3(32'hb848c9e8),
	.w4(32'hb8f1ec05),
	.w5(32'hb9ae7e98),
	.w6(32'hb91516e5),
	.w7(32'hb9bbd152),
	.w8(32'hb9fe66e6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90712ee),
	.w1(32'hb89f6839),
	.w2(32'hb5b13ad4),
	.w3(32'hb8692f19),
	.w4(32'h37c277c5),
	.w5(32'hb8556b7d),
	.w6(32'hb8e40838),
	.w7(32'hb8441463),
	.w8(32'h37efe918),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8920176),
	.w1(32'hb80d4dc8),
	.w2(32'hb81723ad),
	.w3(32'hb8e8257d),
	.w4(32'hb8af3cc9),
	.w5(32'hb7fd9ddd),
	.w6(32'hb940a8d0),
	.w7(32'hb9060f1e),
	.w8(32'hb880e22f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb724a432),
	.w1(32'hb7ea22ba),
	.w2(32'hb86e71cb),
	.w3(32'hb7e7172d),
	.w4(32'hb80eb81d),
	.w5(32'hb862dbf6),
	.w6(32'h370ad32f),
	.w7(32'hb874c5c9),
	.w8(32'hb869173a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3853b2c1),
	.w1(32'h37e285cf),
	.w2(32'hb926ea29),
	.w3(32'hb84f7579),
	.w4(32'hb90b6699),
	.w5(32'hb907bf6f),
	.w6(32'h38d1e4c4),
	.w7(32'hb6a620c0),
	.w8(32'hb8366ee3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb786f7b9),
	.w1(32'hb89479a9),
	.w2(32'hb89b5952),
	.w3(32'hb8a2dc9f),
	.w4(32'h38aeaccc),
	.w5(32'hb8eeb415),
	.w6(32'h386003b0),
	.w7(32'hb8a2b897),
	.w8(32'hb71027d4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910890a),
	.w1(32'hb7b8a9f7),
	.w2(32'h39fc3da7),
	.w3(32'h39951036),
	.w4(32'h38f86eff),
	.w5(32'h391dfaf7),
	.w6(32'h399f0b45),
	.w7(32'h39bc18c6),
	.w8(32'hb7d8945c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398aa20c),
	.w1(32'h39bceb42),
	.w2(32'h3906f0a0),
	.w3(32'h384c710c),
	.w4(32'h387fa99f),
	.w5(32'hb8abdc1e),
	.w6(32'hb9b102a8),
	.w7(32'hb9abdc52),
	.w8(32'hb8173a73),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c669fd),
	.w1(32'hb82e76b9),
	.w2(32'hb85edb42),
	.w3(32'hb8ad46ac),
	.w4(32'hb929b7b3),
	.w5(32'hb7053505),
	.w6(32'hb9451f1a),
	.w7(32'hb89b169a),
	.w8(32'h38823fb9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f9639b),
	.w1(32'h393ce17a),
	.w2(32'h390fc5ba),
	.w3(32'h379890ed),
	.w4(32'h391edb19),
	.w5(32'h38bf4f38),
	.w6(32'h38fe7ea8),
	.w7(32'h388386d1),
	.w8(32'h36803c4f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af2637),
	.w1(32'hb769db38),
	.w2(32'hb84f4f92),
	.w3(32'hb7b86e4c),
	.w4(32'hb74706a3),
	.w5(32'hb7ca7364),
	.w6(32'hb776c788),
	.w7(32'hb8132ba5),
	.w8(32'hb7fccbc3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997efce),
	.w1(32'hb78f9c97),
	.w2(32'h39c5bbdd),
	.w3(32'h363da697),
	.w4(32'h38421ea0),
	.w5(32'h3983c5a6),
	.w6(32'h39b73027),
	.w7(32'h3906347d),
	.w8(32'h36ef5dbf),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385d5779),
	.w1(32'h388cc865),
	.w2(32'h390516a5),
	.w3(32'h380397dc),
	.w4(32'h382421e1),
	.w5(32'h38f7bcdc),
	.w6(32'h392a1ac6),
	.w7(32'h392e9082),
	.w8(32'h390161ea),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a0900c),
	.w1(32'h36571a47),
	.w2(32'h36c3a08a),
	.w3(32'hb6cde3fa),
	.w4(32'hb548e763),
	.w5(32'h3630617e),
	.w6(32'hb6af6138),
	.w7(32'hb6ed8c13),
	.w8(32'hb6a904e3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a297f4),
	.w1(32'hb71a9b9c),
	.w2(32'hb7355cdb),
	.w3(32'hb6ea1f22),
	.w4(32'hb756f66e),
	.w5(32'hb67b6984),
	.w6(32'h35e89094),
	.w7(32'h377a216a),
	.w8(32'h378b3af8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c4480d),
	.w1(32'h3695fd72),
	.w2(32'hb898ef73),
	.w3(32'hb90bbae5),
	.w4(32'hb91def8c),
	.w5(32'hb8ff455d),
	.w6(32'hb84bf742),
	.w7(32'hb8a49d4e),
	.w8(32'hb899970f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b884e),
	.w1(32'hb7f1d434),
	.w2(32'hb7c7440a),
	.w3(32'hb90d62ad),
	.w4(32'hb8c728c2),
	.w5(32'h37e40c28),
	.w6(32'hb900a832),
	.w7(32'hb85d2dda),
	.w8(32'h3829b74a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37334956),
	.w1(32'h38383233),
	.w2(32'h3683a5cc),
	.w3(32'hb7003d7e),
	.w4(32'hb68a9627),
	.w5(32'hb7c106d2),
	.w6(32'hb8a5dd2b),
	.w7(32'hb886b3a1),
	.w8(32'h37f33afc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7852650),
	.w1(32'h38e70ead),
	.w2(32'h37b3cb10),
	.w3(32'hb8a277a5),
	.w4(32'hb755b772),
	.w5(32'hb8e3f3f7),
	.w6(32'hb8ec8790),
	.w7(32'hb8e7316a),
	.w8(32'hb9144fc1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96af3ba),
	.w1(32'hb8e99a1c),
	.w2(32'hb8707e4e),
	.w3(32'hb6326037),
	.w4(32'hb8858c12),
	.w5(32'hb78a1461),
	.w6(32'h386fe451),
	.w7(32'h38ccce89),
	.w8(32'hb7777b52),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37651687),
	.w1(32'hb5d9f590),
	.w2(32'hb8e564c8),
	.w3(32'h3801a027),
	.w4(32'hb83e90a5),
	.w5(32'hb927925f),
	.w6(32'hb94bf9e5),
	.w7(32'hb962f716),
	.w8(32'hb955609c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aed431),
	.w1(32'hb7530e3a),
	.w2(32'hb7bce853),
	.w3(32'hb871d474),
	.w4(32'hb8e18274),
	.w5(32'hb80fbc99),
	.w6(32'hb8d873b0),
	.w7(32'hb8d797d2),
	.w8(32'hb7a242aa),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb635cf7a),
	.w1(32'h36faaeb3),
	.w2(32'h36994ba7),
	.w3(32'hb5a9e487),
	.w4(32'h3776023b),
	.w5(32'h36ac20fe),
	.w6(32'h36b63296),
	.w7(32'h36bad12d),
	.w8(32'h3709cd56),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379c7e07),
	.w1(32'hb69e1875),
	.w2(32'hb6261193),
	.w3(32'hb6984175),
	.w4(32'hb63d7f1f),
	.w5(32'h354d927d),
	.w6(32'hb75cf7d6),
	.w7(32'hb7282352),
	.w8(32'hb6978ecc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5260d11),
	.w1(32'hb5a541e5),
	.w2(32'hb610178c),
	.w3(32'hb5b9d9ce),
	.w4(32'h34f7a69b),
	.w5(32'hb660f929),
	.w6(32'h36306c16),
	.w7(32'h35e5217d),
	.w8(32'h35c8f1ac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c9adbf),
	.w1(32'h36ef298e),
	.w2(32'hb58adb67),
	.w3(32'h3618f4f7),
	.w4(32'hb69633a3),
	.w5(32'hb7227786),
	.w6(32'hb734aa03),
	.w7(32'hb724692c),
	.w8(32'hb6856dc5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8364939),
	.w1(32'hb8160ef3),
	.w2(32'hb841f821),
	.w3(32'hb89cfc15),
	.w4(32'hb8a77546),
	.w5(32'hb7a5581a),
	.w6(32'hb8da4bc3),
	.w7(32'hb88be675),
	.w8(32'h3739201c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a1da92),
	.w1(32'h3785bc8c),
	.w2(32'h38561f78),
	.w3(32'hb823895b),
	.w4(32'h3833cf95),
	.w5(32'h377db899),
	.w6(32'hb85aa0e5),
	.w7(32'hb844b6a0),
	.w8(32'hb6b68f67),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc4fac),
	.w1(32'hb6c6577c),
	.w2(32'hb851789f),
	.w3(32'hb7c3e6db),
	.w4(32'h361faeb6),
	.w5(32'hb86c5d98),
	.w6(32'h38e79c05),
	.w7(32'h3880690e),
	.w8(32'hb7d4081e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d27120),
	.w1(32'hb895f3c0),
	.w2(32'hb839b092),
	.w3(32'hb887326b),
	.w4(32'hb75d2994),
	.w5(32'h37361401),
	.w6(32'hb8a07fe8),
	.w7(32'hb743b2fb),
	.w8(32'hb80ead05),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a1f112),
	.w1(32'h369ae2eb),
	.w2(32'h362ebcb1),
	.w3(32'hb5c9a8f2),
	.w4(32'hb71b6704),
	.w5(32'hb69ef257),
	.w6(32'hb4bda873),
	.w7(32'h35d06db1),
	.w8(32'h36391641),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71e8b8a),
	.w1(32'hb5cabbd7),
	.w2(32'hb6454152),
	.w3(32'hb488ab00),
	.w4(32'h36a03083),
	.w5(32'h348fde4f),
	.w6(32'h378ebc83),
	.w7(32'h37102370),
	.w8(32'h3745ff04),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a7c799),
	.w1(32'h35d7d3fc),
	.w2(32'hb4ac2c82),
	.w3(32'hb6202116),
	.w4(32'h36200b06),
	.w5(32'h34d172df),
	.w6(32'h3699a0c2),
	.w7(32'h348d7d48),
	.w8(32'hb52965fc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb797b7ec),
	.w1(32'hbaf7aded),
	.w2(32'hb9eb30e8),
	.w3(32'hb70582d9),
	.w4(32'hb9ccbefe),
	.w5(32'h3a07cc73),
	.w6(32'hbaa39e96),
	.w7(32'hb9d3f48c),
	.w8(32'h38be229a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ad73e),
	.w1(32'hb8f5b3a8),
	.w2(32'hb99e2f2e),
	.w3(32'h3a773a06),
	.w4(32'hb981594b),
	.w5(32'hb9ee374a),
	.w6(32'h390b137b),
	.w7(32'hb9a2d3ea),
	.w8(32'h3a1a76a0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a461328),
	.w1(32'hb93d5663),
	.w2(32'hb940b65a),
	.w3(32'h3a1e8c31),
	.w4(32'h3949d6c3),
	.w5(32'h3adca802),
	.w6(32'hbb0ec428),
	.w7(32'hbb154b8d),
	.w8(32'hbb45b13a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b609),
	.w1(32'h3a020d88),
	.w2(32'h3a3811b7),
	.w3(32'hb9ccaacc),
	.w4(32'h39f0bfb8),
	.w5(32'h3a287267),
	.w6(32'h3a36486e),
	.w7(32'h39f78fea),
	.w8(32'hb9016140),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a895c1),
	.w1(32'h3a95ebaa),
	.w2(32'h3a875c77),
	.w3(32'hb96e9633),
	.w4(32'hb9e6418d),
	.w5(32'hba5b0308),
	.w6(32'hba001c45),
	.w7(32'hba9477c2),
	.w8(32'hba8a16ed),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986324d),
	.w1(32'hbb606ca4),
	.w2(32'hbba3a1aa),
	.w3(32'hba9e0dc9),
	.w4(32'h3a9537ba),
	.w5(32'hb9bb1d7b),
	.w6(32'h3894eac5),
	.w7(32'hba70a7da),
	.w8(32'hbaf24c41),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e4daa),
	.w1(32'hbb380b1a),
	.w2(32'hb9f16b30),
	.w3(32'hbac46468),
	.w4(32'hbb0609df),
	.w5(32'hb9d99f5c),
	.w6(32'hbab89183),
	.w7(32'hb9af13d3),
	.w8(32'h3af7523d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dbe81),
	.w1(32'h3a38a302),
	.w2(32'h39f1d0c6),
	.w3(32'h3a83886e),
	.w4(32'hba54950f),
	.w5(32'hba9b3ddf),
	.w6(32'h3a82e8c9),
	.w7(32'h3a30a074),
	.w8(32'h3abd63b7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af389e3),
	.w1(32'h398b107d),
	.w2(32'h3a88ae07),
	.w3(32'h37537dc4),
	.w4(32'h39cafb41),
	.w5(32'h3a0fed9e),
	.w6(32'h3a1b150f),
	.w7(32'h3aa075c4),
	.w8(32'h3a27a94e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39def4e0),
	.w1(32'h39be3d3c),
	.w2(32'hb9288daf),
	.w3(32'h3995a3ad),
	.w4(32'h373dc4d5),
	.w5(32'hb9bd53e0),
	.w6(32'h39874581),
	.w7(32'hb9ff2c98),
	.w8(32'h3a14eaf9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a588861),
	.w1(32'hba950cd3),
	.w2(32'hba7c07b8),
	.w3(32'h3a5bd006),
	.w4(32'hba116936),
	.w5(32'hba11f70c),
	.w6(32'hba15ac71),
	.w7(32'hba16c862),
	.w8(32'hb859bbbb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80a3cb),
	.w1(32'h3a7b7a47),
	.w2(32'hb9e2948d),
	.w3(32'hb8bea07e),
	.w4(32'h38ba1daa),
	.w5(32'hbb022c4e),
	.w6(32'h3a9160c9),
	.w7(32'h397d074d),
	.w8(32'hb923dd1a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c6280),
	.w1(32'h3bafad3d),
	.w2(32'h3bace6c0),
	.w3(32'hbb0138db),
	.w4(32'hbaa40229),
	.w5(32'hbaa46282),
	.w6(32'hbad96b5a),
	.w7(32'hb9ddaf51),
	.w8(32'h3a234c12),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b905888),
	.w1(32'hbad5c990),
	.w2(32'hbb498971),
	.w3(32'hbb0d4e6c),
	.w4(32'hbb22c240),
	.w5(32'hbb20d67f),
	.w6(32'hbaba87b1),
	.w7(32'hbb194d79),
	.w8(32'hbac9f5e6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87bf43),
	.w1(32'hb9ece7fc),
	.w2(32'h3a842d35),
	.w3(32'hbaf9738b),
	.w4(32'hb88279b9),
	.w5(32'h3a480ee8),
	.w6(32'hbaa9e5bb),
	.w7(32'hba52cad2),
	.w8(32'hba82b515),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2f5fa),
	.w1(32'h39ee10da),
	.w2(32'hbab92c50),
	.w3(32'h3903850f),
	.w4(32'h3a0f98a4),
	.w5(32'hbab7b875),
	.w6(32'h3933ba18),
	.w7(32'hbac93d2d),
	.w8(32'h3a0974f9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc60b7),
	.w1(32'hbb1b2901),
	.w2(32'hbb641a1b),
	.w3(32'h38ee28d4),
	.w4(32'hbb123772),
	.w5(32'hba82556f),
	.w6(32'hbb25accc),
	.w7(32'hba8c5afd),
	.w8(32'h3ae12805),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9daab2),
	.w1(32'hba53ac6a),
	.w2(32'hba2f72a5),
	.w3(32'h3a555b63),
	.w4(32'hb9f6f2aa),
	.w5(32'hb9cdc4ac),
	.w6(32'hb98a8cc9),
	.w7(32'hb99fe2b4),
	.w8(32'hb9a2927c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49347d),
	.w1(32'h3b8f0d14),
	.w2(32'h3bd49ec2),
	.w3(32'h3777a4e0),
	.w4(32'hbb4b5e01),
	.w5(32'hba9b6981),
	.w6(32'h3ab8995c),
	.w7(32'h3b1786a6),
	.w8(32'h3b448e88),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beed47f),
	.w1(32'h39c205ee),
	.w2(32'hb957ed96),
	.w3(32'h3a69062c),
	.w4(32'h3970c33e),
	.w5(32'hba417e7d),
	.w6(32'h3a065df8),
	.w7(32'h39be2e8e),
	.w8(32'h39a1e455),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b89f5),
	.w1(32'hba00a90e),
	.w2(32'hb90e9fb7),
	.w3(32'hba18acc7),
	.w4(32'hba32e4bd),
	.w5(32'hba689e9e),
	.w6(32'hb9809471),
	.w7(32'hb964c3fe),
	.w8(32'hba54afd2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45420a),
	.w1(32'hba9038aa),
	.w2(32'hbaa4fc14),
	.w3(32'hba41a197),
	.w4(32'hba8b3d97),
	.w5(32'hbaa8bb45),
	.w6(32'hba4e891c),
	.w7(32'hba772e9f),
	.w8(32'hba57176e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91fa9a),
	.w1(32'hb9b7da7e),
	.w2(32'hbb23101f),
	.w3(32'hba3c78dd),
	.w4(32'h3aa37e04),
	.w5(32'hba9590f5),
	.w6(32'h399fd3a2),
	.w7(32'hbafb6699),
	.w8(32'hba1cd37b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afe5aa),
	.w1(32'h3b6e8531),
	.w2(32'hb950cae1),
	.w3(32'h39f6074b),
	.w4(32'h3b03bb91),
	.w5(32'h3a5770ab),
	.w6(32'hb9eae00a),
	.w7(32'hba25cf00),
	.w8(32'hb9d67202),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa236f2),
	.w1(32'h3b00971f),
	.w2(32'h3ae13acc),
	.w3(32'h3a41c648),
	.w4(32'hba9557b2),
	.w5(32'hbb1b579b),
	.w6(32'h3bcafa7d),
	.w7(32'h3bb7c920),
	.w8(32'h3bbf6020),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec2593),
	.w1(32'h390e0135),
	.w2(32'hb9f053d2),
	.w3(32'hbb55e961),
	.w4(32'h39054164),
	.w5(32'hb9898949),
	.w6(32'h398fa945),
	.w7(32'hba0d0a60),
	.w8(32'h38ec0ca9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393503bb),
	.w1(32'hba2d26a7),
	.w2(32'hb9fa37ab),
	.w3(32'h39e25831),
	.w4(32'hb9bc559d),
	.w5(32'hb8adc036),
	.w6(32'hb7c6bd0e),
	.w7(32'hb9be1b3e),
	.w8(32'hba5da110),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cf5a1),
	.w1(32'h3bb97bed),
	.w2(32'h3befc293),
	.w3(32'hba5e0734),
	.w4(32'hbb505371),
	.w5(32'hba95fcac),
	.w6(32'h3b0a3ce2),
	.w7(32'h3b5430d8),
	.w8(32'h3aca6e20),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb63c05),
	.w1(32'hbab0bde6),
	.w2(32'hbaad4764),
	.w3(32'hbae13f9d),
	.w4(32'hba86a4de),
	.w5(32'hba89a7bf),
	.w6(32'hba851392),
	.w7(32'hba427c57),
	.w8(32'hba4328b9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9895af),
	.w1(32'hbb0b7d9c),
	.w2(32'hbb14cfe0),
	.w3(32'hba378960),
	.w4(32'hbb1f2e7a),
	.w5(32'hbab82722),
	.w6(32'hbae9af3b),
	.w7(32'hbaea3b19),
	.w8(32'hbb0f7518),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294493),
	.w1(32'h3b527e4f),
	.w2(32'h3932978c),
	.w3(32'hbb01ace9),
	.w4(32'hba827457),
	.w5(32'hbba97aee),
	.w6(32'h3b1b1431),
	.w7(32'hba22957c),
	.w8(32'h3ab0f2c8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1536ce),
	.w1(32'h3bd2d89c),
	.w2(32'h3b465a4a),
	.w3(32'hbb2dd98a),
	.w4(32'h3ba68262),
	.w5(32'h3b4e7b15),
	.w6(32'h3bb96b74),
	.w7(32'h3afccd15),
	.w8(32'h3b7577fc),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f7270),
	.w1(32'hba130a5e),
	.w2(32'hba85ec3a),
	.w3(32'h3b3de59e),
	.w4(32'h398f7b39),
	.w5(32'hb9df2776),
	.w6(32'hba45274c),
	.w7(32'hbaca4da8),
	.w8(32'hba16c9be),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39076655),
	.w1(32'hb8d18ecf),
	.w2(32'hb688ffe9),
	.w3(32'h3a0b81fd),
	.w4(32'hb98fddee),
	.w5(32'hba0ee33e),
	.w6(32'hb930764e),
	.w7(32'hb992d0f6),
	.w8(32'hb9340bc5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dbe19),
	.w1(32'hbaac3e09),
	.w2(32'hb9ca5fa3),
	.w3(32'hb9163f96),
	.w4(32'hba931861),
	.w5(32'hba530f66),
	.w6(32'hbaf51a33),
	.w7(32'hbac25c1b),
	.w8(32'hbb12af79),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248085),
	.w1(32'hbb44ffb3),
	.w2(32'h3b8a73ca),
	.w3(32'hbb2f48c7),
	.w4(32'hbad724de),
	.w5(32'h3b37a928),
	.w6(32'hbb4f264e),
	.w7(32'h3b5b2dbd),
	.w8(32'hbb350192),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440588),
	.w1(32'h382244c0),
	.w2(32'hb9ca0533),
	.w3(32'hba9b8d29),
	.w4(32'hba4846c4),
	.w5(32'hbab0cf1b),
	.w6(32'hb9e6d171),
	.w7(32'hb9bd60c6),
	.w8(32'hba89ad83),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3760e5),
	.w1(32'hba993366),
	.w2(32'hba8f7cab),
	.w3(32'hbad2e7f0),
	.w4(32'hba38a3a6),
	.w5(32'hba6936f9),
	.w6(32'hba955ef8),
	.w7(32'hba9b4636),
	.w8(32'hba083fa0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af3eb4),
	.w1(32'hb9d5ada1),
	.w2(32'hb9abc2e3),
	.w3(32'hb9faa496),
	.w4(32'h36b6899e),
	.w5(32'hb93d2073),
	.w6(32'h389a5f1d),
	.w7(32'h38963aac),
	.w8(32'h395c868d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954cbf6),
	.w1(32'h3a3238df),
	.w2(32'h3ac22a1c),
	.w3(32'hb9daf902),
	.w4(32'h3a28c23a),
	.w5(32'h3a82cc07),
	.w6(32'h3a15c1f5),
	.w7(32'h3a9b04f6),
	.w8(32'h399de0c9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d058a),
	.w1(32'hb9a64337),
	.w2(32'hba1076f4),
	.w3(32'h3925cd96),
	.w4(32'hb7f3657f),
	.w5(32'hb8f4dd6b),
	.w6(32'hb9091702),
	.w7(32'hba0c40de),
	.w8(32'h38d53c94),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39457f07),
	.w1(32'hb9720c66),
	.w2(32'h39f5c541),
	.w3(32'h3a0fe210),
	.w4(32'hb7ffc42e),
	.w5(32'h39ddd8ad),
	.w6(32'hb938471d),
	.w7(32'h3a03569b),
	.w8(32'h39483851),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8afa36c),
	.w1(32'h3b810dfc),
	.w2(32'h39360a9d),
	.w3(32'h39467622),
	.w4(32'h3ba6479c),
	.w5(32'h3b46f36e),
	.w6(32'h3be134dc),
	.w7(32'h3af34c66),
	.w8(32'h3b6b1b78),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfb175),
	.w1(32'h38d9a3e9),
	.w2(32'hb6be531e),
	.w3(32'h3b0d8e16),
	.w4(32'hba7c8fd2),
	.w5(32'hba4abedc),
	.w6(32'hba508c85),
	.w7(32'hba32bd0c),
	.w8(32'hba4cb15f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1d314),
	.w1(32'hb9d08040),
	.w2(32'h3900d7b3),
	.w3(32'hbaa0c2e3),
	.w4(32'hba1fa00f),
	.w5(32'hb9b687fa),
	.w6(32'hba581730),
	.w7(32'hba4f939c),
	.w8(32'hba8f5f7c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0fd7d),
	.w1(32'h3b45919a),
	.w2(32'h3a28fc21),
	.w3(32'hba22291b),
	.w4(32'h3ad26f4b),
	.w5(32'hba642f61),
	.w6(32'h3b7c4fea),
	.w7(32'h3b092c24),
	.w8(32'h3b3df2b3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad21a22),
	.w1(32'hb930f5d9),
	.w2(32'hbacd1e0b),
	.w3(32'hb9b82ec1),
	.w4(32'h3aa5b1e8),
	.w5(32'hb9a41c5b),
	.w6(32'hb9d180fc),
	.w7(32'hb9436167),
	.w8(32'h38e3e028),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e07b9),
	.w1(32'hbabc92e6),
	.w2(32'hba63b721),
	.w3(32'hba93f2f9),
	.w4(32'hbaab9113),
	.w5(32'hbade5d33),
	.w6(32'hbaab620a),
	.w7(32'hba96df03),
	.w8(32'hbaa2d759),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab54134),
	.w1(32'hbad7d2dd),
	.w2(32'hbb894cfd),
	.w3(32'hbab345ba),
	.w4(32'h3981ca3a),
	.w5(32'h3a5454a8),
	.w6(32'hb9c941ec),
	.w7(32'h3a357df9),
	.w8(32'h3aa1f2d6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6c3a2),
	.w1(32'h3bb77f3a),
	.w2(32'h3b757f79),
	.w3(32'h3b067344),
	.w4(32'hbb125117),
	.w5(32'hbba9f84e),
	.w6(32'h3b13d34b),
	.w7(32'h3a1724b9),
	.w8(32'h3b0126c4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb66cce),
	.w1(32'hb9be6bea),
	.w2(32'h39dd0390),
	.w3(32'hbb331db0),
	.w4(32'hba706a14),
	.w5(32'hba3bf38f),
	.w6(32'hba43e08c),
	.w7(32'hb78b1cd8),
	.w8(32'hba65755a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb2a61),
	.w1(32'h399b8cd8),
	.w2(32'hb9e19acf),
	.w3(32'hba9b1958),
	.w4(32'h39e519c0),
	.w5(32'hb9142a8b),
	.w6(32'h39837989),
	.w7(32'hba271223),
	.w8(32'h39c25e44),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0873ef),
	.w1(32'h39a0cb32),
	.w2(32'hb99dca37),
	.w3(32'h3a809837),
	.w4(32'hb957924a),
	.w5(32'hba89adab),
	.w6(32'h3774a512),
	.w7(32'hba5fe301),
	.w8(32'hb9563760),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ce7b6),
	.w1(32'hb9be4bf1),
	.w2(32'h3a0e6f3b),
	.w3(32'hb9648d32),
	.w4(32'hba704ae7),
	.w5(32'h3aefef96),
	.w6(32'h39971c25),
	.w7(32'hbaa5f1b7),
	.w8(32'hbb3cb21f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13a8db),
	.w1(32'h39ffe1d8),
	.w2(32'hba69c725),
	.w3(32'hba90768c),
	.w4(32'h396a9e2f),
	.w5(32'hba535ce8),
	.w6(32'h3ac470cd),
	.w7(32'hba1cc3bc),
	.w8(32'hba1acf64),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce8e19),
	.w1(32'hbb58afb3),
	.w2(32'h387b578a),
	.w3(32'hba4f1f55),
	.w4(32'hbb24d30d),
	.w5(32'hbabd0841),
	.w6(32'hbae4c07d),
	.w7(32'h38dfb6b4),
	.w8(32'h3abbabac),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c33d2),
	.w1(32'h3a5e1479),
	.w2(32'h3af61a4b),
	.w3(32'hbaa24cc9),
	.w4(32'hb6ac84ea),
	.w5(32'h3a56b9e6),
	.w6(32'h3a357dc6),
	.w7(32'h3adcf295),
	.w8(32'hb99ec6d3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ced667),
	.w1(32'h3b04d3bc),
	.w2(32'hbb9c9191),
	.w3(32'hba630e58),
	.w4(32'h3bdb533d),
	.w5(32'h39f372ae),
	.w6(32'h3bed63ef),
	.w7(32'h3968c72e),
	.w8(32'h3bbbc104),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a787647),
	.w1(32'h3b17ca6b),
	.w2(32'h3ad07ddd),
	.w3(32'h3b87c6ac),
	.w4(32'h3ad0cbbd),
	.w5(32'h3aa497a0),
	.w6(32'h3b0015e8),
	.w7(32'h3aa30ed7),
	.w8(32'h39a34d26),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f2c57),
	.w1(32'hbb874502),
	.w2(32'h39a1f57f),
	.w3(32'h3a1a4019),
	.w4(32'hbb6e9317),
	.w5(32'hba8bfbb5),
	.w6(32'hbb115fa2),
	.w7(32'hba4fc5ef),
	.w8(32'h3a792a68),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91105e1),
	.w1(32'hb9b5de05),
	.w2(32'hb9ac5806),
	.w3(32'h39c8df10),
	.w4(32'h38834b3d),
	.w5(32'h37b99163),
	.w6(32'hb935f690),
	.w7(32'h39b834b1),
	.w8(32'h38f730e2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5bf81),
	.w1(32'hb8c536e8),
	.w2(32'hba0d133d),
	.w3(32'hb937df4d),
	.w4(32'h39633d84),
	.w5(32'hb91f430c),
	.w6(32'h390ba63d),
	.w7(32'hb9d6ecaf),
	.w8(32'hb851d726),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818c9b4),
	.w1(32'hb94c643a),
	.w2(32'h3882c4a1),
	.w3(32'h39a20240),
	.w4(32'hba3cef18),
	.w5(32'hba208ee4),
	.w6(32'hb9d117b6),
	.w7(32'hb9818a91),
	.w8(32'hb9bdcf04),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd7a89),
	.w1(32'h39b59cfd),
	.w2(32'hba1ce0ac),
	.w3(32'hba20bcf0),
	.w4(32'h3acbd668),
	.w5(32'h3a8f9b89),
	.w6(32'hb8c667a9),
	.w7(32'hba832f5e),
	.w8(32'hba086bcf),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99084e9),
	.w1(32'hba15e9be),
	.w2(32'h3a61cffb),
	.w3(32'h3a7357b5),
	.w4(32'hb977a149),
	.w5(32'h3afd5441),
	.w6(32'hbada5bc7),
	.w7(32'hba1676c4),
	.w8(32'hbb3a58a5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7286a5),
	.w1(32'h3ae83b4a),
	.w2(32'h39d1835b),
	.w3(32'hbb63a7a5),
	.w4(32'h3a3675ed),
	.w5(32'hba561cf9),
	.w6(32'h3b14da73),
	.w7(32'h3aa690f8),
	.w8(32'h3ace6d5c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b54e8),
	.w1(32'hba370757),
	.w2(32'hba7aaf8a),
	.w3(32'hba28271e),
	.w4(32'hba1bbd38),
	.w5(32'hbab55828),
	.w6(32'hb9c54284),
	.w7(32'hba52d536),
	.w8(32'hba7960b1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7e656),
	.w1(32'hbb59eab2),
	.w2(32'h3aeb3477),
	.w3(32'hbabe996a),
	.w4(32'hbb32195f),
	.w5(32'h3a7b1b09),
	.w6(32'hbb02992b),
	.w7(32'h388ac90a),
	.w8(32'hb5a495f8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0930a6),
	.w1(32'h3b0f7000),
	.w2(32'h3af593d4),
	.w3(32'h39bcd464),
	.w4(32'h3b71d1db),
	.w5(32'h3b970bd4),
	.w6(32'h3b3cde71),
	.w7(32'h3b2dc294),
	.w8(32'h3b790982),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d4a70),
	.w1(32'h3b5c2eb7),
	.w2(32'h3b7365de),
	.w3(32'h3b8111b3),
	.w4(32'h3b66376e),
	.w5(32'h3b82d16d),
	.w6(32'h3bd8754b),
	.w7(32'h3bbff340),
	.w8(32'h3b442e0a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9c230),
	.w1(32'h39942bba),
	.w2(32'hba3fd989),
	.w3(32'h39e89470),
	.w4(32'h39fd0211),
	.w5(32'h38de3d93),
	.w6(32'h3a3d7739),
	.w7(32'hb98ba983),
	.w8(32'hb965432f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980043e),
	.w1(32'hbb2977c1),
	.w2(32'hba6d628c),
	.w3(32'h39f8e50f),
	.w4(32'hbb1b3143),
	.w5(32'hbb1d4409),
	.w6(32'hbafa0fdb),
	.w7(32'hba8e5f7b),
	.w8(32'hb8d8c254),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ccb96),
	.w1(32'h38f71927),
	.w2(32'hb91bf2ec),
	.w3(32'hba77d54b),
	.w4(32'hb9420647),
	.w5(32'hba2d9986),
	.w6(32'hb93d6106),
	.w7(32'hb98cacd8),
	.w8(32'hb9c71ede),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e4912),
	.w1(32'hb9c00fad),
	.w2(32'hb9ed50de),
	.w3(32'hba23fd84),
	.w4(32'hb880dba6),
	.w5(32'hb87b5af8),
	.w6(32'h380ca80a),
	.w7(32'hb9872e03),
	.w8(32'h3a3c2928),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e552b),
	.w1(32'hb90f5bf4),
	.w2(32'hba036e2d),
	.w3(32'h3a47053d),
	.w4(32'h392a8896),
	.w5(32'hb8a17d79),
	.w6(32'h38a70117),
	.w7(32'hb9e76e1e),
	.w8(32'hb8230495),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384acb23),
	.w1(32'hb8dbaa6c),
	.w2(32'hb9aca245),
	.w3(32'h3a11ea6f),
	.w4(32'hb9d4b8e7),
	.w5(32'hba8d2942),
	.w6(32'hba4d8fe2),
	.w7(32'hbaaf7b17),
	.w8(32'hba578902),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a336949),
	.w1(32'h371930f3),
	.w2(32'hb91c3a03),
	.w3(32'hba13451e),
	.w4(32'hb97a156b),
	.w5(32'hb9b8266a),
	.w6(32'hb78e5fda),
	.w7(32'hb9620324),
	.w8(32'hba260c5d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e198),
	.w1(32'h3ac5612d),
	.w2(32'h3aa25f96),
	.w3(32'hba763782),
	.w4(32'hbab170ef),
	.w5(32'h3af7263f),
	.w6(32'h3a26e10f),
	.w7(32'h3a1f2ac5),
	.w8(32'hb9fe301a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6e23),
	.w1(32'h3a5700ee),
	.w2(32'hba475d83),
	.w3(32'hba27bd4a),
	.w4(32'h3a30413c),
	.w5(32'hba55c51b),
	.w6(32'h3a9e79e3),
	.w7(32'hb9de1507),
	.w8(32'h3ac9ce5c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6126),
	.w1(32'hb9872dac),
	.w2(32'hba31992a),
	.w3(32'h3a94b9bd),
	.w4(32'hba213363),
	.w5(32'hba36419a),
	.w6(32'hba244b6c),
	.w7(32'hba3601c0),
	.w8(32'hba77517e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab43eec),
	.w1(32'h3b28e229),
	.w2(32'h3b94ed67),
	.w3(32'hbaa19b3a),
	.w4(32'hbb4291a0),
	.w5(32'hbac72f4b),
	.w6(32'h39a66a3c),
	.w7(32'h3a97c715),
	.w8(32'hb9e54ef8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05b85c),
	.w1(32'hbacf5b63),
	.w2(32'hbb05fbe6),
	.w3(32'hbb272d3f),
	.w4(32'hb9548c6d),
	.w5(32'hba9670ac),
	.w6(32'hbaafdea7),
	.w7(32'hbb0988f0),
	.w8(32'hb9ad36e1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ef67bc),
	.w1(32'h3a10f6f8),
	.w2(32'hba2c507a),
	.w3(32'h3a23c434),
	.w4(32'h3b435595),
	.w5(32'h3aab6376),
	.w6(32'h3bf3ac28),
	.w7(32'h3bb8cf6d),
	.w8(32'h3bb6160f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8861bd1),
	.w1(32'h3aa69a2d),
	.w2(32'h3a93eb28),
	.w3(32'h3a392d65),
	.w4(32'h3aa51708),
	.w5(32'h3ab668a9),
	.w6(32'h3a1a5b33),
	.w7(32'h39ea297c),
	.w8(32'h39da4180),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20ec05),
	.w1(32'h3a8899c8),
	.w2(32'hb9a4b315),
	.w3(32'h3a3549db),
	.w4(32'h3985a8b3),
	.w5(32'hbab90d49),
	.w6(32'h3ae99fad),
	.w7(32'h3902beb5),
	.w8(32'h3a6f4496),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985458c),
	.w1(32'h3a2ab785),
	.w2(32'h3a295ff9),
	.w3(32'hba8509a2),
	.w4(32'h3a58964c),
	.w5(32'h3a2d5ca3),
	.w6(32'h3a634e99),
	.w7(32'h3a990c2d),
	.w8(32'h39f7dc54),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929e27d),
	.w1(32'h3bc20c5d),
	.w2(32'h3c25562f),
	.w3(32'h3945df26),
	.w4(32'hbb3ab5f3),
	.w5(32'h392eacdf),
	.w6(32'h3aa58710),
	.w7(32'h3bad6895),
	.w8(32'h3b35b224),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf64555),
	.w1(32'h3acaae9c),
	.w2(32'h3a8223aa),
	.w3(32'hbb3d2eaf),
	.w4(32'h3b258bd3),
	.w5(32'h3b2d4e9e),
	.w6(32'h3a96d1bb),
	.w7(32'h39f8e7d2),
	.w8(32'h3a9c8014),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0a107),
	.w1(32'hb92dcb9a),
	.w2(32'hb9e3ff68),
	.w3(32'h3afda911),
	.w4(32'hba42aefb),
	.w5(32'hba9e29b7),
	.w6(32'hba413d24),
	.w7(32'hba98d0fd),
	.w8(32'hba6a738f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84fd098),
	.w1(32'hb96b7015),
	.w2(32'hba8c04ad),
	.w3(32'hba05e1ed),
	.w4(32'h3a0af587),
	.w5(32'hb9edfebd),
	.w6(32'hb9b0b634),
	.w7(32'hbab5376f),
	.w8(32'hba302d8a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b1f50),
	.w1(32'h3a8603d3),
	.w2(32'h3ae30fbd),
	.w3(32'h39b97677),
	.w4(32'h39f09acb),
	.w5(32'h3a966d8e),
	.w6(32'h3ac4b9d7),
	.w7(32'h3b202af8),
	.w8(32'h3a06bb80),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb721dad3),
	.w1(32'hba9ac3e4),
	.w2(32'hbacb6fe1),
	.w3(32'hba146bfc),
	.w4(32'h39cf3a9e),
	.w5(32'hb9dd0b04),
	.w6(32'hb985930a),
	.w7(32'hba5a5539),
	.w8(32'h383fc77b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a24b00),
	.w1(32'h3ac54971),
	.w2(32'h3a0f38fe),
	.w3(32'h3a136527),
	.w4(32'h3a3cf654),
	.w5(32'hb9fccce3),
	.w6(32'h39b63fa1),
	.w7(32'hba68f3a1),
	.w8(32'hba1f3778),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98108a),
	.w1(32'h3a7f6b67),
	.w2(32'h3a4a5c9e),
	.w3(32'h39a8a215),
	.w4(32'h3a93e3c1),
	.w5(32'h38f0b230),
	.w6(32'h3abedc93),
	.w7(32'h3ae0f21e),
	.w8(32'h3a9a179b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39deeed9),
	.w1(32'h3abc985b),
	.w2(32'h3930d1c9),
	.w3(32'hb99fe5a9),
	.w4(32'h39bc1eb6),
	.w5(32'hb9f14f3d),
	.w6(32'h3aec06eb),
	.w7(32'h39a5883e),
	.w8(32'h37c611c4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98432a3),
	.w1(32'hba3533cc),
	.w2(32'hbb3d06b1),
	.w3(32'hbab81af9),
	.w4(32'h3ae7b246),
	.w5(32'hba45f2d8),
	.w6(32'h3bc0f75c),
	.w7(32'h3b364296),
	.w8(32'h3ba097ef),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c6bf5),
	.w1(32'h3a50993a),
	.w2(32'h3a4c8389),
	.w3(32'h38cd45dd),
	.w4(32'hb998243e),
	.w5(32'hb9f58a6e),
	.w6(32'h379b41a4),
	.w7(32'h380abfe3),
	.w8(32'hb9d0784c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39923225),
	.w1(32'h399be619),
	.w2(32'h3abfb000),
	.w3(32'hba793212),
	.w4(32'h393b8324),
	.w5(32'hb9c337a0),
	.w6(32'h393666cb),
	.w7(32'hb9334d7b),
	.w8(32'h39e506b1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0469da),
	.w1(32'hbb135337),
	.w2(32'h3a1e59c8),
	.w3(32'h3a6b93ed),
	.w4(32'hbad9ff04),
	.w5(32'h39fd1d8d),
	.w6(32'h3a33a3d8),
	.w7(32'h3b43c6e1),
	.w8(32'h3a809916),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab38c6b),
	.w1(32'h3a2d2c99),
	.w2(32'h39a5ad35),
	.w3(32'hbb1c8c84),
	.w4(32'hb9df6af5),
	.w5(32'hb9111ba2),
	.w6(32'h3995c526),
	.w7(32'hba1891c9),
	.w8(32'hbb8e9e90),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88c673),
	.w1(32'h3a23040f),
	.w2(32'h3aab3922),
	.w3(32'hbb86633d),
	.w4(32'h39e59531),
	.w5(32'h3a6c3a02),
	.w6(32'h399ec834),
	.w7(32'h3a46ad8a),
	.w8(32'h39431fd3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936ffd4),
	.w1(32'h3a6ce8e8),
	.w2(32'hba52bc44),
	.w3(32'h391a1e5d),
	.w4(32'h3a80b846),
	.w5(32'hba1d6f40),
	.w6(32'h3ad0fafe),
	.w7(32'hb9ea0b68),
	.w8(32'h39831047),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a225fcd),
	.w1(32'hbb596576),
	.w2(32'h3b61aed4),
	.w3(32'h3970bbe2),
	.w4(32'hbb9851ba),
	.w5(32'h39ba5671),
	.w6(32'hbb27514b),
	.w7(32'h3a4f634a),
	.w8(32'hba06e025),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade5c61),
	.w1(32'hbb3d396b),
	.w2(32'h3a8b19a7),
	.w3(32'hbac1da7f),
	.w4(32'hbb146c71),
	.w5(32'hb962ca4b),
	.w6(32'hbac2ea15),
	.w7(32'hba968715),
	.w8(32'h3a1e79e9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5204c7),
	.w1(32'h3aa7e194),
	.w2(32'hba93cf40),
	.w3(32'h3ae33d64),
	.w4(32'h3a9a5c21),
	.w5(32'hbaa1d497),
	.w6(32'h3b17c412),
	.w7(32'hb99c38a3),
	.w8(32'h3b148d09),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adac4eb),
	.w1(32'hbab25fd6),
	.w2(32'hbad2bc94),
	.w3(32'h3aec144d),
	.w4(32'hba185bf2),
	.w5(32'hba15595f),
	.w6(32'hb884be55),
	.w7(32'hb9a36884),
	.w8(32'h3a283fa7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961007a),
	.w1(32'h3a3636fc),
	.w2(32'hba214b91),
	.w3(32'h3a125ad7),
	.w4(32'h3a0a792d),
	.w5(32'hba39207a),
	.w6(32'h3a7d164f),
	.w7(32'hb9bd1f6c),
	.w8(32'h3a8bb6e4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a7630),
	.w1(32'hbaa8e612),
	.w2(32'hbaabc8c1),
	.w3(32'h3a402be0),
	.w4(32'hba65cd65),
	.w5(32'hbaa606f9),
	.w6(32'hba4499b3),
	.w7(32'hba2d03f0),
	.w8(32'hba37eac0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94ee86),
	.w1(32'h3a9672af),
	.w2(32'h3a197160),
	.w3(32'hba24a138),
	.w4(32'hb7fccb08),
	.w5(32'hb9de2131),
	.w6(32'hba06e771),
	.w7(32'hb9e69b6d),
	.w8(32'hba46c43c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c73a8),
	.w1(32'h3a87175c),
	.w2(32'hb9bee953),
	.w3(32'hba8427a3),
	.w4(32'h3ab9c541),
	.w5(32'hb8fb9249),
	.w6(32'h3986135d),
	.w7(32'hbad1a5f0),
	.w8(32'hba50207c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c22dc),
	.w1(32'h3a249588),
	.w2(32'hba225ed7),
	.w3(32'h3a3738e9),
	.w4(32'h3a185362),
	.w5(32'hba2a3431),
	.w6(32'h3a81711e),
	.w7(32'hb98b26ec),
	.w8(32'h3aa05426),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa613),
	.w1(32'hb81b948e),
	.w2(32'hb9d5728f),
	.w3(32'h3a7946e5),
	.w4(32'hb8da261e),
	.w5(32'hba954c5c),
	.w6(32'hb98d20af),
	.w7(32'h3a166b73),
	.w8(32'h385ce504),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba537b06),
	.w1(32'hb9780786),
	.w2(32'hb9eb6254),
	.w3(32'hbb032a92),
	.w4(32'hb9632547),
	.w5(32'hb8de284b),
	.w6(32'h395421ca),
	.w7(32'hba2a1a14),
	.w8(32'hbaa7307c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba110d82),
	.w1(32'hba7bbbb4),
	.w2(32'hb98ea85f),
	.w3(32'hb975a863),
	.w4(32'hb90df129),
	.w5(32'h3b123500),
	.w6(32'hbb05446a),
	.w7(32'hbb1317cb),
	.w8(32'hbb02e853),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fb241),
	.w1(32'hb945d54f),
	.w2(32'hba0c2416),
	.w3(32'hbb29688d),
	.w4(32'hba036e69),
	.w5(32'hb9b177ff),
	.w6(32'hb918b206),
	.w7(32'hba24ed66),
	.w8(32'hba1bfa2d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2da7f),
	.w1(32'hba211021),
	.w2(32'hb71fb905),
	.w3(32'h390c81dd),
	.w4(32'hb9dad96a),
	.w5(32'hb9ca0d04),
	.w6(32'hbacc6b45),
	.w7(32'hba994d76),
	.w8(32'hba267256),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d9ed5),
	.w1(32'hba8a6ad5),
	.w2(32'hb9fc93c1),
	.w3(32'hb7e55eab),
	.w4(32'hba44a47f),
	.w5(32'hba6bf859),
	.w6(32'hba90678b),
	.w7(32'hbadb59d6),
	.w8(32'hbb057d75),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fa568),
	.w1(32'h3a789a56),
	.w2(32'hba6bfeb1),
	.w3(32'hbad4db1b),
	.w4(32'h3a625511),
	.w5(32'hba7576cf),
	.w6(32'h3ac16123),
	.w7(32'hb9dc10a7),
	.w8(32'h3ada975d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fad90),
	.w1(32'h3a1396af),
	.w2(32'hb94a54b2),
	.w3(32'h3aa6fab1),
	.w4(32'h390229af),
	.w5(32'hb9f4e4d8),
	.w6(32'h3a09616a),
	.w7(32'hb9ae69a9),
	.w8(32'h3a3ea0e0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a8337),
	.w1(32'h3a571bac),
	.w2(32'hb982d9ca),
	.w3(32'h3a1a456f),
	.w4(32'h394108d3),
	.w5(32'hba24205a),
	.w6(32'h3a4a1b5d),
	.w7(32'hb9f1e062),
	.w8(32'h3a85e507),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf5dc9),
	.w1(32'h3ab9c531),
	.w2(32'hba065e12),
	.w3(32'h3a5667fe),
	.w4(32'h3a4b23ca),
	.w5(32'h38cf405a),
	.w6(32'hba8cc4c6),
	.w7(32'hbb23e6a9),
	.w8(32'hbb0d4642),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39719b54),
	.w1(32'hbb3f8dc6),
	.w2(32'hb873a70f),
	.w3(32'hb999c319),
	.w4(32'hbb2673e3),
	.w5(32'hbae3fab1),
	.w6(32'hbb0dc751),
	.w7(32'hba2f4251),
	.w8(32'hbb03d4bd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa649a),
	.w1(32'hbae3aa54),
	.w2(32'hba9b3f69),
	.w3(32'hbadc5b8c),
	.w4(32'hbabf8ebb),
	.w5(32'hbaef26fe),
	.w6(32'hbaa8a0d3),
	.w7(32'hba66343f),
	.w8(32'h388904c3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4c720),
	.w1(32'hb9b6ef3c),
	.w2(32'hba726c14),
	.w3(32'hba33df88),
	.w4(32'hb9e0bc5d),
	.w5(32'hbac95317),
	.w6(32'hb9a929dc),
	.w7(32'hbabc5e56),
	.w8(32'hba82be8a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba189447),
	.w1(32'h38d07c2b),
	.w2(32'hb989eea5),
	.w3(32'hba3deed3),
	.w4(32'h398013c9),
	.w5(32'h37bda877),
	.w6(32'h391097c0),
	.w7(32'hb9fd5b6c),
	.w8(32'h396b6bf0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04dadc),
	.w1(32'hba66cf35),
	.w2(32'hbb0385e8),
	.w3(32'h3a679118),
	.w4(32'h39fdd3dd),
	.w5(32'hba277a95),
	.w6(32'hba845184),
	.w7(32'hba915f17),
	.w8(32'hbaea54d1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3989d3),
	.w1(32'h3a0c844a),
	.w2(32'h38c5ef5e),
	.w3(32'hb94a4f92),
	.w4(32'hb97602c7),
	.w5(32'hba879d28),
	.w6(32'h3a9d76d7),
	.w7(32'hb907596c),
	.w8(32'h3a4348b1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3b819),
	.w1(32'hb9c23c09),
	.w2(32'hbab5db67),
	.w3(32'hb922cbfa),
	.w4(32'h3a37495d),
	.w5(32'hba72224f),
	.w6(32'hba71f10e),
	.w7(32'hbb189a19),
	.w8(32'hba72e7df),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965b9e3),
	.w1(32'hbb39eac4),
	.w2(32'hba8a8d85),
	.w3(32'h3a3b745c),
	.w4(32'hbb72bf64),
	.w5(32'hbb1075f4),
	.w6(32'hbb51ca13),
	.w7(32'hbb000162),
	.w8(32'hba8e7f3e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec7549),
	.w1(32'h3b64535e),
	.w2(32'h3b882250),
	.w3(32'hbb3320a1),
	.w4(32'h3b0f251c),
	.w5(32'h3b50c937),
	.w6(32'h3b19b3c3),
	.w7(32'h3b5a7bec),
	.w8(32'h3b4798c5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule