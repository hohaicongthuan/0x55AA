module layer_10_featuremap_172(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd4324),
	.w1(32'h3817891e),
	.w2(32'hb8f4f9f5),
	.w3(32'h38c3686d),
	.w4(32'h39266f4e),
	.w5(32'h38133d98),
	.w6(32'hb8025014),
	.w7(32'hb927bdac),
	.w8(32'hb88a612a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a71e),
	.w1(32'hba134a4b),
	.w2(32'hbb15a625),
	.w3(32'hbbbb224d),
	.w4(32'h3b2f8889),
	.w5(32'h3a62a049),
	.w6(32'hbbd7d6b4),
	.w7(32'h3b1997ee),
	.w8(32'hb9ddca80),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393924b0),
	.w1(32'h38ca01a8),
	.w2(32'h38b7d008),
	.w3(32'h3919e7c0),
	.w4(32'h38474c2a),
	.w5(32'h3896877a),
	.w6(32'h386ecbdb),
	.w7(32'h381d411a),
	.w8(32'h385cd661),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80e616),
	.w1(32'h3a307ec0),
	.w2(32'h3a987d6a),
	.w3(32'h3931fce5),
	.w4(32'hba42b36e),
	.w5(32'h35fe4248),
	.w6(32'hb935e09c),
	.w7(32'h392d5cf5),
	.w8(32'h3891c07e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ece7fb),
	.w1(32'h385a3381),
	.w2(32'h390400bc),
	.w3(32'hb8ea6a6f),
	.w4(32'hb8854afc),
	.w5(32'h3861645d),
	.w6(32'h39409195),
	.w7(32'h37e0aea7),
	.w8(32'h390d4fdd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881826d),
	.w1(32'h387d9a29),
	.w2(32'h388f37bf),
	.w3(32'hb8858303),
	.w4(32'h38b68ec8),
	.w5(32'h38962044),
	.w6(32'h39652e22),
	.w7(32'h38cfe654),
	.w8(32'h394ce26a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e3c6),
	.w1(32'hbbb736f2),
	.w2(32'hbc26dfd9),
	.w3(32'hba1d43de),
	.w4(32'hbbcef42e),
	.w5(32'hbc2c8f94),
	.w6(32'h3b1ab170),
	.w7(32'hbba7b402),
	.w8(32'hbc13b7d7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc147e),
	.w1(32'hbc10081f),
	.w2(32'hbb228aba),
	.w3(32'hbc585c6b),
	.w4(32'hbc0fd0d1),
	.w5(32'hbbafb4b7),
	.w6(32'hbc2473ee),
	.w7(32'hbbee3626),
	.w8(32'hbbc1e41f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1808da),
	.w1(32'h3accfd4f),
	.w2(32'h3a8081ac),
	.w3(32'h3a82252e),
	.w4(32'h3a9729d9),
	.w5(32'h38410845),
	.w6(32'h3a742c78),
	.w7(32'h3a53b3a7),
	.w8(32'hb851a820),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af2ff),
	.w1(32'hb9f8fd0f),
	.w2(32'hbc37ec17),
	.w3(32'hbb811f9e),
	.w4(32'h3becdc22),
	.w5(32'hbb690a9b),
	.w6(32'hbc0fcb20),
	.w7(32'h3b979f95),
	.w8(32'hbbbf91d2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945e302),
	.w1(32'hb9423815),
	.w2(32'hb8a50a13),
	.w3(32'h39295640),
	.w4(32'hb7efbd51),
	.w5(32'hb85c252f),
	.w6(32'hb987fd60),
	.w7(32'hb912b0ea),
	.w8(32'hb980bb5c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c07f2),
	.w1(32'h3ad75099),
	.w2(32'hbbe46617),
	.w3(32'hbb47b6e0),
	.w4(32'hbb45f192),
	.w5(32'hbc23940d),
	.w6(32'h39bec2f7),
	.w7(32'hb8a73f25),
	.w8(32'hbc50ae62),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aabaa),
	.w1(32'hb9f8b2a5),
	.w2(32'hbc4d4687),
	.w3(32'hb9772f4b),
	.w4(32'h3bafd028),
	.w5(32'hbbc33c55),
	.w6(32'hbb60d111),
	.w7(32'h3b45a0f5),
	.w8(32'hbbeab6d3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e33ff),
	.w1(32'hbb73101d),
	.w2(32'hbb501d5c),
	.w3(32'hbb30e88e),
	.w4(32'hba9b1228),
	.w5(32'hbb00b008),
	.w6(32'hbb56bf03),
	.w7(32'hbab42c6f),
	.w8(32'hbb0ae900),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba24c53),
	.w1(32'h3ae2db11),
	.w2(32'hbb8a0852),
	.w3(32'hba82883c),
	.w4(32'h3bf68474),
	.w5(32'h3b07296d),
	.w6(32'hbba6e86b),
	.w7(32'h3b87d4db),
	.w8(32'hb9f29566),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2527b1),
	.w1(32'hbb21bbe5),
	.w2(32'hbc254cdc),
	.w3(32'hbb48b4ab),
	.w4(32'h3b986829),
	.w5(32'hba509f70),
	.w6(32'hbbee71dd),
	.w7(32'hba0a84c9),
	.w8(32'hbbe86721),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e4f2c),
	.w1(32'h391818a6),
	.w2(32'h3995d6e3),
	.w3(32'h39040e35),
	.w4(32'h39287425),
	.w5(32'h396daa22),
	.w6(32'h39bfea33),
	.w7(32'h39936b52),
	.w8(32'h39a049b4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176ff1),
	.w1(32'hbbae6f21),
	.w2(32'hbc32205b),
	.w3(32'hbbc74a66),
	.w4(32'h3a11ff3d),
	.w5(32'hbc2a715a),
	.w6(32'hbc32c2e9),
	.w7(32'hbb948c45),
	.w8(32'hbc486493),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6911),
	.w1(32'hbb4d1e45),
	.w2(32'hbbe8fa7b),
	.w3(32'hbae90de7),
	.w4(32'h3951550a),
	.w5(32'hbb9f397f),
	.w6(32'hbb9b93d1),
	.w7(32'hbb08d33d),
	.w8(32'hbbcb0b13),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b98b9),
	.w1(32'h3995d9ee),
	.w2(32'h38d0dfc8),
	.w3(32'h39505ccc),
	.w4(32'h39b0d140),
	.w5(32'h39430ffd),
	.w6(32'h393198cd),
	.w7(32'h398a6b17),
	.w8(32'h38f23bf9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974b981),
	.w1(32'h38fba071),
	.w2(32'hb6a442b4),
	.w3(32'h397e798e),
	.w4(32'h3864c64b),
	.w5(32'h3865aa2a),
	.w6(32'h39aa3ea8),
	.w7(32'h38394cf3),
	.w8(32'h398c6f62),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c817b4),
	.w1(32'h3b458190),
	.w2(32'hba9065b2),
	.w3(32'h3aa5b774),
	.w4(32'h3b8646a6),
	.w5(32'h3a14ffca),
	.w6(32'h3757b4ab),
	.w7(32'h3b4b50c7),
	.w8(32'hba495e28),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd024e76),
	.w1(32'hbc175a33),
	.w2(32'hbc810dbc),
	.w3(32'hbcb0447c),
	.w4(32'hb90610b0),
	.w5(32'hbc317579),
	.w6(32'hbcc4a864),
	.w7(32'hbbc6952b),
	.w8(32'hbcdcc913),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc225a76),
	.w1(32'h3ad95c0a),
	.w2(32'hbc197d5c),
	.w3(32'hbb54afc6),
	.w4(32'h3c24b69e),
	.w5(32'hbaa133df),
	.w6(32'hbc194456),
	.w7(32'h3bb61c76),
	.w8(32'hbbbfc87b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc876ef5),
	.w1(32'h3ba536b1),
	.w2(32'hbb9cea15),
	.w3(32'hbc1fccc4),
	.w4(32'h3c30ce8e),
	.w5(32'h3b6f6a67),
	.w6(32'hbc835fab),
	.w7(32'h3bf28399),
	.w8(32'hbae777d1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93906d3),
	.w1(32'hba22035a),
	.w2(32'hb95bc9c8),
	.w3(32'hb8b32926),
	.w4(32'hb9ce2276),
	.w5(32'hb9e1e7cd),
	.w6(32'hb8de695c),
	.w7(32'hb9c8cdad),
	.w8(32'hb9d3081b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af9c48),
	.w1(32'h3929fa73),
	.w2(32'h399585f6),
	.w3(32'h39cfe133),
	.w4(32'h382be318),
	.w5(32'h393ba356),
	.w6(32'h39bf17fe),
	.w7(32'h3920c42c),
	.w8(32'h39ade5aa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6058b9),
	.w1(32'h3b9db06f),
	.w2(32'h39e7ccd1),
	.w3(32'hb9a17a39),
	.w4(32'h3bc9bd6a),
	.w5(32'h3c05cea5),
	.w6(32'hba9544d2),
	.w7(32'h3b030f2b),
	.w8(32'h3b17b4ac),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061e4b),
	.w1(32'h39ad012b),
	.w2(32'hbac085fa),
	.w3(32'hbb1b987a),
	.w4(32'hb92e92c5),
	.w5(32'hbaea2aad),
	.w6(32'hbb4fb946),
	.w7(32'hba58ca78),
	.w8(32'hbaed5433),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bf9a9),
	.w1(32'h3bfe691a),
	.w2(32'hba0145e2),
	.w3(32'hbb03138f),
	.w4(32'h3c043e43),
	.w5(32'h3b70a360),
	.w6(32'hbbe6e9f2),
	.w7(32'h3bb13241),
	.w8(32'h3992c4bd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1b14e),
	.w1(32'h3823847b),
	.w2(32'hb7d55876),
	.w3(32'h38d31dd1),
	.w4(32'h37a057ed),
	.w5(32'hb7fc184e),
	.w6(32'h38bfeb7f),
	.w7(32'hb6ad3ea1),
	.w8(32'h37838371),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d5c9e8),
	.w1(32'hb805b17e),
	.w2(32'hb7caab0d),
	.w3(32'h38c637c5),
	.w4(32'hb7fe5da5),
	.w5(32'hb7c7bb0a),
	.w6(32'h38a2ac12),
	.w7(32'hb81d2494),
	.w8(32'h38186cdb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3616ed),
	.w1(32'hb79a36aa),
	.w2(32'hbba881ea),
	.w3(32'hba0dc5b9),
	.w4(32'h3b68616b),
	.w5(32'hbb11b405),
	.w6(32'hbb7df2d7),
	.w7(32'h3a158512),
	.w8(32'hbb8e61f6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d693b),
	.w1(32'h3a84a033),
	.w2(32'hbad70c09),
	.w3(32'hbb4c21df),
	.w4(32'h3b248189),
	.w5(32'h391a2afd),
	.w6(32'hbb82f9d9),
	.w7(32'h3ab321ef),
	.w8(32'hba6acc28),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e5d84),
	.w1(32'h39210f4e),
	.w2(32'h37411500),
	.w3(32'h39a4e9ff),
	.w4(32'h39d1c1f4),
	.w5(32'hb92acbf3),
	.w6(32'h3965bac6),
	.w7(32'hb9b20e92),
	.w8(32'hba0bed04),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a225509),
	.w1(32'hbb2754ed),
	.w2(32'hbbb4f171),
	.w3(32'h3951e7fa),
	.w4(32'hbb146d18),
	.w5(32'hbb94dfc0),
	.w6(32'h3a8f5b7b),
	.w7(32'hbb1c3611),
	.w8(32'hbb89a766),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9180d6),
	.w1(32'h3b9ba753),
	.w2(32'hbc4044aa),
	.w3(32'hbb81e084),
	.w4(32'h3bbdec1f),
	.w5(32'hbab34bef),
	.w6(32'hba86fd23),
	.w7(32'h3bfbb511),
	.w8(32'hbbab0431),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca65a70),
	.w1(32'h3c300828),
	.w2(32'h3ad0909c),
	.w3(32'hbc8d511e),
	.w4(32'h3c5bccde),
	.w5(32'h3c111bc8),
	.w6(32'hbcd041eb),
	.w7(32'h3befd072),
	.w8(32'hbac892fb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dce4e),
	.w1(32'h3c26a9c5),
	.w2(32'h3a5221fd),
	.w3(32'hbc4f6420),
	.w4(32'h3c271825),
	.w5(32'h3b2c3e79),
	.w6(32'hbca944cf),
	.w7(32'h3b050424),
	.w8(32'hbc02d22e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ecfaf),
	.w1(32'h3b05d471),
	.w2(32'h3b08772d),
	.w3(32'hbb03af2c),
	.w4(32'h3b6eab07),
	.w5(32'h3b6ce3cb),
	.w6(32'hbb835f18),
	.w7(32'h3af63b58),
	.w8(32'h3a0d278e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be0d69),
	.w1(32'h38bd6de6),
	.w2(32'h392e68f7),
	.w3(32'h399a278b),
	.w4(32'h38d1ea62),
	.w5(32'h3922488f),
	.w6(32'h39ddf968),
	.w7(32'h38b885f6),
	.w8(32'h39b5b509),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5fe64),
	.w1(32'h38e86757),
	.w2(32'h39bb4e2f),
	.w3(32'h39aac4b6),
	.w4(32'hb8cfedc2),
	.w5(32'h3940799b),
	.w6(32'h39e9ba8e),
	.w7(32'h3986e17e),
	.w8(32'h3a0f5084),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9c61),
	.w1(32'h3a72306b),
	.w2(32'hbae50e0d),
	.w3(32'hbbcca0ec),
	.w4(32'hba954e74),
	.w5(32'hbb3f087d),
	.w6(32'hbba65804),
	.w7(32'hba0d328f),
	.w8(32'hbb4a4736),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48e036),
	.w1(32'hbb39d2dd),
	.w2(32'hbc24f78c),
	.w3(32'hbc0c9a7d),
	.w4(32'h3b0c923c),
	.w5(32'hbb9fceb3),
	.w6(32'hbc5b14a9),
	.w7(32'hbb8fffc9),
	.w8(32'hbc507641),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28234a),
	.w1(32'h3b48c4bf),
	.w2(32'hbc069916),
	.w3(32'hbb60f915),
	.w4(32'h3c2ac464),
	.w5(32'hba260705),
	.w6(32'hbc29ca3d),
	.w7(32'h3bc15957),
	.w8(32'hbba27bd8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc625e31),
	.w1(32'h3ac80aef),
	.w2(32'hbc22a04e),
	.w3(32'hbb8d5c04),
	.w4(32'h3c36c929),
	.w5(32'hba4eb0a5),
	.w6(32'hbc45ee0d),
	.w7(32'h3bd1fdd7),
	.w8(32'hbbc11085),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f9b0a),
	.w1(32'hba1ec09f),
	.w2(32'hbbcaef88),
	.w3(32'hbc1e5ab0),
	.w4(32'h3b69065b),
	.w5(32'hba71e7ce),
	.w6(32'hbc503d94),
	.w7(32'h3a7c3d33),
	.w8(32'hbbd44ea2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82f0c8),
	.w1(32'hbbda0485),
	.w2(32'hbc3b3a59),
	.w3(32'hbbb2647b),
	.w4(32'hbb87d6fd),
	.w5(32'hbc0efeb3),
	.w6(32'hbbbc2160),
	.w7(32'hbba84221),
	.w8(32'hbc4787a1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e925a6),
	.w1(32'hb785d96c),
	.w2(32'h3841a6a8),
	.w3(32'h388829b4),
	.w4(32'hb6d5f0eb),
	.w5(32'h37ce75f7),
	.w6(32'h39072612),
	.w7(32'hb7c70c14),
	.w8(32'h380dbb91),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f46d5),
	.w1(32'h3a04ab5d),
	.w2(32'h3a10bd15),
	.w3(32'h39d1bc19),
	.w4(32'h39f896b0),
	.w5(32'h39d63ad2),
	.w6(32'h39983d66),
	.w7(32'h399bd10c),
	.w8(32'h39187a7c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38334a94),
	.w1(32'h395d0e50),
	.w2(32'h39b95957),
	.w3(32'h381e8b77),
	.w4(32'h396db257),
	.w5(32'h39a625f5),
	.w6(32'h39ce8594),
	.w7(32'h397b01ea),
	.w8(32'h39d98b16),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f981),
	.w1(32'hba79edfa),
	.w2(32'hbbc095ed),
	.w3(32'hbb813dc7),
	.w4(32'h3b96c559),
	.w5(32'hbac945b3),
	.w6(32'hbb9f472e),
	.w7(32'h3b589392),
	.w8(32'hbaccdc4a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15252c),
	.w1(32'hba05458b),
	.w2(32'hbb162814),
	.w3(32'hbaaf9b52),
	.w4(32'h3a0ffef0),
	.w5(32'hbaf1e618),
	.w6(32'hbadadff4),
	.w7(32'h37cdb0e8),
	.w8(32'hbb23e89a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000244),
	.w1(32'hbbe24dec),
	.w2(32'hbc6eefe0),
	.w3(32'hbb5578e2),
	.w4(32'h39545b4a),
	.w5(32'hbbfde08a),
	.w6(32'hbc0570ee),
	.w7(32'hbb274b40),
	.w8(32'hbc2555b5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32706b),
	.w1(32'h391d37c4),
	.w2(32'hb9e79e0f),
	.w3(32'hbb162092),
	.w4(32'hba282d62),
	.w5(32'hbaf913f3),
	.w6(32'hbb0e0bae),
	.w7(32'hba8b8f06),
	.w8(32'hbb39e2c1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d1bcd3),
	.w1(32'hb891a1a5),
	.w2(32'hb8987e0f),
	.w3(32'h3948faca),
	.w4(32'h39538e28),
	.w5(32'h39bf5b90),
	.w6(32'hb9130faa),
	.w7(32'h3880b6a4),
	.w8(32'h399df291),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914e044),
	.w1(32'h394d2c59),
	.w2(32'h39059e4e),
	.w3(32'h39619c55),
	.w4(32'h3931f588),
	.w5(32'h388a94b7),
	.w6(32'h3973f257),
	.w7(32'h3965a606),
	.w8(32'h3966b714),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aeb998),
	.w1(32'h3994b411),
	.w2(32'h370570ea),
	.w3(32'hb816338e),
	.w4(32'hb77cd622),
	.w5(32'h373b9dd1),
	.w6(32'hba022940),
	.w7(32'hb937385f),
	.w8(32'hb81d709a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9295d62),
	.w1(32'h3ad6b64b),
	.w2(32'hb9154a26),
	.w3(32'hb92fbf3b),
	.w4(32'h3ac9a81f),
	.w5(32'h39ae96ce),
	.w6(32'hba9167f2),
	.w7(32'h39acf5f0),
	.w8(32'hba01948c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9957bf6),
	.w1(32'hb91fe84b),
	.w2(32'hb8cff5dd),
	.w3(32'h39dc31f3),
	.w4(32'hb8fdbaaf),
	.w5(32'hb95c08de),
	.w6(32'hb9cd9b44),
	.w7(32'hba6a2c78),
	.w8(32'hba2fa8a7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86157b),
	.w1(32'hbac95723),
	.w2(32'hbb9fec47),
	.w3(32'hbafa6d43),
	.w4(32'h3a045f47),
	.w5(32'hbb508849),
	.w6(32'hbaef3e34),
	.w7(32'hb921078f),
	.w8(32'hbba54f30),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02dfcf),
	.w1(32'hbb0fceb8),
	.w2(32'hbb36092b),
	.w3(32'hbba97efb),
	.w4(32'hbb1b84e6),
	.w5(32'hbb08b25f),
	.w6(32'hbb9fce01),
	.w7(32'hbb5d4aa0),
	.w8(32'hbbab0098),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fb862f),
	.w1(32'h37d94538),
	.w2(32'h3799bf82),
	.w3(32'hb77d8dd1),
	.w4(32'hb6d68bd8),
	.w5(32'hb86916be),
	.w6(32'h36c0fc92),
	.w7(32'hb948b859),
	.w8(32'h395e436c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b50fc7),
	.w1(32'h399db84c),
	.w2(32'h39a98dfb),
	.w3(32'hb7819e66),
	.w4(32'h398efeac),
	.w5(32'h399a09cf),
	.w6(32'h39fadb73),
	.w7(32'h39ba8747),
	.w8(32'h39ed91fe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a10774),
	.w1(32'h387bec5e),
	.w2(32'h37c5360b),
	.w3(32'h39c8f851),
	.w4(32'h38bf8daf),
	.w5(32'h3829a2f5),
	.w6(32'h3944b4aa),
	.w7(32'h38831fdb),
	.w8(32'h392e357d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f0862),
	.w1(32'hb909b72f),
	.w2(32'hb5d02352),
	.w3(32'h398f8eaa),
	.w4(32'hb8fdba2a),
	.w5(32'hb90fc856),
	.w6(32'h39687125),
	.w7(32'hb8ce632b),
	.w8(32'h39833cd9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09febf),
	.w1(32'hbc00e69f),
	.w2(32'hbc231bce),
	.w3(32'hbb9deffd),
	.w4(32'hbb8056c3),
	.w5(32'hbad5c4cf),
	.w6(32'hbc1ce772),
	.w7(32'hbbe7227d),
	.w8(32'hbc03f8bd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b8f12),
	.w1(32'hbabf2261),
	.w2(32'hbc4f19e9),
	.w3(32'hbba5fecc),
	.w4(32'h3b9457ea),
	.w5(32'hbc18e606),
	.w6(32'hbc265474),
	.w7(32'hb934b983),
	.w8(32'hbc705abb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c8f5b),
	.w1(32'h3acb8554),
	.w2(32'hbbfa04b9),
	.w3(32'hbc134976),
	.w4(32'h3ba6d39e),
	.w5(32'hbbd36048),
	.w6(32'hbc3d5329),
	.w7(32'hbb0d76ac),
	.w8(32'hbc561856),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71e8e5),
	.w1(32'h3c7d0140),
	.w2(32'hbbb0e3a0),
	.w3(32'hbbb616a5),
	.w4(32'h3cc92d61),
	.w5(32'h3c0533f5),
	.w6(32'hbca42b5f),
	.w7(32'h3c80c942),
	.w8(32'hbb1b9ab5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395dca62),
	.w1(32'h3937c3d3),
	.w2(32'h398cffba),
	.w3(32'h39818b53),
	.w4(32'h3906ab44),
	.w5(32'h3953d253),
	.w6(32'h39f27ad0),
	.w7(32'h397f6569),
	.w8(32'h39da5881),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13bbcd),
	.w1(32'h3758aa78),
	.w2(32'h394cbb42),
	.w3(32'h39fbae78),
	.w4(32'hb819644e),
	.w5(32'h3946e69f),
	.w6(32'h39e30e8d),
	.w7(32'h39015de8),
	.w8(32'h39db6ede),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b89d0b),
	.w1(32'hb76c2f71),
	.w2(32'h3925f1b4),
	.w3(32'h39b42ef1),
	.w4(32'hb8b31541),
	.w5(32'h39182046),
	.w6(32'h39fb8a96),
	.w7(32'h3873c5c2),
	.w8(32'h39aedfcd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9955395),
	.w1(32'hb9158d2c),
	.w2(32'hba8dd803),
	.w3(32'hb99d9e9f),
	.w4(32'h3950c250),
	.w5(32'hbabe1413),
	.w6(32'hba6cda9e),
	.w7(32'hb9e13106),
	.w8(32'hbadc7f89),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a37f9),
	.w1(32'h380eeef8),
	.w2(32'h39175f81),
	.w3(32'h3937f267),
	.w4(32'hb8816555),
	.w5(32'h385b615b),
	.w6(32'h39a3c08e),
	.w7(32'h38789e30),
	.w8(32'h3986e50b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3350ac),
	.w1(32'hbbb03789),
	.w2(32'hbb7bf287),
	.w3(32'hbb8a76df),
	.w4(32'hbbae56ac),
	.w5(32'hbb70d7a3),
	.w6(32'hbb41bcb3),
	.w7(32'hbb434198),
	.w8(32'hbb78716c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcddab6),
	.w1(32'hbb08d8c4),
	.w2(32'hbc001cfa),
	.w3(32'hbb9c10c3),
	.w4(32'h3a73a19a),
	.w5(32'hbb3ba5b9),
	.w6(32'hbbf8700e),
	.w7(32'hbb8478d8),
	.w8(32'hbbf2c2c5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19734e),
	.w1(32'h39e0efcc),
	.w2(32'hbbc4a243),
	.w3(32'hbb8527c0),
	.w4(32'h3c06f672),
	.w5(32'h3b41eac8),
	.w6(32'hbbcd1fa4),
	.w7(32'h3bf10c50),
	.w8(32'h3b1ecfdf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895fc5),
	.w1(32'hb9f72022),
	.w2(32'hbb92790e),
	.w3(32'hbb26f49b),
	.w4(32'h3b18290e),
	.w5(32'hbaca82a8),
	.w6(32'hbba9128f),
	.w7(32'hb8e2ab9f),
	.w8(32'hbb7f2670),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab16684),
	.w1(32'hb9cde17e),
	.w2(32'hbb9e44fa),
	.w3(32'h398967cf),
	.w4(32'h3aeab9d0),
	.w5(32'hb9d0fdc2),
	.w6(32'hba967997),
	.w7(32'h3aece1a8),
	.w8(32'hba8ab13f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8092b3),
	.w1(32'h37408b58),
	.w2(32'hbb82ebff),
	.w3(32'hbac845f4),
	.w4(32'h3b1bec4b),
	.w5(32'hba83e0bb),
	.w6(32'hbb5b2942),
	.w7(32'h3a894f26),
	.w8(32'hbb199df8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ce09f),
	.w1(32'hbb3e7fee),
	.w2(32'hbbc9716f),
	.w3(32'hbb2199ec),
	.w4(32'hbb06f537),
	.w5(32'hbba0575c),
	.w6(32'hbb343dfc),
	.w7(32'hba9bb00a),
	.w8(32'hbb91f6fb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3867e353),
	.w1(32'h388e269c),
	.w2(32'h381ca763),
	.w3(32'h38119728),
	.w4(32'h3857b564),
	.w5(32'h36175da6),
	.w6(32'h390c8559),
	.w7(32'h384adfe0),
	.w8(32'h39021ffb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa7cf8),
	.w1(32'h38d4a545),
	.w2(32'h38e31bfc),
	.w3(32'h39043e1f),
	.w4(32'h38c50a88),
	.w5(32'h39062c41),
	.w6(32'h39058892),
	.w7(32'h38d2ff8b),
	.w8(32'h39020896),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906fff0),
	.w1(32'h39626273),
	.w2(32'h39a2e68f),
	.w3(32'hb866ecb7),
	.w4(32'h38e15bb3),
	.w5(32'h3901a2e8),
	.w6(32'h36f5ca3b),
	.w7(32'h382179c1),
	.w8(32'hb7dfe412),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a989e),
	.w1(32'h3a1c0539),
	.w2(32'h3a3ba685),
	.w3(32'hb8b85aed),
	.w4(32'h3a10cd53),
	.w5(32'h3a4aa5b4),
	.w6(32'hba0916cc),
	.w7(32'h39db8b8e),
	.w8(32'h39da61ae),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d1a41),
	.w1(32'h3b2f93b1),
	.w2(32'h3a23a9b5),
	.w3(32'hbc292662),
	.w4(32'h3b6f5f0c),
	.w5(32'h3b4db7e2),
	.w6(32'hbc47d2d3),
	.w7(32'h3b79eeca),
	.w8(32'h3a0017f8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8539e),
	.w1(32'h3ad68e7b),
	.w2(32'hb81d3c52),
	.w3(32'h3aae64a3),
	.w4(32'h3b33451e),
	.w5(32'h3a25295c),
	.w6(32'hba69576c),
	.w7(32'h3a2c60cb),
	.w8(32'hb9fb568e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4c581),
	.w1(32'hbaabbb37),
	.w2(32'hbba9dd89),
	.w3(32'hbb036151),
	.w4(32'h3b334c3a),
	.w5(32'hbaa91be5),
	.w6(32'hbbc88dfe),
	.w7(32'h3ac2dc73),
	.w8(32'hbb3cca2d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc530537),
	.w1(32'hbbbd2690),
	.w2(32'hbbad16c1),
	.w3(32'hbc65e54e),
	.w4(32'hbb3c741e),
	.w5(32'hbbaf89ad),
	.w6(32'hbc97caf3),
	.w7(32'hbc0814ea),
	.w8(32'hbc31058d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963c9c),
	.w1(32'h3b8dc7ab),
	.w2(32'hba550d80),
	.w3(32'hbba9ca44),
	.w4(32'h3b478317),
	.w5(32'h3a870e61),
	.w6(32'hbbe1afc9),
	.w7(32'h3b02ec4e),
	.w8(32'hbb0a84de),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f7c6b),
	.w1(32'hbb2ebc65),
	.w2(32'hbbd0b672),
	.w3(32'hbbf7313e),
	.w4(32'h39015904),
	.w5(32'hbb0a456f),
	.w6(32'hbb9b3396),
	.w7(32'hba7a68d8),
	.w8(32'hbc0cf8aa),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2cbb),
	.w1(32'h3be267d8),
	.w2(32'h3b207eed),
	.w3(32'hb9c6b4bd),
	.w4(32'h3c04edf1),
	.w5(32'h3b8c681c),
	.w6(32'hbb3481ed),
	.w7(32'h3be06684),
	.w8(32'h3b58b4dc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e170e),
	.w1(32'hba777131),
	.w2(32'hbbd964c1),
	.w3(32'hbbd55a82),
	.w4(32'h3b91e16d),
	.w5(32'h39586566),
	.w6(32'hbc5e8aaa),
	.w7(32'hbb220322),
	.w8(32'hbbf46592),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01b784),
	.w1(32'h385eea09),
	.w2(32'hbb6136bb),
	.w3(32'hbbb56f46),
	.w4(32'h3b21bbe7),
	.w5(32'h3aaf5d66),
	.w6(32'hbbb2026a),
	.w7(32'h3b62644f),
	.w8(32'hbaa6a07e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb3b2),
	.w1(32'h3b93c8a1),
	.w2(32'hba08d3cc),
	.w3(32'hbbb43cba),
	.w4(32'h3c1e4ea8),
	.w5(32'h3b8a4b88),
	.w6(32'hbc2425ea),
	.w7(32'h3bd7dbde),
	.w8(32'h3abe254c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce18c3),
	.w1(32'h398d5808),
	.w2(32'h39b01bca),
	.w3(32'h39ae8ca8),
	.w4(32'h3820db37),
	.w5(32'h3958dc7e),
	.w6(32'h3988a388),
	.w7(32'hb84ad853),
	.w8(32'h3930dc9d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19a5d7),
	.w1(32'hba93ac4c),
	.w2(32'hbc261de0),
	.w3(32'hbb9da403),
	.w4(32'h3bdcc994),
	.w5(32'hbb7e049a),
	.w6(32'hbc372c41),
	.w7(32'hba866a54),
	.w8(32'hbc2529de),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0251),
	.w1(32'hbaf3636b),
	.w2(32'hbbd6109a),
	.w3(32'hbb61a247),
	.w4(32'h3a0d7faa),
	.w5(32'hbb640d4e),
	.w6(32'hbb79163d),
	.w7(32'hb682d5d0),
	.w8(32'hbbed7fc1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6869e8),
	.w1(32'hbb99ad42),
	.w2(32'hbc8b0a91),
	.w3(32'hbb9ea0d6),
	.w4(32'h3b61c69c),
	.w5(32'hbba997e7),
	.w6(32'hb94d709f),
	.w7(32'h3b4da508),
	.w8(32'hbc44b1b4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7fac3),
	.w1(32'h3bcb77b7),
	.w2(32'h3b8a330a),
	.w3(32'hbca47562),
	.w4(32'h3c0252da),
	.w5(32'h3bfed4ab),
	.w6(32'hbcbc1dbf),
	.w7(32'h3b006741),
	.w8(32'hbafac6b6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe984d5),
	.w1(32'h3bae0c92),
	.w2(32'hbbbc90e0),
	.w3(32'hbad34e1a),
	.w4(32'h3c49011d),
	.w5(32'h3af02a27),
	.w6(32'hbc0a7e79),
	.w7(32'h3c0aba88),
	.w8(32'hba973f23),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebc8e4),
	.w1(32'hbb87ea5c),
	.w2(32'hbc1b7701),
	.w3(32'hbbbece4e),
	.w4(32'hbb49b2de),
	.w5(32'hbb7f46bf),
	.w6(32'hbb2721af),
	.w7(32'h398d8da5),
	.w8(32'hbc036dc4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b665ce),
	.w1(32'hb867c109),
	.w2(32'h38f6625c),
	.w3(32'h390022f2),
	.w4(32'hb90aa174),
	.w5(32'h3811a045),
	.w6(32'h399f97aa),
	.w7(32'hb64c235f),
	.w8(32'h398557ed),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc824275),
	.w1(32'hbc5be621),
	.w2(32'hbc8b37ff),
	.w3(32'hbbed72c0),
	.w4(32'hba8f160a),
	.w5(32'hbb949abe),
	.w6(32'h3951e69d),
	.w7(32'h3bfc0ce4),
	.w8(32'hb8efcc5c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a0a1a),
	.w1(32'h3b96c4d3),
	.w2(32'hbb64c1f9),
	.w3(32'hba0ee4e2),
	.w4(32'h3b0fdb13),
	.w5(32'hbb82b044),
	.w6(32'hb92b5208),
	.w7(32'h3ba5c667),
	.w8(32'hbb9ce155),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef5441),
	.w1(32'h39516718),
	.w2(32'hb869e4e1),
	.w3(32'h383bade9),
	.w4(32'h39edae11),
	.w5(32'h3984d024),
	.w6(32'h387d07d3),
	.w7(32'h39f8c1c8),
	.w8(32'h39808937),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d4f7c),
	.w1(32'hba6866d8),
	.w2(32'hbac04bcc),
	.w3(32'hbab947b2),
	.w4(32'hb9298b86),
	.w5(32'hb9bd8423),
	.w6(32'hbb45c698),
	.w7(32'hba5f3d59),
	.w8(32'hba5e486d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd412f3),
	.w1(32'hbacffec9),
	.w2(32'hbb8be4dd),
	.w3(32'hbb998995),
	.w4(32'h3aefe5c1),
	.w5(32'hbaf2ff9e),
	.w6(32'hbc02cfd1),
	.w7(32'hbb03a5ad),
	.w8(32'hbbc27315),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6266a9),
	.w1(32'h3b5595cb),
	.w2(32'hbb20b42d),
	.w3(32'hba7a40a6),
	.w4(32'h3c034eb0),
	.w5(32'h3b0e3e5f),
	.w6(32'hbb8e3ddb),
	.w7(32'h3be1ebc2),
	.w8(32'h3a6fdca9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda49b),
	.w1(32'h3a24ae99),
	.w2(32'hbaccd758),
	.w3(32'hbb5e2c8c),
	.w4(32'h3b33ffcc),
	.w5(32'h3a35c3ad),
	.w6(32'hbc14c6f2),
	.w7(32'hb95d4047),
	.w8(32'hbb3fd309),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbef1ae),
	.w1(32'h3a47a7c2),
	.w2(32'hbad9ac37),
	.w3(32'hbb29ca70),
	.w4(32'h3b8cff79),
	.w5(32'h3a87425b),
	.w6(32'hbbbbedb2),
	.w7(32'h3b28a49c),
	.w8(32'hbaa1d7de),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33b2ca),
	.w1(32'h3aee04ec),
	.w2(32'hbb5be989),
	.w3(32'hbb7e59e6),
	.w4(32'h3a058e7d),
	.w5(32'hbb52056a),
	.w6(32'hbb97cfc0),
	.w7(32'hbad040fa),
	.w8(32'hbbd06a93),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca91a9),
	.w1(32'hbb138c4d),
	.w2(32'hbbe2aa38),
	.w3(32'hba676a36),
	.w4(32'h3b5ff804),
	.w5(32'h3a43211e),
	.w6(32'hbb930926),
	.w7(32'h3abdc4c9),
	.w8(32'hbb43b9a9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eca8d),
	.w1(32'h3ac181f7),
	.w2(32'hbb0ef8a1),
	.w3(32'hbb08ce60),
	.w4(32'h3b68ebfd),
	.w5(32'hb9b9288e),
	.w6(32'hbbae9d87),
	.w7(32'h3abd9454),
	.w8(32'hbb311934),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957c4d5),
	.w1(32'hb97d949a),
	.w2(32'hb9b51dc8),
	.w3(32'hb9770160),
	.w4(32'hb8fadb3d),
	.w5(32'hb913cbc9),
	.w6(32'hb8ebc298),
	.w7(32'hb95b7d2c),
	.w8(32'hb8478a73),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bea39),
	.w1(32'hb9d86748),
	.w2(32'hb9f74876),
	.w3(32'hb7bd6f2e),
	.w4(32'h396a5df6),
	.w5(32'h382bec01),
	.w6(32'hba2b464a),
	.w7(32'hb63cbc0b),
	.w8(32'hb911b94b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3852f289),
	.w1(32'h383fdc9b),
	.w2(32'hb85db1dc),
	.w3(32'hb8ad1a5b),
	.w4(32'h37fca327),
	.w5(32'hb85a7a33),
	.w6(32'hb7428778),
	.w7(32'hb87a8eb3),
	.w8(32'hb707488b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39081279),
	.w1(32'hb8c0a454),
	.w2(32'hb8b056cb),
	.w3(32'h38e8dcfe),
	.w4(32'hb87ef05b),
	.w5(32'h3927af0b),
	.w6(32'h38f0c3c3),
	.w7(32'hb940dfb1),
	.w8(32'h3715064a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a8bd),
	.w1(32'h3b2886e0),
	.w2(32'hbb8cbcf1),
	.w3(32'hba9f831c),
	.w4(32'h3bdd9936),
	.w5(32'h3918a448),
	.w6(32'hbba6f555),
	.w7(32'h3b814bf4),
	.w8(32'hbb0f9eee),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14c2e9),
	.w1(32'hb9ea8806),
	.w2(32'hba3c1cd1),
	.w3(32'hb953880c),
	.w4(32'hb943db90),
	.w5(32'hb9d856a8),
	.w6(32'hba15a87a),
	.w7(32'hb9a308fd),
	.w8(32'hba25cfb9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7822c0a),
	.w1(32'hbaafec9d),
	.w2(32'hbb8f07da),
	.w3(32'hba9e6e83),
	.w4(32'hba928909),
	.w5(32'hbb1ba1b3),
	.w6(32'h39c5d48c),
	.w7(32'hba8acd90),
	.w8(32'hbb87273c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc600561),
	.w1(32'h3a485b24),
	.w2(32'hbb306626),
	.w3(32'hbc0c85f6),
	.w4(32'h3bb36a6e),
	.w5(32'h3a8ed42b),
	.w6(32'hbc3ebe1f),
	.w7(32'h3b3a5e61),
	.w8(32'hbab7accd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925de0f),
	.w1(32'h39004599),
	.w2(32'h38d8bfd7),
	.w3(32'h3992cd7a),
	.w4(32'h397e524b),
	.w5(32'h39783cb3),
	.w6(32'h39acea66),
	.w7(32'h398ca2ff),
	.w8(32'hb79a4a07),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396289f3),
	.w1(32'h39700484),
	.w2(32'hb8fc93e5),
	.w3(32'h3a2aaab5),
	.w4(32'h3a2e4a43),
	.w5(32'h394462fd),
	.w6(32'h3959a648),
	.w7(32'h3920094e),
	.w8(32'hb836a226),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396dfa5b),
	.w1(32'h37bdd034),
	.w2(32'hb8471902),
	.w3(32'h39528770),
	.w4(32'hb70033b7),
	.w5(32'hb855a10f),
	.w6(32'h38af6823),
	.w7(32'hb837dc40),
	.w8(32'h37dd0c45),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3a7d8),
	.w1(32'hbcb7e688),
	.w2(32'hbc311dbc),
	.w3(32'hbad64db7),
	.w4(32'hbc13feb4),
	.w5(32'hbc8b80b8),
	.w6(32'hbc6881d2),
	.w7(32'hbc6bc5e5),
	.w8(32'hbb932ebc),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908b7eb),
	.w1(32'hbcd7ffdd),
	.w2(32'h399b0f25),
	.w3(32'hbb6cae62),
	.w4(32'hbc1c7a39),
	.w5(32'hbc780478),
	.w6(32'hbb0f8b5f),
	.w7(32'hbb823dcc),
	.w8(32'hbb8b7aab),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb175fa),
	.w1(32'h3c87b202),
	.w2(32'hbcaf83f8),
	.w3(32'hbbf6b849),
	.w4(32'h3c39d6f6),
	.w5(32'hbc8fe817),
	.w6(32'hbbed7536),
	.w7(32'hbb8ad6ac),
	.w8(32'h3b59083a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c377448),
	.w1(32'h3d4016fb),
	.w2(32'hbc3fc09e),
	.w3(32'hbc87dd7c),
	.w4(32'h3c8490da),
	.w5(32'h3ba0b047),
	.w6(32'h3c250f0d),
	.w7(32'hbbffc10a),
	.w8(32'hbc9f391a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00cfeb),
	.w1(32'h3cf9f863),
	.w2(32'hbbec2886),
	.w3(32'hbbd55895),
	.w4(32'h3bfb1e2b),
	.w5(32'hb9925d13),
	.w6(32'h3ad6219a),
	.w7(32'hbc58debf),
	.w8(32'hbca15716),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e5b51),
	.w1(32'h38c60b75),
	.w2(32'h39e6a840),
	.w3(32'hbbabc487),
	.w4(32'h3bb6dd86),
	.w5(32'h3c32e194),
	.w6(32'h3c0cc064),
	.w7(32'h3b5cfa91),
	.w8(32'h3c5c584c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dc101),
	.w1(32'hbbe6ed6e),
	.w2(32'h3b9f1ffb),
	.w3(32'h3b9afced),
	.w4(32'h3a6ffd1e),
	.w5(32'hbb2b0241),
	.w6(32'h3b991cac),
	.w7(32'h3b5ea334),
	.w8(32'hba93f2f7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c7a55),
	.w1(32'hbcb1fc76),
	.w2(32'h3b80e2ab),
	.w3(32'hbc0dded8),
	.w4(32'h3b23b752),
	.w5(32'h3b6365d4),
	.w6(32'hbbc0a1c4),
	.w7(32'hba5b8956),
	.w8(32'h3bfa92a4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c996404),
	.w1(32'h3d4f60f8),
	.w2(32'hbc860209),
	.w3(32'h3ba48627),
	.w4(32'h3c8c247b),
	.w5(32'h3a3d53d4),
	.w6(32'h3bffe5cd),
	.w7(32'hbc169760),
	.w8(32'hbd0d7cce),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2cdf94),
	.w1(32'hbcf6c4e0),
	.w2(32'h3c097dc4),
	.w3(32'hbc515066),
	.w4(32'hbbab3eed),
	.w5(32'hbc136762),
	.w6(32'hbc820777),
	.w7(32'h3b304781),
	.w8(32'hb9f1d25c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba91cd),
	.w1(32'hbc4123bd),
	.w2(32'hbc3419f6),
	.w3(32'hbc894230),
	.w4(32'hba077712),
	.w5(32'hbc5564e2),
	.w6(32'hbc101bdb),
	.w7(32'hbc675ddd),
	.w8(32'hbca4d48d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1daff),
	.w1(32'h3d87dcf1),
	.w2(32'hbd0a85f1),
	.w3(32'hbcca78d4),
	.w4(32'h3c908928),
	.w5(32'hbbae83f3),
	.w6(32'h3c519320),
	.w7(32'hbc780ea2),
	.w8(32'hbce648e4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd362f04),
	.w1(32'h3b4775a1),
	.w2(32'hbb1877e2),
	.w3(32'hbbc40bcc),
	.w4(32'h3bb0c592),
	.w5(32'h39676c0a),
	.w6(32'hbb2605e0),
	.w7(32'h3b972ed7),
	.w8(32'h3b631d89),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9134a1),
	.w1(32'hbbd1a29d),
	.w2(32'hbbccff71),
	.w3(32'hbc135b36),
	.w4(32'hbb22a749),
	.w5(32'hbc07d5c3),
	.w6(32'hbc28d8cc),
	.w7(32'h3ab934eb),
	.w8(32'hbb8bf236),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e58dd),
	.w1(32'hbc0b53de),
	.w2(32'hbb6ba539),
	.w3(32'hbc483e6c),
	.w4(32'hba8335a7),
	.w5(32'hbb8b09dc),
	.w6(32'hba290ede),
	.w7(32'h3a01ace9),
	.w8(32'h3b2e6c62),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1023c6),
	.w1(32'hbc805a2a),
	.w2(32'h3cf0fac7),
	.w3(32'hbbaedf9f),
	.w4(32'h3c47212e),
	.w5(32'h3b8513ea),
	.w6(32'hbbceecb6),
	.w7(32'h3caa4881),
	.w8(32'h3c62ad14),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca142bc),
	.w1(32'h3bdd757b),
	.w2(32'h3b5abfe8),
	.w3(32'hbc1f1066),
	.w4(32'h3aebd8bf),
	.w5(32'hbc0fbcd3),
	.w6(32'hba15f319),
	.w7(32'h3c154e8a),
	.w8(32'h3c0ed0f3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaad15),
	.w1(32'hbc10fc24),
	.w2(32'h3ac0472a),
	.w3(32'hbc3dd066),
	.w4(32'hbacf5b5b),
	.w5(32'hbbb88995),
	.w6(32'hbbafad4c),
	.w7(32'hbbf507ea),
	.w8(32'hbc65afb9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49d1dc),
	.w1(32'h3b3c065b),
	.w2(32'hbad84384),
	.w3(32'hbc8b85e7),
	.w4(32'h3b80ef6d),
	.w5(32'h3b5129a7),
	.w6(32'h3b6b6010),
	.w7(32'hbaf3c707),
	.w8(32'h3a9f7322),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8949b6),
	.w1(32'h3d950a75),
	.w2(32'hbc7e6a75),
	.w3(32'h39d077ce),
	.w4(32'h3caa4550),
	.w5(32'h3ba64ec0),
	.w6(32'h3c87e03d),
	.w7(32'hbc17af0c),
	.w8(32'hbceedd02),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd508ee0),
	.w1(32'h3cb17a3b),
	.w2(32'hbc4a26a7),
	.w3(32'hbc1e426c),
	.w4(32'h3c0080ff),
	.w5(32'h3bb60b97),
	.w6(32'hbc67b3fb),
	.w7(32'hbbd2683e),
	.w8(32'hbc72530f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd31e0d),
	.w1(32'hbbbcf4ff),
	.w2(32'hbc8035a3),
	.w3(32'hbc119563),
	.w4(32'h3b87bfe0),
	.w5(32'hbc39db82),
	.w6(32'hbc0a7c35),
	.w7(32'hbbea2341),
	.w8(32'hbc6d6c8b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9f5e),
	.w1(32'hbcb64f0c),
	.w2(32'h3c20f4bc),
	.w3(32'hbc42ac35),
	.w4(32'hbc2d1773),
	.w5(32'hbb069756),
	.w6(32'hbc184fd1),
	.w7(32'hb90493bd),
	.w8(32'h3c00a3b1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0eb543),
	.w1(32'h3cd91515),
	.w2(32'hbb86ea32),
	.w3(32'hbb615bbc),
	.w4(32'h3c4481e7),
	.w5(32'hbaa6332a),
	.w6(32'hb983d9b9),
	.w7(32'h3c84eebe),
	.w8(32'hbb8a9856),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb4cbf),
	.w1(32'hbba8ed5a),
	.w2(32'hba51fca4),
	.w3(32'hbc803362),
	.w4(32'h3a8ac4bf),
	.w5(32'h3b272850),
	.w6(32'hbbba9bb5),
	.w7(32'h3b902c04),
	.w8(32'h3bbc0f72),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac98c8),
	.w1(32'hbd08c61e),
	.w2(32'hb8cc9a3b),
	.w3(32'h3ac02869),
	.w4(32'hbc14abc2),
	.w5(32'hbc6cb0c9),
	.w6(32'hbbd93e83),
	.w7(32'h3ad55bcf),
	.w8(32'hbbf2522e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7fb8e),
	.w1(32'h3c4df259),
	.w2(32'hbc0a67e1),
	.w3(32'hbc6b5c71),
	.w4(32'h3c5a043c),
	.w5(32'h3be50349),
	.w6(32'h3a22a4a8),
	.w7(32'h3bdafaa4),
	.w8(32'h3a400a9e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf987e2),
	.w1(32'hbb856611),
	.w2(32'h3b1cc40a),
	.w3(32'hba3a1f92),
	.w4(32'h3bd549b7),
	.w5(32'h3b603a0a),
	.w6(32'hbb1e1457),
	.w7(32'h39a9873a),
	.w8(32'h3a92b36e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c679d10),
	.w1(32'hbc14b2b3),
	.w2(32'hbb6c3500),
	.w3(32'hba852f09),
	.w4(32'hbb38a66f),
	.w5(32'hbc0471c6),
	.w6(32'hbb834946),
	.w7(32'hbbfbfc26),
	.w8(32'hbc1c5d37),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3757f5),
	.w1(32'h3c562d67),
	.w2(32'hbc84a93e),
	.w3(32'hbc6cfb9e),
	.w4(32'h3a642189),
	.w5(32'hbbb654ca),
	.w6(32'hba764eba),
	.w7(32'h3b14f3d5),
	.w8(32'h3b0ee3ff),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a2e0),
	.w1(32'hbb898cb1),
	.w2(32'hbc9bbe68),
	.w3(32'hbbdd8fc6),
	.w4(32'h3abcab26),
	.w5(32'hbc824442),
	.w6(32'hbc16ff32),
	.w7(32'hbc8a9791),
	.w8(32'hbbbe63a7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74fa86),
	.w1(32'h3b44465e),
	.w2(32'hbb874ca1),
	.w3(32'hbb0ca0f8),
	.w4(32'h3bcf03eb),
	.w5(32'h3abe7f61),
	.w6(32'hbc0bba7e),
	.w7(32'hbbb2f844),
	.w8(32'hba9421c8),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897aa97),
	.w1(32'hbc6fa989),
	.w2(32'hbaa4389a),
	.w3(32'h3b2fa484),
	.w4(32'hbc072538),
	.w5(32'hbbd3f28d),
	.w6(32'hbbc2fc88),
	.w7(32'hbb8ac635),
	.w8(32'hba57310f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13c0cf),
	.w1(32'hbc47e7c3),
	.w2(32'hb94fab88),
	.w3(32'hbb874569),
	.w4(32'hbb6b95b9),
	.w5(32'hbba7eb6a),
	.w6(32'hbb8f8a0d),
	.w7(32'hbad79433),
	.w8(32'hba7cec53),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd10a9),
	.w1(32'hbbc32b15),
	.w2(32'hbd022fc6),
	.w3(32'hbc1641c0),
	.w4(32'h3aa4d1ee),
	.w5(32'hbc50f5b1),
	.w6(32'hbc757abe),
	.w7(32'hbc9c8ace),
	.w8(32'hbc0984ec),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d99c),
	.w1(32'hbca43d59),
	.w2(32'hbc5d3754),
	.w3(32'hbb782031),
	.w4(32'hbb88eb81),
	.w5(32'hbc241dcc),
	.w6(32'hbc4fa9e9),
	.w7(32'hbb9b16eb),
	.w8(32'hbb8b23c3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf20d),
	.w1(32'h3d7684de),
	.w2(32'hbcb8e250),
	.w3(32'hbbc975b2),
	.w4(32'h3c9c9665),
	.w5(32'hba8c158a),
	.w6(32'h3bebcc1e),
	.w7(32'hbc2f35ac),
	.w8(32'hbcbb7d98),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1378a6),
	.w1(32'hbc224014),
	.w2(32'hbb004411),
	.w3(32'hbc052b17),
	.w4(32'hbba3b250),
	.w5(32'hbc18f9be),
	.w6(32'hbb1843f9),
	.w7(32'h3a895459),
	.w8(32'hbaad092b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dce64),
	.w1(32'h3d365af0),
	.w2(32'hbb1aa43c),
	.w3(32'hbc290399),
	.w4(32'h3c52c7a1),
	.w5(32'h3c03da3c),
	.w6(32'h3c16dca1),
	.w7(32'h3a7e1805),
	.w8(32'hbc9c5b29),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc946c0),
	.w1(32'h3d513bc2),
	.w2(32'hbbfcaf5a),
	.w3(32'h3ba14b57),
	.w4(32'h3c965bf6),
	.w5(32'h3bd14ef3),
	.w6(32'h3c5f224b),
	.w7(32'hbbd1feb7),
	.w8(32'hbca56e80),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf9d9fb),
	.w1(32'hbcb319cc),
	.w2(32'h3c1c0012),
	.w3(32'hbba5c894),
	.w4(32'hbbaa2b66),
	.w5(32'hbbd8b710),
	.w6(32'hbb684f1d),
	.w7(32'h3a24f784),
	.w8(32'hbb0c9df8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40a4d6),
	.w1(32'h3cdfdbe9),
	.w2(32'hbbad90a1),
	.w3(32'hbc96c4f2),
	.w4(32'h3b8aaf83),
	.w5(32'h3bb42056),
	.w6(32'hbba723a4),
	.w7(32'h3a3c5388),
	.w8(32'hbc78593c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18b253),
	.w1(32'hbba7e666),
	.w2(32'hbc329ef6),
	.w3(32'hbc8fb34b),
	.w4(32'hba3b146f),
	.w5(32'hbc1ac1ed),
	.w6(32'hbc9d8aa7),
	.w7(32'hbbc6aa00),
	.w8(32'hbc5b9b86),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5b0d2),
	.w1(32'h3cf3dad4),
	.w2(32'hbae6e5a5),
	.w3(32'h3bcdd327),
	.w4(32'h3bbc71c8),
	.w5(32'h3bfc054c),
	.w6(32'h3bc97a52),
	.w7(32'h3b02ffd4),
	.w8(32'hbc4fe791),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc574a2),
	.w1(32'hbc16404a),
	.w2(32'hbb054928),
	.w3(32'hba856426),
	.w4(32'h3b74ced6),
	.w5(32'hbb0be728),
	.w6(32'hbc27a84b),
	.w7(32'h3b4bc5ec),
	.w8(32'h3ab8413c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9d3bc),
	.w1(32'h3dc57396),
	.w2(32'hbcb4fa13),
	.w3(32'hbb85e5f4),
	.w4(32'h3cfb5cee),
	.w5(32'h3ba209cd),
	.w6(32'h3d047d80),
	.w7(32'hbc3f6428),
	.w8(32'hbcb42550),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a9dd6),
	.w1(32'h3d2c5b9e),
	.w2(32'hbcc7ab9e),
	.w3(32'h39e9ee79),
	.w4(32'h3cd3544c),
	.w5(32'hbc3662f3),
	.w6(32'h3bef3bb6),
	.w7(32'hbbf1c893),
	.w8(32'hbccb4542),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d26bb),
	.w1(32'h3d1dd97f),
	.w2(32'hbc9a6ad6),
	.w3(32'hbc74f3d7),
	.w4(32'h3c881020),
	.w5(32'hba8705d5),
	.w6(32'hb9cb2510),
	.w7(32'hbc08a32f),
	.w8(32'hbcc67cc3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef5985),
	.w1(32'h3bcb20f7),
	.w2(32'hbbe1e71f),
	.w3(32'hbc4504af),
	.w4(32'h3bad9dce),
	.w5(32'hbb9fda12),
	.w6(32'hbad3c852),
	.w7(32'h3bb9306d),
	.w8(32'hbc2c4946),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0f5de),
	.w1(32'h3a9cb9e2),
	.w2(32'hbc033e81),
	.w3(32'hbc41fcbd),
	.w4(32'hba0f7d15),
	.w5(32'hbb6eefd1),
	.w6(32'h3b68a550),
	.w7(32'hbbe6c500),
	.w8(32'h3a4d4b94),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01b0a6),
	.w1(32'hbc46e3b4),
	.w2(32'hbbfa085f),
	.w3(32'hbadf987a),
	.w4(32'hbac2fcb8),
	.w5(32'hbba8ec1f),
	.w6(32'hbbbcd41e),
	.w7(32'hbb4ada62),
	.w8(32'hbb926697),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dedc7a),
	.w1(32'hbcb0d668),
	.w2(32'h3c93dc73),
	.w3(32'hbbab4a2e),
	.w4(32'hbb6ea963),
	.w5(32'hbad82a7f),
	.w6(32'hb9a74393),
	.w7(32'h3bfa4ab4),
	.w8(32'h3b6147e0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3540dd),
	.w1(32'h3d4fbf51),
	.w2(32'hbc92ed10),
	.w3(32'hbbeecabf),
	.w4(32'h3ca3fcc1),
	.w5(32'hb98fc8f8),
	.w6(32'h3cb075e3),
	.w7(32'hbbf0b1b6),
	.w8(32'hbcba8262),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd08eaf5),
	.w1(32'h3c14e4b3),
	.w2(32'hbc8f1924),
	.w3(32'hbc174570),
	.w4(32'h3b961b1e),
	.w5(32'hbb03a5f3),
	.w6(32'hbbc6fc31),
	.w7(32'h39a3a533),
	.w8(32'h3af78aab),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae353a5),
	.w1(32'hbb771d92),
	.w2(32'h3b91e999),
	.w3(32'h3b82f8f9),
	.w4(32'h3c105d7c),
	.w5(32'h3bb76e3f),
	.w6(32'hbbac10a3),
	.w7(32'hbac9b021),
	.w8(32'hbc05c09d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dcd29),
	.w1(32'hbb80a060),
	.w2(32'hbb880822),
	.w3(32'hb9a8c432),
	.w4(32'hbad09585),
	.w5(32'hbba895bf),
	.w6(32'hbb24c41b),
	.w7(32'hbb4c78ad),
	.w8(32'h3bba52ba),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd53e7),
	.w1(32'h3b9f5fdc),
	.w2(32'hbbe61e70),
	.w3(32'h3ac1ee98),
	.w4(32'hba54a453),
	.w5(32'h37c4a590),
	.w6(32'hbb2b3c34),
	.w7(32'hbb834fcf),
	.w8(32'hbbd031e5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bab8f),
	.w1(32'hbbc17fcf),
	.w2(32'hba4314f5),
	.w3(32'h3b297c3f),
	.w4(32'hbbc0c3ed),
	.w5(32'h3a811b3f),
	.w6(32'hbc7c0be9),
	.w7(32'hbbc30371),
	.w8(32'h3b194ba8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99c9a4),
	.w1(32'h3c80826d),
	.w2(32'hbbdbd437),
	.w3(32'hba766cd2),
	.w4(32'h3c093ab2),
	.w5(32'h3c16583c),
	.w6(32'h3b0a61e7),
	.w7(32'h39c58065),
	.w8(32'hbc1f3139),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79fe8a),
	.w1(32'h3c170227),
	.w2(32'hbcd22b17),
	.w3(32'hba0440ad),
	.w4(32'h3c05f4cd),
	.w5(32'hbc40836c),
	.w6(32'h3bd749d3),
	.w7(32'h3b745140),
	.w8(32'h3c4f2f47),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9a46a),
	.w1(32'h3d5834e3),
	.w2(32'hbc97e597),
	.w3(32'hbb70e3b5),
	.w4(32'h3c7801c4),
	.w5(32'hbbb43406),
	.w6(32'h3c8a9343),
	.w7(32'hbc1e65c9),
	.w8(32'hbca0d2d1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd169492),
	.w1(32'hbce246e3),
	.w2(32'hbc282ea8),
	.w3(32'hbbd5b945),
	.w4(32'hbb70ad24),
	.w5(32'hbc855c85),
	.w6(32'hbba76a4f),
	.w7(32'h3af4767c),
	.w8(32'hbc651134),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54a513),
	.w1(32'h3cdac6f9),
	.w2(32'hbc57af4a),
	.w3(32'hbcdfd85a),
	.w4(32'h3b97295b),
	.w5(32'h3b8f1f6f),
	.w6(32'hbcab3cce),
	.w7(32'hbb325233),
	.w8(32'hbce20b93),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0e1266),
	.w1(32'hbc123a1b),
	.w2(32'h3c7b1d59),
	.w3(32'hbc0be558),
	.w4(32'hbba951ff),
	.w5(32'h3a173f4a),
	.w6(32'h3bba15ab),
	.w7(32'h3bf39915),
	.w8(32'hba528e3e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74f6ab),
	.w1(32'hbbd267c9),
	.w2(32'hbd24b374),
	.w3(32'hbbb23c00),
	.w4(32'hbbcc6f32),
	.w5(32'hbd0337b3),
	.w6(32'hbc135c9b),
	.w7(32'hbc9c0b3a),
	.w8(32'h394cc9e4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7520a2),
	.w1(32'h3d85e7a1),
	.w2(32'hbc96ed62),
	.w3(32'hbb8de61a),
	.w4(32'h3c9f477f),
	.w5(32'h3b011b60),
	.w6(32'h3ca83b67),
	.w7(32'hbc2c1649),
	.w8(32'hbc8c8a5c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbd32c),
	.w1(32'h3c584c18),
	.w2(32'hbba660ad),
	.w3(32'h3b4155be),
	.w4(32'h3ac1e8ae),
	.w5(32'hba1d774b),
	.w6(32'h374caa15),
	.w7(32'hbbd8e6b3),
	.w8(32'hbc6b23ba),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9301d7),
	.w1(32'hbb1ba9eb),
	.w2(32'hbcb13c45),
	.w3(32'hbbdddebc),
	.w4(32'hb9612ced),
	.w5(32'hbbe7fd78),
	.w6(32'h39d7f9da),
	.w7(32'hbbc1fe00),
	.w8(32'hb8b6f4d2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133883),
	.w1(32'hbba1a0be),
	.w2(32'hbbb7c573),
	.w3(32'h3b7461e0),
	.w4(32'h3a4150bd),
	.w5(32'h3bba01be),
	.w6(32'hbc6af43f),
	.w7(32'hba310093),
	.w8(32'hbaa3eb49),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba987f49),
	.w1(32'hbbbb2052),
	.w2(32'hbbeb8d8e),
	.w3(32'h3c1e60cf),
	.w4(32'h3b77f629),
	.w5(32'hba290390),
	.w6(32'hbc4ea01d),
	.w7(32'h3b089abd),
	.w8(32'h3b858b25),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bb058),
	.w1(32'hbc07cc68),
	.w2(32'h3c5e82ec),
	.w3(32'h3b85377a),
	.w4(32'h3ba01a4c),
	.w5(32'h39c543e7),
	.w6(32'hbb46650d),
	.w7(32'h39a928d9),
	.w8(32'hbc37be24),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31dd12),
	.w1(32'h3c8f6b3f),
	.w2(32'hbcc1ad0e),
	.w3(32'hbc8a9b5a),
	.w4(32'h3c0a114d),
	.w5(32'hbc5ec9dc),
	.w6(32'h3ad69c9f),
	.w7(32'hbb32fe6a),
	.w8(32'hbc6362d3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ae127),
	.w1(32'h3d60baaa),
	.w2(32'hbc70b64d),
	.w3(32'hbc104214),
	.w4(32'h3c9b9262),
	.w5(32'h3ad0a0ef),
	.w6(32'h3c68de47),
	.w7(32'hbc156d19),
	.w8(32'hbcac91aa),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce29b99),
	.w1(32'hbc724501),
	.w2(32'h3b7d3241),
	.w3(32'h3923fb51),
	.w4(32'hbb7235d2),
	.w5(32'hbc196b3f),
	.w6(32'h39e1b380),
	.w7(32'hbaab6eba),
	.w8(32'hbbe82512),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b3c47),
	.w1(32'hbca8d611),
	.w2(32'h3c20a857),
	.w3(32'hbc62db70),
	.w4(32'hbbb0db05),
	.w5(32'hbba7e26a),
	.w6(32'hbb2b1da2),
	.w7(32'h3b3ad253),
	.w8(32'hbabcddf4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8111d3),
	.w1(32'hbc5bbefb),
	.w2(32'h3b2f9b70),
	.w3(32'hbc44d69b),
	.w4(32'hbb08d7af),
	.w5(32'hbb83c01a),
	.w6(32'hbb7205ab),
	.w7(32'h3a196ae0),
	.w8(32'h3ad458b6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e370),
	.w1(32'h3d186f07),
	.w2(32'hbc7f1fb5),
	.w3(32'hbc601f12),
	.w4(32'h3c72a25d),
	.w5(32'h3b148759),
	.w6(32'h3b9b47f0),
	.w7(32'h3847493e),
	.w8(32'hbc8504b1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05f494),
	.w1(32'h3c9db994),
	.w2(32'hbc335aa2),
	.w3(32'hbbfd0c05),
	.w4(32'h3ba5d717),
	.w5(32'h3c49a249),
	.w6(32'hbc3dac25),
	.w7(32'hb91385f7),
	.w8(32'hbc5fb249),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e511e),
	.w1(32'hbd14af87),
	.w2(32'h3c6855bd),
	.w3(32'hbb9fea1e),
	.w4(32'hbb84075c),
	.w5(32'hbc12169d),
	.w6(32'hbc3c082d),
	.w7(32'h3b775240),
	.w8(32'h3c18b200),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea9686),
	.w1(32'h3cd73352),
	.w2(32'hbc8c7d7a),
	.w3(32'hbb8aa71c),
	.w4(32'h3aa59c86),
	.w5(32'hbb91359e),
	.w6(32'h3a329fea),
	.w7(32'hbc22afc8),
	.w8(32'hbbd580ee),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf0104f),
	.w1(32'hbb236fe8),
	.w2(32'hbc371d1d),
	.w3(32'h3b296113),
	.w4(32'h3ba83195),
	.w5(32'h3baca623),
	.w6(32'hbc4dc5b4),
	.w7(32'hbac7a60b),
	.w8(32'h3bd20f03),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc96eea),
	.w1(32'hbcba7489),
	.w2(32'hbbd8063f),
	.w3(32'h3bcf2e72),
	.w4(32'hbbf4f5ad),
	.w5(32'hbc61a1b1),
	.w6(32'hbc84756d),
	.w7(32'hbc41ff59),
	.w8(32'hbbe7b3cc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc63c7),
	.w1(32'hbb5a6574),
	.w2(32'hbbd418e0),
	.w3(32'hbc24b08e),
	.w4(32'h3b6fd0d2),
	.w5(32'h3a429938),
	.w6(32'hbc44bfe3),
	.w7(32'h3b83f0aa),
	.w8(32'hbafbb372),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d7a00),
	.w1(32'h3d20f199),
	.w2(32'h3bd9a0a8),
	.w3(32'h3bf836f4),
	.w4(32'h3c54eb48),
	.w5(32'h3c5c8e57),
	.w6(32'h3c6386c4),
	.w7(32'h3bffc0a3),
	.w8(32'hbc08ad84),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0bff8),
	.w1(32'h3b430358),
	.w2(32'hbb61726f),
	.w3(32'h3a42475e),
	.w4(32'h3af56256),
	.w5(32'h3b20c149),
	.w6(32'h3b972626),
	.w7(32'h382a1db6),
	.w8(32'h3b24e2a4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc142236),
	.w1(32'h3d199881),
	.w2(32'hbc3eb6c9),
	.w3(32'h3ad83ef0),
	.w4(32'h3c1fbb08),
	.w5(32'hbb2d8f5a),
	.w6(32'h3a3bf671),
	.w7(32'hbb1a9f91),
	.w8(32'hbce0324f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2764aa),
	.w1(32'hbc114ba4),
	.w2(32'hbc177f5e),
	.w3(32'hbc79747f),
	.w4(32'h3b326667),
	.w5(32'hbbb2a9a0),
	.w6(32'hbc0ec165),
	.w7(32'h3be3e00c),
	.w8(32'hbc7b3c28),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca27053),
	.w1(32'h3caa1269),
	.w2(32'hbbd155e1),
	.w3(32'hbbf8dc1f),
	.w4(32'h3c8bcf3f),
	.w5(32'h3c433906),
	.w6(32'hbac3296c),
	.w7(32'h3ba79ddf),
	.w8(32'hbbc9a2f6),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4185),
	.w1(32'h3c79fb61),
	.w2(32'hbcb7b149),
	.w3(32'h3b74c9dd),
	.w4(32'h3bd2c465),
	.w5(32'hbbb2781c),
	.w6(32'h3a19fc42),
	.w7(32'hbc052150),
	.w8(32'hbb96790f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf809f),
	.w1(32'hbc472652),
	.w2(32'h3b793bd8),
	.w3(32'h3be4d036),
	.w4(32'hbb8ab0fa),
	.w5(32'hbaf7508c),
	.w6(32'hbb9b08b6),
	.w7(32'hba9dbd18),
	.w8(32'h3abdf902),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d43d9),
	.w1(32'h3bbe1e7d),
	.w2(32'hbbd8e337),
	.w3(32'hbb4d4b69),
	.w4(32'hba4d2f6e),
	.w5(32'h39f71f0b),
	.w6(32'hbad62c92),
	.w7(32'hbb1a9ab5),
	.w8(32'hbbb3d7d4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42ac7),
	.w1(32'hbc736806),
	.w2(32'hbb00e94e),
	.w3(32'h3a873751),
	.w4(32'hbc4006fd),
	.w5(32'hbc83b7dc),
	.w6(32'hbbfbc35b),
	.w7(32'hbb8c91c5),
	.w8(32'hbbed05a4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dea68),
	.w1(32'hbc82eed3),
	.w2(32'hbb89406e),
	.w3(32'hbbf58357),
	.w4(32'hbb096826),
	.w5(32'hbba5154a),
	.w6(32'hbba92843),
	.w7(32'h3bb2e4b5),
	.w8(32'h3ae65c3b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5ed2),
	.w1(32'h3d466c35),
	.w2(32'hbc8b1889),
	.w3(32'hbb9728e4),
	.w4(32'h3c78f91c),
	.w5(32'h3b91f93e),
	.w6(32'h3c43c994),
	.w7(32'hbc4b97f9),
	.w8(32'hbd0a9e36),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3e381f),
	.w1(32'h3cfc36d2),
	.w2(32'h3bdee055),
	.w3(32'hbc05598f),
	.w4(32'h3c911fa1),
	.w5(32'h3c6a7d67),
	.w6(32'hbbe370fe),
	.w7(32'h3b6b8dc4),
	.w8(32'hbbd1615f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc987b08),
	.w1(32'hbc2b23fd),
	.w2(32'hbbc884f7),
	.w3(32'h39f3dee8),
	.w4(32'hbaeadfdf),
	.w5(32'hbb0615c5),
	.w6(32'hbca14450),
	.w7(32'hbba00a76),
	.w8(32'hbb3d5b71),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8df12e),
	.w1(32'h3d022244),
	.w2(32'h3a2a16df),
	.w3(32'h3b19bf9a),
	.w4(32'h3c023de1),
	.w5(32'h3b4b6a4b),
	.w6(32'h3bd0ac38),
	.w7(32'hbba5675f),
	.w8(32'hbc5a5dd5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68727f),
	.w1(32'hbb5760a5),
	.w2(32'h3a2c29e5),
	.w3(32'hbbd744f4),
	.w4(32'h3a9167e9),
	.w5(32'h3b42e6d7),
	.w6(32'hbaf846ef),
	.w7(32'hbbd24ec0),
	.w8(32'h3af5fd22),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dc9e7),
	.w1(32'hbb95bc23),
	.w2(32'hbb0cfbd5),
	.w3(32'h3b9d607b),
	.w4(32'hbc031a8b),
	.w5(32'hbb9409cc),
	.w6(32'hbb0aa85b),
	.w7(32'hba5be212),
	.w8(32'hbae03c46),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49b712),
	.w1(32'h39bfb2f5),
	.w2(32'hbcd9d067),
	.w3(32'h3c1892e1),
	.w4(32'h3b279470),
	.w5(32'hbc60d9e5),
	.w6(32'hbb77d7bc),
	.w7(32'hbc3f6e38),
	.w8(32'h3c63af5f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa0fc9),
	.w1(32'h3cea9954),
	.w2(32'hbb1a4f37),
	.w3(32'h3c66b1be),
	.w4(32'hbb992553),
	.w5(32'h3b8a8288),
	.w6(32'h38b4a332),
	.w7(32'hbb07c053),
	.w8(32'hbcb9a25f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd350303),
	.w1(32'h3b70ccaa),
	.w2(32'hba11ef2c),
	.w3(32'hbc28328e),
	.w4(32'h3c0d1740),
	.w5(32'h3b96454e),
	.w6(32'hbbabda07),
	.w7(32'hbaeef540),
	.w8(32'hbba8da2d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933f0c),
	.w1(32'h3bd425f9),
	.w2(32'hbc8df5ff),
	.w3(32'h3bca1010),
	.w4(32'h3b4eea17),
	.w5(32'hbbafa8b6),
	.w6(32'hbc06badb),
	.w7(32'hbbb405a8),
	.w8(32'h3a0e0262),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46556e),
	.w1(32'h3b568d46),
	.w2(32'h3b7b2bac),
	.w3(32'h3c042531),
	.w4(32'h3b8316c4),
	.w5(32'h3b37af5b),
	.w6(32'h3c205783),
	.w7(32'hbbb811e5),
	.w8(32'hbbff4156),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3c907),
	.w1(32'hbd6da993),
	.w2(32'h3c7a1528),
	.w3(32'hb845b63b),
	.w4(32'hbc4f7885),
	.w5(32'hbcab6d62),
	.w6(32'hbb500544),
	.w7(32'h3bbd9c8b),
	.w8(32'h3c3e904f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d333d65),
	.w1(32'hbc675c1a),
	.w2(32'h3acc2cc8),
	.w3(32'hbb89a98f),
	.w4(32'h3a8a7989),
	.w5(32'hbc28a755),
	.w6(32'h39e52dde),
	.w7(32'hbb9416e5),
	.w8(32'hbc1aafbd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a4ff),
	.w1(32'hbcef17d7),
	.w2(32'h3c56e08e),
	.w3(32'hbc42d327),
	.w4(32'hbbf1898d),
	.w5(32'hbbf2849e),
	.w6(32'hbb3a008e),
	.w7(32'h3ab121cf),
	.w8(32'h3c2bd956),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb937f5),
	.w1(32'hbc141dc4),
	.w2(32'hbc29f868),
	.w3(32'hbb4ee855),
	.w4(32'hbbb117d9),
	.w5(32'hbc48a43c),
	.w6(32'hbbafdca6),
	.w7(32'hbc2e86b0),
	.w8(32'hbc35aa79),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c499a),
	.w1(32'h3d09b16d),
	.w2(32'h3a815755),
	.w3(32'hbc09162e),
	.w4(32'h3bcff406),
	.w5(32'hb9afbdd4),
	.w6(32'h3c12fd9d),
	.w7(32'hbad22f41),
	.w8(32'hbc8abb72),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc792da),
	.w1(32'hbc798097),
	.w2(32'h3c330dd0),
	.w3(32'hbc2db537),
	.w4(32'hbb9e1dfc),
	.w5(32'h3b65a886),
	.w6(32'hbb42bdcf),
	.w7(32'h3be31e4b),
	.w8(32'h3c4aa04f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71f09f),
	.w1(32'hbcf0570c),
	.w2(32'h3c75b602),
	.w3(32'h3b1d9889),
	.w4(32'hbbd2d304),
	.w5(32'hbbc86fad),
	.w6(32'hba508a7f),
	.w7(32'h3b53b8b8),
	.w8(32'h3c34546e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc44d30),
	.w1(32'h3d5ba4e4),
	.w2(32'hbc40a8ab),
	.w3(32'hbac27abb),
	.w4(32'h3c98223b),
	.w5(32'hbab93bad),
	.w6(32'h3ce09f8e),
	.w7(32'hbb717c2f),
	.w8(32'hbc89ddc1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f3604),
	.w1(32'hbc487003),
	.w2(32'h3c3a5ebc),
	.w3(32'hbc40bb1c),
	.w4(32'h3a9a559f),
	.w5(32'h3adb560c),
	.w6(32'hbbdaecde),
	.w7(32'h3bb7e14a),
	.w8(32'h381c8fa1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bc245),
	.w1(32'hb9b86763),
	.w2(32'hbc8d292c),
	.w3(32'hbc460ab9),
	.w4(32'hba19a048),
	.w5(32'hbc86caa0),
	.w6(32'hbc046ca3),
	.w7(32'hbbbbed6f),
	.w8(32'hbbf8d3bc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45c77d),
	.w1(32'hbc328ce7),
	.w2(32'h3b0dd01b),
	.w3(32'hbbde23c1),
	.w4(32'h3b617195),
	.w5(32'hbbe94958),
	.w6(32'hbbc4fced),
	.w7(32'h3a66dc70),
	.w8(32'hbbd7f072),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb018db3),
	.w1(32'h3d2ae2cd),
	.w2(32'hbccd2cbc),
	.w3(32'hbc61b0f4),
	.w4(32'h3c6af853),
	.w5(32'hbb1f5310),
	.w6(32'h3c11d0b0),
	.w7(32'hbbfb6b6d),
	.w8(32'hbc88e81b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bc4aa),
	.w1(32'h3992ea54),
	.w2(32'h3c3fe05f),
	.w3(32'h3b664458),
	.w4(32'h3c0fd27d),
	.w5(32'h3c3f720c),
	.w6(32'h3c030ecc),
	.w7(32'h3b589027),
	.w8(32'h3bcc59d5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59ffe5),
	.w1(32'hbd2f0b8a),
	.w2(32'h3ca508c6),
	.w3(32'h3b3d36c5),
	.w4(32'hbc226305),
	.w5(32'hbc21e4d6),
	.w6(32'hbb0ec42b),
	.w7(32'h3b4d65e3),
	.w8(32'h3c806fcd),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e0b3a),
	.w1(32'hbce25b39),
	.w2(32'h3c177ca0),
	.w3(32'hbb189dd6),
	.w4(32'hbbf7daf5),
	.w5(32'hbc01346d),
	.w6(32'hbbe2b397),
	.w7(32'hb94221fb),
	.w8(32'h3b6e8132),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65f617),
	.w1(32'hbd004871),
	.w2(32'h3c2c4cf0),
	.w3(32'hbb9694ff),
	.w4(32'hbc175931),
	.w5(32'hbc02c59d),
	.w6(32'hbc1123e0),
	.w7(32'hba94abcd),
	.w8(32'h3bd164ec),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb0b2d),
	.w1(32'hbb267ff8),
	.w2(32'hbbb18f4c),
	.w3(32'hbbdcd24e),
	.w4(32'hbb45ea93),
	.w5(32'hbbda20c4),
	.w6(32'hbb9260ca),
	.w7(32'h3ba4ac3b),
	.w8(32'h3b341ed7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd7d86),
	.w1(32'h3cea40f3),
	.w2(32'hbc8d5f5a),
	.w3(32'hbab87d0c),
	.w4(32'h3c1d4ac1),
	.w5(32'h3c0be0f9),
	.w6(32'hbb8c06c9),
	.w7(32'hbc10d355),
	.w8(32'hbbeb9222),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc351a08),
	.w1(32'hbabfd2ed),
	.w2(32'hb9a29fb7),
	.w3(32'hba905d00),
	.w4(32'h3c058e02),
	.w5(32'hbb4b65c2),
	.w6(32'h3b45923f),
	.w7(32'hbb2eb5fb),
	.w8(32'hbace6133),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f37b3),
	.w1(32'hbbb939a8),
	.w2(32'hbb0a8f37),
	.w3(32'hbb999a90),
	.w4(32'hba9231eb),
	.w5(32'hba4e1215),
	.w6(32'hbb379b4e),
	.w7(32'hbb8ef1d1),
	.w8(32'hba825971),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc5e6d),
	.w1(32'hbcdfc10f),
	.w2(32'h3c2a190b),
	.w3(32'hbc19dda1),
	.w4(32'hbc08e69f),
	.w5(32'hbc16be42),
	.w6(32'hbbb0e398),
	.w7(32'h394eb059),
	.w8(32'hbb071052),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1955bf),
	.w1(32'h3a87f99a),
	.w2(32'hba81de78),
	.w3(32'hbc8699b1),
	.w4(32'hba1918d6),
	.w5(32'h3b543f1e),
	.w6(32'h39c62180),
	.w7(32'h3ba45cc8),
	.w8(32'hbb618fde),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6ca3),
	.w1(32'hbc1c7ce6),
	.w2(32'h3c1f46d7),
	.w3(32'h3b28d891),
	.w4(32'h3b749a0b),
	.w5(32'h3bb9854e),
	.w6(32'hbb2ce8e6),
	.w7(32'hbc14bfbb),
	.w8(32'hba68b354),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985da58),
	.w1(32'hbcd2c01c),
	.w2(32'hbc59f898),
	.w3(32'h3b170ed9),
	.w4(32'hbc34512c),
	.w5(32'hbc4e6720),
	.w6(32'hbca4f4ca),
	.w7(32'hbc573ba8),
	.w8(32'hbc1dc0fd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62c9d0),
	.w1(32'hb8c9e6ec),
	.w2(32'hb8033eaf),
	.w3(32'hbc33dc2b),
	.w4(32'hb902c9fa),
	.w5(32'hb8293978),
	.w6(32'h38112048),
	.w7(32'hb8d71816),
	.w8(32'h37914179),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacaa86),
	.w1(32'h3b843d77),
	.w2(32'h3b9ed537),
	.w3(32'hbb94bf59),
	.w4(32'h3b4f5eab),
	.w5(32'h3b48f434),
	.w6(32'hbc27fcbe),
	.w7(32'hbb5101a5),
	.w8(32'hbb2dabc6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule