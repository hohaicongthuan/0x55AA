module layer_10_featuremap_285(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa25874),
	.w1(32'hbc0d8b1f),
	.w2(32'hbc28ff61),
	.w3(32'hbb68d76f),
	.w4(32'h3ae37aa6),
	.w5(32'h3b0cc10a),
	.w6(32'h3c075560),
	.w7(32'hba8b1e15),
	.w8(32'hbb014c1d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231c83),
	.w1(32'hbb984828),
	.w2(32'hba988c78),
	.w3(32'h3b8132c4),
	.w4(32'hbb9d41b6),
	.w5(32'hbc076190),
	.w6(32'h3b8f842f),
	.w7(32'h3b77e0c1),
	.w8(32'hbb4eb634),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26dd20),
	.w1(32'hba35b62f),
	.w2(32'hbb8fd656),
	.w3(32'hbc3a8e3d),
	.w4(32'hbbd84635),
	.w5(32'h3b4819e4),
	.w6(32'hbb895526),
	.w7(32'hbaca591d),
	.w8(32'hba97387a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7e06),
	.w1(32'h3abfaa0c),
	.w2(32'h3b96819f),
	.w3(32'h3b8f9270),
	.w4(32'h3b9a5828),
	.w5(32'hbbcf8cc1),
	.w6(32'hba0a676d),
	.w7(32'h3b822521),
	.w8(32'hbb9a73ec),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee3f3),
	.w1(32'h38e86c73),
	.w2(32'hbb04ab45),
	.w3(32'hbb8fcb94),
	.w4(32'hbc106c17),
	.w5(32'h3ba639a9),
	.w6(32'hbba61a7a),
	.w7(32'hbb875069),
	.w8(32'h3b3805ed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c826e),
	.w1(32'hbb72d0c5),
	.w2(32'h3b3a068c),
	.w3(32'h3c2f8b48),
	.w4(32'h3bed32da),
	.w5(32'h3be9c4d5),
	.w6(32'h3b8827d3),
	.w7(32'h3bcdf952),
	.w8(32'hb9ea8e6d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f5982),
	.w1(32'hbb177595),
	.w2(32'h3aafbd07),
	.w3(32'h3bdf01d6),
	.w4(32'h3c038e2b),
	.w5(32'hbab6993b),
	.w6(32'hb9783acc),
	.w7(32'h3bb8af98),
	.w8(32'h3ac51b56),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc15e8b),
	.w1(32'h3a8c9d9b),
	.w2(32'h3bc60275),
	.w3(32'hbc13e719),
	.w4(32'hbb219624),
	.w5(32'h3c19dc60),
	.w6(32'hbb423815),
	.w7(32'hbabc65fd),
	.w8(32'h3bd457cf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d7e62),
	.w1(32'hba685c3a),
	.w2(32'h3ad6cd36),
	.w3(32'h3b51c89b),
	.w4(32'h3af38895),
	.w5(32'h3bc3a966),
	.w6(32'h3b63b8bb),
	.w7(32'h3b8d5cdd),
	.w8(32'hb9e918de),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcef9e),
	.w1(32'hbc3ad007),
	.w2(32'hba50bd69),
	.w3(32'h3baef9c5),
	.w4(32'h3b47444a),
	.w5(32'hba5c626c),
	.w6(32'h3ba068c7),
	.w7(32'h3bc7fcf0),
	.w8(32'h399aa5a2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e3360),
	.w1(32'hbbbd326b),
	.w2(32'h3a593cb8),
	.w3(32'h3ba94c01),
	.w4(32'h3b6fa0ce),
	.w5(32'hbba423a3),
	.w6(32'h3b26bda9),
	.w7(32'h3b88106b),
	.w8(32'hbb88aad6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f6a6c),
	.w1(32'hb80d5977),
	.w2(32'hbbd1c6c3),
	.w3(32'h3ae39bc9),
	.w4(32'hb98f3186),
	.w5(32'hbad39f36),
	.w6(32'hbbea4e0f),
	.w7(32'hbb365af4),
	.w8(32'h3b3b1939),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2901fb),
	.w1(32'hbba7bd2e),
	.w2(32'h3b9cc905),
	.w3(32'hbb6da808),
	.w4(32'hbbe1eb17),
	.w5(32'hba649817),
	.w6(32'h3b96006d),
	.w7(32'hba9cd16a),
	.w8(32'h3af23a79),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04126a),
	.w1(32'hbbd9bde4),
	.w2(32'hba0011d0),
	.w3(32'hbbc8d350),
	.w4(32'hbc046198),
	.w5(32'h3b6e97ae),
	.w6(32'hbbb1708d),
	.w7(32'hba928f0e),
	.w8(32'hbaa11519),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e9bad),
	.w1(32'hbba88871),
	.w2(32'h3b90d8e6),
	.w3(32'h3bf01adf),
	.w4(32'h3bc01efa),
	.w5(32'h3ad19b6c),
	.w6(32'hbb4eb873),
	.w7(32'h3aa923e3),
	.w8(32'h3a63d43f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0899c),
	.w1(32'hbc33db6b),
	.w2(32'hbbaa694e),
	.w3(32'hbb4e58fb),
	.w4(32'hbb36acd4),
	.w5(32'h3b4f0789),
	.w6(32'hbc0f9b12),
	.w7(32'hbadd44aa),
	.w8(32'h3b889155),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87fe57),
	.w1(32'h399edf43),
	.w2(32'h3b8ec03d),
	.w3(32'h3b4f480d),
	.w4(32'h3aad9343),
	.w5(32'h3a053c3e),
	.w6(32'h3bc91fd5),
	.w7(32'h3b4516f4),
	.w8(32'h3a62838a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0b2a5),
	.w1(32'hbc427db7),
	.w2(32'hbb1179b1),
	.w3(32'hbacf201c),
	.w4(32'hbb89c12e),
	.w5(32'hba049c5d),
	.w6(32'h3b95b9e3),
	.w7(32'h3b9237aa),
	.w8(32'h3bb4315b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9ab89),
	.w1(32'hbc118c1f),
	.w2(32'hbb0e5216),
	.w3(32'hb9cabd01),
	.w4(32'hbb2d2c8b),
	.w5(32'h3b833f92),
	.w6(32'h3b42e1de),
	.w7(32'h3a96bd49),
	.w8(32'hbb95dd80),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1388),
	.w1(32'h3abccebc),
	.w2(32'hbb06a9b3),
	.w3(32'h3b54596b),
	.w4(32'hbb3740d9),
	.w5(32'h3b8428a0),
	.w6(32'h3b3f1ebf),
	.w7(32'h3aeae8a0),
	.w8(32'h3bffebfb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb882d1),
	.w1(32'hbc077fa6),
	.w2(32'hbc028d67),
	.w3(32'hbbf64980),
	.w4(32'hbbbf1c6b),
	.w5(32'hb9c2711e),
	.w6(32'hbbe41de0),
	.w7(32'hbbdbbf53),
	.w8(32'hbb071e15),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7b4b4),
	.w1(32'h3bba3a19),
	.w2(32'h3c088014),
	.w3(32'hbb27e0f6),
	.w4(32'h3adf04c3),
	.w5(32'hb98cc9a1),
	.w6(32'hbb0bbabf),
	.w7(32'h3b7a3880),
	.w8(32'hbb44de0a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04cda5),
	.w1(32'hbc35c772),
	.w2(32'h3aed420f),
	.w3(32'h394300c2),
	.w4(32'hbc01f857),
	.w5(32'hbb15079f),
	.w6(32'hbb76f9b9),
	.w7(32'hb9e8a4d0),
	.w8(32'h3bd21d18),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082f9f),
	.w1(32'hbc5b0ccc),
	.w2(32'hbac43064),
	.w3(32'hba9b79a5),
	.w4(32'hbbfea9d8),
	.w5(32'hbba5e500),
	.w6(32'hbc0bef11),
	.w7(32'hbc09f363),
	.w8(32'hb9dee1a5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5b213),
	.w1(32'hbb6455fb),
	.w2(32'h3a86b24c),
	.w3(32'hbb8a58a2),
	.w4(32'hbadd4183),
	.w5(32'h3afb2c2a),
	.w6(32'h393b9c90),
	.w7(32'h39dc079e),
	.w8(32'h3a004c1a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73e1c0),
	.w1(32'hbbc99e9f),
	.w2(32'hbb14426d),
	.w3(32'h39b658db),
	.w4(32'h3b9e914b),
	.w5(32'hbb49f606),
	.w6(32'hb911b484),
	.w7(32'hbb2a3a34),
	.w8(32'hbaade818),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4ab5b),
	.w1(32'hb8ee0564),
	.w2(32'hba56f2b6),
	.w3(32'hbb18a1f9),
	.w4(32'h38dd4a55),
	.w5(32'h3bbb5744),
	.w6(32'hbb59fe17),
	.w7(32'hba0b181d),
	.w8(32'h3bd9580e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7ce2f),
	.w1(32'hbbb16779),
	.w2(32'hbbb44f55),
	.w3(32'h3b7ba635),
	.w4(32'h3b5c8085),
	.w5(32'h3bb18cae),
	.w6(32'h3c0738c5),
	.w7(32'h3af28572),
	.w8(32'hbb93bb96),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5cf3c),
	.w1(32'hbb056a5a),
	.w2(32'hbaecc56b),
	.w3(32'h3a767c0e),
	.w4(32'hba25cb5b),
	.w5(32'hbb3a96d5),
	.w6(32'h3ac7060c),
	.w7(32'hba39ef44),
	.w8(32'hbc2094f2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0286),
	.w1(32'h3b53815b),
	.w2(32'h3acb0ad1),
	.w3(32'h3ac41860),
	.w4(32'hbbb10d5b),
	.w5(32'h3c3f39af),
	.w6(32'h3bb8c2e5),
	.w7(32'hbb089912),
	.w8(32'h3baef583),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd30b78),
	.w1(32'hbabba120),
	.w2(32'h3ba2fada),
	.w3(32'h3baa6839),
	.w4(32'h3b80d72f),
	.w5(32'h3a4fbad7),
	.w6(32'h3bc1c7cb),
	.w7(32'h3b4cf180),
	.w8(32'h3b8a128d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf5893),
	.w1(32'hba1a8639),
	.w2(32'hbb29dc58),
	.w3(32'hbba61a33),
	.w4(32'hbb13486e),
	.w5(32'hbb9fcf17),
	.w6(32'hbaf6c545),
	.w7(32'hbb07979a),
	.w8(32'hbb98b70c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca07dd),
	.w1(32'hbb10a248),
	.w2(32'hbb0bef38),
	.w3(32'hba19746b),
	.w4(32'hb9fac79d),
	.w5(32'h3b3cec7a),
	.w6(32'h3aa61acb),
	.w7(32'h3a8cfa18),
	.w8(32'h3a5d0d7c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10a49),
	.w1(32'hbb85d2b3),
	.w2(32'h39f70022),
	.w3(32'h3bcd58c6),
	.w4(32'h3b2eebd7),
	.w5(32'h39d4518b),
	.w6(32'hba48868c),
	.w7(32'h3b722c90),
	.w8(32'hbb1d5713),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393087d0),
	.w1(32'hbb5d9554),
	.w2(32'hbb0c1940),
	.w3(32'hbb524c2e),
	.w4(32'hbb858769),
	.w5(32'h3be17699),
	.w6(32'hbb60ad6d),
	.w7(32'hbbe1a52c),
	.w8(32'h3bab4de5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef0938),
	.w1(32'hbc4948b7),
	.w2(32'hbb66ce19),
	.w3(32'hb71b5544),
	.w4(32'hbb0bc9e7),
	.w5(32'h3bb67391),
	.w6(32'h3c0cd4ea),
	.w7(32'hb8bbf56f),
	.w8(32'hba85bccc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf0b32),
	.w1(32'hbb89b950),
	.w2(32'hbb025bf1),
	.w3(32'h3c0404bd),
	.w4(32'h3ab4a33e),
	.w5(32'h3b0f89dd),
	.w6(32'h3bba8588),
	.w7(32'h3af688d0),
	.w8(32'h3b855fc7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6c86),
	.w1(32'h3966a05e),
	.w2(32'hbb82c194),
	.w3(32'h3c257989),
	.w4(32'h3c47ae55),
	.w5(32'h3af67674),
	.w6(32'h3bba29a9),
	.w7(32'h3c1f6268),
	.w8(32'hbc254024),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a14f),
	.w1(32'hbc1e937f),
	.w2(32'h3924b069),
	.w3(32'hbb6806d0),
	.w4(32'hba4b6389),
	.w5(32'hba8bc16a),
	.w6(32'hbb4f362d),
	.w7(32'hbbc35be5),
	.w8(32'hbb3c5bec),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7240de),
	.w1(32'h3c0807a4),
	.w2(32'h3c145fd9),
	.w3(32'hba418b64),
	.w4(32'h3c1cf34e),
	.w5(32'hbb5cea10),
	.w6(32'h3b0dadf7),
	.w7(32'h3c11e8fc),
	.w8(32'hbb1d8ee5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8b23b),
	.w1(32'h3b43ed23),
	.w2(32'h3aea6119),
	.w3(32'hba4dd5fe),
	.w4(32'hbbb6d0e6),
	.w5(32'hbaf0973d),
	.w6(32'hbb2c3edc),
	.w7(32'hbb8dfd9e),
	.w8(32'hbbf1d0a4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4131b7),
	.w1(32'hbbad97dc),
	.w2(32'hbafb3490),
	.w3(32'hbb31e892),
	.w4(32'h3a4a9233),
	.w5(32'hba9a5c23),
	.w6(32'hbc1499af),
	.w7(32'hbb8e3da3),
	.w8(32'hbb4bfae0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d540e),
	.w1(32'hbc1c9450),
	.w2(32'hbc2cd0de),
	.w3(32'h3a15f857),
	.w4(32'hba5570df),
	.w5(32'hbac7c439),
	.w6(32'hbba97f01),
	.w7(32'hbbeb4175),
	.w8(32'h3b042c36),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9c133),
	.w1(32'hbc048a63),
	.w2(32'hbb435504),
	.w3(32'hbac220ea),
	.w4(32'hbb75e387),
	.w5(32'h3ae87c99),
	.w6(32'h3b37af02),
	.w7(32'h3bdd172a),
	.w8(32'h3a43e701),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80a104),
	.w1(32'hb991064b),
	.w2(32'hba191ced),
	.w3(32'h3b9211ec),
	.w4(32'h3b8ded1d),
	.w5(32'hbb3aefec),
	.w6(32'h3acc8134),
	.w7(32'h3b21aa16),
	.w8(32'hbae9884b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6faf79),
	.w1(32'hbc3c8e8e),
	.w2(32'hbbdf612f),
	.w3(32'hbbd223e3),
	.w4(32'hbb363efe),
	.w5(32'hbb6a3908),
	.w6(32'hbba5bead),
	.w7(32'hbb9c430a),
	.w8(32'hba3cb934),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d86d7),
	.w1(32'hbb2a567f),
	.w2(32'hbbb0c266),
	.w3(32'hbbb11076),
	.w4(32'hbb699bc4),
	.w5(32'h3b95c4a1),
	.w6(32'hba836aa1),
	.w7(32'hbb363bdd),
	.w8(32'h3b4a5625),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc5de),
	.w1(32'hbc5d38bb),
	.w2(32'h3b65c754),
	.w3(32'hbbc6161e),
	.w4(32'hbc135a12),
	.w5(32'hb8756915),
	.w6(32'h3af70c23),
	.w7(32'h3abebd81),
	.w8(32'h3bc77eb4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae9ce4),
	.w1(32'hbbbffe74),
	.w2(32'hbb07d76b),
	.w3(32'h3a6354d4),
	.w4(32'hbb1a383d),
	.w5(32'hbafc3599),
	.w6(32'h3b695ef5),
	.w7(32'hb982821e),
	.w8(32'hbb87a300),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdf2a1),
	.w1(32'h3b4dbb1c),
	.w2(32'h3ba29dcc),
	.w3(32'hbb0a8afe),
	.w4(32'h3b2c0b32),
	.w5(32'hbb922633),
	.w6(32'hbbaa58a9),
	.w7(32'h3b3563b7),
	.w8(32'h3b917b2a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c107424),
	.w1(32'hba78bfb6),
	.w2(32'hbb8458a8),
	.w3(32'hbb84559a),
	.w4(32'hbaad2613),
	.w5(32'h3b0e420d),
	.w6(32'hbbb481ac),
	.w7(32'hbb8f6a3f),
	.w8(32'h3b91b568),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896262),
	.w1(32'hbaa79ac4),
	.w2(32'hbb85bafe),
	.w3(32'hbad58ef5),
	.w4(32'hbad21b6b),
	.w5(32'hbb627cfa),
	.w6(32'h3bed4a31),
	.w7(32'h3b2e3283),
	.w8(32'hbb4af697),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5fc2f),
	.w1(32'hbbbd29e9),
	.w2(32'h3b3e4328),
	.w3(32'hbb25b74d),
	.w4(32'hba95b511),
	.w5(32'hbb4c15af),
	.w6(32'hbc0b8e74),
	.w7(32'hbbb95c9f),
	.w8(32'hbbd7dcbd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e50ec),
	.w1(32'hbc157b25),
	.w2(32'hbb87fb94),
	.w3(32'h3b8eb6d5),
	.w4(32'hba71c554),
	.w5(32'h3b01933f),
	.w6(32'h3b284430),
	.w7(32'h3b6f8575),
	.w8(32'h3a8a3702),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1618c2),
	.w1(32'hb9983244),
	.w2(32'hba9359dd),
	.w3(32'h377bb978),
	.w4(32'hbab89604),
	.w5(32'hbadac20c),
	.w6(32'h3aa42d4b),
	.w7(32'h3a9f3c69),
	.w8(32'hbb04e049),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ced7e),
	.w1(32'hbbc0987c),
	.w2(32'hbb994291),
	.w3(32'hbbe87004),
	.w4(32'hbb584b99),
	.w5(32'h3ad4dad8),
	.w6(32'hbb3eb2b8),
	.w7(32'hbb0ce53a),
	.w8(32'h3b6b0aff),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd05d),
	.w1(32'h3b83c08a),
	.w2(32'h3b5335af),
	.w3(32'hbaafcf34),
	.w4(32'hbb1cc89c),
	.w5(32'h3a6c4d77),
	.w6(32'h3bc7459a),
	.w7(32'h3b1b40bc),
	.w8(32'hbb95a4e5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ebff2),
	.w1(32'hbbb0b3f3),
	.w2(32'h3b8f5f74),
	.w3(32'hba249cff),
	.w4(32'h3a8bcb38),
	.w5(32'hba61f195),
	.w6(32'hbbcad412),
	.w7(32'h3964a12f),
	.w8(32'hbb1d3e52),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad631e),
	.w1(32'h3ae66324),
	.w2(32'h3b28144a),
	.w3(32'hbb67cf6e),
	.w4(32'h3b6a2f78),
	.w5(32'hbb56cd5d),
	.w6(32'hbbf78fd3),
	.w7(32'hbaaf4d5f),
	.w8(32'hbbd968bc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7052d1),
	.w1(32'h3c31b94e),
	.w2(32'hbb88760b),
	.w3(32'hbb39684f),
	.w4(32'hbbd8dd25),
	.w5(32'h3ab6c048),
	.w6(32'hbb2a7f7d),
	.w7(32'hbbe4a380),
	.w8(32'hbc5d7991),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ac51c),
	.w1(32'hbc31514b),
	.w2(32'hbadc2549),
	.w3(32'hbb97965f),
	.w4(32'hbb5a5c42),
	.w5(32'h3b131326),
	.w6(32'hbc08d372),
	.w7(32'hbb349116),
	.w8(32'hbbca31c0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99c67b),
	.w1(32'hbb7ca0fc),
	.w2(32'hbb2e7038),
	.w3(32'h3a7f2e7f),
	.w4(32'h3b7cb515),
	.w5(32'hbba7d640),
	.w6(32'h3b252032),
	.w7(32'hbb160e50),
	.w8(32'hb8bac6bd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b159f55),
	.w1(32'h3affe38c),
	.w2(32'h3abb75b2),
	.w3(32'hbb67d7be),
	.w4(32'hbb96e98b),
	.w5(32'hbabf0591),
	.w6(32'hbb517127),
	.w7(32'hbba3d0d3),
	.w8(32'hbaa54a63),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad67a81),
	.w1(32'hba0f4c7c),
	.w2(32'h393ea012),
	.w3(32'hbb2e10f0),
	.w4(32'hbb2f1ccd),
	.w5(32'h3b43237a),
	.w6(32'hbb04caea),
	.w7(32'hba9a29be),
	.w8(32'hb9c319ab),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71bf19),
	.w1(32'h3ad6ac3c),
	.w2(32'h3b58e33d),
	.w3(32'h3b50702c),
	.w4(32'h3b5f5e5e),
	.w5(32'hbbb5a87e),
	.w6(32'h3b2dadef),
	.w7(32'h3bc8135d),
	.w8(32'h3a31027d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ad724),
	.w1(32'hb782ba58),
	.w2(32'hbb817ee9),
	.w3(32'hbaa0b9ae),
	.w4(32'hbadc479a),
	.w5(32'hbb4eae28),
	.w6(32'h3aa8f488),
	.w7(32'hbaa8c224),
	.w8(32'h39dbada5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cc865),
	.w1(32'hbb91f96b),
	.w2(32'hba53f610),
	.w3(32'h37667904),
	.w4(32'hb9818ec3),
	.w5(32'h3c0a500e),
	.w6(32'hbb8b568a),
	.w7(32'hba012820),
	.w8(32'h3c2ee36d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb803cd9a),
	.w1(32'h3b66b022),
	.w2(32'h3ba3e758),
	.w3(32'h3a22268f),
	.w4(32'hbaa0cc5c),
	.w5(32'hbb932883),
	.w6(32'h3acd5520),
	.w7(32'h3bf359f4),
	.w8(32'hbb1bc604),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1787a),
	.w1(32'hbb1147d2),
	.w2(32'hbac09711),
	.w3(32'hbbfb90f7),
	.w4(32'hb9ca4b80),
	.w5(32'hbb9d5338),
	.w6(32'hbc15f2e4),
	.w7(32'hbb02036e),
	.w8(32'hb8a4fdbc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7e550),
	.w1(32'hbbeeeb02),
	.w2(32'hbba6fa40),
	.w3(32'hbb58e159),
	.w4(32'h3a75499b),
	.w5(32'hba1da02d),
	.w6(32'h3a8bd87a),
	.w7(32'h3b0694eb),
	.w8(32'h3a3cc4f1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9090af),
	.w1(32'hbb09497f),
	.w2(32'hbabb7f58),
	.w3(32'hb9dc0d83),
	.w4(32'h3a0915a0),
	.w5(32'h3be582c2),
	.w6(32'h399f5fa8),
	.w7(32'hbab6f0da),
	.w8(32'hbc2f3dac),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e33b9),
	.w1(32'hbb94ccda),
	.w2(32'hb9d1adae),
	.w3(32'hbc4c10e0),
	.w4(32'h3bb0551d),
	.w5(32'h3ba361f6),
	.w6(32'h3c3121ff),
	.w7(32'h3b5cc6a8),
	.w8(32'h3bf9c4a2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45bf90),
	.w1(32'hbc89f9df),
	.w2(32'hbc29dc95),
	.w3(32'hbc78aa41),
	.w4(32'h3aa9f733),
	.w5(32'h3ba5568a),
	.w6(32'h3cf00b7b),
	.w7(32'h3b94f39c),
	.w8(32'hbb3bd824),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2e063),
	.w1(32'hba06dec2),
	.w2(32'hbb39633c),
	.w3(32'h3bef368e),
	.w4(32'hba721f1a),
	.w5(32'hbb5eee3d),
	.w6(32'h3b3472cf),
	.w7(32'h3b3ae994),
	.w8(32'hbb1661ed),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04f60c),
	.w1(32'hbb4b574f),
	.w2(32'hbb08cd9f),
	.w3(32'h3c12ec2f),
	.w4(32'h3b56d67f),
	.w5(32'hba3c197c),
	.w6(32'h39fc94a4),
	.w7(32'h3b666064),
	.w8(32'h3b706a57),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981ffe),
	.w1(32'hbb9b25c5),
	.w2(32'hbb4995ad),
	.w3(32'hbaf13f88),
	.w4(32'hbb913f14),
	.w5(32'hbaf56206),
	.w6(32'h3b878552),
	.w7(32'h3ac44f81),
	.w8(32'hb9ef5cc5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc256238),
	.w1(32'hbb30c6b3),
	.w2(32'h3b95f8ae),
	.w3(32'h3a68c24e),
	.w4(32'hbaaa2984),
	.w5(32'hb9104d04),
	.w6(32'hba457924),
	.w7(32'h3ad19467),
	.w8(32'h3a39bd07),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeacd0),
	.w1(32'hbc09c482),
	.w2(32'hbb264f18),
	.w3(32'hbbe8339e),
	.w4(32'hbbc4ceb9),
	.w5(32'h3b80584b),
	.w6(32'hbb3723c7),
	.w7(32'hb9f02cef),
	.w8(32'h3be913af),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0715cd),
	.w1(32'hb99cbddd),
	.w2(32'h3b47edee),
	.w3(32'hbaf3e2b6),
	.w4(32'hbac7f0f6),
	.w5(32'h3bb6b2f3),
	.w6(32'h3be2d238),
	.w7(32'h3b759089),
	.w8(32'h3b2f957c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba191183),
	.w1(32'hbc16713b),
	.w2(32'h3baf8263),
	.w3(32'h3c105261),
	.w4(32'h3b76bbd2),
	.w5(32'hbc37ad73),
	.w6(32'h3bfd6bc8),
	.w7(32'h3c1668db),
	.w8(32'hbbdf626e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a704),
	.w1(32'h3bca61c1),
	.w2(32'h3a77e5b4),
	.w3(32'hbc644660),
	.w4(32'hbbe63bd2),
	.w5(32'h3b7e360e),
	.w6(32'hbc0e1d0f),
	.w7(32'hbbae2fe2),
	.w8(32'h3b2ada91),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a6a2),
	.w1(32'hbba1100a),
	.w2(32'hbb2434bc),
	.w3(32'h3a9df645),
	.w4(32'hb80d4ef4),
	.w5(32'hbbdd8200),
	.w6(32'hb9da108f),
	.w7(32'hbb134a20),
	.w8(32'hbb9dde8f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05a6c4),
	.w1(32'h3b8df8b2),
	.w2(32'h3c2b60a5),
	.w3(32'hbb74e07d),
	.w4(32'h3b0e1b5c),
	.w5(32'h3a098569),
	.w6(32'hbb612f4d),
	.w7(32'h3b628b62),
	.w8(32'h3b056d37),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684c01),
	.w1(32'h3beef3f8),
	.w2(32'h3bfb1dce),
	.w3(32'h3bd0d171),
	.w4(32'h3ae1eff0),
	.w5(32'hbaf00960),
	.w6(32'h3b424542),
	.w7(32'h3baa9d94),
	.w8(32'hbb6829b6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515e62),
	.w1(32'hbaafafa1),
	.w2(32'h3b1361d0),
	.w3(32'hbb78d2fc),
	.w4(32'hbb501134),
	.w5(32'hbb94bf09),
	.w6(32'hbb35f219),
	.w7(32'hbab8c375),
	.w8(32'h3b9a79af),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60c9be),
	.w1(32'hbc1d6ba1),
	.w2(32'hbb6cefe5),
	.w3(32'hbb82d0a3),
	.w4(32'h3899b673),
	.w5(32'hbacc012a),
	.w6(32'hbb072f33),
	.w7(32'hba87da4b),
	.w8(32'hbbdd753f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0a50e),
	.w1(32'h3b97a7ef),
	.w2(32'hbb12e920),
	.w3(32'h3ac42d5f),
	.w4(32'h3c11b6b9),
	.w5(32'hbb2c72ae),
	.w6(32'hbb589a17),
	.w7(32'h3b097c93),
	.w8(32'hbbb663c9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b72975),
	.w1(32'h3a5d4bcd),
	.w2(32'h3a68e004),
	.w3(32'hba730b78),
	.w4(32'hbb88ef2d),
	.w5(32'h3bb4e8ad),
	.w6(32'hbb1c0d72),
	.w7(32'hb79ad895),
	.w8(32'h3a5c7cd8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d053c),
	.w1(32'hbb94f356),
	.w2(32'h3ae71fa1),
	.w3(32'h3c0f30ac),
	.w4(32'h3bc4776c),
	.w5(32'hbbfbcd42),
	.w6(32'h3b3f1f4d),
	.w7(32'h3bac4a38),
	.w8(32'hbafd3ddf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1009),
	.w1(32'hb94b1f80),
	.w2(32'h3aa63d00),
	.w3(32'hba582cd4),
	.w4(32'hbbbf8d3a),
	.w5(32'hbb3e637b),
	.w6(32'h3c30cf94),
	.w7(32'hbbe5c76a),
	.w8(32'hb980806c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5a74b),
	.w1(32'hbbe888aa),
	.w2(32'h3c05ec21),
	.w3(32'h3bc9c03b),
	.w4(32'h3a6ca908),
	.w5(32'hbbb6b999),
	.w6(32'hbbaacae5),
	.w7(32'h3c6ad8aa),
	.w8(32'hbbbb6875),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c3d9),
	.w1(32'h3abb20a2),
	.w2(32'hbb159620),
	.w3(32'hbba5b643),
	.w4(32'hbbda8ce9),
	.w5(32'hbbadc4d7),
	.w6(32'hbb2c105b),
	.w7(32'hbba5bc0e),
	.w8(32'hbb9c73f3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231529),
	.w1(32'h3b87ad91),
	.w2(32'h3a9784d4),
	.w3(32'h3b571211),
	.w4(32'hbb28e421),
	.w5(32'hbafaa05d),
	.w6(32'hbb4667a5),
	.w7(32'h3b557b40),
	.w8(32'h3a3ee08a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa445a3),
	.w1(32'hbbba1451),
	.w2(32'hbbbd88ca),
	.w3(32'hbb820896),
	.w4(32'hbb5c14ba),
	.w5(32'hba67590b),
	.w6(32'hbb01a74f),
	.w7(32'h39af1e4e),
	.w8(32'hbbf423f9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9a825),
	.w1(32'hbb64e5e8),
	.w2(32'hbc37cfa9),
	.w3(32'h3bd407c7),
	.w4(32'hbb0ed5dc),
	.w5(32'hbbd435bc),
	.w6(32'h3c25a233),
	.w7(32'h3bbad6c2),
	.w8(32'hbba6d714),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc180e7),
	.w1(32'hbbb8ba5b),
	.w2(32'hbc50d180),
	.w3(32'hbb51937c),
	.w4(32'hb9b35b67),
	.w5(32'hbae635bf),
	.w6(32'hb9f28b03),
	.w7(32'hbb0c027a),
	.w8(32'h37bf2523),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5519),
	.w1(32'h3b6658ae),
	.w2(32'h3b9d7031),
	.w3(32'hbb3b60ca),
	.w4(32'h3aacdb44),
	.w5(32'h3a7d4600),
	.w6(32'hba4877a6),
	.w7(32'h397734e3),
	.w8(32'h3b314bbb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119bc1),
	.w1(32'hbb7ab3a8),
	.w2(32'h3bb5da19),
	.w3(32'h3c0de84b),
	.w4(32'hbaf4863c),
	.w5(32'hbb403196),
	.w6(32'h3a527d05),
	.w7(32'hba80fa5f),
	.w8(32'h398994df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084b43),
	.w1(32'hbb116110),
	.w2(32'hbbec0a01),
	.w3(32'h3b9b4d3d),
	.w4(32'h3a393df9),
	.w5(32'hb96db0c0),
	.w6(32'hbb105dda),
	.w7(32'h3b32eb16),
	.w8(32'h3b939160),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e023cb),
	.w1(32'hbb3ac61a),
	.w2(32'hbc46cea8),
	.w3(32'h3a54eeaa),
	.w4(32'hbbbbe001),
	.w5(32'h3b05d3c0),
	.w6(32'h3bf58ea5),
	.w7(32'h3ae94b79),
	.w8(32'h3ca454b9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75b0bf),
	.w1(32'h3c310655),
	.w2(32'hbc495be6),
	.w3(32'h3c34685c),
	.w4(32'h3b86454e),
	.w5(32'h3a351ed9),
	.w6(32'h3b581728),
	.w7(32'hbbfb4857),
	.w8(32'h3c82f0c4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3c06),
	.w1(32'hba5243fe),
	.w2(32'hbb30fb97),
	.w3(32'h3beb0b03),
	.w4(32'hb920ddd8),
	.w5(32'h3ba90749),
	.w6(32'h3c4930fb),
	.w7(32'h3bcd4015),
	.w8(32'h3b661c3f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13448d),
	.w1(32'hbb1731be),
	.w2(32'hbbf57ee9),
	.w3(32'h3ae7e9cb),
	.w4(32'hbbee037a),
	.w5(32'hbc81b86e),
	.w6(32'h3c0d4298),
	.w7(32'h39412fe3),
	.w8(32'hbc81f4c0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d3e41),
	.w1(32'h3bbc34f3),
	.w2(32'h3c9ec10c),
	.w3(32'h3b5d7a41),
	.w4(32'h3c7d4286),
	.w5(32'h3be9abcf),
	.w6(32'h3b8efe2a),
	.w7(32'h3ce8aad7),
	.w8(32'h3c5f5240),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ecaf6),
	.w1(32'hbb8ccf61),
	.w2(32'hbbac2d4a),
	.w3(32'hbbc6226e),
	.w4(32'hbbda79ab),
	.w5(32'h3abe0238),
	.w6(32'h3b6f41de),
	.w7(32'hbc1db133),
	.w8(32'h3aef1f65),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e524c),
	.w1(32'hba85158c),
	.w2(32'hbbcace46),
	.w3(32'h3b27876b),
	.w4(32'h3a89f41e),
	.w5(32'hbb649145),
	.w6(32'hb8274e21),
	.w7(32'hbb44c82a),
	.w8(32'h3b3ec34b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3812),
	.w1(32'hbc3aa5de),
	.w2(32'hbb8cfa27),
	.w3(32'hbc284004),
	.w4(32'hbb32691d),
	.w5(32'h3c1168c3),
	.w6(32'hbc11134f),
	.w7(32'hbc3d505f),
	.w8(32'h3c26ab49),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf22a7c),
	.w1(32'hbb2067ff),
	.w2(32'hbbefd7d9),
	.w3(32'hbad57985),
	.w4(32'hbb827a5f),
	.w5(32'h3b906e71),
	.w6(32'hba361765),
	.w7(32'hbbe139bb),
	.w8(32'h3bfd667e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac92d1f),
	.w1(32'hbba4cbad),
	.w2(32'hbb83de35),
	.w3(32'hbb048333),
	.w4(32'hbbdbbeea),
	.w5(32'hb98db388),
	.w6(32'hbbc71d37),
	.w7(32'hbbce096b),
	.w8(32'h3a8d8961),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb867498),
	.w1(32'hbbbb04ab),
	.w2(32'hbb0b81bd),
	.w3(32'hba7e8841),
	.w4(32'hbabd51ef),
	.w5(32'hbaefdaa0),
	.w6(32'hbb99f477),
	.w7(32'hbb2323bd),
	.w8(32'h3ab87f7a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a823875),
	.w1(32'h3a2825af),
	.w2(32'hbbba5e49),
	.w3(32'h3bd5e175),
	.w4(32'h3b47c223),
	.w5(32'h3b45a1fd),
	.w6(32'h3bdf26d3),
	.w7(32'hbb13a3d4),
	.w8(32'h3a093e5a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58d7ea),
	.w1(32'hbb49c223),
	.w2(32'hbba93da0),
	.w3(32'h39878e3f),
	.w4(32'hba48b10c),
	.w5(32'hbbc01be5),
	.w6(32'h3c3c0f40),
	.w7(32'hb9e25e86),
	.w8(32'hbbccb26f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe8297),
	.w1(32'hbc021464),
	.w2(32'hbc0d8e80),
	.w3(32'hbb265e04),
	.w4(32'hbbf702cd),
	.w5(32'hbbd949f8),
	.w6(32'hbbdd368c),
	.w7(32'hbc2d8ec3),
	.w8(32'hb8d349e1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fbdf6),
	.w1(32'hbb97f11f),
	.w2(32'hbb1180e3),
	.w3(32'hbc0818cc),
	.w4(32'hbc26493e),
	.w5(32'h3acdc8b5),
	.w6(32'hbba00487),
	.w7(32'hbb7ee354),
	.w8(32'h3c373fbf),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b2faf),
	.w1(32'h3c53863d),
	.w2(32'hbb67c8c2),
	.w3(32'hbb39b54c),
	.w4(32'hbb1c45fd),
	.w5(32'hba35ccc9),
	.w6(32'h3c329d2b),
	.w7(32'hbb880b16),
	.w8(32'hbba71609),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9559c0e),
	.w1(32'h3b6ab5eb),
	.w2(32'hbb8f1a5d),
	.w3(32'h3b833c68),
	.w4(32'h3bb41799),
	.w5(32'hbadee571),
	.w6(32'h3bce44fc),
	.w7(32'h3b577fda),
	.w8(32'hbad8273f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dca3a9),
	.w1(32'hbb5fbdbf),
	.w2(32'hbbb2958e),
	.w3(32'hbb5fdc26),
	.w4(32'hbbb1f548),
	.w5(32'h3ab14395),
	.w6(32'hbbc68006),
	.w7(32'hbbd9ef22),
	.w8(32'h3c2be080),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06aa8f),
	.w1(32'h3b8ef538),
	.w2(32'hbc0b4f86),
	.w3(32'hbbf8042f),
	.w4(32'h3b2d55dc),
	.w5(32'h396dfd3d),
	.w6(32'hbbcb1a9e),
	.w7(32'hbc4e4097),
	.w8(32'h3aceecd5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910a766),
	.w1(32'h3a574006),
	.w2(32'h3b020dc8),
	.w3(32'h3b1acff7),
	.w4(32'h3a4b0225),
	.w5(32'hbc24eb4e),
	.w6(32'hbaf9e340),
	.w7(32'h3b18e031),
	.w8(32'hbbf22b79),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b7f65),
	.w1(32'hbb8e1b72),
	.w2(32'hba2e9876),
	.w3(32'hbbafed2f),
	.w4(32'h3bb872d0),
	.w5(32'h3bd163fb),
	.w6(32'hbc587f18),
	.w7(32'hbb02343a),
	.w8(32'hbb2afce9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9389d55),
	.w1(32'hbb9749bc),
	.w2(32'hba52c0ad),
	.w3(32'h3a54ebce),
	.w4(32'hbb966b75),
	.w5(32'h3ab78bb3),
	.w6(32'hbba5680b),
	.w7(32'h3a1b0d9f),
	.w8(32'hbb625cf0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc839),
	.w1(32'hbbaf9fb5),
	.w2(32'h3a4a7f91),
	.w3(32'hbae909cd),
	.w4(32'h3944c2de),
	.w5(32'hbb945171),
	.w6(32'h39babf90),
	.w7(32'h3c316cba),
	.w8(32'hbbd8ace8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe376aa),
	.w1(32'hbb7f3320),
	.w2(32'hbb20ed24),
	.w3(32'h3beaea68),
	.w4(32'h3bca4c75),
	.w5(32'hbb61441d),
	.w6(32'h3b64c3b6),
	.w7(32'h3b4582d2),
	.w8(32'hbbb2bf13),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959240e),
	.w1(32'hbba2dd9c),
	.w2(32'hb8a628f2),
	.w3(32'hbb03be93),
	.w4(32'hba27f3bd),
	.w5(32'hbb622747),
	.w6(32'hbb3fc804),
	.w7(32'hbac14f6d),
	.w8(32'hbc09a9fb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc41eb),
	.w1(32'h3ac3d1e7),
	.w2(32'hbaf03902),
	.w3(32'hbb5f8e5b),
	.w4(32'hbb5c305c),
	.w5(32'hbac48309),
	.w6(32'h3bf0cd7a),
	.w7(32'h3be19224),
	.w8(32'hbb48701c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba335),
	.w1(32'hbbeba86e),
	.w2(32'hbba05389),
	.w3(32'hbb6bad4f),
	.w4(32'h3a540260),
	.w5(32'h3b837cf1),
	.w6(32'h3ab6d015),
	.w7(32'hbb416c86),
	.w8(32'h3bc07999),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81f486),
	.w1(32'hbb753130),
	.w2(32'hbbaecc1d),
	.w3(32'hbb0f6861),
	.w4(32'hbbde182e),
	.w5(32'h3ab3c0e7),
	.w6(32'hbb0216e6),
	.w7(32'hbb925469),
	.w8(32'h3bd33ff1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a940005),
	.w1(32'hbb312823),
	.w2(32'h39ff1e21),
	.w3(32'hbb87db53),
	.w4(32'hbaaf3684),
	.w5(32'hbbfc1a53),
	.w6(32'h3bece3ad),
	.w7(32'hbb13eed6),
	.w8(32'hbbc96c8e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2908df),
	.w1(32'hbc1900d7),
	.w2(32'hbbff943a),
	.w3(32'hbb2a1590),
	.w4(32'hbbefe78b),
	.w5(32'h3b5b6710),
	.w6(32'h3ab4e3c1),
	.w7(32'hbac7ed8e),
	.w8(32'h3b137605),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab88a92),
	.w1(32'hba5e2123),
	.w2(32'hbb842d5b),
	.w3(32'hbb54b123),
	.w4(32'hbb80dd31),
	.w5(32'hbae9a7c1),
	.w6(32'h3b25bae1),
	.w7(32'hbc039a37),
	.w8(32'hbb6bf793),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7ee9),
	.w1(32'h3b97e445),
	.w2(32'hbb9a5905),
	.w3(32'hbb124d28),
	.w4(32'h39650a15),
	.w5(32'h3ae053d8),
	.w6(32'hb9977a79),
	.w7(32'hbaa10c03),
	.w8(32'h3bb49ee0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e2fa9),
	.w1(32'hbb0b50ee),
	.w2(32'hbb865498),
	.w3(32'hbb1d5545),
	.w4(32'hbb391b06),
	.w5(32'hbc41d99f),
	.w6(32'hbb5e040a),
	.w7(32'hbb0920b0),
	.w8(32'hbc0b27bd),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61c78c),
	.w1(32'h3b90751e),
	.w2(32'h3bbc8732),
	.w3(32'hb808e870),
	.w4(32'h3a0f1f73),
	.w5(32'h3b05fe1d),
	.w6(32'h3ba9dfd8),
	.w7(32'h3c0a2da7),
	.w8(32'h3b28c9f6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab01f8c),
	.w1(32'hbb88ec74),
	.w2(32'hbbb9d883),
	.w3(32'h3a61e15c),
	.w4(32'hbb6cba83),
	.w5(32'hbb112672),
	.w6(32'hbb35c444),
	.w7(32'hbb36f84f),
	.w8(32'hb9910072),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b794),
	.w1(32'hbb5d7b32),
	.w2(32'hbc0ac8e9),
	.w3(32'hbc026e9d),
	.w4(32'hbc3c18a3),
	.w5(32'hbb8153e0),
	.w6(32'hbb2c9e13),
	.w7(32'hbb9676d0),
	.w8(32'h3b453820),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf04b84),
	.w1(32'hbc21747b),
	.w2(32'hbba37ab1),
	.w3(32'h3b15fa8f),
	.w4(32'hbb1fcc89),
	.w5(32'hba0f9e9e),
	.w6(32'hbb0682be),
	.w7(32'hba16e932),
	.w8(32'hba931300),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88d959),
	.w1(32'hbbfb0082),
	.w2(32'hbbf08e2d),
	.w3(32'hbb9a4113),
	.w4(32'hbc183f4e),
	.w5(32'h39f8a950),
	.w6(32'hbbc64a1b),
	.w7(32'hbbb972f3),
	.w8(32'h3b591a83),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9ee81),
	.w1(32'hbbc02452),
	.w2(32'hbb8addf5),
	.w3(32'h3a629de0),
	.w4(32'hbaa77e45),
	.w5(32'h3a9498a6),
	.w6(32'hb96aaea1),
	.w7(32'h3a75bcd7),
	.w8(32'h3b1feca3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8175e7),
	.w1(32'hbbb08866),
	.w2(32'hbbd06009),
	.w3(32'hbb35396c),
	.w4(32'hbbb37f06),
	.w5(32'h3acf1b3f),
	.w6(32'hbba5e3c1),
	.w7(32'hbb510fd1),
	.w8(32'h3bc1f87a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d34fc4),
	.w1(32'hbbcdec71),
	.w2(32'hba7e4517),
	.w3(32'h3a85ac6c),
	.w4(32'hbc02d32d),
	.w5(32'hbb8b56f7),
	.w6(32'hbb8c90b8),
	.w7(32'hbb61c5f0),
	.w8(32'hbc1e49ab),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50d14a),
	.w1(32'hbbf4f275),
	.w2(32'h3b260f92),
	.w3(32'hbb6f7d0b),
	.w4(32'h3ae2ddec),
	.w5(32'hb993fe74),
	.w6(32'hbba19e1d),
	.w7(32'h3bd66f12),
	.w8(32'h39e5d78f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b0e9),
	.w1(32'hbbeacea6),
	.w2(32'hba992e9a),
	.w3(32'hbb5bae17),
	.w4(32'hbaedfd70),
	.w5(32'h3b64400e),
	.w6(32'h3c2d99ad),
	.w7(32'h3b3d5675),
	.w8(32'h3b7b3eca),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baacbc6),
	.w1(32'h3b228676),
	.w2(32'hbbdf8124),
	.w3(32'h3c0501be),
	.w4(32'h3b93c5a0),
	.w5(32'hbbee44f3),
	.w6(32'h3bd5872f),
	.w7(32'h3a6befc8),
	.w8(32'hbb68501e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64396c),
	.w1(32'hbbbf4235),
	.w2(32'hbb8a4713),
	.w3(32'hbabfacb9),
	.w4(32'hbb879238),
	.w5(32'h3c16ef1b),
	.w6(32'h3a08745b),
	.w7(32'hbb5d4b02),
	.w8(32'h3c4cb54b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf28899),
	.w1(32'hb83026a7),
	.w2(32'hbbec66cc),
	.w3(32'h3a1e91ca),
	.w4(32'hbb926009),
	.w5(32'hbc0b9ff1),
	.w6(32'h3aa5b1ea),
	.w7(32'hbc3a9fab),
	.w8(32'hbc213769),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fca17),
	.w1(32'hbba84cdc),
	.w2(32'hba505254),
	.w3(32'hbba987bf),
	.w4(32'h3b088bdc),
	.w5(32'hbc06f880),
	.w6(32'hbc27c758),
	.w7(32'h3bad62c8),
	.w8(32'hbab1d9fa),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c52ac),
	.w1(32'h3a53290d),
	.w2(32'hbaa73a90),
	.w3(32'h3c18c279),
	.w4(32'h3b9e1154),
	.w5(32'h3a55bd6a),
	.w6(32'h3c0e374f),
	.w7(32'h3bab8ee9),
	.w8(32'hbbb24dc0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77a39d),
	.w1(32'hbc6c24ac),
	.w2(32'hbc0ac11a),
	.w3(32'hbc393ef7),
	.w4(32'hbc061694),
	.w5(32'hb9acea08),
	.w6(32'h3baaa6ab),
	.w7(32'hbb8d2a38),
	.w8(32'h3adcae21),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ece36),
	.w1(32'hbbbebd41),
	.w2(32'hbb8b0c53),
	.w3(32'hbba1e6fe),
	.w4(32'hbb6d15fe),
	.w5(32'h3b8f2f68),
	.w6(32'h3b0b2ef2),
	.w7(32'h399fa7bc),
	.w8(32'h3b68a742),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2a925),
	.w1(32'hbb973889),
	.w2(32'hbbba38c6),
	.w3(32'hbb4e42cb),
	.w4(32'hbc19855b),
	.w5(32'h3a93d3b9),
	.w6(32'hbbd3ea5b),
	.w7(32'hbbd8d41c),
	.w8(32'h3a68e05e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb36858),
	.w1(32'h38b0e516),
	.w2(32'hbaca24c8),
	.w3(32'hbac1b858),
	.w4(32'hbb9d7562),
	.w5(32'hbba1c30a),
	.w6(32'h3bdb1462),
	.w7(32'h3b8ad802),
	.w8(32'hbb87d7b6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d3372),
	.w1(32'hbc942a29),
	.w2(32'hbb5dfe0f),
	.w3(32'hbc67dad1),
	.w4(32'hbc054420),
	.w5(32'hbbae156a),
	.w6(32'hbbe9569d),
	.w7(32'h3b48abda),
	.w8(32'hbb69a1d6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082d2c),
	.w1(32'hbbb3758b),
	.w2(32'hbbaec736),
	.w3(32'hbad79773),
	.w4(32'h3b50706f),
	.w5(32'h3b88fc06),
	.w6(32'hbbebee20),
	.w7(32'h390dfa31),
	.w8(32'h3c67db55),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55a4e0),
	.w1(32'h3bd87db1),
	.w2(32'hbc26c2ae),
	.w3(32'h3c3daf2d),
	.w4(32'h3a9a00ca),
	.w5(32'h3b921954),
	.w6(32'h3bbd1662),
	.w7(32'hbbcbeed9),
	.w8(32'h3c465bdd),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a7f81),
	.w1(32'hbb561466),
	.w2(32'hbba85e3b),
	.w3(32'hba84f60c),
	.w4(32'hbbc195b4),
	.w5(32'hbb90b6a2),
	.w6(32'hbb464de6),
	.w7(32'hbc32c731),
	.w8(32'hbb9cd96d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdba6e7),
	.w1(32'hbbecf99f),
	.w2(32'hbb287a5e),
	.w3(32'hbbb4572a),
	.w4(32'hbb68844d),
	.w5(32'h3b41590a),
	.w6(32'hbc14801a),
	.w7(32'hbbd315ed),
	.w8(32'h3bc1821e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026895),
	.w1(32'h3b34eac2),
	.w2(32'hbc20c621),
	.w3(32'h3be35ebf),
	.w4(32'h3c2a91e3),
	.w5(32'h3b2519ed),
	.w6(32'h3c88baab),
	.w7(32'h3c0aa64b),
	.w8(32'h3bc0194c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b693a13),
	.w1(32'h3b968a9c),
	.w2(32'hbad745e9),
	.w3(32'h3b7721e0),
	.w4(32'h3b4212e9),
	.w5(32'h3b12e96d),
	.w6(32'h3bdd2e99),
	.w7(32'h3b00f46f),
	.w8(32'h3bb3ef6b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399976b1),
	.w1(32'hbaa818cf),
	.w2(32'hbb2b4aef),
	.w3(32'h3b7a29b1),
	.w4(32'hbab5efcb),
	.w5(32'hbbba7276),
	.w6(32'hb9880af2),
	.w7(32'hbb4456ac),
	.w8(32'h3c31d1af),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb4b7),
	.w1(32'h3ba9e3bd),
	.w2(32'hb9015f99),
	.w3(32'hbbf918fe),
	.w4(32'hbb8e1012),
	.w5(32'h3aa324bd),
	.w6(32'h3958eeab),
	.w7(32'hbbdbeae1),
	.w8(32'h3c8ce44c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85322e),
	.w1(32'hbb3cd099),
	.w2(32'hbb2af6b6),
	.w3(32'h3c4da0a6),
	.w4(32'hbc0f11be),
	.w5(32'hbc18f455),
	.w6(32'h3c470f27),
	.w7(32'hbc14ec4e),
	.w8(32'hbc0edd33),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8eab2),
	.w1(32'hbba4533b),
	.w2(32'hbbbd88ac),
	.w3(32'hbbdc620e),
	.w4(32'hba2685cd),
	.w5(32'hbb139230),
	.w6(32'hbc3d4431),
	.w7(32'h3abc0b54),
	.w8(32'h3b073162),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09ff92),
	.w1(32'h3ac63f0b),
	.w2(32'h39cba84d),
	.w3(32'hbb81306e),
	.w4(32'hbaa10af5),
	.w5(32'hbb3c89f9),
	.w6(32'h3b4f1b75),
	.w7(32'h35c92b1d),
	.w8(32'h38e2f6af),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a945ee5),
	.w1(32'h3b86d087),
	.w2(32'hb9e3e4ab),
	.w3(32'h3964c026),
	.w4(32'hb99b5dee),
	.w5(32'h3a7ead8b),
	.w6(32'h3b403d71),
	.w7(32'h38e184b1),
	.w8(32'h3c1ae9fb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1361d3),
	.w1(32'hbaede72e),
	.w2(32'hbbb6524a),
	.w3(32'hbbb00956),
	.w4(32'h3b9a3222),
	.w5(32'h3bb11706),
	.w6(32'hbc177216),
	.w7(32'hbc1cc533),
	.w8(32'h3bcef384),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b366ece),
	.w1(32'h3b186e06),
	.w2(32'hbae642ea),
	.w3(32'h3b8b6680),
	.w4(32'hbad58e24),
	.w5(32'hbb1c6e62),
	.w6(32'h3a8175b6),
	.w7(32'hbb112469),
	.w8(32'hbbb7c595),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61e8e),
	.w1(32'h3b947047),
	.w2(32'h3b68b627),
	.w3(32'hba8a419b),
	.w4(32'hbb162c4d),
	.w5(32'hbc0f969f),
	.w6(32'h3ab4a313),
	.w7(32'h3b9fa37a),
	.w8(32'hbc011a74),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd99e05),
	.w1(32'h3b3b0f78),
	.w2(32'h3b9c44f6),
	.w3(32'h3a814ad6),
	.w4(32'hbb0d13d7),
	.w5(32'hbb054395),
	.w6(32'h3b408a03),
	.w7(32'h3bf61bcd),
	.w8(32'hbbe11876),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6929c),
	.w1(32'hba906311),
	.w2(32'hba6e5758),
	.w3(32'hbb93b9cd),
	.w4(32'hba55d4cf),
	.w5(32'h3b2b9f91),
	.w6(32'h3b5124d7),
	.w7(32'h3ae86c8c),
	.w8(32'h3c1c016f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3b6d4),
	.w1(32'h3ab5740b),
	.w2(32'hbbd7643e),
	.w3(32'hba97689f),
	.w4(32'hbbd5e1e2),
	.w5(32'hbb5412c9),
	.w6(32'hbbbcd366),
	.w7(32'hbc18c992),
	.w8(32'hbabfed72),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3495ff37),
	.w1(32'hbc04a9bc),
	.w2(32'hbba06c26),
	.w3(32'hbbea2a9b),
	.w4(32'hba84fba4),
	.w5(32'h3c88c273),
	.w6(32'hbbcb6f9f),
	.w7(32'hbbce7ecd),
	.w8(32'h3cf4254d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fdbfa),
	.w1(32'h3b821607),
	.w2(32'hbca6bd50),
	.w3(32'hbb737b8f),
	.w4(32'hbc0bb91a),
	.w5(32'hbb7c8e56),
	.w6(32'h3c002b8b),
	.w7(32'hbcb82da9),
	.w8(32'h3bca1d72),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58567),
	.w1(32'hbc4c567b),
	.w2(32'hbc3147f2),
	.w3(32'hbc074240),
	.w4(32'hbbc8740d),
	.w5(32'h3b0aefb0),
	.w6(32'hbbf1991f),
	.w7(32'hbab5e310),
	.w8(32'h3bfa48a3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ff890),
	.w1(32'hbbd9cdd2),
	.w2(32'hbbb8fdbe),
	.w3(32'hb9d64fe6),
	.w4(32'h3ab9afe6),
	.w5(32'h3bdea9b0),
	.w6(32'hbb326250),
	.w7(32'hbb875154),
	.w8(32'h3c1b6f1e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830254),
	.w1(32'hbbb4423c),
	.w2(32'hbba02389),
	.w3(32'hbb9d53cd),
	.w4(32'hbb39a356),
	.w5(32'h3b6c6c20),
	.w6(32'hbba576b6),
	.w7(32'hbbae4aed),
	.w8(32'h3b3238df),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d0e5e),
	.w1(32'hbae256a7),
	.w2(32'hbb03ec0e),
	.w3(32'h3b48b6eb),
	.w4(32'hbb75b855),
	.w5(32'hbaed4f00),
	.w6(32'h390a5b48),
	.w7(32'hbb591dee),
	.w8(32'hbbfc41f0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81db61),
	.w1(32'hbbbdc041),
	.w2(32'hbbb3fa1a),
	.w3(32'hbaaf9700),
	.w4(32'hbafadc62),
	.w5(32'hb96aed76),
	.w6(32'hbad016dc),
	.w7(32'h3bc50b5a),
	.w8(32'h3b55821c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2162d),
	.w1(32'h3a6e1569),
	.w2(32'hbbb31f8c),
	.w3(32'h3a154516),
	.w4(32'hbbe848f4),
	.w5(32'hbbacb7a4),
	.w6(32'hbb9bf9fe),
	.w7(32'hbc004b15),
	.w8(32'hbc124f00),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb620f5f),
	.w1(32'hbb861e06),
	.w2(32'h3b4bc61d),
	.w3(32'hbbdb2fd8),
	.w4(32'h3b8faae3),
	.w5(32'hba722e65),
	.w6(32'hba4b9d00),
	.w7(32'h3c1d6de6),
	.w8(32'h3afaec07),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a379),
	.w1(32'h3b98d7f6),
	.w2(32'hbacf4a72),
	.w3(32'hbad792f0),
	.w4(32'h3b568825),
	.w5(32'h3bf202da),
	.w6(32'hbb7966f3),
	.w7(32'hba3602c2),
	.w8(32'h3ad93a3b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb736eec),
	.w1(32'hbbf09899),
	.w2(32'hbb722655),
	.w3(32'hbc19a7db),
	.w4(32'hbc423135),
	.w5(32'hbb6a8151),
	.w6(32'hbb5eb4ae),
	.w7(32'h3a1bb28d),
	.w8(32'hbbce2c44),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc3218),
	.w1(32'hbc018781),
	.w2(32'hbb868965),
	.w3(32'hbb8b6538),
	.w4(32'hbb5e2c42),
	.w5(32'h3baab894),
	.w6(32'hbac3c33f),
	.w7(32'hbb66972a),
	.w8(32'hbb205dcd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a1ce),
	.w1(32'h3a069a05),
	.w2(32'hbaa8380b),
	.w3(32'h3ab5aee5),
	.w4(32'h3a2e3ee4),
	.w5(32'hbb1e73f6),
	.w6(32'h3c3a6ab3),
	.w7(32'hb9a114c4),
	.w8(32'h3a5014bd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71d8cb),
	.w1(32'h3b395320),
	.w2(32'h3af4cd54),
	.w3(32'hba2b5320),
	.w4(32'h3b19303c),
	.w5(32'h3b12dc3f),
	.w6(32'h3bc0b214),
	.w7(32'h3aba8a1f),
	.w8(32'hba91edcc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabde2b6),
	.w1(32'hbb5f28cb),
	.w2(32'hb9c5176e),
	.w3(32'h3b4a1dd9),
	.w4(32'h3b038e11),
	.w5(32'h3aa2b051),
	.w6(32'h3b5a0da8),
	.w7(32'h3b1b5024),
	.w8(32'h3aa59222),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96e3f1),
	.w1(32'hba247859),
	.w2(32'hbbcdaca8),
	.w3(32'hbb3b3015),
	.w4(32'hbb984f2f),
	.w5(32'h3a00993f),
	.w6(32'h3be2991b),
	.w7(32'hbc0b42a8),
	.w8(32'h3b9656f3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b857c12),
	.w1(32'hb9bd1479),
	.w2(32'hbbe01066),
	.w3(32'h3aa57fc6),
	.w4(32'hbbce82bb),
	.w5(32'hbbc05c3b),
	.w6(32'hbbbde5d0),
	.w7(32'hbbed11a0),
	.w8(32'hbbbca706),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc740ec),
	.w1(32'hbcc7d181),
	.w2(32'hbb8d413b),
	.w3(32'hbca066b3),
	.w4(32'hbc832804),
	.w5(32'h3b675de9),
	.w6(32'hbcc148b1),
	.w7(32'hbacb8158),
	.w8(32'h3b61a92f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a41fa1),
	.w1(32'h3bad7c5c),
	.w2(32'hbc220049),
	.w3(32'h3b516feb),
	.w4(32'hbaca1ea9),
	.w5(32'hbb914069),
	.w6(32'h3ba8cbc1),
	.w7(32'hb816c92a),
	.w8(32'h3ac3727c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b56a5),
	.w1(32'hba44f804),
	.w2(32'hbbdaaa10),
	.w3(32'hba7b59f3),
	.w4(32'hbb92b54b),
	.w5(32'hbb612cbc),
	.w6(32'hbb767748),
	.w7(32'hbc058624),
	.w8(32'hbad28277),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba542ed3),
	.w1(32'h3aaa876d),
	.w2(32'h3900bb55),
	.w3(32'h3b470182),
	.w4(32'h3b9857df),
	.w5(32'h3b1a6cff),
	.w6(32'h3b51e089),
	.w7(32'hba2cec64),
	.w8(32'hbb06a824),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d099a),
	.w1(32'h3c0a15ff),
	.w2(32'h3b09b4e2),
	.w3(32'h3ba03760),
	.w4(32'h3c129821),
	.w5(32'hba2849f1),
	.w6(32'h3c422705),
	.w7(32'h3ba5d7ab),
	.w8(32'h39312f10),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00ebbb),
	.w1(32'hb98410e6),
	.w2(32'h3aedf383),
	.w3(32'hbb866bcf),
	.w4(32'h3add75e4),
	.w5(32'hb980f172),
	.w6(32'h3c09d0cb),
	.w7(32'h3b3986df),
	.w8(32'hbb0bf244),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffc2fb),
	.w1(32'hbb924880),
	.w2(32'hbb1d2f58),
	.w3(32'h3b81178e),
	.w4(32'hba1eb109),
	.w5(32'hbae6dbc6),
	.w6(32'h3ab91b1c),
	.w7(32'h3aac304f),
	.w8(32'h39b23ef2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0ac55),
	.w1(32'h39c6d07b),
	.w2(32'hbc0af50d),
	.w3(32'h3b8702c3),
	.w4(32'hbb3e6c35),
	.w5(32'h3b1cf116),
	.w6(32'h3bb8d7df),
	.w7(32'h3b14922d),
	.w8(32'h3b21cf2f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61ffce),
	.w1(32'hbc5f6973),
	.w2(32'hbbb68482),
	.w3(32'hbb9fd3fb),
	.w4(32'hbb873f60),
	.w5(32'hbb3fdd87),
	.w6(32'hbbf79bc7),
	.w7(32'hbbc2cf1f),
	.w8(32'h3977abd7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bb8da),
	.w1(32'hbc8b43da),
	.w2(32'hbbb5859b),
	.w3(32'hbc3ca9ab),
	.w4(32'hbb649cf9),
	.w5(32'h3c2ff445),
	.w6(32'h3aa6bdf0),
	.w7(32'hbb179026),
	.w8(32'h3c9e961e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9394cc),
	.w1(32'hbbd01346),
	.w2(32'hbc3b556c),
	.w3(32'hbbaf59fc),
	.w4(32'hbc105c9b),
	.w5(32'h3aaab499),
	.w6(32'hbc2ab1c5),
	.w7(32'hbc8a40fd),
	.w8(32'h3c33a060),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa9219),
	.w1(32'hbb8caaee),
	.w2(32'hbbd5be2d),
	.w3(32'h35bc75d0),
	.w4(32'hbb23ad86),
	.w5(32'h3a6f26d1),
	.w6(32'hbbffd989),
	.w7(32'hbc28ddb1),
	.w8(32'h3b64abd6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf6972),
	.w1(32'h3b89d63a),
	.w2(32'h3bb4465d),
	.w3(32'h3bb0b298),
	.w4(32'h3aea3a73),
	.w5(32'hbbb4a6d8),
	.w6(32'h3c013754),
	.w7(32'h39637401),
	.w8(32'hbb83ed55),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574ae0),
	.w1(32'h3b65d1f8),
	.w2(32'h3bc0b1d8),
	.w3(32'h3a83c5b2),
	.w4(32'h3aa83139),
	.w5(32'hbbae83e2),
	.w6(32'hba62950a),
	.w7(32'h3b182436),
	.w8(32'hbbb271b4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883209),
	.w1(32'hb9f8ee4d),
	.w2(32'hbbb10072),
	.w3(32'hbb16aa91),
	.w4(32'h3b4b1ef6),
	.w5(32'hba9d4e72),
	.w6(32'hba6e4eb2),
	.w7(32'hba167a78),
	.w8(32'hba2f4f0b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf104ae),
	.w1(32'hbb9b90a7),
	.w2(32'hbbe98ebc),
	.w3(32'hbb4c7e85),
	.w4(32'hbbb58f41),
	.w5(32'hbc2716c7),
	.w6(32'h3a0255f1),
	.w7(32'hbbdf28f2),
	.w8(32'hbc8e5c1c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15fae8),
	.w1(32'h3b0ab4a7),
	.w2(32'h392806f4),
	.w3(32'h3b65e45f),
	.w4(32'h3c5a4513),
	.w5(32'hbb7a2c6d),
	.w6(32'h3b6c5262),
	.w7(32'h3c8f5b4c),
	.w8(32'hbbaa6366),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cbe53),
	.w1(32'hbb01f0b6),
	.w2(32'hbb6407f5),
	.w3(32'hbbadc723),
	.w4(32'hbbaf9f45),
	.w5(32'hbae55476),
	.w6(32'h3a06da23),
	.w7(32'hb9b4fffd),
	.w8(32'h3c0f2c9b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af51e9a),
	.w1(32'h3af28694),
	.w2(32'h3b379220),
	.w3(32'hbaee2195),
	.w4(32'h3aece06a),
	.w5(32'hbc254ac2),
	.w6(32'hbb6b7bb1),
	.w7(32'h3973c54f),
	.w8(32'hbc56230c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8878c2),
	.w1(32'hba5a2b44),
	.w2(32'h3c1e0a43),
	.w3(32'h3b8e4f2a),
	.w4(32'h3c14fa6c),
	.w5(32'h3acb5f8b),
	.w6(32'h3c00c7be),
	.w7(32'h3cd01524),
	.w8(32'h3b35f77b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb217dbc),
	.w1(32'hbbe6869c),
	.w2(32'hbc2b4696),
	.w3(32'hbb87f8fe),
	.w4(32'hbc1b3bd6),
	.w5(32'hbb99cdbf),
	.w6(32'hbb550e1f),
	.w7(32'hbc1f6910),
	.w8(32'hbbcc273e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912701),
	.w1(32'hbc438a09),
	.w2(32'hbbc9ab82),
	.w3(32'hbbbccb3c),
	.w4(32'hbb3fe819),
	.w5(32'hba29ed31),
	.w6(32'hbbe4e4a7),
	.w7(32'hb80749d6),
	.w8(32'hbb14f7a7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97afbd),
	.w1(32'h3abc9fba),
	.w2(32'h3aabe464),
	.w3(32'hb90a51f0),
	.w4(32'h3b41806a),
	.w5(32'h39a9beb3),
	.w6(32'hbb4dbf74),
	.w7(32'h3c057dcf),
	.w8(32'h3a025f4a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f2d9a),
	.w1(32'hbb883b38),
	.w2(32'hbb218bf2),
	.w3(32'hbb0aba0f),
	.w4(32'hb99cdb2c),
	.w5(32'h3bbd475e),
	.w6(32'h3b1338f3),
	.w7(32'h3bc6714e),
	.w8(32'h3b82a8fc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6b24),
	.w1(32'hb9d1e74a),
	.w2(32'h3afd1f6b),
	.w3(32'h3b5ea92c),
	.w4(32'h3ba84733),
	.w5(32'hbb1e04d1),
	.w6(32'h3b8a2660),
	.w7(32'h3bee9392),
	.w8(32'hbb0a7c0c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe86145),
	.w1(32'hbaf4e3de),
	.w2(32'hb9b51ec8),
	.w3(32'hbb8fb409),
	.w4(32'hbb14357c),
	.w5(32'h3b4118a9),
	.w6(32'h3ae427f4),
	.w7(32'h3b45dcfc),
	.w8(32'h3c098be3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf7ee),
	.w1(32'hbb09c2c5),
	.w2(32'hbc715dd7),
	.w3(32'hbac618c3),
	.w4(32'hbc151d8a),
	.w5(32'h3b1e7c8a),
	.w6(32'h3b1c70b5),
	.w7(32'hbb124e21),
	.w8(32'h3b6b9e37),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9732a2),
	.w1(32'hbba74772),
	.w2(32'hbbd0292d),
	.w3(32'hbad60b86),
	.w4(32'hbb857e3a),
	.w5(32'hbb20bf08),
	.w6(32'h3abd16bf),
	.w7(32'hbc31953d),
	.w8(32'hbb68e61c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbade4a1),
	.w1(32'hbbca6e07),
	.w2(32'hbb7b09b0),
	.w3(32'hbabbc0af),
	.w4(32'hb8ee6ca3),
	.w5(32'h3b75b1d4),
	.w6(32'h3afd0dd1),
	.w7(32'hbb01c61a),
	.w8(32'h3b9e1ada),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51ddae),
	.w1(32'hb9032e0e),
	.w2(32'hbbed9804),
	.w3(32'hbb1cdf6f),
	.w4(32'hbbd14e7f),
	.w5(32'hbb19838f),
	.w6(32'hbb4d9d55),
	.w7(32'hbc0427e0),
	.w8(32'hbb10e04f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafed54b),
	.w1(32'hbb8f2c11),
	.w2(32'h3ad57caf),
	.w3(32'hba400877),
	.w4(32'hba1c6b03),
	.w5(32'hbbae6031),
	.w6(32'hbb3a1e93),
	.w7(32'h3a1ad3d5),
	.w8(32'hbc0070a7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b6802),
	.w1(32'hbae37466),
	.w2(32'h3b49bd3b),
	.w3(32'hbbb0968b),
	.w4(32'h3bd8af06),
	.w5(32'h3bddcd6a),
	.w6(32'h3bbed687),
	.w7(32'h3c36aa95),
	.w8(32'h3c88982e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b606322),
	.w1(32'hbb9f256b),
	.w2(32'hbbfc9cb8),
	.w3(32'hbbc7cdab),
	.w4(32'hbc2d8b9d),
	.w5(32'hbb6ae402),
	.w6(32'h3b616e07),
	.w7(32'hbadec540),
	.w8(32'h3c832772),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce1ecf),
	.w1(32'h3bc8f753),
	.w2(32'hbc3a82a6),
	.w3(32'hbab1aa2e),
	.w4(32'h3b2438e4),
	.w5(32'hbb0c547f),
	.w6(32'h3c360a31),
	.w7(32'hbbd3b450),
	.w8(32'hbaee709c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c0ca),
	.w1(32'hbbc9d145),
	.w2(32'h3ad43073),
	.w3(32'hbbfd5d11),
	.w4(32'h3b8b1e16),
	.w5(32'hba944033),
	.w6(32'hbc20e499),
	.w7(32'hb91f65c1),
	.w8(32'h3b70da8e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba556c4c),
	.w1(32'hba4b212c),
	.w2(32'h39cc35c7),
	.w3(32'h3ad37fec),
	.w4(32'h3ab53ab7),
	.w5(32'h3b5cdbe2),
	.w6(32'hb8dd4ded),
	.w7(32'h3af6394d),
	.w8(32'h3c07778d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8858b92),
	.w1(32'hb9e12f5e),
	.w2(32'h3ae3ea4a),
	.w3(32'h3a0198bc),
	.w4(32'hbb83fecc),
	.w5(32'hbc8e63a7),
	.w6(32'hba94f4cf),
	.w7(32'hbafd853b),
	.w8(32'hbcd57a79),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9086b),
	.w1(32'hbaa85b6b),
	.w2(32'h3c8c10b4),
	.w3(32'h3b4e2b12),
	.w4(32'h3c543819),
	.w5(32'h3a286456),
	.w6(32'h3b639d4f),
	.w7(32'h3cf066e3),
	.w8(32'h3baa7b46),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91ade9),
	.w1(32'hbbd9a3b0),
	.w2(32'hbb8e14f6),
	.w3(32'h39830776),
	.w4(32'hba566c74),
	.w5(32'hb7bffe64),
	.w6(32'h3c0047e4),
	.w7(32'hbb9a3acc),
	.w8(32'hba392303),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada8fdb),
	.w1(32'h39eaab64),
	.w2(32'h3a1e7f33),
	.w3(32'hb9652e0b),
	.w4(32'h3a9fc2da),
	.w5(32'hbb0f84bb),
	.w6(32'hb95d2e73),
	.w7(32'h3a24db3e),
	.w8(32'hbb455244),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a210),
	.w1(32'hbbf27749),
	.w2(32'hbbb25a4c),
	.w3(32'hbba494fe),
	.w4(32'hbb936c13),
	.w5(32'hbb152d07),
	.w6(32'hbbaa2a7c),
	.w7(32'hbb5d28f8),
	.w8(32'hbabb398f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6eb2e),
	.w1(32'hbbcad514),
	.w2(32'hbb5f3504),
	.w3(32'hbb31b354),
	.w4(32'hbb642842),
	.w5(32'h35ff6232),
	.w6(32'hbb2ba2fa),
	.w7(32'hbb3939c9),
	.w8(32'h3aa786bf),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b9cc6),
	.w1(32'h3bb5c59d),
	.w2(32'h3bb3756f),
	.w3(32'h39bcfc17),
	.w4(32'hb9396f6d),
	.w5(32'h3b71eada),
	.w6(32'h3aeaaa37),
	.w7(32'h3b9a2870),
	.w8(32'h3b26c437),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b6945),
	.w1(32'hbbe2c2f3),
	.w2(32'hbbb9f0c1),
	.w3(32'h3ac144c4),
	.w4(32'hbb7749c8),
	.w5(32'hbb5ea50a),
	.w6(32'h3b0bba94),
	.w7(32'hba5d3441),
	.w8(32'h3a3bbe5e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb126b18),
	.w1(32'hbba3afd7),
	.w2(32'hbba03401),
	.w3(32'hba67c8b1),
	.w4(32'hbab3a5a6),
	.w5(32'h3b8dabec),
	.w6(32'hbb13c0e5),
	.w7(32'hbb6b17ce),
	.w8(32'h3ab80cb6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a512ded),
	.w1(32'h3b3c657a),
	.w2(32'h3b818955),
	.w3(32'h3b8f1893),
	.w4(32'h3b9a6dda),
	.w5(32'hbac75553),
	.w6(32'h394cf4f6),
	.w7(32'h3b6badd3),
	.w8(32'hba937755),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cfb4e),
	.w1(32'hbb83605c),
	.w2(32'hbb5a932e),
	.w3(32'hbb2fb6b3),
	.w4(32'hbb888578),
	.w5(32'h3a5a1a54),
	.w6(32'hba2b3cb2),
	.w7(32'hbaecb038),
	.w8(32'hbac2b34f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825802),
	.w1(32'hbb6cf8f1),
	.w2(32'hbbaba8d3),
	.w3(32'h3b0d3649),
	.w4(32'hb9e51ad5),
	.w5(32'h3ab20168),
	.w6(32'hbb0e6911),
	.w7(32'hbb386e05),
	.w8(32'h38733f4c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b1239),
	.w1(32'hba462c93),
	.w2(32'hbb4243a9),
	.w3(32'h3a781902),
	.w4(32'hbaea548a),
	.w5(32'hba0b7f04),
	.w6(32'h3abd3d54),
	.w7(32'hbb557352),
	.w8(32'hba4fbb9b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bb61e),
	.w1(32'hb7b604e7),
	.w2(32'h3b1442f8),
	.w3(32'hb94821dd),
	.w4(32'h3b19ceb1),
	.w5(32'h3b4715ed),
	.w6(32'h39b18c26),
	.w7(32'h3b1f614a),
	.w8(32'h3a9e5a87),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad40c11),
	.w1(32'h3a72b0e7),
	.w2(32'h3b372182),
	.w3(32'h3b10cd85),
	.w4(32'h3b0e68cc),
	.w5(32'hba8973a9),
	.w6(32'h3a7b549c),
	.w7(32'h3ab45481),
	.w8(32'hbaa3ccff),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c7a18),
	.w1(32'hbb190991),
	.w2(32'hb9a882d2),
	.w3(32'h3a60086c),
	.w4(32'h3a5d661b),
	.w5(32'h39f85b97),
	.w6(32'h39c7aa6c),
	.w7(32'h39d1096e),
	.w8(32'h3b62b82d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3898ffd7),
	.w1(32'hbacf6cc7),
	.w2(32'h3b5e854c),
	.w3(32'hbac7a5df),
	.w4(32'h3b56f7f5),
	.w5(32'hba37a684),
	.w6(32'h3a747b3e),
	.w7(32'h3c14aac0),
	.w8(32'h3a40ebbc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368640d4),
	.w1(32'h3a4950c8),
	.w2(32'h3b75fbc5),
	.w3(32'hba2bf325),
	.w4(32'hba13a8b5),
	.w5(32'h3b0cb8aa),
	.w6(32'h3b048e26),
	.w7(32'h3b5468fb),
	.w8(32'h3b5ef318),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffe65e),
	.w1(32'hbaf2eaed),
	.w2(32'h3b53c14b),
	.w3(32'h3ac27c2a),
	.w4(32'h3b1ffe51),
	.w5(32'h3948c361),
	.w6(32'h3ade1521),
	.w7(32'h3b14ecd3),
	.w8(32'h3a2e492a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfb9e6),
	.w1(32'hbaf6f70a),
	.w2(32'hba9cbd49),
	.w3(32'hbaedc8f9),
	.w4(32'h3a8af2b0),
	.w5(32'hbae7cc46),
	.w6(32'hbb278221),
	.w7(32'hba6a8cec),
	.w8(32'h3ab1c604),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3afb1),
	.w1(32'h3b22c9ad),
	.w2(32'h3bae239d),
	.w3(32'hba2e6efb),
	.w4(32'h3b12f92d),
	.w5(32'h39c371e1),
	.w6(32'h3946dee8),
	.w7(32'h3be6e14e),
	.w8(32'h3ac6949d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b192ec7),
	.w1(32'h3b651c8f),
	.w2(32'h3b878b69),
	.w3(32'h3a615769),
	.w4(32'h3b493aa9),
	.w5(32'h39b777c4),
	.w6(32'h3ad5861b),
	.w7(32'h3b1ce65d),
	.w8(32'h38b35a6f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff5a96),
	.w1(32'hba445c9f),
	.w2(32'hbb78481b),
	.w3(32'hbb0c8eb4),
	.w4(32'hbaf75c89),
	.w5(32'h3977e24c),
	.w6(32'hbaa3431e),
	.w7(32'hba9c2940),
	.w8(32'hba07188d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb4896),
	.w1(32'hbb35afa8),
	.w2(32'hbb60f7d4),
	.w3(32'h3af1dfe7),
	.w4(32'h39e8f72a),
	.w5(32'h3abf5d74),
	.w6(32'h3b4f569d),
	.w7(32'h3a718357),
	.w8(32'h3a6de2db),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba472df7),
	.w1(32'hba76b464),
	.w2(32'hbab0eff3),
	.w3(32'h3b38f2e3),
	.w4(32'h3b01a365),
	.w5(32'hb9f701e5),
	.w6(32'h3b10b90c),
	.w7(32'hbac3f34a),
	.w8(32'h3a20336a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a3e56),
	.w1(32'h3b18e94e),
	.w2(32'h39f9d865),
	.w3(32'hbb447edb),
	.w4(32'hba961aea),
	.w5(32'hbb8888cd),
	.w6(32'hbb0be181),
	.w7(32'h391691d8),
	.w8(32'hbb4e9f86),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae235bd),
	.w1(32'hbb5864bf),
	.w2(32'hbab4e754),
	.w3(32'hba634971),
	.w4(32'h3a165c68),
	.w5(32'h3ade856a),
	.w6(32'hbb33e67d),
	.w7(32'h386f857b),
	.w8(32'hbaa34740),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacfeb5),
	.w1(32'h3a4941d5),
	.w2(32'h39985113),
	.w3(32'hba989fe1),
	.w4(32'hbb417030),
	.w5(32'hbba10e47),
	.w6(32'h39b1a962),
	.w7(32'h39f12160),
	.w8(32'hbb7e226a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd03d25),
	.w1(32'hbbc04f79),
	.w2(32'hbb1a2d0c),
	.w3(32'hbb925435),
	.w4(32'hbb8883e4),
	.w5(32'h3b36aab9),
	.w6(32'hbabbbcb5),
	.w7(32'hbae72210),
	.w8(32'h3afc570f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97c4cc),
	.w1(32'h3b0e935e),
	.w2(32'h3b1a6e93),
	.w3(32'h3ac3de8e),
	.w4(32'h3a95b709),
	.w5(32'h3b45e164),
	.w6(32'h3b15e787),
	.w7(32'h3ac768a9),
	.w8(32'h3b042c69),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dfeb48),
	.w1(32'hba699b93),
	.w2(32'hbaea8c30),
	.w3(32'hba3f6536),
	.w4(32'hba3355af),
	.w5(32'hba3307d5),
	.w6(32'hbb0c4227),
	.w7(32'h3992a0c9),
	.w8(32'hbab1499e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af76033),
	.w1(32'h3ac35412),
	.w2(32'h3b572953),
	.w3(32'h3a45e44d),
	.w4(32'h3b25705c),
	.w5(32'hb9939ea6),
	.w6(32'hba93e531),
	.w7(32'h3a040c48),
	.w8(32'h388bf7c7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8725e7),
	.w1(32'hbac37c04),
	.w2(32'hbb700ac0),
	.w3(32'h3adde1f9),
	.w4(32'h3b95a5d7),
	.w5(32'h3b6787b6),
	.w6(32'hb9e937b9),
	.w7(32'h3b53c2cb),
	.w8(32'h3b877ff4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule