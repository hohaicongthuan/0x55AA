module layer_10_featuremap_84(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398929b5),
	.w1(32'hbaf54864),
	.w2(32'hbb33c223),
	.w3(32'hba9e1ea0),
	.w4(32'h3b0d8ab2),
	.w5(32'h3b8bb413),
	.w6(32'hbcdab1c5),
	.w7(32'h3b6aac21),
	.w8(32'h3ac34c14),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcceb8f1),
	.w1(32'h3bb7ef64),
	.w2(32'h3c1be309),
	.w3(32'h3ba3a50c),
	.w4(32'h3baea512),
	.w5(32'h3c172a9f),
	.w6(32'hba9aa5df),
	.w7(32'hbb802df7),
	.w8(32'h3b3e49d2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909c2b),
	.w1(32'h39d0bf78),
	.w2(32'h3b05c69d),
	.w3(32'h3ab558d6),
	.w4(32'hbb8ade9c),
	.w5(32'hba66bb9c),
	.w6(32'hbb3a26b9),
	.w7(32'hb990750e),
	.w8(32'hba83d6b1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb822d),
	.w1(32'hba38e0c8),
	.w2(32'h3ac02b89),
	.w3(32'hba9ab802),
	.w4(32'h3b56bcc8),
	.w5(32'hb9d2e0e3),
	.w6(32'h3a7c9217),
	.w7(32'h3b338c4a),
	.w8(32'hbb60c5c2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0738da),
	.w1(32'hbae7d09a),
	.w2(32'h3aa0b91b),
	.w3(32'hbb0e9a43),
	.w4(32'hbb517e6c),
	.w5(32'hba4bc68f),
	.w6(32'h3b0ceabe),
	.w7(32'hbac7a59c),
	.w8(32'hbb7f21c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b6ed),
	.w1(32'hbafc5ba1),
	.w2(32'h3b94ce7a),
	.w3(32'h3a650b33),
	.w4(32'hbb3041bf),
	.w5(32'h3b9ef7ff),
	.w6(32'hbc54fe27),
	.w7(32'hbb22c276),
	.w8(32'h3a75830f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4880b5),
	.w1(32'hbc01fdf0),
	.w2(32'hbc97706b),
	.w3(32'h3c077aca),
	.w4(32'hbbde1ff0),
	.w5(32'hbcc61956),
	.w6(32'hbc2fc15e),
	.w7(32'hbc0597dd),
	.w8(32'hb8899db0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1fb530),
	.w1(32'hbc68b6f2),
	.w2(32'hbc46b754),
	.w3(32'hbc105588),
	.w4(32'hbc088b4d),
	.w5(32'hb901bfbd),
	.w6(32'h3bcc15cb),
	.w7(32'h3c31feb8),
	.w8(32'h3b357426),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59569),
	.w1(32'h3c01a844),
	.w2(32'hbbf5f54f),
	.w3(32'h3b85578d),
	.w4(32'h386f2ef8),
	.w5(32'h3ae7445e),
	.w6(32'hbb3db97b),
	.w7(32'hb9a9c41f),
	.w8(32'hb8c60834),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc74fac),
	.w1(32'hbb97a050),
	.w2(32'hbc06be55),
	.w3(32'hbb36e6b9),
	.w4(32'hbbe327e6),
	.w5(32'hbc5a26c8),
	.w6(32'hbb8fc118),
	.w7(32'hbbb0af7e),
	.w8(32'hbbf4473a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ed2e9),
	.w1(32'hb9c38888),
	.w2(32'hb848decb),
	.w3(32'h3b42cb23),
	.w4(32'h3c57fc89),
	.w5(32'hbd0131ac),
	.w6(32'h3af1c31c),
	.w7(32'hb931c475),
	.w8(32'h3990ef05),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a7215),
	.w1(32'h3a8a069f),
	.w2(32'hbccd1643),
	.w3(32'h3bc2b28e),
	.w4(32'h3bb78f24),
	.w5(32'hbccde4e6),
	.w6(32'hbbc29ba0),
	.w7(32'hbbaa5652),
	.w8(32'hbc0039aa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46109a),
	.w1(32'hbc3e9493),
	.w2(32'hbc374563),
	.w3(32'hbbdc2689),
	.w4(32'hbc0a918a),
	.w5(32'hbc09dcf8),
	.w6(32'hbaf57907),
	.w7(32'h3b0133b5),
	.w8(32'hbb2fb3d5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c556b32),
	.w1(32'hbc218524),
	.w2(32'hbbb0e897),
	.w3(32'hbc12573e),
	.w4(32'hbc4796e5),
	.w5(32'hbb71009e),
	.w6(32'h3b090554),
	.w7(32'h3cd42194),
	.w8(32'hbb15a943),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f9a67),
	.w1(32'h3b9d0875),
	.w2(32'h3baf312c),
	.w3(32'h3b824f1f),
	.w4(32'h3c20667c),
	.w5(32'h3bffd589),
	.w6(32'h3b0c9184),
	.w7(32'hbaad6512),
	.w8(32'hbb6421e7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c83d5),
	.w1(32'hbbe843a9),
	.w2(32'h3c31adea),
	.w3(32'hbc2b4bc6),
	.w4(32'hbb0f27fb),
	.w5(32'h3bd2e472),
	.w6(32'h3b4dadb0),
	.w7(32'hbb124cc4),
	.w8(32'h3ca82b29),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfadf9),
	.w1(32'h3cce8c6d),
	.w2(32'hb9c519e0),
	.w3(32'hba497aa1),
	.w4(32'h38961364),
	.w5(32'hbbe970a9),
	.w6(32'h3b8180e1),
	.w7(32'hba976ab1),
	.w8(32'h3b1dfc52),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d442f),
	.w1(32'hbd2c0be8),
	.w2(32'hbcd6e129),
	.w3(32'hbbcfb538),
	.w4(32'hbc67b479),
	.w5(32'hbc1b34a0),
	.w6(32'h3abb7a78),
	.w7(32'hbbc3ee13),
	.w8(32'h3bd3a092),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67048a),
	.w1(32'hbccdfef6),
	.w2(32'hbb8d5cbe),
	.w3(32'hbb35d162),
	.w4(32'hbb2d6c92),
	.w5(32'hbbe8be54),
	.w6(32'h3aa4255f),
	.w7(32'hbb70d38a),
	.w8(32'hb986a63b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb6b5d),
	.w1(32'h3a42264f),
	.w2(32'h3b23dce0),
	.w3(32'h3b34d172),
	.w4(32'h3bf30567),
	.w5(32'h3aaf6da4),
	.w6(32'h3a32be54),
	.w7(32'hbaea0e6b),
	.w8(32'hbb0861c7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0516da),
	.w1(32'hba27f7e6),
	.w2(32'h3b1c756d),
	.w3(32'h3a878e12),
	.w4(32'h3a43f8a4),
	.w5(32'hba69d4d6),
	.w6(32'hbc5c9c04),
	.w7(32'hbac5207e),
	.w8(32'h3a60418d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5a092),
	.w1(32'h3b788565),
	.w2(32'h3b4f55be),
	.w3(32'hb9ccb4df),
	.w4(32'h3b1b5c0a),
	.w5(32'h3b635dab),
	.w6(32'hbb49f40c),
	.w7(32'hba99140d),
	.w8(32'h3af348d1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85f26b),
	.w1(32'h3c074ea4),
	.w2(32'hbcb7d6ce),
	.w3(32'h3bca5cfd),
	.w4(32'h3b4877c0),
	.w5(32'hbd0d7040),
	.w6(32'hbc112165),
	.w7(32'hbaa30df6),
	.w8(32'hbc4b8951),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81eded),
	.w1(32'hba470d83),
	.w2(32'hbb212d3f),
	.w3(32'h3b884933),
	.w4(32'h3b54c825),
	.w5(32'h390f3640),
	.w6(32'h3ba712eb),
	.w7(32'hba99c035),
	.w8(32'hbb2a6275),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92dd08a),
	.w1(32'h3bdfb8ca),
	.w2(32'h3c1bd288),
	.w3(32'h3991d1ef),
	.w4(32'h3c28fa16),
	.w5(32'h3c9c6dde),
	.w6(32'hbbacf008),
	.w7(32'hbb49f738),
	.w8(32'hbbd2e081),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0023bb),
	.w1(32'hbb8cd699),
	.w2(32'h3bcb04d3),
	.w3(32'hb92b9a13),
	.w4(32'hbc11005c),
	.w5(32'h3a04d55e),
	.w6(32'h3c06f7ce),
	.w7(32'hba218752),
	.w8(32'hb9aa5b92),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b10e7),
	.w1(32'h3a777639),
	.w2(32'hba87c339),
	.w3(32'hbb106403),
	.w4(32'h3b817ec2),
	.w5(32'hbad9cfe1),
	.w6(32'h3ad671b5),
	.w7(32'h3a175bd4),
	.w8(32'h3b88a9b0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8fcd),
	.w1(32'hbd090a52),
	.w2(32'hbc41c799),
	.w3(32'h3a6127f8),
	.w4(32'hbc934800),
	.w5(32'hbcdb466c),
	.w6(32'h3b27982c),
	.w7(32'h3da21c2b),
	.w8(32'hbcb7e8d3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8b0d8),
	.w1(32'h3b758945),
	.w2(32'hb9d355aa),
	.w3(32'hbb881217),
	.w4(32'h3b3952a8),
	.w5(32'h3a1dbaba),
	.w6(32'h3bf270c6),
	.w7(32'hbb5f7596),
	.w8(32'h3adfbce0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1e1bd),
	.w1(32'hbb260500),
	.w2(32'h3b4116ac),
	.w3(32'h3b500547),
	.w4(32'hbbb4f446),
	.w5(32'h3a1466ed),
	.w6(32'h3be9fd24),
	.w7(32'hbc1c0613),
	.w8(32'hbc9c36bb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f6583),
	.w1(32'h3b4b5e32),
	.w2(32'hbbdd7612),
	.w3(32'hbb96b930),
	.w4(32'h3b7bafbc),
	.w5(32'h3b4763b8),
	.w6(32'hbb4c9d9f),
	.w7(32'h3c1de055),
	.w8(32'h3b156d98),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03a486),
	.w1(32'h3b628262),
	.w2(32'h3a7f986b),
	.w3(32'hbc11989f),
	.w4(32'hbb0611a8),
	.w5(32'h3b800886),
	.w6(32'h3b054407),
	.w7(32'hbb64add1),
	.w8(32'h3b13836a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b725b),
	.w1(32'hbb8bcf19),
	.w2(32'hbb5b3926),
	.w3(32'h3bac6c11),
	.w4(32'h3c0786da),
	.w5(32'hbb2532a5),
	.w6(32'h3b81cbad),
	.w7(32'hbc2f94fc),
	.w8(32'hbb0fcc15),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d339c),
	.w1(32'hbc4949a9),
	.w2(32'h3c95b2d3),
	.w3(32'h3bbc8d2a),
	.w4(32'hbaa0fc04),
	.w5(32'h3ba03be0),
	.w6(32'hbb7116ed),
	.w7(32'hbb3056d8),
	.w8(32'hbbb3e4e9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82099c),
	.w1(32'hbb0849d5),
	.w2(32'hbac1e7eb),
	.w3(32'hbadf78bc),
	.w4(32'hbaa7a481),
	.w5(32'hbbbbfea9),
	.w6(32'h3b92cc88),
	.w7(32'hbb8a0aae),
	.w8(32'h3bc507b0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3406f9),
	.w1(32'h3caefddb),
	.w2(32'hbbb134d1),
	.w3(32'h3ab8b3d2),
	.w4(32'hbb7821e6),
	.w5(32'hbbad2a3e),
	.w6(32'hbd8641b1),
	.w7(32'h3c2975c2),
	.w8(32'h39e0a17f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128e4c),
	.w1(32'h3d79ea19),
	.w2(32'hbc874082),
	.w3(32'h3d19f312),
	.w4(32'h3d8a1f21),
	.w5(32'hbdc01030),
	.w6(32'hbad73451),
	.w7(32'h3b9bfed4),
	.w8(32'hbca1cb5d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42af6c),
	.w1(32'hbb860666),
	.w2(32'h3c93f4e7),
	.w3(32'hb88b00d2),
	.w4(32'h3b4512dd),
	.w5(32'h3c92d9a5),
	.w6(32'hbc5cfb18),
	.w7(32'hbcb79b85),
	.w8(32'hbc404934),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f8bf3),
	.w1(32'hbc8eedac),
	.w2(32'h3b487de2),
	.w3(32'hbc428766),
	.w4(32'hbcc4074d),
	.w5(32'h3baf8406),
	.w6(32'hbbb157ed),
	.w7(32'hbc83a37e),
	.w8(32'h3c68bd8a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160f07),
	.w1(32'hba88d579),
	.w2(32'h3b372a86),
	.w3(32'hba8b0f8c),
	.w4(32'h3bd0dfe0),
	.w5(32'h3bd0fd01),
	.w6(32'h3c7728c3),
	.w7(32'hbaa2f7a6),
	.w8(32'h3c9f8782),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872b528),
	.w1(32'h3c298e32),
	.w2(32'hbb7f0e47),
	.w3(32'hbb262a7a),
	.w4(32'h3bea9782),
	.w5(32'hbb90d06c),
	.w6(32'hb9f243b8),
	.w7(32'h3b314668),
	.w8(32'h3bc2ff82),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a582d28),
	.w1(32'hbb73a256),
	.w2(32'hbb538526),
	.w3(32'h3c371f3a),
	.w4(32'hbd10119c),
	.w5(32'hb9df779a),
	.w6(32'h3c784036),
	.w7(32'h3b12e99a),
	.w8(32'hbcec1bb5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4af08a),
	.w1(32'h3be0fe39),
	.w2(32'hbad71125),
	.w3(32'hbb5bf85d),
	.w4(32'hbb9bf40c),
	.w5(32'hb7ad545c),
	.w6(32'hbb4fd726),
	.w7(32'h3a85be00),
	.w8(32'h3b8030a7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c22ec),
	.w1(32'hbcef2e19),
	.w2(32'hbc33d2d4),
	.w3(32'hbb9099c6),
	.w4(32'hbc3fbeac),
	.w5(32'hbbce51d7),
	.w6(32'h3afe7ff1),
	.w7(32'hbd719762),
	.w8(32'hb90d6fd7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e4d6),
	.w1(32'hbd0142b3),
	.w2(32'h3bcf8595),
	.w3(32'h3c0e18bc),
	.w4(32'h3a35bc15),
	.w5(32'hbd041b9e),
	.w6(32'hb8d21dbf),
	.w7(32'h3bdbf5db),
	.w8(32'hbbb35074),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987e09),
	.w1(32'h3bbaa77a),
	.w2(32'h3a4373c1),
	.w3(32'h3b806e67),
	.w4(32'h3bacdda8),
	.w5(32'h3c2a8573),
	.w6(32'h3d255701),
	.w7(32'h3c0e3618),
	.w8(32'hbb334b7e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35073d),
	.w1(32'h3b4f9bfe),
	.w2(32'h3bc5dc9c),
	.w3(32'h3c9558d9),
	.w4(32'h3c27b131),
	.w5(32'hbcc99649),
	.w6(32'h3af2ebd7),
	.w7(32'h3b3f369c),
	.w8(32'h3c06c30b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81888e),
	.w1(32'hbc4eca7b),
	.w2(32'hbc3e843d),
	.w3(32'hbb918d05),
	.w4(32'hbcbb03b2),
	.w5(32'hbccfbf77),
	.w6(32'h3ac1ca23),
	.w7(32'hbbe886ac),
	.w8(32'h39f1383d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398856d9),
	.w1(32'hbbffcc33),
	.w2(32'hbd0bc5fb),
	.w3(32'h3b30f827),
	.w4(32'h3ab066e3),
	.w5(32'hbb7f0ea2),
	.w6(32'hba7f1bec),
	.w7(32'hbb8d47f1),
	.w8(32'hbb7cf889),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeba693),
	.w1(32'h3c155d6a),
	.w2(32'hbbbe540c),
	.w3(32'hbb47914e),
	.w4(32'h3c99e54d),
	.w5(32'hbc00f4b8),
	.w6(32'h3a77166c),
	.w7(32'h3a21fee9),
	.w8(32'hb9e0d90a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15addd),
	.w1(32'h3a74975d),
	.w2(32'h3a68069f),
	.w3(32'h3aaf7168),
	.w4(32'hb954ba4e),
	.w5(32'h3a16c33b),
	.w6(32'h3a0b219c),
	.w7(32'h3b0e349e),
	.w8(32'h3b46162c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805416),
	.w1(32'hbc47182c),
	.w2(32'hbc0da0fa),
	.w3(32'hbcb3a60a),
	.w4(32'hbb46aa60),
	.w5(32'hbbae971f),
	.w6(32'hbba132bb),
	.w7(32'hba9b03c4),
	.w8(32'hbaf72851),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f8fe2),
	.w1(32'hbb97857f),
	.w2(32'h3ae1ff89),
	.w3(32'hbb8d1488),
	.w4(32'h3b09e948),
	.w5(32'hbb9b73eb),
	.w6(32'h3c180e5b),
	.w7(32'h3b8719f9),
	.w8(32'h3b1f62dc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ef50c),
	.w1(32'hbbff4d81),
	.w2(32'hb986d10c),
	.w3(32'h3b5351f0),
	.w4(32'h3c289df2),
	.w5(32'hbc9f1615),
	.w6(32'h3ba8b01a),
	.w7(32'hba1a7bf1),
	.w8(32'hbc1faff1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d8d1c),
	.w1(32'hba507a8d),
	.w2(32'hbae008c2),
	.w3(32'h3ba14333),
	.w4(32'hbbd315aa),
	.w5(32'hbb66fe5d),
	.w6(32'h3adaa243),
	.w7(32'h3b3935ed),
	.w8(32'h3b2f5e83),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a260296),
	.w1(32'hbb273c14),
	.w2(32'h3bd5b955),
	.w3(32'hbaafe368),
	.w4(32'h3ab148d3),
	.w5(32'hbc3bdbe2),
	.w6(32'hbafb84eb),
	.w7(32'hb9bf0f8e),
	.w8(32'h3ba42f00),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadc6e5),
	.w1(32'hbb45a81b),
	.w2(32'h3ba905af),
	.w3(32'h3c11dfd4),
	.w4(32'hba90063f),
	.w5(32'hbb7bb9cb),
	.w6(32'h3b587c63),
	.w7(32'hbbd47249),
	.w8(32'hbad8e352),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70553b),
	.w1(32'h3b5f64c8),
	.w2(32'h3b9433eb),
	.w3(32'hbc690b57),
	.w4(32'hbad731df),
	.w5(32'h3be7b47e),
	.w6(32'hb98ed929),
	.w7(32'h39f0fe44),
	.w8(32'h392ce197),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbb21b),
	.w1(32'hbb96c90c),
	.w2(32'hbb09823a),
	.w3(32'hbba2457c),
	.w4(32'h3c2ae618),
	.w5(32'h3b4a7b1e),
	.w6(32'h3c1167b3),
	.w7(32'h3a954c4f),
	.w8(32'h3b658c1d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ac101),
	.w1(32'h3c19330e),
	.w2(32'hbb494a4c),
	.w3(32'hbd1f8697),
	.w4(32'h3a9eab1b),
	.w5(32'hba9ea58f),
	.w6(32'hbbc7635a),
	.w7(32'hbbfa9768),
	.w8(32'hbbdf5579),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2c9a1),
	.w1(32'h3baa4a3a),
	.w2(32'hbc0b9a0c),
	.w3(32'hbb9684b2),
	.w4(32'hbaa0d46f),
	.w5(32'hbb57bbb1),
	.w6(32'hbc009489),
	.w7(32'hb9f90f1b),
	.w8(32'h3bc62683),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37c9b7),
	.w1(32'hbcab04d1),
	.w2(32'h3a77c696),
	.w3(32'h3acde3a9),
	.w4(32'hbb969375),
	.w5(32'h3d8de9e3),
	.w6(32'hbbc6a02b),
	.w7(32'hbc20d8cb),
	.w8(32'hb91d50c1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b650241),
	.w1(32'hbae73f15),
	.w2(32'h3bf9fab7),
	.w3(32'h3a6acb18),
	.w4(32'hbb85b2fd),
	.w5(32'h3c391174),
	.w6(32'hbb88cff5),
	.w7(32'hbb30bc82),
	.w8(32'hbb609752),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4204),
	.w1(32'hbd8f56aa),
	.w2(32'h3c0e1ec7),
	.w3(32'h3b52340f),
	.w4(32'hbb88afa4),
	.w5(32'hbc13386a),
	.w6(32'hbb453cab),
	.w7(32'hbba9ef09),
	.w8(32'hbc1aada8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7012f),
	.w1(32'h3c057219),
	.w2(32'hbb9699b3),
	.w3(32'hbb8ee4fc),
	.w4(32'h3a8314f5),
	.w5(32'hbbe85109),
	.w6(32'h3b4f4d5c),
	.w7(32'hbb90258a),
	.w8(32'h3bcbbd86),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38430c),
	.w1(32'hbb90f673),
	.w2(32'hbb2aa0f5),
	.w3(32'hba71cb9f),
	.w4(32'h3bcab857),
	.w5(32'h38aa3629),
	.w6(32'h3b43f862),
	.w7(32'hbc1ebb97),
	.w8(32'h3c4021f1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97a9e4),
	.w1(32'h3bce6bb3),
	.w2(32'h3c7e1152),
	.w3(32'h3b878312),
	.w4(32'hbcd7247b),
	.w5(32'hbb94f36f),
	.w6(32'h3c3edd28),
	.w7(32'hbc2216a3),
	.w8(32'hbb444832),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb118b),
	.w1(32'hbc9e3fb4),
	.w2(32'hbc76237b),
	.w3(32'h3c6d02c5),
	.w4(32'h3bd59de1),
	.w5(32'hbb5afeb1),
	.w6(32'h3cc488d5),
	.w7(32'h3cc9f184),
	.w8(32'h3c6a0ffc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf6aa),
	.w1(32'hbc7807c2),
	.w2(32'hbbd31453),
	.w3(32'hbc0ae400),
	.w4(32'h3af2fae1),
	.w5(32'h3a31533a),
	.w6(32'h3b92d666),
	.w7(32'h3d1dfe92),
	.w8(32'hba43cf50),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09ffc1),
	.w1(32'hbba66b9a),
	.w2(32'h3c5bdbbc),
	.w3(32'h3c3dbd6c),
	.w4(32'h3cadc65e),
	.w5(32'h3cb56408),
	.w6(32'hbac91dce),
	.w7(32'hbc1ba84c),
	.w8(32'hbc8f9a65),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318edb),
	.w1(32'hbd532a43),
	.w2(32'hbb675d4b),
	.w3(32'hbc4b958a),
	.w4(32'h3a3b4af4),
	.w5(32'hbc1186ca),
	.w6(32'h3c937a95),
	.w7(32'hbba7655e),
	.w8(32'hbbec9eed),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7bfd9),
	.w1(32'hbc44f622),
	.w2(32'h3bcac0b3),
	.w3(32'h3a06df99),
	.w4(32'h3b5737df),
	.w5(32'h3ba3ded1),
	.w6(32'hbbc0e2b0),
	.w7(32'h39a265fd),
	.w8(32'h3c68dce4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c152504),
	.w1(32'hba7688a7),
	.w2(32'hbc0b1e03),
	.w3(32'h3b8acf2f),
	.w4(32'h397e832a),
	.w5(32'hbafb4193),
	.w6(32'h3b844613),
	.w7(32'h3ad7dac4),
	.w8(32'h398e5bab),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89603f),
	.w1(32'hbb491c4e),
	.w2(32'hbc2d5dc4),
	.w3(32'h3b5081e9),
	.w4(32'hbbe71c31),
	.w5(32'h3abef814),
	.w6(32'hbb6e49ce),
	.w7(32'h3b8c7608),
	.w8(32'hba31df1a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d73ae),
	.w1(32'hbc27b787),
	.w2(32'h3a0c0363),
	.w3(32'h3bfa6b81),
	.w4(32'h3d59bb37),
	.w5(32'h3bbe06e4),
	.w6(32'h3c060049),
	.w7(32'hbc760956),
	.w8(32'hbc132209),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbdb4a),
	.w1(32'hbbb4d10d),
	.w2(32'hba3f7175),
	.w3(32'h3b823581),
	.w4(32'hbc32c5db),
	.w5(32'hbbc5db7c),
	.w6(32'h3ba1b7a4),
	.w7(32'h3b9b97df),
	.w8(32'hbba057d6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c8a2b),
	.w1(32'hbd76b78f),
	.w2(32'hbbca1e4f),
	.w3(32'hbb4d9c06),
	.w4(32'h3c2658a0),
	.w5(32'hbca59c8a),
	.w6(32'h3c435a40),
	.w7(32'h3c1a8abe),
	.w8(32'hbc2d59f4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02bb45),
	.w1(32'h39340609),
	.w2(32'hbb4db1d0),
	.w3(32'h3c4e8095),
	.w4(32'hb984dd21),
	.w5(32'hbaf96df0),
	.w6(32'hbc69b3f4),
	.w7(32'hbd87f871),
	.w8(32'hbd46ffc3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92cf2c),
	.w1(32'hbb4e22c9),
	.w2(32'h3a99f288),
	.w3(32'h3bcd705a),
	.w4(32'h3947e68e),
	.w5(32'hbb25de70),
	.w6(32'h3bc6aa66),
	.w7(32'h3ba621de),
	.w8(32'h3c1ddb82),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75ad8),
	.w1(32'hbb2d1645),
	.w2(32'h3c6b829f),
	.w3(32'hbb2deb2c),
	.w4(32'hbb9500a5),
	.w5(32'hbd06fc76),
	.w6(32'h3b319c09),
	.w7(32'hbca63a85),
	.w8(32'hbb2ba1a2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba92dd7),
	.w1(32'hbbb2d5db),
	.w2(32'h3b4ac570),
	.w3(32'hbb93b97f),
	.w4(32'hba91d9ed),
	.w5(32'h39abdd89),
	.w6(32'hbc04a0ca),
	.w7(32'hbb8e1e8e),
	.w8(32'h388c459c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc709c),
	.w1(32'hbd0e8c24),
	.w2(32'hbc36eea2),
	.w3(32'h3b462eb0),
	.w4(32'h3a1ec1ce),
	.w5(32'hbb655dc5),
	.w6(32'hbc4c361c),
	.w7(32'hbc159bdc),
	.w8(32'hbca26688),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10dd94),
	.w1(32'hbc3b1a8b),
	.w2(32'hbaccc063),
	.w3(32'h39ca0c2e),
	.w4(32'hba251778),
	.w5(32'h3aca3958),
	.w6(32'h3bc14e70),
	.w7(32'h3b77bbb1),
	.w8(32'hbb654b80),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14634d),
	.w1(32'h3958fc1a),
	.w2(32'h3bd9fe34),
	.w3(32'hb9e0398d),
	.w4(32'h39d940d0),
	.w5(32'hbb94adc2),
	.w6(32'h3b4af41c),
	.w7(32'h3c215a69),
	.w8(32'hbb111742),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57023f),
	.w1(32'hbaa41338),
	.w2(32'h3b13d916),
	.w3(32'hbb3c0f8c),
	.w4(32'hbd0ea18a),
	.w5(32'hbb60507e),
	.w6(32'hbb82345a),
	.w7(32'hbb7b32ea),
	.w8(32'h3b9092eb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140f78),
	.w1(32'hbb367f92),
	.w2(32'hbb1b26a4),
	.w3(32'hbb250434),
	.w4(32'hbb451e82),
	.w5(32'h3c12c06c),
	.w6(32'h3b7af618),
	.w7(32'h3afd22b6),
	.w8(32'h3b38bf41),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd89eed),
	.w1(32'h3cdbadc5),
	.w2(32'hbb4d7d6e),
	.w3(32'h3c0b3b00),
	.w4(32'h3c68951c),
	.w5(32'h3aba806f),
	.w6(32'hbbc73dfb),
	.w7(32'hbb994ce4),
	.w8(32'hbb75ded0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9dbb2),
	.w1(32'hbb300886),
	.w2(32'hbb7f289b),
	.w3(32'h3add1bdf),
	.w4(32'h3bb5bb5b),
	.w5(32'h3b7eb0aa),
	.w6(32'hbbaa5533),
	.w7(32'hbc9012cc),
	.w8(32'h3b8117be),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c194274),
	.w1(32'h3c17129c),
	.w2(32'hba4fa6ab),
	.w3(32'h3b805d70),
	.w4(32'h3c88b47b),
	.w5(32'h3b30c4d1),
	.w6(32'h3bdeb2fc),
	.w7(32'h3b730cf1),
	.w8(32'h3bca3d33),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5198e),
	.w1(32'hbb967df0),
	.w2(32'hba4ef53b),
	.w3(32'hbbaa0704),
	.w4(32'hbc27dae1),
	.w5(32'hbc86275d),
	.w6(32'h3babed1c),
	.w7(32'hbbda4125),
	.w8(32'h3b58673a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0369df),
	.w1(32'hbbdfa9f1),
	.w2(32'hbb7f7110),
	.w3(32'hbb7d4080),
	.w4(32'hbb72a91d),
	.w5(32'hb9d0d828),
	.w6(32'hbc15f59f),
	.w7(32'h3beda6bc),
	.w8(32'hbbd0edb7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e1ea5),
	.w1(32'h3b85b11c),
	.w2(32'hbc412d21),
	.w3(32'h3c8858b5),
	.w4(32'hbc02491a),
	.w5(32'hbcdfd3c5),
	.w6(32'h3b479f1c),
	.w7(32'hbc5eb0f1),
	.w8(32'hbc1fe5df),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7630fb),
	.w1(32'hbc005acc),
	.w2(32'h3bbbd49c),
	.w3(32'h3d97a8d7),
	.w4(32'hbc1dffb4),
	.w5(32'hbb02790e),
	.w6(32'hbc15fa41),
	.w7(32'hbbd4183e),
	.w8(32'hbba996d4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdabaa5),
	.w1(32'hbbcdedbe),
	.w2(32'h3d2f21ff),
	.w3(32'h3c4e111b),
	.w4(32'h3c168bc8),
	.w5(32'h3c1ab105),
	.w6(32'h3c627a3d),
	.w7(32'h3bb4504e),
	.w8(32'h3b9ad08f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc43338),
	.w1(32'hba9c842e),
	.w2(32'h3c093fdd),
	.w3(32'h3bfdae60),
	.w4(32'h3b8b2acc),
	.w5(32'h3b1b801c),
	.w6(32'h3b6ed11e),
	.w7(32'hbb3bf92a),
	.w8(32'hbcc6372d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1dfb7),
	.w1(32'hb9b65167),
	.w2(32'h3c03f2a0),
	.w3(32'hbb90ed80),
	.w4(32'h3bb63c6c),
	.w5(32'hbc528cca),
	.w6(32'hbb0f136e),
	.w7(32'hbbbe44e5),
	.w8(32'h3b91e716),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6737),
	.w1(32'h3b3015bc),
	.w2(32'hbb83edb8),
	.w3(32'h3a6a5f66),
	.w4(32'h3b6580a1),
	.w5(32'h3b055f0d),
	.w6(32'h3982bbe6),
	.w7(32'hb89c1e4a),
	.w8(32'h3953ffc5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c607de8),
	.w1(32'hbb4dcfd1),
	.w2(32'hbc0ae76a),
	.w3(32'h3b092a69),
	.w4(32'hbaee1286),
	.w5(32'hbbdef606),
	.w6(32'h3b808aa9),
	.w7(32'h3b87a7fa),
	.w8(32'hbb8b04ac),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d26db),
	.w1(32'h3bb0ce68),
	.w2(32'hbc853029),
	.w3(32'h3bdfe56b),
	.w4(32'hbbf7c06b),
	.w5(32'hbc7d09a8),
	.w6(32'h3a39f91c),
	.w7(32'hbc3dcc08),
	.w8(32'hbccd432d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b7fcf),
	.w1(32'h3d0b0b6e),
	.w2(32'hbce4e7a9),
	.w3(32'h3bb7e787),
	.w4(32'h3cd710ae),
	.w5(32'hbc9b2231),
	.w6(32'hbc17cb51),
	.w7(32'h3c1d96a2),
	.w8(32'h3ca4798c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41754f),
	.w1(32'h399a73a7),
	.w2(32'h3bbf0740),
	.w3(32'h3b386ca0),
	.w4(32'h3dad52a7),
	.w5(32'h3c73e607),
	.w6(32'h392e8bde),
	.w7(32'h3bcdbcf3),
	.w8(32'h3c06be85),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6b78),
	.w1(32'h3bb2d5c0),
	.w2(32'h3d0012ca),
	.w3(32'hba0843f2),
	.w4(32'h3c2dee91),
	.w5(32'h3bd8b5ac),
	.w6(32'h3bac689f),
	.w7(32'hbb27faef),
	.w8(32'hbba3a2d5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70c98b),
	.w1(32'h3c36b2b5),
	.w2(32'hba9f448c),
	.w3(32'hbca390b5),
	.w4(32'h3c95b392),
	.w5(32'hbc8b717f),
	.w6(32'h3b752ecf),
	.w7(32'h3a5dc48e),
	.w8(32'h3c0b71ec),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20695),
	.w1(32'h3c702b14),
	.w2(32'h3c63f631),
	.w3(32'h3aca6494),
	.w4(32'h3b487e76),
	.w5(32'hbb3f1994),
	.w6(32'hbbd8d089),
	.w7(32'hbb14b875),
	.w8(32'h3ae57723),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb82e79),
	.w1(32'h3cf21d93),
	.w2(32'hbc8d677b),
	.w3(32'h3c4c64c5),
	.w4(32'h3c67d210),
	.w5(32'hbcf84aae),
	.w6(32'hbbae4902),
	.w7(32'hb994eb57),
	.w8(32'hb9a83e81),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22762a),
	.w1(32'hbbac3757),
	.w2(32'hbca23400),
	.w3(32'h392eda0e),
	.w4(32'hbc1e1a3a),
	.w5(32'hbcb125bd),
	.w6(32'hbc5216d0),
	.w7(32'h3cfd26f4),
	.w8(32'hbc1e7a94),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca36f27),
	.w1(32'hb9b7616b),
	.w2(32'h3a995866),
	.w3(32'h3a884200),
	.w4(32'hb747128e),
	.w5(32'h3b84a907),
	.w6(32'hbaa2f243),
	.w7(32'h3b3d6de6),
	.w8(32'h392f428f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8ee93),
	.w1(32'h3b243085),
	.w2(32'h3a39d6c9),
	.w3(32'hba7cac8a),
	.w4(32'h3b8e2f3a),
	.w5(32'h3bc2f515),
	.w6(32'hbbded45f),
	.w7(32'hbb5f4d38),
	.w8(32'hbba3e314),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae65b4),
	.w1(32'hbbdfeaa0),
	.w2(32'hbc4b1fb0),
	.w3(32'hbcb639bd),
	.w4(32'hbc0f67bf),
	.w5(32'hbc741148),
	.w6(32'hba015fd3),
	.w7(32'hbbe5f4dd),
	.w8(32'hbabbc666),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76eeda),
	.w1(32'hbb198e5b),
	.w2(32'h3aa41a59),
	.w3(32'h3a43319a),
	.w4(32'h3b8b2223),
	.w5(32'h3ba6cdf5),
	.w6(32'hbb30700b),
	.w7(32'hbb0ac623),
	.w8(32'hbb3a8aba),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba03328),
	.w1(32'hbbfd2b5d),
	.w2(32'h3abfc8b6),
	.w3(32'hbb3067cc),
	.w4(32'hbca1c643),
	.w5(32'hbbada7f3),
	.w6(32'hbc0f226e),
	.w7(32'hbd12b01f),
	.w8(32'hbaae0afc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b08ca),
	.w1(32'h3c24a36e),
	.w2(32'h3c0c897c),
	.w3(32'h3afc661c),
	.w4(32'h3b53ac7e),
	.w5(32'h3a367281),
	.w6(32'hbb01ccc6),
	.w7(32'hbac286aa),
	.w8(32'hbad7f07d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad767c),
	.w1(32'hbae7c999),
	.w2(32'hbbc4cc96),
	.w3(32'h3bea6a14),
	.w4(32'h3c3b841e),
	.w5(32'h3bbe4c05),
	.w6(32'h3aa301f6),
	.w7(32'h3c5fe34f),
	.w8(32'hbc7f050c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce3defc),
	.w1(32'hbb3b9d10),
	.w2(32'h3c2424b4),
	.w3(32'hbc6826fa),
	.w4(32'hbc239fbf),
	.w5(32'h3bba6672),
	.w6(32'hbb14c3e3),
	.w7(32'hbbd28469),
	.w8(32'h3aa533ab),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f0288),
	.w1(32'h3bad1590),
	.w2(32'hba033944),
	.w3(32'hb94ad0fb),
	.w4(32'h3b3ada4b),
	.w5(32'h3bbfa2df),
	.w6(32'h3ac6d7aa),
	.w7(32'hbc259cd7),
	.w8(32'h3a35d8b4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bcc59),
	.w1(32'hbc225a61),
	.w2(32'hbb5a5c67),
	.w3(32'hbbafb607),
	.w4(32'h3a007353),
	.w5(32'hbae0bd9f),
	.w6(32'h3c03f6ad),
	.w7(32'hbab778d5),
	.w8(32'h39351d7a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af28c),
	.w1(32'h39624634),
	.w2(32'hbb7fe441),
	.w3(32'h3a0d5f7e),
	.w4(32'hbbaedf2b),
	.w5(32'h3b46910d),
	.w6(32'hbbf29c99),
	.w7(32'h3af03e2b),
	.w8(32'h38f97469),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e387b),
	.w1(32'hbb952774),
	.w2(32'h3c287fbb),
	.w3(32'h3b1e5693),
	.w4(32'h38a6013c),
	.w5(32'h3ac1c350),
	.w6(32'hbaa10f78),
	.w7(32'hbaf73379),
	.w8(32'hbbee4d2e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d6551),
	.w1(32'h3a397282),
	.w2(32'hbd40a035),
	.w3(32'hbb524873),
	.w4(32'h3b8f5e93),
	.w5(32'h3b597129),
	.w6(32'hbb5e1cc0),
	.w7(32'hbacb7d89),
	.w8(32'h3c3a79c3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc85c44),
	.w1(32'hba230f0a),
	.w2(32'hb9f64adb),
	.w3(32'hbaabf327),
	.w4(32'h3b915e53),
	.w5(32'hba9a5ac0),
	.w6(32'h3bb3488f),
	.w7(32'hbbb61b8e),
	.w8(32'hbb2a0be7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adff906),
	.w1(32'h3bc4ee25),
	.w2(32'hbc966692),
	.w3(32'hb9ecbbce),
	.w4(32'h3b737615),
	.w5(32'h3acf7343),
	.w6(32'h3cb75c94),
	.w7(32'h3c8d4aca),
	.w8(32'hbb648fde),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aef3b),
	.w1(32'hbba1e1af),
	.w2(32'hbc30cfed),
	.w3(32'hbad6c4f1),
	.w4(32'hbb75121b),
	.w5(32'hbc432c02),
	.w6(32'h3be994bc),
	.w7(32'hba103598),
	.w8(32'hbc25d9a6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb178157),
	.w1(32'h3b740aea),
	.w2(32'h3c36836e),
	.w3(32'h3b1ff8e9),
	.w4(32'h3b6b8a7c),
	.w5(32'h3ca138e6),
	.w6(32'hbb17e76f),
	.w7(32'hbc3e133d),
	.w8(32'hbbaaa77d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0229),
	.w1(32'hbc7f738b),
	.w2(32'hbbb2b6d1),
	.w3(32'h39bb5de1),
	.w4(32'hbc3b84b0),
	.w5(32'hbb8cb946),
	.w6(32'hbb041b1f),
	.w7(32'h3c2904a0),
	.w8(32'hbb9133e4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0041),
	.w1(32'h3b87c055),
	.w2(32'h3bb072d2),
	.w3(32'h3ae480fc),
	.w4(32'h3c252d69),
	.w5(32'h3c1b528d),
	.w6(32'hbcce9b27),
	.w7(32'h3c6c0a59),
	.w8(32'hbad5a766),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29bd2d),
	.w1(32'h369a19c6),
	.w2(32'h3b2ca16b),
	.w3(32'h3b52f61b),
	.w4(32'hbc5c8513),
	.w5(32'h3ad480e1),
	.w6(32'hbb90544a),
	.w7(32'h3a00824b),
	.w8(32'hbae2040c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238828),
	.w1(32'hbac77139),
	.w2(32'h39da0d64),
	.w3(32'h3b91a809),
	.w4(32'hbc2e388a),
	.w5(32'h3bc31152),
	.w6(32'hbb1121b2),
	.w7(32'hbb11b6fe),
	.w8(32'h3b865c6a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c121525),
	.w1(32'hbc999c25),
	.w2(32'hbc80c59a),
	.w3(32'h3c1bfab3),
	.w4(32'hbc25b2d8),
	.w5(32'hbc8ea518),
	.w6(32'h3b94b4de),
	.w7(32'h3cf134b6),
	.w8(32'h3c09ef62),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2186e),
	.w1(32'hbb76536e),
	.w2(32'h3bb30cf4),
	.w3(32'h3a5463a5),
	.w4(32'hbc49878b),
	.w5(32'hbc88100b),
	.w6(32'hbb1b07f0),
	.w7(32'hbb8dd445),
	.w8(32'h3c4bbae1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fb165),
	.w1(32'h3ae0d0a9),
	.w2(32'h3bcaf386),
	.w3(32'hbad135e6),
	.w4(32'hbbabae47),
	.w5(32'hbbc43c0a),
	.w6(32'hba9c46bd),
	.w7(32'hbb5a7f2c),
	.w8(32'hbb705262),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da19fe),
	.w1(32'hbc1c06b8),
	.w2(32'hb98f33d7),
	.w3(32'hbb7792ee),
	.w4(32'h3bbb3b7a),
	.w5(32'hbb49a9ff),
	.w6(32'h3a6c7fa2),
	.w7(32'hbac2d29c),
	.w8(32'h3bf8cf64),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064c3d),
	.w1(32'hbd519bb7),
	.w2(32'hbbc1a666),
	.w3(32'hbb0cf745),
	.w4(32'h3b37af21),
	.w5(32'hb951c5e7),
	.w6(32'hbac42600),
	.w7(32'hb9eff644),
	.w8(32'h3a069e07),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb2862),
	.w1(32'h3a98f56c),
	.w2(32'hbb830da6),
	.w3(32'h3cd412c5),
	.w4(32'h3b45f8cb),
	.w5(32'h3c843870),
	.w6(32'h3bc741b4),
	.w7(32'h3c65974b),
	.w8(32'hb9e098f2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ff471),
	.w1(32'hbb98c902),
	.w2(32'h3b859147),
	.w3(32'h3b61afae),
	.w4(32'hbb0e12dd),
	.w5(32'hbbc89b12),
	.w6(32'h3d0d877f),
	.w7(32'hbb907d0c),
	.w8(32'h3a7092a2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca153c6),
	.w1(32'hbc1b63c4),
	.w2(32'hbc76cd02),
	.w3(32'h3a2f0973),
	.w4(32'h3cf59d08),
	.w5(32'hbd158b7b),
	.w6(32'hbc1ec058),
	.w7(32'hbb2f1bbc),
	.w8(32'hbbdbb112),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98059d0),
	.w1(32'h3b44a103),
	.w2(32'hbb731ca7),
	.w3(32'h3afce0a3),
	.w4(32'h3b65b785),
	.w5(32'h39e381cb),
	.w6(32'hbb100d16),
	.w7(32'hbace7caf),
	.w8(32'h3b53a403),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9378d3),
	.w1(32'hbb8d4091),
	.w2(32'hbbc39b44),
	.w3(32'h3a7a610a),
	.w4(32'h3c1a0bff),
	.w5(32'hbc4dc540),
	.w6(32'h3a6d7161),
	.w7(32'h3c0c9364),
	.w8(32'h3b7c7305),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021f1a),
	.w1(32'hba950533),
	.w2(32'hbc5d2370),
	.w3(32'h3bcddb37),
	.w4(32'h3c10d6a8),
	.w5(32'hbbc47f85),
	.w6(32'h3b8ee2f4),
	.w7(32'h3b046f81),
	.w8(32'h3c2aece4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ad585),
	.w1(32'h3c25c987),
	.w2(32'hbc9cb642),
	.w3(32'h3c0cdf01),
	.w4(32'h3c6e8993),
	.w5(32'h3c05b9e1),
	.w6(32'hbadf5112),
	.w7(32'hb94bad7d),
	.w8(32'h3b727b38),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf10cb9),
	.w1(32'hbb3e4927),
	.w2(32'hbb890e39),
	.w3(32'h3c3acc8f),
	.w4(32'hbaec7888),
	.w5(32'h3b92c2ce),
	.w6(32'hbc2520d2),
	.w7(32'h3b834efa),
	.w8(32'hbb1aaa43),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa516c8),
	.w1(32'hbba1788e),
	.w2(32'hbaac4841),
	.w3(32'h3acb3a81),
	.w4(32'h3b676845),
	.w5(32'hbb7fa474),
	.w6(32'h3b09eade),
	.w7(32'h38d940ab),
	.w8(32'h3b8994fa),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0cd8),
	.w1(32'hbcd0756e),
	.w2(32'h3a51e7e7),
	.w3(32'h3c119096),
	.w4(32'hbc9bad12),
	.w5(32'h3bf56b51),
	.w6(32'h3a7af14c),
	.w7(32'hbc5e095e),
	.w8(32'hbb91e0f0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aa198),
	.w1(32'h39a0ee9c),
	.w2(32'h3b34bee7),
	.w3(32'h3b2ae8fb),
	.w4(32'h3c81c9b1),
	.w5(32'hb97f8ef1),
	.w6(32'h3ae53bfe),
	.w7(32'h3b13d92b),
	.w8(32'h38020de7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06ffee),
	.w1(32'h39697aa3),
	.w2(32'hbb6a1bc8),
	.w3(32'h3b8a815f),
	.w4(32'hbad7185f),
	.w5(32'h3ab0762e),
	.w6(32'h3b8f4636),
	.w7(32'hbb582a99),
	.w8(32'hba73a316),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b651d3b),
	.w1(32'hbb2c319d),
	.w2(32'h3c0ca251),
	.w3(32'hbaabbfdf),
	.w4(32'hbbe853ef),
	.w5(32'h3a8de711),
	.w6(32'hbbe06ef6),
	.w7(32'h3bba8afe),
	.w8(32'hbad476e8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b75ce),
	.w1(32'h3b614d6a),
	.w2(32'hbb29bf81),
	.w3(32'h3ab4b949),
	.w4(32'hb9e07a42),
	.w5(32'hba1c8914),
	.w6(32'h3c14254e),
	.w7(32'hbb2d5f27),
	.w8(32'hbb047721),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14793f),
	.w1(32'h3bdfc63b),
	.w2(32'h3a34c5c5),
	.w3(32'h3b9e4358),
	.w4(32'h3c317cef),
	.w5(32'h3a5aeae8),
	.w6(32'h3b1c9d8d),
	.w7(32'h3b0b5ff7),
	.w8(32'hbb82fa02),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0dc85),
	.w1(32'h3956f582),
	.w2(32'hbc47e3ae),
	.w3(32'hbc7c46d3),
	.w4(32'h3c877180),
	.w5(32'hbbc20e8a),
	.w6(32'hbbfe40c2),
	.w7(32'hbb6f5ce7),
	.w8(32'hbb87140b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b2bc),
	.w1(32'hbba05f11),
	.w2(32'h3b4f0c4a),
	.w3(32'h3b1ce9c7),
	.w4(32'hb99df257),
	.w5(32'h3b2069f0),
	.w6(32'h39a821e6),
	.w7(32'hbbd47158),
	.w8(32'h3b6a246e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900fb71),
	.w1(32'hbb8082e5),
	.w2(32'hbb2da7e8),
	.w3(32'hbbe657a7),
	.w4(32'hbb1aa5a9),
	.w5(32'hbbee0317),
	.w6(32'hbb95aa39),
	.w7(32'hbaac2a3a),
	.w8(32'h3c7dbf88),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16b037),
	.w1(32'h3b49ee61),
	.w2(32'hbbaf788c),
	.w3(32'h3adeee05),
	.w4(32'hbb60e7f1),
	.w5(32'hbb9a8f69),
	.w6(32'h3bbf2718),
	.w7(32'h3b3805cb),
	.w8(32'h3d14b346),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf21db),
	.w1(32'h3a3f1289),
	.w2(32'hbbebb5f3),
	.w3(32'h3c2c7100),
	.w4(32'h39370038),
	.w5(32'hbbf61c10),
	.w6(32'h3c2d4a9f),
	.w7(32'hba425e11),
	.w8(32'hbb4abc57),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c237c),
	.w1(32'hbc69ed43),
	.w2(32'hbc5c74ee),
	.w3(32'h3ab2ac54),
	.w4(32'hbbb2dc13),
	.w5(32'hbbe6b970),
	.w6(32'hb7e02216),
	.w7(32'hbc977056),
	.w8(32'hbca6db37),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be11622),
	.w1(32'h3bac42bd),
	.w2(32'hbafe82e7),
	.w3(32'h3b23a3f0),
	.w4(32'h3b9197d1),
	.w5(32'h3b87171e),
	.w6(32'h3b8e15a4),
	.w7(32'hbb72a2f4),
	.w8(32'hbb87d730),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f27a0),
	.w1(32'hba85276e),
	.w2(32'h3a05840b),
	.w3(32'h3adf1dad),
	.w4(32'hb98490e0),
	.w5(32'h3a7bd514),
	.w6(32'hba867cf0),
	.w7(32'h39f3b963),
	.w8(32'h3ba139d0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fca07),
	.w1(32'h396870a6),
	.w2(32'h3b30dcd7),
	.w3(32'h3b2d84a2),
	.w4(32'h3b05a476),
	.w5(32'hbbfb5f2c),
	.w6(32'h3b372e50),
	.w7(32'hba1a096e),
	.w8(32'h3b8903e4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451fe0),
	.w1(32'h3a7f3a38),
	.w2(32'h3b906340),
	.w3(32'h3b00ff1c),
	.w4(32'h3b444da8),
	.w5(32'h3bd2bbab),
	.w6(32'hb9a8db19),
	.w7(32'hbb102e48),
	.w8(32'hbb708422),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bed37),
	.w1(32'hbbc098a1),
	.w2(32'h3b9a2548),
	.w3(32'h38657046),
	.w4(32'h3c12b5c8),
	.w5(32'h3c256a6b),
	.w6(32'h3a10edeb),
	.w7(32'h382e2baa),
	.w8(32'h3adea10c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c080fa0),
	.w1(32'hba098919),
	.w2(32'hbb411f9d),
	.w3(32'h3b337b3a),
	.w4(32'hbac4520d),
	.w5(32'hbb3212f5),
	.w6(32'h38e49be9),
	.w7(32'hbbef3f33),
	.w8(32'hbba51843),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd889a7),
	.w1(32'h3a8023dc),
	.w2(32'hba4c8a17),
	.w3(32'hba6e08ea),
	.w4(32'h3b611b6d),
	.w5(32'h3b852c55),
	.w6(32'hbb2ba363),
	.w7(32'h3c0469ef),
	.w8(32'h3cb2107f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c30d2),
	.w1(32'h3b2c5fea),
	.w2(32'hbb8bc5ae),
	.w3(32'h3a3c9777),
	.w4(32'hbbfe5d28),
	.w5(32'hbc055084),
	.w6(32'h3b8005ac),
	.w7(32'h3c6ca54b),
	.w8(32'hbbeba580),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d9c68),
	.w1(32'hb9ba17ae),
	.w2(32'hbc691640),
	.w3(32'h3b3453cf),
	.w4(32'hb9e8b0e6),
	.w5(32'hbb898402),
	.w6(32'h3c6bd0ca),
	.w7(32'h3a7b8788),
	.w8(32'hbb26a392),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba365c2),
	.w1(32'hbb438a36),
	.w2(32'h39aa7563),
	.w3(32'hbb8da5ef),
	.w4(32'h3bfbbe65),
	.w5(32'h3b2050a6),
	.w6(32'h3b86aacd),
	.w7(32'h3ba1d45f),
	.w8(32'hbbd8dae2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2964),
	.w1(32'hb6b6df17),
	.w2(32'h3b15b532),
	.w3(32'hbb067e55),
	.w4(32'hb8c2acca),
	.w5(32'h380452e7),
	.w6(32'h383256e4),
	.w7(32'h3af9fba2),
	.w8(32'h3bbbb4b4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1a2af),
	.w1(32'hbb9e0dca),
	.w2(32'hbabc1f38),
	.w3(32'hb9f5041a),
	.w4(32'hbb23818a),
	.w5(32'hbc3706ee),
	.w6(32'h3b5d13f4),
	.w7(32'hba9d6be8),
	.w8(32'h3bd2a722),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9586780),
	.w1(32'h3a7fa327),
	.w2(32'h3ab25107),
	.w3(32'hba9816f6),
	.w4(32'hb99ff84d),
	.w5(32'h3a2a5269),
	.w6(32'h3bca69ce),
	.w7(32'hbb8b0526),
	.w8(32'hbb26efc6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b1b3a),
	.w1(32'hb75cd5d3),
	.w2(32'h3a008c57),
	.w3(32'h3bac2c49),
	.w4(32'hb96379d4),
	.w5(32'hbae8f3f0),
	.w6(32'h39bb7cf2),
	.w7(32'h3ba506ea),
	.w8(32'h3af35ed1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa17b65),
	.w1(32'h3b4dec38),
	.w2(32'h3b566a39),
	.w3(32'hbb04b6a6),
	.w4(32'hbb9dd7d1),
	.w5(32'h3ba342bb),
	.w6(32'h3c62e782),
	.w7(32'h3ababf4a),
	.w8(32'h3b240881),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c446706),
	.w1(32'hba964b56),
	.w2(32'hbc91eb6e),
	.w3(32'h3c104813),
	.w4(32'h3b01e3c0),
	.w5(32'hbc7e533b),
	.w6(32'h3be712fd),
	.w7(32'h3c06cdc7),
	.w8(32'h3beabe53),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3db96d),
	.w1(32'hbb83b166),
	.w2(32'hbb778955),
	.w3(32'h3b4747c5),
	.w4(32'h3b6ea3a7),
	.w5(32'h3b0ac4cc),
	.w6(32'h3b9e5a01),
	.w7(32'h3c33ba1d),
	.w8(32'hbb8cc34c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c574837),
	.w1(32'h3bb23a86),
	.w2(32'h3b173abe),
	.w3(32'h3bf3e3fc),
	.w4(32'hbb53dba8),
	.w5(32'h3ab48b46),
	.w6(32'h3b40e8bc),
	.w7(32'h3c178150),
	.w8(32'hbbd311e3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f48d9),
	.w1(32'h3b77f603),
	.w2(32'hbc0c508f),
	.w3(32'hbb22289a),
	.w4(32'h3b9f6cb3),
	.w5(32'hbbe4e8bf),
	.w6(32'hbc32a6e9),
	.w7(32'hbaaccf4a),
	.w8(32'hbca44d2f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8e0d8),
	.w1(32'hbc94dfe1),
	.w2(32'hbc0f4b40),
	.w3(32'hbbbe6504),
	.w4(32'hbc0d8074),
	.w5(32'hbb4044c4),
	.w6(32'hbc833e96),
	.w7(32'hbc57bdf7),
	.w8(32'h3c06e4e4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc1aa7),
	.w1(32'h3b953f9e),
	.w2(32'hbc0183e8),
	.w3(32'hbc4d1843),
	.w4(32'h3b89ece1),
	.w5(32'hbc6572cc),
	.w6(32'h3ba4db05),
	.w7(32'hbac1cedb),
	.w8(32'hbb7880b4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c72b9),
	.w1(32'hbb57574c),
	.w2(32'h3b61286f),
	.w3(32'hbb11ff92),
	.w4(32'hbb8ea026),
	.w5(32'hbaf5f4eb),
	.w6(32'hbbed4df1),
	.w7(32'h3c06cb98),
	.w8(32'hbc185d3f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ed08),
	.w1(32'hbc0508d1),
	.w2(32'hbb606890),
	.w3(32'hb82471f1),
	.w4(32'h3a3d46b2),
	.w5(32'h3a6fae8d),
	.w6(32'h3bb6ac64),
	.w7(32'h3cf02dc7),
	.w8(32'h3bdade26),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c904151),
	.w1(32'hbc0bb548),
	.w2(32'h3bd047ae),
	.w3(32'h3bd2f3fb),
	.w4(32'hba9b3eae),
	.w5(32'h3b344a95),
	.w6(32'h3b4b36cd),
	.w7(32'hbbbbde03),
	.w8(32'h3b9f9ad4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5eae),
	.w1(32'hbbbeda28),
	.w2(32'hbb2ca901),
	.w3(32'h3b6a9b80),
	.w4(32'hb9e1cf0b),
	.w5(32'hbbe165e6),
	.w6(32'hbb628343),
	.w7(32'hbabbbeb7),
	.w8(32'h3c57e94d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc35d84),
	.w1(32'hbbde2ce7),
	.w2(32'hbaeaa34d),
	.w3(32'h3b7ddca1),
	.w4(32'hbb1197ec),
	.w5(32'h3955f21f),
	.w6(32'h3b9a8202),
	.w7(32'hbbd2130b),
	.w8(32'h3ae5c724),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fe86f),
	.w1(32'h3b287852),
	.w2(32'h3c097100),
	.w3(32'hbbb93afc),
	.w4(32'h3b47f164),
	.w5(32'hb9c4bce9),
	.w6(32'hbbc181d9),
	.w7(32'hba0d8821),
	.w8(32'hbc573675),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c6c5),
	.w1(32'hbba6ef05),
	.w2(32'h3bc0db2a),
	.w3(32'hbc3d7062),
	.w4(32'hbac304f3),
	.w5(32'h3c531cfb),
	.w6(32'hbbada809),
	.w7(32'h3b9dd158),
	.w8(32'h3b7d14dc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c6bfb),
	.w1(32'h3b2638b4),
	.w2(32'hbb8d4ef1),
	.w3(32'h3a9cf4f0),
	.w4(32'hbaadb9e0),
	.w5(32'h38c4c839),
	.w6(32'hb8ed762e),
	.w7(32'hbb4a4ba2),
	.w8(32'h3a666db0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d3167),
	.w1(32'h3c241b66),
	.w2(32'h3bd514e4),
	.w3(32'h3b975703),
	.w4(32'h3861f4f4),
	.w5(32'hbb48d0bd),
	.w6(32'h38218e33),
	.w7(32'h390fe059),
	.w8(32'hba10585e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ea3c),
	.w1(32'h3a3f6219),
	.w2(32'h3c069303),
	.w3(32'h3acded43),
	.w4(32'h3b5caca3),
	.w5(32'h3c142191),
	.w6(32'hbb03a623),
	.w7(32'hbb4539ab),
	.w8(32'hbac54994),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad24a15),
	.w1(32'hbbe9e9a5),
	.w2(32'hba8b6662),
	.w3(32'h3c05817d),
	.w4(32'h3bd37fcd),
	.w5(32'hba841735),
	.w6(32'hbaf8975c),
	.w7(32'h3c9a4609),
	.w8(32'hbc80ff5b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad17648),
	.w1(32'h3c5761c0),
	.w2(32'hbb99863d),
	.w3(32'h3bca6f0f),
	.w4(32'h3c924c56),
	.w5(32'hbcdaa1df),
	.w6(32'h3a7e48a4),
	.w7(32'hbadb9b2b),
	.w8(32'hbca4db2f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3e6e2),
	.w1(32'hbb85c0ae),
	.w2(32'h3aba1296),
	.w3(32'hbbe79ce7),
	.w4(32'hbb56f632),
	.w5(32'h3bc2e3ce),
	.w6(32'h3b5089ca),
	.w7(32'hbafe784d),
	.w8(32'h3b1224f1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ea2f),
	.w1(32'hbc6d46b4),
	.w2(32'hbc384ad9),
	.w3(32'hbc14fcd1),
	.w4(32'hbb96b420),
	.w5(32'hb9a8f212),
	.w6(32'h3c296366),
	.w7(32'h3c2de51c),
	.w8(32'h3c0d8ce6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f97ab),
	.w1(32'hbc404652),
	.w2(32'h3cff4554),
	.w3(32'hbb2bc177),
	.w4(32'h38d27b1c),
	.w5(32'hbab0dbcb),
	.w6(32'h3b482666),
	.w7(32'hbbf20536),
	.w8(32'h3bba7d94),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ae01b),
	.w1(32'h38ff722d),
	.w2(32'hbc168d89),
	.w3(32'hbb8cb1fe),
	.w4(32'hbbb274c6),
	.w5(32'hbc3e7616),
	.w6(32'h3c80c0b1),
	.w7(32'h3a60a319),
	.w8(32'h3b81e224),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567edc),
	.w1(32'h3c768c4c),
	.w2(32'hbbc0243c),
	.w3(32'h3ac4c47a),
	.w4(32'hbbd3a025),
	.w5(32'h3b5c9604),
	.w6(32'h39b184ce),
	.w7(32'h385a4e11),
	.w8(32'hba2b9988),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b952),
	.w1(32'hbadb5cba),
	.w2(32'hbbd66b75),
	.w3(32'h3b729ded),
	.w4(32'h3bb836c5),
	.w5(32'h3795fffe),
	.w6(32'hbbb30fa0),
	.w7(32'h3c12b2b8),
	.w8(32'h3af6f80a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7984d),
	.w1(32'hb6fa0d60),
	.w2(32'hba4f6b69),
	.w3(32'h397b5874),
	.w4(32'hba9ce997),
	.w5(32'h3c0dc6da),
	.w6(32'hb8c3597c),
	.w7(32'h3b6ddc36),
	.w8(32'h3c3b55b2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0eef2),
	.w1(32'hbbf5f8ef),
	.w2(32'h3b467cbc),
	.w3(32'h3b4ff30a),
	.w4(32'h3c6e279b),
	.w5(32'hbc6bed62),
	.w6(32'hbc11b2a6),
	.w7(32'h3c75ab5e),
	.w8(32'hbbf2619e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade88c1),
	.w1(32'h3caaeec3),
	.w2(32'hbb554540),
	.w3(32'h3bca4535),
	.w4(32'hba832882),
	.w5(32'h3b6eedc8),
	.w6(32'h3bc0991d),
	.w7(32'hbb86df5c),
	.w8(32'h3b5819c7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c4b3),
	.w1(32'h3c0981d3),
	.w2(32'hbba07943),
	.w3(32'h3b247d05),
	.w4(32'h3c13e58c),
	.w5(32'hbb332de7),
	.w6(32'hbc004000),
	.w7(32'hbb743a4f),
	.w8(32'hbacf1c33),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf060ee),
	.w1(32'hbaa8468a),
	.w2(32'hbc035721),
	.w3(32'hbbaa1a94),
	.w4(32'h3c6ab7af),
	.w5(32'h39d0619f),
	.w6(32'h3c6d84ca),
	.w7(32'h3b23a679),
	.w8(32'h3cb2ed65),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fe754),
	.w1(32'hbb360646),
	.w2(32'hbcae737d),
	.w3(32'hbaffd1a4),
	.w4(32'hbbbc8917),
	.w5(32'hbc15f869),
	.w6(32'h3bc1c13c),
	.w7(32'h3a0862e1),
	.w8(32'hbb214c40),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac54972),
	.w1(32'hbc1fe929),
	.w2(32'hbb8bcbf1),
	.w3(32'hbb926c4e),
	.w4(32'h3c0ddb78),
	.w5(32'hbc048720),
	.w6(32'h3d3b09a7),
	.w7(32'hbc1f7045),
	.w8(32'hbc876ae8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc302f45),
	.w1(32'h3c053753),
	.w2(32'h3aadfb07),
	.w3(32'hbb937ed7),
	.w4(32'hbbffd727),
	.w5(32'h3bcc9cbe),
	.w6(32'hbb722025),
	.w7(32'h3b9622de),
	.w8(32'h3bed6e8d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bcf88),
	.w1(32'hbb4717b7),
	.w2(32'h3bc8e787),
	.w3(32'hb9a9e238),
	.w4(32'hbb9e2aa8),
	.w5(32'hbb2fde87),
	.w6(32'hb9ae8881),
	.w7(32'hbb9718ae),
	.w8(32'h3a4219c5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98b613),
	.w1(32'hbc3a831b),
	.w2(32'h3b1dab92),
	.w3(32'hbba67e0b),
	.w4(32'hb9e87750),
	.w5(32'hbc256332),
	.w6(32'h3c27d7ff),
	.w7(32'h3b94e94f),
	.w8(32'h3bbd2dc5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58c32b),
	.w1(32'h3b6dbbe0),
	.w2(32'hbb2c45e9),
	.w3(32'h3bbfa04c),
	.w4(32'hbc226711),
	.w5(32'hbbeaf143),
	.w6(32'hbc1e264f),
	.w7(32'hbc08ecb9),
	.w8(32'hbad4075a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f4afb),
	.w1(32'h3a7b8f5b),
	.w2(32'h3c5c6626),
	.w3(32'h3b8efbde),
	.w4(32'h3c9d4c93),
	.w5(32'h3ab7babc),
	.w6(32'hbbd0fb13),
	.w7(32'hbc3d1f56),
	.w8(32'hbbec96c5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70e130),
	.w1(32'h3b8f5d54),
	.w2(32'hbb731f97),
	.w3(32'hba8062e4),
	.w4(32'h3bb9658a),
	.w5(32'hbbb7a959),
	.w6(32'hbbcf1d16),
	.w7(32'hbb8f5a98),
	.w8(32'hbbdecf12),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5426d8),
	.w1(32'hb9060869),
	.w2(32'hbc1abeb1),
	.w3(32'h3b78e740),
	.w4(32'hb8c587e8),
	.w5(32'h3b23ee7b),
	.w6(32'hbc835a57),
	.w7(32'h3bf2c9c9),
	.w8(32'hbd0e0bc0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d228cef),
	.w1(32'hbaca441e),
	.w2(32'h3bd60bc6),
	.w3(32'hbc32d890),
	.w4(32'h3c59f78d),
	.w5(32'h3cae5544),
	.w6(32'hbb8f849f),
	.w7(32'hbc134b40),
	.w8(32'hbb1fcc18),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba61bb6),
	.w1(32'hbbbf2542),
	.w2(32'hbac90c54),
	.w3(32'h3bf3d564),
	.w4(32'hbb9c50d5),
	.w5(32'h3c597f2f),
	.w6(32'h3b6fddaf),
	.w7(32'hbbdf5843),
	.w8(32'hba7dd057),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb292d),
	.w1(32'hbc1d648c),
	.w2(32'h3c973723),
	.w3(32'hbc00d447),
	.w4(32'hbbb5d42a),
	.w5(32'hbb87fe3d),
	.w6(32'hba84870d),
	.w7(32'hbbf8d7a8),
	.w8(32'hbc847ace),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cf7a2),
	.w1(32'h3b087f68),
	.w2(32'h3b6df9e6),
	.w3(32'hbb1be06c),
	.w4(32'h3ae0cae5),
	.w5(32'hbb9898ff),
	.w6(32'h3bb176fc),
	.w7(32'h3c6e31cc),
	.w8(32'hbc146d39),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1943f),
	.w1(32'h3acb355f),
	.w2(32'hb7c595ba),
	.w3(32'h3c08aed1),
	.w4(32'hbab41e9a),
	.w5(32'hbad6ac1c),
	.w6(32'hbba6298c),
	.w7(32'h3c7150ac),
	.w8(32'hb9bfb91a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64419f),
	.w1(32'hbc78fb4b),
	.w2(32'hbcbf1823),
	.w3(32'h3bf85442),
	.w4(32'h3a311dcd),
	.w5(32'hbc0a4ddc),
	.w6(32'h3ca29abf),
	.w7(32'h3ba6bce6),
	.w8(32'hbaa21374),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c8fe),
	.w1(32'hbc8dfead),
	.w2(32'hbc8398de),
	.w3(32'h3bd0ea4f),
	.w4(32'h3a887885),
	.w5(32'hbc298f3f),
	.w6(32'hbc25c557),
	.w7(32'h3c49c20b),
	.w8(32'hba4bd8d9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b901299),
	.w1(32'h3c2eac4f),
	.w2(32'h3badc10a),
	.w3(32'h39780ccb),
	.w4(32'h3c569f39),
	.w5(32'h3b83eaad),
	.w6(32'h3c13ebd2),
	.w7(32'h3b3a1028),
	.w8(32'hbb0bc690),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae61bca),
	.w1(32'h3add9bb8),
	.w2(32'hbb2e23d3),
	.w3(32'h3a57dd0f),
	.w4(32'hbbce6d24),
	.w5(32'hba018e98),
	.w6(32'hbd30f63c),
	.w7(32'hbc4222c5),
	.w8(32'hbc5d8aa5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfba8ba),
	.w1(32'h3b0ff28c),
	.w2(32'h3b7c5481),
	.w3(32'hb9f5c497),
	.w4(32'hbb0705b6),
	.w5(32'hbbfab181),
	.w6(32'h3b584ee7),
	.w7(32'h3a30ca9d),
	.w8(32'h3c2931ac),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0824f2),
	.w1(32'hbab30022),
	.w2(32'hbbc78a84),
	.w3(32'hbbd2ba50),
	.w4(32'h3b85707e),
	.w5(32'h3cab8150),
	.w6(32'h3a34835f),
	.w7(32'hba1c5d6c),
	.w8(32'h3b054308),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7da31),
	.w1(32'h3bed5e42),
	.w2(32'hbd30cc89),
	.w3(32'h3ba2e157),
	.w4(32'h39d50034),
	.w5(32'hbd47bbed),
	.w6(32'hba65d3ef),
	.w7(32'hbc2c5ca6),
	.w8(32'hbcce8ef4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994587),
	.w1(32'hbc23a6d6),
	.w2(32'hbc235317),
	.w3(32'h389f13c8),
	.w4(32'hbbd3ba80),
	.w5(32'hbbde2cb6),
	.w6(32'hbb1bc3c4),
	.w7(32'h3c612220),
	.w8(32'h3b8a6ba5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00bbd9),
	.w1(32'hbc1af55b),
	.w2(32'hbbdf15f7),
	.w3(32'h3c35cc1c),
	.w4(32'h3b634682),
	.w5(32'hbc867c35),
	.w6(32'hbb17a2dc),
	.w7(32'h3bb9b2ec),
	.w8(32'h3bc23d62),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2cbb),
	.w1(32'hbbf6411b),
	.w2(32'h3a819fd4),
	.w3(32'h3d3d9de4),
	.w4(32'h3c2aa42c),
	.w5(32'h3bad78b8),
	.w6(32'hbbced4ab),
	.w7(32'hbc179688),
	.w8(32'hbb29908c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284f64),
	.w1(32'h3b926ded),
	.w2(32'h3bd8e4b6),
	.w3(32'h38a834b9),
	.w4(32'h3bc5d453),
	.w5(32'hbb52599f),
	.w6(32'hbbd23521),
	.w7(32'hbc26ac79),
	.w8(32'hbd03a87d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a9bc),
	.w1(32'h3996cf41),
	.w2(32'hbbcfc6f3),
	.w3(32'h3b267210),
	.w4(32'hbbbfc3bc),
	.w5(32'hbabdd75f),
	.w6(32'h3b9b86dd),
	.w7(32'hbb660bcf),
	.w8(32'h3b02b314),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0875c),
	.w1(32'h3b96565f),
	.w2(32'hba9fcf28),
	.w3(32'h3b7dc642),
	.w4(32'h3b19fa50),
	.w5(32'h3bb46f90),
	.w6(32'h3b459812),
	.w7(32'hbbdf7652),
	.w8(32'h3babb1f9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53df3b),
	.w1(32'h3b35ef4a),
	.w2(32'h3ad6913b),
	.w3(32'h3cc60a68),
	.w4(32'hbc2dcb45),
	.w5(32'h3c50e99a),
	.w6(32'h3b002c51),
	.w7(32'hbbb301bf),
	.w8(32'h3a3a04c7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcccd0b),
	.w1(32'hbb1b0d1a),
	.w2(32'hba2b43f0),
	.w3(32'hbb167a99),
	.w4(32'hbb316629),
	.w5(32'hbb823ba4),
	.w6(32'h3afa2402),
	.w7(32'hbbbda065),
	.w8(32'hbad891f2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ce955),
	.w1(32'hbc20188d),
	.w2(32'hbca7cb81),
	.w3(32'hba8ed90c),
	.w4(32'hbc50f1cd),
	.w5(32'hbcb91c08),
	.w6(32'hba8641da),
	.w7(32'h3b4f033a),
	.w8(32'h3c52471e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd19873),
	.w1(32'hbc11cd33),
	.w2(32'hbc4f81c6),
	.w3(32'h3b95d354),
	.w4(32'h3bb2217e),
	.w5(32'h3b0825c8),
	.w6(32'hb9cc78b4),
	.w7(32'h3bfd184d),
	.w8(32'h3b31995e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc0fd8),
	.w1(32'hbab2837e),
	.w2(32'h3ba7b3c4),
	.w3(32'h39c4de42),
	.w4(32'h3c1c36a2),
	.w5(32'h3c251601),
	.w6(32'h3bc657e8),
	.w7(32'h3b9945d0),
	.w8(32'hbc57b8a9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10e52b),
	.w1(32'hbb79fc26),
	.w2(32'hbb238c20),
	.w3(32'hbc3a00a3),
	.w4(32'h3a88016c),
	.w5(32'hbc7264f4),
	.w6(32'h3a647550),
	.w7(32'h3b724e13),
	.w8(32'hbb7dfc9d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43746a),
	.w1(32'h3abbffca),
	.w2(32'hbca547fc),
	.w3(32'h3c56d5db),
	.w4(32'h3b7a350b),
	.w5(32'hbc6031d9),
	.w6(32'h3a5ba630),
	.w7(32'hbb9b52a1),
	.w8(32'hbc460ecc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b57c2),
	.w1(32'h3b100868),
	.w2(32'hbc910347),
	.w3(32'h3b78aa58),
	.w4(32'hbb2d5648),
	.w5(32'hbab4f85c),
	.w6(32'hb9cc65aa),
	.w7(32'h3b80daab),
	.w8(32'hbbcc0f07),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25ff5f),
	.w1(32'hb9e9eec5),
	.w2(32'h3b3acf0a),
	.w3(32'hba225300),
	.w4(32'hbd6799f1),
	.w5(32'hbb710e7f),
	.w6(32'hbc2d2724),
	.w7(32'h3b626624),
	.w8(32'h39f2c982),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf50218),
	.w1(32'h3bcd2a00),
	.w2(32'h3b4a50e4),
	.w3(32'hbb1066ed),
	.w4(32'hbb86811c),
	.w5(32'hbaa192a0),
	.w6(32'h3ba38e0c),
	.w7(32'hbbc46710),
	.w8(32'hb980a1ff),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57e9b9),
	.w1(32'h3bb5ce5c),
	.w2(32'h3bc37f91),
	.w3(32'h3c0be349),
	.w4(32'h3c5f112b),
	.w5(32'hbae83956),
	.w6(32'hba9463a4),
	.w7(32'h3c314fca),
	.w8(32'hbbc9f357),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde07da),
	.w1(32'hb8f78261),
	.w2(32'hbbe37031),
	.w3(32'h3aa2dd15),
	.w4(32'hbbb91fe6),
	.w5(32'hbaee07ca),
	.w6(32'hbb5a4618),
	.w7(32'h3bc9b5ab),
	.w8(32'h3b538dea),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed4a6),
	.w1(32'hbb0302b9),
	.w2(32'hbab8a72c),
	.w3(32'h3a835231),
	.w4(32'h38ce12d4),
	.w5(32'hbce1cea3),
	.w6(32'hbcbeff6c),
	.w7(32'hbc1627ab),
	.w8(32'hb80c2b62),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d331),
	.w1(32'h3ac3c771),
	.w2(32'hbba76be0),
	.w3(32'h3b83076c),
	.w4(32'hbc8b80f0),
	.w5(32'h3b0797a1),
	.w6(32'h3b0d7955),
	.w7(32'hbc2918d5),
	.w8(32'hbb89fceb),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52c86f),
	.w1(32'h3ada5329),
	.w2(32'hbb490e49),
	.w3(32'hbba5eafd),
	.w4(32'h3b463543),
	.w5(32'hbb01bace),
	.w6(32'hbb2bf761),
	.w7(32'hb7dcca0e),
	.w8(32'h3bd656cf),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce5cba5),
	.w1(32'hbb440e5c),
	.w2(32'hbb8c4478),
	.w3(32'h3a77535e),
	.w4(32'hba32df42),
	.w5(32'h3b4c7874),
	.w6(32'h3a661ad3),
	.w7(32'hbc3d681d),
	.w8(32'hbc1483a8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a7f9),
	.w1(32'h3ba8262f),
	.w2(32'hbb3b5cf6),
	.w3(32'hbbb57cae),
	.w4(32'hbb93dd01),
	.w5(32'hbc1d03ca),
	.w6(32'h3b7a0e75),
	.w7(32'h3a61253c),
	.w8(32'h3c361188),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7c16),
	.w1(32'hbbbe6013),
	.w2(32'hbb10d7ac),
	.w3(32'h3bce7a91),
	.w4(32'hbbe68e16),
	.w5(32'hbc81eca8),
	.w6(32'h3c088cea),
	.w7(32'hbbcf1694),
	.w8(32'hbad34673),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506423),
	.w1(32'hbb5c3b9f),
	.w2(32'hbbb1a5a3),
	.w3(32'hbc23e381),
	.w4(32'hbb654f56),
	.w5(32'h3b2d0958),
	.w6(32'hbbd23ce9),
	.w7(32'hbb69f4f6),
	.w8(32'hbb10eaf7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac02c18),
	.w1(32'h3b546742),
	.w2(32'hbb006861),
	.w3(32'hbb4b559a),
	.w4(32'hbcc2b795),
	.w5(32'h3a09aa16),
	.w6(32'h3ac35788),
	.w7(32'hbbb56226),
	.w8(32'h3c640c42),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d8c0ef),
	.w1(32'h3a8451eb),
	.w2(32'h3b9990d0),
	.w3(32'hbb5c5708),
	.w4(32'hbb766e9c),
	.w5(32'hbb32a94b),
	.w6(32'h3b4387c5),
	.w7(32'hbbd1e0b6),
	.w8(32'h3cbe7039),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda193a),
	.w1(32'hba6cb1a4),
	.w2(32'h3be4ac70),
	.w3(32'hbd6be1b6),
	.w4(32'h3a609794),
	.w5(32'hbbcb790b),
	.w6(32'hbb7e376f),
	.w7(32'hbbb2927b),
	.w8(32'hbcd3006b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20ea2e),
	.w1(32'hbc3da177),
	.w2(32'h3ae21e88),
	.w3(32'h3c626004),
	.w4(32'hba3b4fb2),
	.w5(32'hba27f525),
	.w6(32'h3bd7a139),
	.w7(32'h3bc181f1),
	.w8(32'h3c134477),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ffff0),
	.w1(32'hbb38382c),
	.w2(32'h3b748fc1),
	.w3(32'h3b6ced9e),
	.w4(32'h3b2c8d40),
	.w5(32'hbc1d50f9),
	.w6(32'hbc54b1d8),
	.w7(32'hb98ef4c9),
	.w8(32'hbb8f9657),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60803d),
	.w1(32'hb9cf6311),
	.w2(32'hba3f4c6d),
	.w3(32'h3b07ed47),
	.w4(32'h3bb91544),
	.w5(32'hbbe18fa3),
	.w6(32'h3cf5ebb1),
	.w7(32'hbb61eede),
	.w8(32'h3bb181e7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42754c),
	.w1(32'hbbb6e1ed),
	.w2(32'hbc134d2b),
	.w3(32'hbb02a85c),
	.w4(32'h3b523ec2),
	.w5(32'h3a339ff5),
	.w6(32'h3b3a2395),
	.w7(32'hbb9bb019),
	.w8(32'h3a94d106),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eea0f),
	.w1(32'h3c257579),
	.w2(32'hbaf8b97c),
	.w3(32'hbb2f2d5b),
	.w4(32'h3aaa9a1b),
	.w5(32'hbb8b834a),
	.w6(32'hbd9241e0),
	.w7(32'hbc292517),
	.w8(32'hbb02e382),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082d6c),
	.w1(32'hba23a6b6),
	.w2(32'hbc23e026),
	.w3(32'hbc8a1e57),
	.w4(32'h3c2e7c4b),
	.w5(32'hbba8bb28),
	.w6(32'h39e0e692),
	.w7(32'h3b1e1e08),
	.w8(32'hbab80838),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c744730),
	.w1(32'hbb2f0b4a),
	.w2(32'h3b7b22a7),
	.w3(32'h3aac474d),
	.w4(32'hbc468c91),
	.w5(32'h3be0c581),
	.w6(32'hbb852e3a),
	.w7(32'hbc8b16e9),
	.w8(32'h3b6ed16e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750c17),
	.w1(32'hbc7c7e35),
	.w2(32'h3ca7ecc3),
	.w3(32'hbb76fbfc),
	.w4(32'hbc090a49),
	.w5(32'h3b42aa8d),
	.w6(32'h3c0da9bb),
	.w7(32'h3b232d02),
	.w8(32'h3c865a12),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1082c5),
	.w1(32'h3a41d0ed),
	.w2(32'hb76c1731),
	.w3(32'hba7db65c),
	.w4(32'hbb8a5150),
	.w5(32'h3b3308dd),
	.w6(32'hbb00d0f8),
	.w7(32'h39e90f1d),
	.w8(32'hbc1670e4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38766d05),
	.w1(32'hbc7e656d),
	.w2(32'hbbfccb86),
	.w3(32'h3cbe8461),
	.w4(32'h3bf78a88),
	.w5(32'h39830e64),
	.w6(32'hbb58acbf),
	.w7(32'h3b5f5f5b),
	.w8(32'h398f4dc2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule