module layer_10_featuremap_497(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39020ae4),
	.w1(32'h3a8db83f),
	.w2(32'h3a4ac3eb),
	.w3(32'hb959f057),
	.w4(32'h3b692403),
	.w5(32'hbb09d580),
	.w6(32'h3a38b80f),
	.w7(32'h3be76965),
	.w8(32'h3a2b64bf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6438a),
	.w1(32'hb8bb6598),
	.w2(32'hbae92b99),
	.w3(32'h39cdadac),
	.w4(32'h3959aceb),
	.w5(32'hbb091887),
	.w6(32'hbb44db6e),
	.w7(32'hbba4ad5f),
	.w8(32'hbbae2b84),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfab6e6),
	.w1(32'hb9e88a05),
	.w2(32'hbb65b47a),
	.w3(32'hba5d92b0),
	.w4(32'h3bc84e81),
	.w5(32'h3a4ccd4d),
	.w6(32'h3a85ca49),
	.w7(32'hbc12732a),
	.w8(32'hbc2cee98),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03178d),
	.w1(32'hbc26c0a5),
	.w2(32'hbb392154),
	.w3(32'h3ac27b84),
	.w4(32'hbb8867f5),
	.w5(32'h3ce665e3),
	.w6(32'hbb37ce5b),
	.w7(32'h3b0035fb),
	.w8(32'h3c03d030),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409539),
	.w1(32'h3ab74ce4),
	.w2(32'hbb05fe3c),
	.w3(32'hba027b94),
	.w4(32'h3ab54445),
	.w5(32'hbbda1c70),
	.w6(32'h3b124bf1),
	.w7(32'hb9b73a15),
	.w8(32'hbb82888f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3762b),
	.w1(32'h3b22791d),
	.w2(32'hbbd7259f),
	.w3(32'hbbc0a0df),
	.w4(32'hbbf63355),
	.w5(32'hbbc387da),
	.w6(32'hba28ef4e),
	.w7(32'hbb9081ce),
	.w8(32'hbb9e7ac9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc73f04),
	.w1(32'h3ba45909),
	.w2(32'h3c321b1c),
	.w3(32'hb9b290bf),
	.w4(32'h3c9c36a6),
	.w5(32'h3cb85a1a),
	.w6(32'h3b6ae87e),
	.w7(32'h39a6efe8),
	.w8(32'h3b2fa4f3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051a17),
	.w1(32'h3b0f5ea1),
	.w2(32'h3b8c0b5a),
	.w3(32'h3c9b79b6),
	.w4(32'h3bb94065),
	.w5(32'hbbccecd8),
	.w6(32'hba4431bc),
	.w7(32'h3b6a99b5),
	.w8(32'hbb5b27ac),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87127),
	.w1(32'hbb80e642),
	.w2(32'h3b815bda),
	.w3(32'h3b6665eb),
	.w4(32'hbc37f51f),
	.w5(32'h3c55d7e8),
	.w6(32'h3b98ffde),
	.w7(32'hbb46f83a),
	.w8(32'h3b8e5b93),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb710fe),
	.w1(32'h3b210243),
	.w2(32'h3bcdccf5),
	.w3(32'hbbc8c070),
	.w4(32'h3c67f2ec),
	.w5(32'h3cc2870f),
	.w6(32'hbc3287f4),
	.w7(32'h3b9473b4),
	.w8(32'h3bf54c56),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b7b82),
	.w1(32'hbb5f2ef0),
	.w2(32'h3aa9c248),
	.w3(32'h3c0f787f),
	.w4(32'h3ae890f0),
	.w5(32'h39d6edab),
	.w6(32'h3c12b532),
	.w7(32'hbb04eabf),
	.w8(32'hbaad2f55),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4c7e),
	.w1(32'h3bb82d28),
	.w2(32'h3bd8414d),
	.w3(32'hbb30e971),
	.w4(32'hba142830),
	.w5(32'h3a64c8d4),
	.w6(32'hbb01f6bf),
	.w7(32'hbc288964),
	.w8(32'hbbb24ab2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e528),
	.w1(32'h3c7e1f4d),
	.w2(32'hbbaec684),
	.w3(32'hbbf70832),
	.w4(32'hbb204181),
	.w5(32'hbbaf2adb),
	.w6(32'hbc30145f),
	.w7(32'hbb8273d4),
	.w8(32'hbbf90652),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b02c0),
	.w1(32'h3c26c6d3),
	.w2(32'hbae6aebb),
	.w3(32'h3b8e35e4),
	.w4(32'h3bc725b4),
	.w5(32'h39e1fbae),
	.w6(32'h3be4cf86),
	.w7(32'h3c39aade),
	.w8(32'h3b98cd9d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86f346),
	.w1(32'hbb1030a5),
	.w2(32'hbc0e9455),
	.w3(32'h3bb9ff0c),
	.w4(32'h3b8e7128),
	.w5(32'hbc41fd30),
	.w6(32'h3a214a2f),
	.w7(32'h3aa08c77),
	.w8(32'hbc231eea),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ab4b6),
	.w1(32'h3c40ad26),
	.w2(32'hbb939a47),
	.w3(32'h3b791466),
	.w4(32'h3c2935d6),
	.w5(32'hbc53a43b),
	.w6(32'hbb762574),
	.w7(32'h3b09fb0f),
	.w8(32'hbc47a944),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10f474),
	.w1(32'h3bf37859),
	.w2(32'h3b93aece),
	.w3(32'hbb8fd156),
	.w4(32'h3b99f1c8),
	.w5(32'hbb16f525),
	.w6(32'h39ae71be),
	.w7(32'hbc5b0894),
	.w8(32'hbbe7ae7e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae37ff7),
	.w1(32'hbab07708),
	.w2(32'h3c79d633),
	.w3(32'hbb30c08a),
	.w4(32'hbbaa9403),
	.w5(32'h3b448023),
	.w6(32'hbc0be83f),
	.w7(32'hbad92021),
	.w8(32'h3b1f4c55),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86565b),
	.w1(32'h3c8f6106),
	.w2(32'h3c36acb3),
	.w3(32'hbc3ce1e8),
	.w4(32'h3b22fb1d),
	.w5(32'hbac73a89),
	.w6(32'hbc09641b),
	.w7(32'hbbb711d3),
	.w8(32'hba7a21ce),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd47a),
	.w1(32'h3ba2810d),
	.w2(32'hbb9ca00e),
	.w3(32'hba33da93),
	.w4(32'h3bd229f4),
	.w5(32'hbc35a410),
	.w6(32'hbb88be35),
	.w7(32'hbc001e03),
	.w8(32'hbc9f208e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd12b9c),
	.w1(32'h3b849fa3),
	.w2(32'hbb72e95f),
	.w3(32'hbbb29fd2),
	.w4(32'hbbb9548d),
	.w5(32'hbbcf46fa),
	.w6(32'hbc0adb66),
	.w7(32'hbc0f7925),
	.w8(32'hbaff5749),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e9ba8),
	.w1(32'h3ba9f59d),
	.w2(32'hbc7fa51e),
	.w3(32'h3b85c8ad),
	.w4(32'h3a1e4931),
	.w5(32'hbc67c1f3),
	.w6(32'h39f459ac),
	.w7(32'h3b774a07),
	.w8(32'hbc305555),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16fff7),
	.w1(32'h3aa2f8f9),
	.w2(32'h3bdded35),
	.w3(32'hbbaf51ad),
	.w4(32'h3bea39d3),
	.w5(32'h3d025ec3),
	.w6(32'hbb74bc50),
	.w7(32'h3b01c9e2),
	.w8(32'h3c6f21b7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7348d9),
	.w1(32'h3bd5e136),
	.w2(32'hbbbe95a9),
	.w3(32'h3c9b517b),
	.w4(32'hbb8b9de8),
	.w5(32'hbc188b70),
	.w6(32'hbbc48fbc),
	.w7(32'h3a54ed91),
	.w8(32'hbb3f59fb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4c046),
	.w1(32'hbbc30694),
	.w2(32'h3c90c7c4),
	.w3(32'h3a8e82f3),
	.w4(32'hbbbaaa20),
	.w5(32'h3c055c73),
	.w6(32'h39e463af),
	.w7(32'h3c36b451),
	.w8(32'h3a8bb623),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99936be),
	.w1(32'hbb4cb3aa),
	.w2(32'hbc07f16f),
	.w3(32'hba0084d9),
	.w4(32'hbbaf9094),
	.w5(32'hbc22f673),
	.w6(32'h3a4a7f10),
	.w7(32'h3afdca4c),
	.w8(32'h3a3fc80c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d21be2),
	.w1(32'hbb287681),
	.w2(32'hbb3e5242),
	.w3(32'h3b8508f7),
	.w4(32'hbb8176a0),
	.w5(32'h3c4ec5c3),
	.w6(32'h3c87c0e5),
	.w7(32'h39a96339),
	.w8(32'hba39d365),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb63f00),
	.w1(32'h3adfc94b),
	.w2(32'h3c335d08),
	.w3(32'h3bf585a1),
	.w4(32'hbb2be869),
	.w5(32'h3c20ecb4),
	.w6(32'h3b0d5b0f),
	.w7(32'hbb19c519),
	.w8(32'h3c5c6bb1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4122f5),
	.w1(32'h3b42478e),
	.w2(32'h3d41769e),
	.w3(32'h3c94760d),
	.w4(32'h3d206c81),
	.w5(32'h3d098e33),
	.w6(32'h3c189e54),
	.w7(32'h3c7da4f6),
	.w8(32'h3c1e9b3a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81377c),
	.w1(32'h399af71e),
	.w2(32'hbba3f8a2),
	.w3(32'h3c4566ef),
	.w4(32'h3a817317),
	.w5(32'hb9403040),
	.w6(32'h3bcf63f5),
	.w7(32'hbba5de90),
	.w8(32'hbbc1c842),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ea30),
	.w1(32'hbae3cd49),
	.w2(32'h3bdcd7a9),
	.w3(32'h3c06b370),
	.w4(32'h3c0aaae1),
	.w5(32'hbb5d0e8c),
	.w6(32'hba354993),
	.w7(32'hbb6b2f84),
	.w8(32'hbb998eba),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13a46f),
	.w1(32'hbb3a6188),
	.w2(32'hbbae471a),
	.w3(32'h3c35b1b0),
	.w4(32'hbba67a77),
	.w5(32'hbba94008),
	.w6(32'hbbac23f9),
	.w7(32'hbba17851),
	.w8(32'h3a137650),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd29e49),
	.w1(32'h3bc2efd9),
	.w2(32'hbaea1ab9),
	.w3(32'hbb2ecc2e),
	.w4(32'h3b2c73e6),
	.w5(32'hba186e6a),
	.w6(32'h3b327d48),
	.w7(32'hb9c5712d),
	.w8(32'h3b760798),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b58928),
	.w1(32'hbb5bf49d),
	.w2(32'hbb2e4289),
	.w3(32'h3b81c703),
	.w4(32'hbc2bb046),
	.w5(32'hbb7c4c19),
	.w6(32'h39797532),
	.w7(32'h3b4a1b3d),
	.w8(32'h3c2cea37),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc3acc),
	.w1(32'h3b8b324a),
	.w2(32'hbbd08bf5),
	.w3(32'h3c7fc588),
	.w4(32'hbbabbc0c),
	.w5(32'hbcca2314),
	.w6(32'h3a45e81f),
	.w7(32'h3a9181b8),
	.w8(32'hbb075cc5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6ca3a),
	.w1(32'hbc5e4f10),
	.w2(32'hbb27c791),
	.w3(32'h3b3f5ac6),
	.w4(32'hbc11a9cc),
	.w5(32'h3bbcd701),
	.w6(32'h3c0904df),
	.w7(32'hbb3e8ca9),
	.w8(32'h3b3b93ad),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dd0c21),
	.w1(32'hbc225271),
	.w2(32'h3c016862),
	.w3(32'h38ba0a77),
	.w4(32'hbc048a07),
	.w5(32'h3c91c322),
	.w6(32'hbad7d6d7),
	.w7(32'hbbe21b2c),
	.w8(32'hba8acbb4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c470847),
	.w1(32'h3ab5aedb),
	.w2(32'hbb8d59c1),
	.w3(32'hbb9d76a9),
	.w4(32'hbbc90097),
	.w5(32'hbba0544e),
	.w6(32'hbc4ef51c),
	.w7(32'hbc75c151),
	.w8(32'hbc4a3193),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae684b5),
	.w1(32'hb9ae0331),
	.w2(32'h3be3d65a),
	.w3(32'hbba5e59f),
	.w4(32'h3bba0665),
	.w5(32'hbada8e8d),
	.w6(32'hbb38e133),
	.w7(32'h3a93af32),
	.w8(32'hba25da1b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092885),
	.w1(32'hbb053fc1),
	.w2(32'hbb668850),
	.w3(32'h3b7620f8),
	.w4(32'hbb283d85),
	.w5(32'h3b8f4f8e),
	.w6(32'h3bdaf7bc),
	.w7(32'h3a38d558),
	.w8(32'h3aef1dc5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0d2d7),
	.w1(32'h3c31b56b),
	.w2(32'hbba7446b),
	.w3(32'h3b26ece4),
	.w4(32'h3c0b2a07),
	.w5(32'h3b6ef94a),
	.w6(32'h3b49294e),
	.w7(32'hba96493d),
	.w8(32'h3b5532f4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3269b5),
	.w1(32'h3a0873c9),
	.w2(32'hbb655a2f),
	.w3(32'h3b45ad24),
	.w4(32'hbb6f8e26),
	.w5(32'h3c283e0e),
	.w6(32'hbb8aaf8a),
	.w7(32'hbb9a1967),
	.w8(32'hbaaad5e0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32a3fa),
	.w1(32'hbc0274b2),
	.w2(32'hbb7eec00),
	.w3(32'hbb28e8a4),
	.w4(32'hbb16a8d2),
	.w5(32'h3c977ca5),
	.w6(32'hbb86152d),
	.w7(32'hbb8abc3e),
	.w8(32'hbbc36067),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d40ad),
	.w1(32'h3c75b570),
	.w2(32'h3ce01d67),
	.w3(32'hbc97f909),
	.w4(32'h3c03edfa),
	.w5(32'h3c9d79e6),
	.w6(32'hbc3ea6b6),
	.w7(32'h3c192ac7),
	.w8(32'h3cf8737f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c310536),
	.w1(32'h3c04ed4f),
	.w2(32'h3ab8c5c9),
	.w3(32'h3c580ad8),
	.w4(32'h3b829cc2),
	.w5(32'h3c16d569),
	.w6(32'h3c173b04),
	.w7(32'hbbab73fb),
	.w8(32'hba98e373),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94777f),
	.w1(32'h3c2c6dc6),
	.w2(32'hbb8ff255),
	.w3(32'h3b8dc2aa),
	.w4(32'hbab892d6),
	.w5(32'hbc43aae8),
	.w6(32'h3ab4f870),
	.w7(32'hba248ee2),
	.w8(32'hbb23a9c1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ab100),
	.w1(32'h3c262a47),
	.w2(32'h396af5cb),
	.w3(32'hba6a3bff),
	.w4(32'hbb6f4fa2),
	.w5(32'h3b42d4c8),
	.w6(32'h3be90c39),
	.w7(32'hbbbb3d3e),
	.w8(32'hb9f9e4a8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e5d24),
	.w1(32'h3accdd01),
	.w2(32'h3c38c149),
	.w3(32'hbb8b670b),
	.w4(32'hba4bb899),
	.w5(32'h3ba31edc),
	.w6(32'h3bceafe0),
	.w7(32'h3ba31c38),
	.w8(32'h3c2aa240),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7ae64),
	.w1(32'hb767e641),
	.w2(32'h3c06e3ae),
	.w3(32'h3b5d41d3),
	.w4(32'h3b030d48),
	.w5(32'hbb8cb11c),
	.w6(32'h3ba1601d),
	.w7(32'h3bd3ba67),
	.w8(32'hbb6ddfeb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2110),
	.w1(32'hb9d1691b),
	.w2(32'hbbbbe9bb),
	.w3(32'hbb5b81b1),
	.w4(32'h3b2cbbe0),
	.w5(32'hbba76d7c),
	.w6(32'hb8cbbcd8),
	.w7(32'hb9bfe88f),
	.w8(32'hba56f241),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc138a74),
	.w1(32'h3c980c39),
	.w2(32'h3c35748d),
	.w3(32'hbbc5be44),
	.w4(32'h3c77f4f5),
	.w5(32'hbb92e519),
	.w6(32'h3b4d4342),
	.w7(32'h3c260d50),
	.w8(32'hbb950357),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab73bc8),
	.w1(32'h3ae1d47a),
	.w2(32'hbbef12ba),
	.w3(32'hbc042f86),
	.w4(32'hbb75ba29),
	.w5(32'h3993cee8),
	.w6(32'hbafdce46),
	.w7(32'hbb9f2727),
	.w8(32'h3b4b16d0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb598b25),
	.w1(32'hbbc87cd7),
	.w2(32'hbb8a15c6),
	.w3(32'hbc199b11),
	.w4(32'hbbbfe97d),
	.w5(32'h3b6fd26c),
	.w6(32'hbbf5cacf),
	.w7(32'hbbfdb011),
	.w8(32'hbb8f6ff0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6139),
	.w1(32'h3c09e700),
	.w2(32'hbada15c7),
	.w3(32'hbb417381),
	.w4(32'h3bcc6783),
	.w5(32'hbba1838d),
	.w6(32'hbbe1977b),
	.w7(32'h3bd9b804),
	.w8(32'h3c190bf9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf1756),
	.w1(32'hbb316011),
	.w2(32'h3b4b6dd6),
	.w3(32'h3b9be5d3),
	.w4(32'hbbe99235),
	.w5(32'h3a334e50),
	.w6(32'h3be725d4),
	.w7(32'hbc2afc36),
	.w8(32'hba07fed2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0d21),
	.w1(32'h3ad3fbc2),
	.w2(32'hbb0a7afe),
	.w3(32'hbba2fa60),
	.w4(32'hb9844bf1),
	.w5(32'h3b20852c),
	.w6(32'hbbcc1008),
	.w7(32'h3b95300b),
	.w8(32'h39e3c060),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecef23),
	.w1(32'h3c0e345c),
	.w2(32'h3b2c17ec),
	.w3(32'hba50c1ae),
	.w4(32'h3a25fe28),
	.w5(32'h3b8fdb15),
	.w6(32'hbb147978),
	.w7(32'hb91db28c),
	.w8(32'h3b1bf9c0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1975),
	.w1(32'hbbeccffd),
	.w2(32'hbc46ec09),
	.w3(32'hbb925e7c),
	.w4(32'hbc815560),
	.w5(32'hbbb875cb),
	.w6(32'hb92ac410),
	.w7(32'hbc106912),
	.w8(32'hbc24cae8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc388a5b),
	.w1(32'hbb0ff993),
	.w2(32'hb8c399ed),
	.w3(32'hbbec4af9),
	.w4(32'hbbda6086),
	.w5(32'hb9dd7b34),
	.w6(32'hbc1500e1),
	.w7(32'hbc028c84),
	.w8(32'hbc2bcc2d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19f054),
	.w1(32'hbbd7863d),
	.w2(32'hbba55e9b),
	.w3(32'h3ad81132),
	.w4(32'hbbec5fcf),
	.w5(32'hbc70124a),
	.w6(32'h3a999cfd),
	.w7(32'hbc2f6038),
	.w8(32'hbc41e798),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4a1ba),
	.w1(32'hbbec0905),
	.w2(32'hbbe78a27),
	.w3(32'hbbb045e5),
	.w4(32'hbc1ad8ce),
	.w5(32'hbb0f55e5),
	.w6(32'hbba7d703),
	.w7(32'hbbd74db8),
	.w8(32'hbbc3844f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8b25c),
	.w1(32'h3b4af77f),
	.w2(32'h3ba7b482),
	.w3(32'h3b91126f),
	.w4(32'h3b58e103),
	.w5(32'h3b98eb2f),
	.w6(32'h3b7a7446),
	.w7(32'hbbbe6d22),
	.w8(32'h3afaad09),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399498dd),
	.w1(32'hbb97ddff),
	.w2(32'h3b187d1f),
	.w3(32'hbaa9e46e),
	.w4(32'h3a9a7ba4),
	.w5(32'h3c7c4611),
	.w6(32'hbba2309c),
	.w7(32'h3afe9759),
	.w8(32'h3a105394),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd82d0),
	.w1(32'h3c760de7),
	.w2(32'h3bc958de),
	.w3(32'hbc1a415f),
	.w4(32'h3b7832f9),
	.w5(32'hbb9ae1d5),
	.w6(32'hbb90fe0c),
	.w7(32'hbb072fdf),
	.w8(32'hbbfb7c0d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39fcf3),
	.w1(32'h3c9a4a9c),
	.w2(32'h377bcdc1),
	.w3(32'hbc370e3f),
	.w4(32'h3c0c3fc7),
	.w5(32'hbc2c52c2),
	.w6(32'h3a75c1ce),
	.w7(32'h3c3e1657),
	.w8(32'hbaeb6731),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e9bda),
	.w1(32'hbc886fb9),
	.w2(32'hbc05b189),
	.w3(32'h3b5be13b),
	.w4(32'hbbec81ba),
	.w5(32'h3c32f7cb),
	.w6(32'h3bf51c65),
	.w7(32'hbae6711b),
	.w8(32'hbb7e2206),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e8bfe),
	.w1(32'h3ae6a7c6),
	.w2(32'h3b4bf661),
	.w3(32'hbc7019b6),
	.w4(32'hbbd2e6c4),
	.w5(32'h3b477b36),
	.w6(32'hbc5254a1),
	.w7(32'h39dc257b),
	.w8(32'h3ab2c185),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768aea),
	.w1(32'hba803a3e),
	.w2(32'h3c43c282),
	.w3(32'h3bf3445f),
	.w4(32'hbc124923),
	.w5(32'hbbd7717b),
	.w6(32'h3b3c5a7e),
	.w7(32'h3c34b0ac),
	.w8(32'hbb97d0f5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd450ac),
	.w1(32'h3c4cceee),
	.w2(32'h3cd26725),
	.w3(32'hbbd08212),
	.w4(32'h3cb5e849),
	.w5(32'h3b9e083b),
	.w6(32'hbbc08f35),
	.w7(32'h3c48586d),
	.w8(32'h3c75bedb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16c2cc),
	.w1(32'h3b397180),
	.w2(32'h3a3a2b78),
	.w3(32'hbbded5ef),
	.w4(32'h3a296e06),
	.w5(32'hbb1129fd),
	.w6(32'hbb2ede98),
	.w7(32'hba313f2f),
	.w8(32'hbb34d75d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3a962),
	.w1(32'hb95b9453),
	.w2(32'hb928f65d),
	.w3(32'h39628a21),
	.w4(32'hb7b1ca42),
	.w5(32'hb809f555),
	.w6(32'hb8aaaad8),
	.w7(32'h394ad688),
	.w8(32'h39c80dce),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd57f0),
	.w1(32'h39971c37),
	.w2(32'hb9d6b35f),
	.w3(32'hb8fd8213),
	.w4(32'h379b4713),
	.w5(32'h398aee00),
	.w6(32'h396555f3),
	.w7(32'hb93c5077),
	.w8(32'hb91bb6a0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92dcc51),
	.w1(32'hba1781e5),
	.w2(32'hb91e0cf3),
	.w3(32'h3962791a),
	.w4(32'hba1cc143),
	.w5(32'hb873dfbd),
	.w6(32'h38ad9506),
	.w7(32'hba1f62f6),
	.w8(32'hba62590d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba279758),
	.w1(32'hb700bcd9),
	.w2(32'h3a2545f3),
	.w3(32'hba764140),
	.w4(32'hba5a5251),
	.w5(32'hb8bb07d7),
	.w6(32'hba1a7176),
	.w7(32'hb97638cd),
	.w8(32'h39c73d4b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aab3ec),
	.w1(32'hb93bd551),
	.w2(32'hb943a7a6),
	.w3(32'hb942f23e),
	.w4(32'hb8d0b3ff),
	.w5(32'h391a938b),
	.w6(32'hb90b6cee),
	.w7(32'h390d3148),
	.w8(32'h3a0ddbcc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6887a9),
	.w1(32'h395f1ca6),
	.w2(32'h3ab63953),
	.w3(32'hba8aae24),
	.w4(32'hba7fc7ea),
	.w5(32'h37895954),
	.w6(32'hbaad1c45),
	.w7(32'hba79b045),
	.w8(32'hb8196ff2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d2a6),
	.w1(32'hba46d5ce),
	.w2(32'h3b5ce3d6),
	.w3(32'hbaf22e0d),
	.w4(32'hbb0e6821),
	.w5(32'h3a8b1a0d),
	.w6(32'h3a9627b7),
	.w7(32'h39cc13f7),
	.w8(32'h3ab2ee59),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49b2db),
	.w1(32'h3af5600f),
	.w2(32'h3ac239d5),
	.w3(32'h3a8939d9),
	.w4(32'h3a0c6b44),
	.w5(32'hb8e2d3fb),
	.w6(32'hba9c4b07),
	.w7(32'hba411fce),
	.w8(32'hba84777e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eec84c),
	.w1(32'h39d4fe9b),
	.w2(32'h3ae58378),
	.w3(32'hba535ad9),
	.w4(32'hb9a7596b),
	.w5(32'h3a84c1f2),
	.w6(32'hb97224ed),
	.w7(32'h397fda27),
	.w8(32'h3ab1769b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a8551),
	.w1(32'h39f737f6),
	.w2(32'h3b17d24f),
	.w3(32'hba987fb7),
	.w4(32'h38ea350c),
	.w5(32'h3b1e4bed),
	.w6(32'hbb25bdac),
	.w7(32'hba9f2655),
	.w8(32'hb8f496fc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d9761),
	.w1(32'h3a43bd3f),
	.w2(32'h3a8d3a21),
	.w3(32'h38aa42ef),
	.w4(32'hb972d4ef),
	.w5(32'h38860759),
	.w6(32'hba5645e8),
	.w7(32'hba49ec48),
	.w8(32'hb972189a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c53af8),
	.w1(32'h39a9cf1c),
	.w2(32'h3a9ed847),
	.w3(32'hba870f31),
	.w4(32'hba9b88f6),
	.w5(32'hb9c09670),
	.w6(32'hba6bc3ca),
	.w7(32'hba055dc2),
	.w8(32'h398548ac),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374d8887),
	.w1(32'h3923db19),
	.w2(32'h387333f2),
	.w3(32'hb81147a6),
	.w4(32'h38dc4309),
	.w5(32'h39083f6f),
	.w6(32'hb927c227),
	.w7(32'h368d76d7),
	.w8(32'h384ce8ab),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf4683),
	.w1(32'hb9de410d),
	.w2(32'h3900a681),
	.w3(32'h39eafbad),
	.w4(32'hb9218b7b),
	.w5(32'h3a01ded2),
	.w6(32'h399045a0),
	.w7(32'hb8e61852),
	.w8(32'hb9931b36),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a41b78),
	.w1(32'h38ce7b30),
	.w2(32'h39903d29),
	.w3(32'hb887feb3),
	.w4(32'h393b3912),
	.w5(32'hb8b6adab),
	.w6(32'h3843df0b),
	.w7(32'h38663615),
	.w8(32'hb7b5cb3a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c5a0c),
	.w1(32'hba971c25),
	.w2(32'hba130461),
	.w3(32'h398c7e3f),
	.w4(32'hb98571af),
	.w5(32'hba1e8d0d),
	.w6(32'h398c3e44),
	.w7(32'hb8416705),
	.w8(32'hb8efdaa7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada0da4),
	.w1(32'hb87000fd),
	.w2(32'hb9ba0bc1),
	.w3(32'h39dec8d0),
	.w4(32'h38949ce5),
	.w5(32'hba8f4492),
	.w6(32'hba631b12),
	.w7(32'hba4b5811),
	.w8(32'hbaec1a0e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ffce65),
	.w1(32'hb928f776),
	.w2(32'h399f408a),
	.w3(32'h38cafb8b),
	.w4(32'h3927bb28),
	.w5(32'h3a277a13),
	.w6(32'h39b97af6),
	.w7(32'hb8a98e96),
	.w8(32'h39a68919),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaee69),
	.w1(32'h3abd6eb7),
	.w2(32'h3acac538),
	.w3(32'h3a8fbc7a),
	.w4(32'hb9ceae50),
	.w5(32'hb984786b),
	.w6(32'h3a9963a2),
	.w7(32'h3a0a2abf),
	.w8(32'h3a1282fb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d42d),
	.w1(32'h39a88f4d),
	.w2(32'h3b0fa0ee),
	.w3(32'hbb7778d5),
	.w4(32'hbb4c0f95),
	.w5(32'hba808ed8),
	.w6(32'hbb0063a6),
	.w7(32'hbaa26991),
	.w8(32'hb937df1f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e78c4),
	.w1(32'h396a3c6b),
	.w2(32'hbb231fa5),
	.w3(32'h3a583cc2),
	.w4(32'hb997d4c7),
	.w5(32'hbb5206f9),
	.w6(32'hb9d8899e),
	.w7(32'hbb36cee4),
	.w8(32'hbb9a42f5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc2a06),
	.w1(32'h3a692116),
	.w2(32'h3bb284b7),
	.w3(32'hba66ee02),
	.w4(32'hb8aded8b),
	.w5(32'h3b7e06db),
	.w6(32'hbb381b0f),
	.w7(32'hbb3bab8f),
	.w8(32'h3ac70f88),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d24b13),
	.w1(32'hba93e0ec),
	.w2(32'hbb3aa7fc),
	.w3(32'hb88fe7ad),
	.w4(32'hbb148d70),
	.w5(32'hbb80792a),
	.w6(32'hb969f9db),
	.w7(32'hbb356fe5),
	.w8(32'hbb8a08d8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f53c9),
	.w1(32'h3b3df924),
	.w2(32'h3be49a9f),
	.w3(32'hbb2cf41e),
	.w4(32'h397093bc),
	.w5(32'h3b9104d8),
	.w6(32'hba80c174),
	.w7(32'h3ac83c33),
	.w8(32'h3b92e61e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a529680),
	.w1(32'h3aa1653c),
	.w2(32'h3abd8f99),
	.w3(32'hba3c7c94),
	.w4(32'h3a52e342),
	.w5(32'h3a39c133),
	.w6(32'hbaba37d6),
	.w7(32'hba06abe6),
	.w8(32'hba67a4f4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98be39),
	.w1(32'hb8cc9efc),
	.w2(32'hbaf34afa),
	.w3(32'hba8beedd),
	.w4(32'hba23646f),
	.w5(32'hbb6fa996),
	.w6(32'hbab51a79),
	.w7(32'hbb0d0c8c),
	.w8(32'hbb98c999),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8baacac),
	.w1(32'h38f62ecc),
	.w2(32'h3900135f),
	.w3(32'h39c880d3),
	.w4(32'h39731b9d),
	.w5(32'hb7e97499),
	.w6(32'h3a0aa5cb),
	.w7(32'h398c330d),
	.w8(32'h39cc31b6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabcb7b),
	.w1(32'h3b37ddae),
	.w2(32'h3b918c8c),
	.w3(32'hba608eb9),
	.w4(32'hb981ff1b),
	.w5(32'h3b050047),
	.w6(32'h39616f05),
	.w7(32'h388eff40),
	.w8(32'h3b3cbb45),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7d4f2),
	.w1(32'h3a4d52b4),
	.w2(32'h3b035eed),
	.w3(32'hbaaf8527),
	.w4(32'hb9e045f2),
	.w5(32'h3a7897d6),
	.w6(32'hbb8d559b),
	.w7(32'hbb749420),
	.w8(32'hbaf227fb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b4d68),
	.w1(32'hbb490db9),
	.w2(32'h3b0c6eae),
	.w3(32'h3bedeb4a),
	.w4(32'hbb1e891a),
	.w5(32'hba9683bb),
	.w6(32'h3bdf5fbd),
	.w7(32'h3b8567fa),
	.w8(32'h3b80f3f9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0df60),
	.w1(32'hbb460ac2),
	.w2(32'hbb873264),
	.w3(32'h3aab5589),
	.w4(32'hbb842383),
	.w5(32'hbbad39bc),
	.w6(32'hb8ea3262),
	.w7(32'hbbe3f141),
	.w8(32'hbc0e4460),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663990),
	.w1(32'h3b0b09c9),
	.w2(32'h3b07421e),
	.w3(32'h39a80079),
	.w4(32'hb8161a34),
	.w5(32'hba18c549),
	.w6(32'hba7ebabe),
	.w7(32'hb942d8bd),
	.w8(32'hb9c80a90),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca1c78),
	.w1(32'hba139421),
	.w2(32'h3b70fb81),
	.w3(32'hb83af447),
	.w4(32'hbad2d6ba),
	.w5(32'h3a45fab2),
	.w6(32'hba9bb3ce),
	.w7(32'hbb074454),
	.w8(32'hba86da6c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc196d),
	.w1(32'hba0ed584),
	.w2(32'hb7c407d9),
	.w3(32'h3a5facfa),
	.w4(32'hba52a4ef),
	.w5(32'hb9ac903d),
	.w6(32'h3a0fbdde),
	.w7(32'hb9701312),
	.w8(32'hba19730c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8441cf),
	.w1(32'h39f42525),
	.w2(32'h3b33ae35),
	.w3(32'h3c0b6004),
	.w4(32'h3b0e307c),
	.w5(32'h3ad630dc),
	.w6(32'h3bf70a80),
	.w7(32'h3bcb4e4d),
	.w8(32'h39f48735),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a373301),
	.w1(32'hbabb5df9),
	.w2(32'h3a78c619),
	.w3(32'hba5c6339),
	.w4(32'hbafbf77c),
	.w5(32'h39840836),
	.w6(32'hbaff25b8),
	.w7(32'hbb2522a1),
	.w8(32'hb932beb7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3508313d),
	.w1(32'hb9ed707b),
	.w2(32'hb972d900),
	.w3(32'hb8a38e3d),
	.w4(32'hb9b89329),
	.w5(32'hb97d03fe),
	.w6(32'hb98dbd18),
	.w7(32'hba04b2bd),
	.w8(32'hb9d1d883),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e5dce),
	.w1(32'h3a681cc5),
	.w2(32'h3a7a0e9f),
	.w3(32'h38456deb),
	.w4(32'h39df3bab),
	.w5(32'h39dfba8c),
	.w6(32'h39851298),
	.w7(32'h3a242470),
	.w8(32'h3a4b2bcd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c4c0),
	.w1(32'h3b1b640c),
	.w2(32'h3b758edd),
	.w3(32'hbab38c4b),
	.w4(32'hba9197c3),
	.w5(32'h3a87e7a5),
	.w6(32'hbad6f503),
	.w7(32'hba2700a8),
	.w8(32'h3a978a5b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd1b2),
	.w1(32'h3a8dfa18),
	.w2(32'h3a8ce2d9),
	.w3(32'h38ed06ef),
	.w4(32'hb8f17944),
	.w5(32'hb9fd8283),
	.w6(32'hba8220df),
	.w7(32'hb9559593),
	.w8(32'hba56a9dd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacfc75),
	.w1(32'h39925f2b),
	.w2(32'hbacfa1e1),
	.w3(32'hb98ed275),
	.w4(32'hba311987),
	.w5(32'hbb1ddbf8),
	.w6(32'hbb1db3df),
	.w7(32'hbb1d37f5),
	.w8(32'hbb757209),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa489ee),
	.w1(32'h3a1bf8ca),
	.w2(32'h3a0cb1c4),
	.w3(32'h3839e0b2),
	.w4(32'hb9962ceb),
	.w5(32'hba35d7d8),
	.w6(32'hb98479e5),
	.w7(32'hb9b674d3),
	.w8(32'hba61c2a4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98444f0),
	.w1(32'hba8d5b40),
	.w2(32'h3a9bf4ef),
	.w3(32'h399df3c9),
	.w4(32'hbb04a16d),
	.w5(32'hba2089fb),
	.w6(32'h3b6a63e5),
	.w7(32'h3ac69267),
	.w8(32'h3b01963e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcfe15),
	.w1(32'h3b7cb7dd),
	.w2(32'h3b9b5a9e),
	.w3(32'h3ad0929d),
	.w4(32'h3b3e8943),
	.w5(32'h3b7255f3),
	.w6(32'hb992fed9),
	.w7(32'h3ace9060),
	.w8(32'h3b43e73f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbbf3f),
	.w1(32'h3a8849f3),
	.w2(32'h3a4e8942),
	.w3(32'hba1490fd),
	.w4(32'hba00c464),
	.w5(32'hb93bf16b),
	.w6(32'hba2612e4),
	.w7(32'hba0f96d8),
	.w8(32'hb9c86535),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916cdee),
	.w1(32'h370816c5),
	.w2(32'hb94fdd40),
	.w3(32'hb8795317),
	.w4(32'h3889d302),
	.w5(32'hb7ae4b5b),
	.w6(32'hb8eb929f),
	.w7(32'h393181ac),
	.w8(32'h377bf53c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c921fd),
	.w1(32'h3a6d9473),
	.w2(32'h3aaca6be),
	.w3(32'h39ea43a8),
	.w4(32'h3a7d2b95),
	.w5(32'h39acc384),
	.w6(32'h39499bfa),
	.w7(32'h3a7a5b51),
	.w8(32'h39913d88),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b2e30),
	.w1(32'h3a2b2758),
	.w2(32'h3a1273a2),
	.w3(32'hb95999be),
	.w4(32'h395c396a),
	.w5(32'h3932e5e9),
	.w6(32'h36f8c1aa),
	.w7(32'h39816561),
	.w8(32'hb65574b8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ccdc3),
	.w1(32'hb94793c7),
	.w2(32'hb9bbe8e1),
	.w3(32'h38d60747),
	.w4(32'hb905de36),
	.w5(32'h393b3f8c),
	.w6(32'hb99c5ab6),
	.w7(32'hb90e867a),
	.w8(32'h39ccf1b8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6da32),
	.w1(32'h3a9c3871),
	.w2(32'h3a9897ac),
	.w3(32'hb81c8d8e),
	.w4(32'hba20bda8),
	.w5(32'hba7d9a7a),
	.w6(32'hba49f45e),
	.w7(32'hb9e5f608),
	.w8(32'hb95c44e9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce8f37),
	.w1(32'hb993909b),
	.w2(32'hb9adfef6),
	.w3(32'h391043c2),
	.w4(32'hb960b0ce),
	.w5(32'hb97a6910),
	.w6(32'h3994c89c),
	.w7(32'hb8e9795a),
	.w8(32'hb8c623c2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8743e),
	.w1(32'hba57de0e),
	.w2(32'h3a19ccdf),
	.w3(32'hba40a97f),
	.w4(32'hba8c0651),
	.w5(32'hb72cfd60),
	.w6(32'hb9817e64),
	.w7(32'hb9c62888),
	.w8(32'h394ee7b7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a814002),
	.w1(32'h3ac27424),
	.w2(32'hb98fbc4a),
	.w3(32'hb99513a3),
	.w4(32'h3acccd12),
	.w5(32'hbac991d8),
	.w6(32'hba8c06af),
	.w7(32'h39b5a92e),
	.w8(32'hbb09efc6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d9cab),
	.w1(32'hba0649a1),
	.w2(32'hb84215d3),
	.w3(32'h392d328e),
	.w4(32'hb8974193),
	.w5(32'hba14ae60),
	.w6(32'h3a0f6052),
	.w7(32'h36dab122),
	.w8(32'hb9e4d2ff),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9750165),
	.w1(32'h3920b813),
	.w2(32'h39f246ab),
	.w3(32'hb703eb70),
	.w4(32'hb92005ba),
	.w5(32'h3923ed02),
	.w6(32'h394a48de),
	.w7(32'h38bec636),
	.w8(32'h39a26b6c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2fb5e),
	.w1(32'h39046840),
	.w2(32'hb90a5a01),
	.w3(32'h382e5ede),
	.w4(32'hb914e77c),
	.w5(32'h39dd92dd),
	.w6(32'h39027d3b),
	.w7(32'h38f5c1de),
	.w8(32'h398f7f6c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963aabc),
	.w1(32'hb987ea38),
	.w2(32'hb8291496),
	.w3(32'h3864b471),
	.w4(32'h394abbe4),
	.w5(32'h3a1019a8),
	.w6(32'hb7a63aa4),
	.w7(32'h3907f2e7),
	.w8(32'h3a2600e9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae87383),
	.w1(32'h38afb73d),
	.w2(32'h3b95dcaf),
	.w3(32'hbb114096),
	.w4(32'hba67be08),
	.w5(32'h3b2d1618),
	.w6(32'h3afe5c6a),
	.w7(32'h3ab420d1),
	.w8(32'h3b5ed8fa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70e5d9),
	.w1(32'h3afdc0df),
	.w2(32'h3b62d904),
	.w3(32'hbb2aa8b7),
	.w4(32'hba15c0e1),
	.w5(32'h3b1cb190),
	.w6(32'hbacec0bc),
	.w7(32'hba1aa9d1),
	.w8(32'h3b1b3d56),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd671e),
	.w1(32'hb9a9212b),
	.w2(32'h3888cb2d),
	.w3(32'hb9ec510d),
	.w4(32'hb9b8eeb2),
	.w5(32'hb9b94589),
	.w6(32'hba41d53e),
	.w7(32'hb9c0c0fc),
	.w8(32'hba1c5f09),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a398a3),
	.w1(32'h3a643074),
	.w2(32'h3b09e2f2),
	.w3(32'h39926baf),
	.w4(32'h398f8fd7),
	.w5(32'h3ae47d8a),
	.w6(32'h3a10d006),
	.w7(32'h3a95b324),
	.w8(32'h3ac79a92),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d13a6c),
	.w1(32'h398f5d7c),
	.w2(32'hb9aadf85),
	.w3(32'h395d6af3),
	.w4(32'hb9e0d44e),
	.w5(32'hba865adb),
	.w6(32'hba1a7c45),
	.w7(32'hb9a5b167),
	.w8(32'hba3d581d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c45111),
	.w1(32'h3ab4cc7c),
	.w2(32'h3b0a9acc),
	.w3(32'hb8882f89),
	.w4(32'h39265db8),
	.w5(32'h3aa62624),
	.w6(32'h39aa8b5f),
	.w7(32'h3a8b45b0),
	.w8(32'h3abb08a9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2a209),
	.w1(32'h3ae5b337),
	.w2(32'h3ab7169c),
	.w3(32'h392e1084),
	.w4(32'h3abee0a8),
	.w5(32'h3ab99cfd),
	.w6(32'hb9eb4b74),
	.w7(32'h39c12343),
	.w8(32'h3a09f344),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b9a57),
	.w1(32'h3a9b2352),
	.w2(32'h3b6d22e8),
	.w3(32'hbad696b3),
	.w4(32'hbaae0701),
	.w5(32'h3afa286b),
	.w6(32'hbabba709),
	.w7(32'hbaf798f0),
	.w8(32'h3ade497d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a251d92),
	.w1(32'h3a072d21),
	.w2(32'h39518ee6),
	.w3(32'hb8772f0a),
	.w4(32'hb7393a31),
	.w5(32'hba29345e),
	.w6(32'hba114f22),
	.w7(32'hba978593),
	.w8(32'hbabe0c04),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a681f00),
	.w1(32'h3a013feb),
	.w2(32'h3afe14fa),
	.w3(32'hb81f427c),
	.w4(32'hba5eae75),
	.w5(32'h393e6061),
	.w6(32'hba777c6c),
	.w7(32'hba3322db),
	.w8(32'h384a1de1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9993c5),
	.w1(32'h3a4959c9),
	.w2(32'h3b031424),
	.w3(32'hbaf42989),
	.w4(32'hbad84208),
	.w5(32'h39aa1da8),
	.w6(32'hbacfb91b),
	.w7(32'hbaa44f6c),
	.w8(32'hb9bb4f27),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa57cef),
	.w1(32'hb8bdd111),
	.w2(32'h393eb156),
	.w3(32'h392a78be),
	.w4(32'hba0b46c3),
	.w5(32'hbaa49674),
	.w6(32'h39ef377d),
	.w7(32'h3a007825),
	.w8(32'hba411777),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83d124c),
	.w1(32'h3aa1bc71),
	.w2(32'h3b4db3d7),
	.w3(32'hba6d5523),
	.w4(32'hb90f7e7d),
	.w5(32'h3afc5462),
	.w6(32'hbaf8466d),
	.w7(32'hbaaf695c),
	.w8(32'h3a8019b1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39968255),
	.w1(32'h3999145d),
	.w2(32'h39b588ea),
	.w3(32'hb94379bd),
	.w4(32'hb91f97eb),
	.w5(32'hb96dc12f),
	.w6(32'hb9521b4b),
	.w7(32'hb8c248b3),
	.w8(32'hb937a00a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e668),
	.w1(32'h39d20f29),
	.w2(32'hbaf7a57b),
	.w3(32'hbaa5f1c7),
	.w4(32'hba3c0c4a),
	.w5(32'hbb7422ad),
	.w6(32'hbaed5009),
	.w7(32'hbb0499c8),
	.w8(32'hbbb712e9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11005a),
	.w1(32'hb9ac6f7b),
	.w2(32'h39e633ba),
	.w3(32'hba4b9b13),
	.w4(32'hba4bcda5),
	.w5(32'hba9af571),
	.w6(32'h38a4f0e9),
	.w7(32'hb9b9cb3c),
	.w8(32'hba60a225),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39888ec4),
	.w1(32'hb9a4d737),
	.w2(32'h3884de74),
	.w3(32'h399b2da9),
	.w4(32'hb9a72835),
	.w5(32'h3a0bb457),
	.w6(32'h39052467),
	.w7(32'hb88c07a9),
	.w8(32'h3978a548),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9054c58),
	.w1(32'h39a2c67d),
	.w2(32'h3903223d),
	.w3(32'h3932b3a9),
	.w4(32'h38adc3e7),
	.w5(32'h38d18b26),
	.w6(32'h38b304e9),
	.w7(32'hb9558c08),
	.w8(32'hb98d0e8a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e452d),
	.w1(32'hb95105dc),
	.w2(32'hb9bf4d92),
	.w3(32'h39849605),
	.w4(32'hb7084c25),
	.w5(32'h39936dc4),
	.w6(32'hb9674ea0),
	.w7(32'hb9234d0f),
	.w8(32'hba0f03ea),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c6b1e),
	.w1(32'hb891c453),
	.w2(32'hb94e1099),
	.w3(32'hb9c99069),
	.w4(32'hba904aca),
	.w5(32'hbb1eabba),
	.w6(32'hba7c1ad4),
	.w7(32'hbab3666b),
	.w8(32'hbb517a16),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0fdb9),
	.w1(32'h3b08fbf4),
	.w2(32'h3b176aff),
	.w3(32'hb9c5dcc6),
	.w4(32'hba258230),
	.w5(32'h3a08a97f),
	.w6(32'hb99ac0d7),
	.w7(32'hb96a3e5f),
	.w8(32'h3a836ca3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38435517),
	.w1(32'hb98e0c46),
	.w2(32'hb9c06329),
	.w3(32'hb84c6e16),
	.w4(32'h395f65e0),
	.w5(32'hb9bcdcf4),
	.w6(32'hb97ca9ce),
	.w7(32'hb91de029),
	.w8(32'hb98ca016),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be190),
	.w1(32'h3b3fb40d),
	.w2(32'h3b9cafea),
	.w3(32'hba6bd4ed),
	.w4(32'h396ae58c),
	.w5(32'h3b3f70e2),
	.w6(32'hba9ee25a),
	.w7(32'hba66773c),
	.w8(32'h3af1e417),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b048b91),
	.w1(32'h3aef38b1),
	.w2(32'h3ac0f75a),
	.w3(32'h3a10aaa1),
	.w4(32'hb945d6cb),
	.w5(32'h398c4e7c),
	.w6(32'h37cf0c46),
	.w7(32'h38d0a08a),
	.w8(32'h395be87f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3690fd),
	.w1(32'h38e4a519),
	.w2(32'h3b3c3e1a),
	.w3(32'hbac7026c),
	.w4(32'hba7fc63b),
	.w5(32'h3ab28223),
	.w6(32'hba893a46),
	.w7(32'hba4f16e0),
	.w8(32'h3aa15437),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ca802),
	.w1(32'h3ae8d108),
	.w2(32'hba455dfe),
	.w3(32'h39d6f62f),
	.w4(32'hb910371b),
	.w5(32'hbac0fb7c),
	.w6(32'hba9891c6),
	.w7(32'hba9f083b),
	.w8(32'hbb25db6b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a036801),
	.w1(32'h3a8d3150),
	.w2(32'h3aef0745),
	.w3(32'h3a220c8b),
	.w4(32'h3a8fb028),
	.w5(32'h3a7524e8),
	.w6(32'h39b00184),
	.w7(32'h3a4e71fa),
	.w8(32'h3a458bc6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39698215),
	.w1(32'hb9ceece5),
	.w2(32'hb8af7bde),
	.w3(32'h39f6ae33),
	.w4(32'h38c813f2),
	.w5(32'h38e401ce),
	.w6(32'h3a096f43),
	.w7(32'hb90aa280),
	.w8(32'h39bd3a3a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac06d50),
	.w1(32'h3a2ceece),
	.w2(32'hb9a78966),
	.w3(32'h39a3f489),
	.w4(32'hba170008),
	.w5(32'hbad60090),
	.w6(32'h3867fbfc),
	.w7(32'hba04d6a0),
	.w8(32'hbaac69e5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21649b),
	.w1(32'hb9bcef1d),
	.w2(32'hba40f42e),
	.w3(32'hba6c55b7),
	.w4(32'hba00a455),
	.w5(32'hba99c76c),
	.w6(32'hba6e52e4),
	.w7(32'hbad02c57),
	.w8(32'hbb496b59),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a330afc),
	.w1(32'hb9c8f80b),
	.w2(32'hbab4213e),
	.w3(32'h3a27d1e5),
	.w4(32'hb9bdfe8c),
	.w5(32'hbada6969),
	.w6(32'h39db95c6),
	.w7(32'hba17c1f4),
	.w8(32'hbac8111d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f4cfb),
	.w1(32'h39cfff78),
	.w2(32'h3a3ef5e6),
	.w3(32'hba38fae0),
	.w4(32'h38a4effe),
	.w5(32'h3a2ee393),
	.w6(32'hba3c6126),
	.w7(32'hb9df0308),
	.w8(32'hb8bb3f9d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39659b5c),
	.w1(32'h3912720f),
	.w2(32'h39a49e86),
	.w3(32'hb902b9c6),
	.w4(32'h3929213b),
	.w5(32'hb94fade4),
	.w6(32'hb9e63224),
	.w7(32'h39615bf1),
	.w8(32'hb78bdde5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e0a0a7),
	.w1(32'h3aa0a805),
	.w2(32'h3b5809e8),
	.w3(32'hba903137),
	.w4(32'hba65b838),
	.w5(32'h3a7ad319),
	.w6(32'hba282366),
	.w7(32'hb8f9dacb),
	.w8(32'h3a599bc2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958abb2),
	.w1(32'hba1e29b3),
	.w2(32'h39b78524),
	.w3(32'hba4da64e),
	.w4(32'hba05deba),
	.w5(32'hb94e5224),
	.w6(32'hba311e99),
	.w7(32'hba811507),
	.w8(32'hba8a6664),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57b4f9),
	.w1(32'h3a65ee78),
	.w2(32'h3a8e747d),
	.w3(32'hba4880e8),
	.w4(32'h39694270),
	.w5(32'h39667ec2),
	.w6(32'hb925d16f),
	.w7(32'h39d0173b),
	.w8(32'h3a765ae5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e2cf9),
	.w1(32'hb9b5afb7),
	.w2(32'hb9fd510e),
	.w3(32'h3aa5110b),
	.w4(32'hb8b90b4c),
	.w5(32'hb97d7d60),
	.w6(32'h3a014d75),
	.w7(32'h35661156),
	.w8(32'hb98a0981),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378883cd),
	.w1(32'h3a44ef9a),
	.w2(32'h3aa88e05),
	.w3(32'hb8cef98c),
	.w4(32'h3a112b52),
	.w5(32'h39e3488b),
	.w6(32'h3a593b53),
	.w7(32'h3ac3cf8d),
	.w8(32'h3a2b620c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9441caf),
	.w1(32'h3855e9bb),
	.w2(32'h376bfeec),
	.w3(32'h382d5454),
	.w4(32'h3819b53b),
	.w5(32'hb9cf97d9),
	.w6(32'hb8314e68),
	.w7(32'hb8e95f63),
	.w8(32'hb9e64037),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ef126),
	.w1(32'h38281963),
	.w2(32'h39556146),
	.w3(32'hb780b037),
	.w4(32'h3880298e),
	.w5(32'hba273686),
	.w6(32'hb7ba4509),
	.w7(32'h387c9279),
	.w8(32'hb9417e2b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9fc32),
	.w1(32'h3994db67),
	.w2(32'h38efc620),
	.w3(32'hba3c1787),
	.w4(32'hb9f8a27e),
	.w5(32'hba605a18),
	.w6(32'hba928c39),
	.w7(32'hba9497a5),
	.w8(32'hba93888e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02a68d),
	.w1(32'hb74e5c53),
	.w2(32'h3b432f93),
	.w3(32'hbac66077),
	.w4(32'hbb7174ba),
	.w5(32'hba4c974c),
	.w6(32'hb9cf184c),
	.w7(32'hba92bf70),
	.w8(32'h3a2cd569),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e1e70),
	.w1(32'hba07f727),
	.w2(32'hb96f97d7),
	.w3(32'h3a2da9e5),
	.w4(32'h39076a4b),
	.w5(32'hba0d4459),
	.w6(32'h3a279fab),
	.w7(32'hb936a5f9),
	.w8(32'h37d48daf),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab109a1),
	.w1(32'h3a8ff1b6),
	.w2(32'h3999512c),
	.w3(32'hba04aef9),
	.w4(32'hba2c0ce0),
	.w5(32'hb99c8bbf),
	.w6(32'hbaf30e10),
	.w7(32'hbab9e3b3),
	.w8(32'hba6faeaa),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaea092),
	.w1(32'h38d37af6),
	.w2(32'h3878fe26),
	.w3(32'hba0437dd),
	.w4(32'h380fc733),
	.w5(32'hb7e9cc3c),
	.w6(32'hba937f49),
	.w7(32'hba379e37),
	.w8(32'hb9901193),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb11cb),
	.w1(32'h3ab14837),
	.w2(32'h3b2a2cd5),
	.w3(32'h3914e7c4),
	.w4(32'hba52c00f),
	.w5(32'h3a838236),
	.w6(32'hb9318576),
	.w7(32'hba95b300),
	.w8(32'h3b0303a6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ec6bb),
	.w1(32'h3a9c0746),
	.w2(32'h3b1d13be),
	.w3(32'hba14e000),
	.w4(32'hb8da85fc),
	.w5(32'h3afc8bcd),
	.w6(32'hba70dcbd),
	.w7(32'hb9c43d7e),
	.w8(32'h3a08c516),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900d163),
	.w1(32'h3afaf199),
	.w2(32'h3b3e0e23),
	.w3(32'hba9cd721),
	.w4(32'hba1b3dd2),
	.w5(32'h3aefcfe9),
	.w6(32'hba1c7104),
	.w7(32'hba441e0b),
	.w8(32'h3ad22247),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e82982),
	.w1(32'hb9e74dab),
	.w2(32'hb9872779),
	.w3(32'h393bd023),
	.w4(32'hb9d5a200),
	.w5(32'hb9ea2dff),
	.w6(32'hb968dd9e),
	.w7(32'hb9d48189),
	.w8(32'hba06da1b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce1724),
	.w1(32'h3a7ef874),
	.w2(32'h3aed65f9),
	.w3(32'hb9efaa4f),
	.w4(32'h3a02c089),
	.w5(32'h3a8bbc04),
	.w6(32'hba7b4b03),
	.w7(32'hb99ea511),
	.w8(32'h394e0d94),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b95f43),
	.w1(32'hb9ab550a),
	.w2(32'hba0bd86a),
	.w3(32'h37d8192a),
	.w4(32'h39cc5c7e),
	.w5(32'hb97568fc),
	.w6(32'h39d20977),
	.w7(32'h3966a46c),
	.w8(32'h38b8e6ab),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2ba10),
	.w1(32'h3980972c),
	.w2(32'hb9465740),
	.w3(32'h3874a217),
	.w4(32'h37f1a7ce),
	.w5(32'h39dd31c7),
	.w6(32'h39b91c93),
	.w7(32'h38b492f6),
	.w8(32'h39465aeb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb840574a),
	.w1(32'h391da09b),
	.w2(32'h3a555326),
	.w3(32'h39715fed),
	.w4(32'hb9845472),
	.w5(32'h39bd6650),
	.w6(32'h39b5f048),
	.w7(32'h379c80c8),
	.w8(32'h39d71e75),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4957d),
	.w1(32'h3b1bd879),
	.w2(32'h3b39f22d),
	.w3(32'h39faee21),
	.w4(32'h3acfe278),
	.w5(32'h3b06be99),
	.w6(32'h39b07234),
	.w7(32'h3a5948ec),
	.w8(32'h3adcdc59),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a9b1e),
	.w1(32'h3913fde3),
	.w2(32'h3984e23f),
	.w3(32'h38bbde93),
	.w4(32'h39203d18),
	.w5(32'h3804ff1a),
	.w6(32'hb886b05a),
	.w7(32'hb95cca0c),
	.w8(32'hb8f0df25),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38bc3d),
	.w1(32'hb60e839f),
	.w2(32'hb9a5e6dd),
	.w3(32'h39a30160),
	.w4(32'h3983cab7),
	.w5(32'hb621ce38),
	.w6(32'h39ebc0c0),
	.w7(32'h399676a4),
	.w8(32'h38ee2bff),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8736d2a),
	.w1(32'h3a118a83),
	.w2(32'hb9303782),
	.w3(32'h398be686),
	.w4(32'h39bcb431),
	.w5(32'hba82539b),
	.w6(32'h3864fb97),
	.w7(32'h3a519dc8),
	.w8(32'hb9ceab0a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6596),
	.w1(32'h3af15780),
	.w2(32'h3b264c17),
	.w3(32'hb8b74af3),
	.w4(32'h3a5cb977),
	.w5(32'h3b180d3a),
	.w6(32'hb9c267a2),
	.w7(32'h3a4f7c4e),
	.w8(32'h3af3ea31),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b40d3),
	.w1(32'hba8db325),
	.w2(32'h3aa1e1af),
	.w3(32'h3b965bac),
	.w4(32'hba235052),
	.w5(32'h39411340),
	.w6(32'h3b55cdc4),
	.w7(32'h3a82d2f0),
	.w8(32'hb944e953),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38722630),
	.w1(32'h39dbea5e),
	.w2(32'hb91865f2),
	.w3(32'h38ea7da1),
	.w4(32'h39314f42),
	.w5(32'h390c302d),
	.w6(32'h3959361b),
	.w7(32'hb69d314d),
	.w8(32'h36d78288),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b368933),
	.w1(32'h3b887401),
	.w2(32'h3bb9df17),
	.w3(32'hb9e69607),
	.w4(32'h3a9a42cc),
	.w5(32'h3b7007d7),
	.w6(32'h39cdac7d),
	.w7(32'h3b0f8111),
	.w8(32'h3bcaca12),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d23306),
	.w1(32'h3aa12658),
	.w2(32'h3a1c828a),
	.w3(32'h3a002abf),
	.w4(32'hb8d57d20),
	.w5(32'hb9c5725a),
	.w6(32'hbb38d1e8),
	.w7(32'hbba1d9fc),
	.w8(32'hbb9041a2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f1261),
	.w1(32'hb9b1df63),
	.w2(32'h3a98f7e4),
	.w3(32'hb930af46),
	.w4(32'hba55a320),
	.w5(32'h378a946e),
	.w6(32'h381b4c2a),
	.w7(32'hba405c53),
	.w8(32'hb9c25155),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980b162),
	.w1(32'h385c7efb),
	.w2(32'hb9a3a9eb),
	.w3(32'h39b30440),
	.w4(32'hb963905f),
	.w5(32'h342c53bc),
	.w6(32'h3887f368),
	.w7(32'h38d4c55e),
	.w8(32'h398653cf),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949b60b),
	.w1(32'h39085d4d),
	.w2(32'hb78dcc41),
	.w3(32'h3967a087),
	.w4(32'h38c3618f),
	.w5(32'h3a000b1d),
	.w6(32'h38b0b979),
	.w7(32'h391aaa5a),
	.w8(32'h397f8807),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ff197),
	.w1(32'hb887b84e),
	.w2(32'h3816f919),
	.w3(32'hb89ad560),
	.w4(32'hb8b82065),
	.w5(32'hb93ab783),
	.w6(32'hb98cac24),
	.w7(32'hb8f37de0),
	.w8(32'hb9023fc2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9981ab4),
	.w1(32'hbaa439d6),
	.w2(32'h3aa29aaf),
	.w3(32'hb953a408),
	.w4(32'hba8d3bfc),
	.w5(32'h39bc5232),
	.w6(32'h39666693),
	.w7(32'hba621159),
	.w8(32'h39ac0b00),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00b187),
	.w1(32'hba1b5533),
	.w2(32'hb93320bf),
	.w3(32'hba919e84),
	.w4(32'hbad7fc01),
	.w5(32'hbad22137),
	.w6(32'h36bf381a),
	.w7(32'hba82ed6a),
	.w8(32'hba8bd511),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b066ef9),
	.w1(32'h3b08ffb4),
	.w2(32'h3a98896b),
	.w3(32'h3a974914),
	.w4(32'h3a98e67d),
	.w5(32'hb9f55608),
	.w6(32'hb90ac925),
	.w7(32'h3a3019c4),
	.w8(32'hba694eea),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09ed3c),
	.w1(32'h3a3d7154),
	.w2(32'h3992017c),
	.w3(32'h39d267a7),
	.w4(32'h398816bf),
	.w5(32'hb916661c),
	.w6(32'hb9457fae),
	.w7(32'h39cff9ec),
	.w8(32'hb8979b29),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8faa5),
	.w1(32'hbb73ecd0),
	.w2(32'hbb928f47),
	.w3(32'hb96ba777),
	.w4(32'hbaabccb6),
	.w5(32'h3b06bc42),
	.w6(32'hba363037),
	.w7(32'h3a5bd4f5),
	.w8(32'h3c0a4ddd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5cfd4),
	.w1(32'h3bd0fb3f),
	.w2(32'h3b7a5fff),
	.w3(32'h3b1954de),
	.w4(32'hba6cef4c),
	.w5(32'hbbf89d64),
	.w6(32'h3bac02e5),
	.w7(32'h3abcf2cf),
	.w8(32'h3aa2576a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad81fa),
	.w1(32'h3bf9708c),
	.w2(32'h3c2aef83),
	.w3(32'hbb590be1),
	.w4(32'h3b490ed7),
	.w5(32'hbbb863f5),
	.w6(32'hbb86758f),
	.w7(32'hbaba2392),
	.w8(32'hba8e4fff),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd87c6d),
	.w1(32'h3bdc6c71),
	.w2(32'h3baaa3c6),
	.w3(32'h3bd71391),
	.w4(32'h3c1e6aca),
	.w5(32'h3b5563c7),
	.w6(32'h3b294552),
	.w7(32'h3bd49e53),
	.w8(32'h3c01b424),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba15156),
	.w1(32'hbbe55eb2),
	.w2(32'h3b0e218d),
	.w3(32'hb9abd762),
	.w4(32'hbae55d80),
	.w5(32'hb971ce91),
	.w6(32'h3af34fc8),
	.w7(32'hbabd6211),
	.w8(32'hba8e3fa3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39909c70),
	.w1(32'h3a5f54ff),
	.w2(32'h3b91b2e3),
	.w3(32'hbaf0d5d1),
	.w4(32'hbbb53eb9),
	.w5(32'h3933afbb),
	.w6(32'h398b532e),
	.w7(32'hbb453562),
	.w8(32'hbb209442),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d5240),
	.w1(32'hbb03bbcd),
	.w2(32'h3c0289e3),
	.w3(32'hbba6b5b5),
	.w4(32'h3b0d5e13),
	.w5(32'h3aaad814),
	.w6(32'hbb23af32),
	.w7(32'hbb0ea0d5),
	.w8(32'hbb9858cb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89feaf),
	.w1(32'hbb71e751),
	.w2(32'hbbc363ac),
	.w3(32'h3bc63596),
	.w4(32'hbb12fa96),
	.w5(32'hb82a2d36),
	.w6(32'h3ac62d33),
	.w7(32'hbb953d0f),
	.w8(32'hb9b07100),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe204a9),
	.w1(32'h3b00f25f),
	.w2(32'h3a0a0d09),
	.w3(32'h3979bcb1),
	.w4(32'hba63d7c3),
	.w5(32'hbba949d6),
	.w6(32'h3b616cd4),
	.w7(32'h3a82447a),
	.w8(32'h37f24c15),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beabd2b),
	.w1(32'h3b0f79fa),
	.w2(32'h3b6aee18),
	.w3(32'hb9e36d30),
	.w4(32'h3b1d1735),
	.w5(32'h3a1a4f5d),
	.w6(32'hbbcb8817),
	.w7(32'h3b2f51d6),
	.w8(32'hba8823c6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be58057),
	.w1(32'h39f31e45),
	.w2(32'h3bed8474),
	.w3(32'h3b6de316),
	.w4(32'hbb25b716),
	.w5(32'h3a0f62ff),
	.w6(32'hbb01cc09),
	.w7(32'h38836858),
	.w8(32'h3b061183),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc8237),
	.w1(32'hbc0ff29e),
	.w2(32'hbbc3c431),
	.w3(32'h3afbb268),
	.w4(32'hbb594683),
	.w5(32'h3b755346),
	.w6(32'h3bed5f79),
	.w7(32'hbb2dff07),
	.w8(32'h3bd70bad),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf39bd3),
	.w1(32'h3a076bb4),
	.w2(32'hba5c14b7),
	.w3(32'h3adf8630),
	.w4(32'hbae87547),
	.w5(32'hbaefd4f6),
	.w6(32'h3bc4cf42),
	.w7(32'hbb1ac0ec),
	.w8(32'hbb98c1c7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f25a9),
	.w1(32'hbb72a4db),
	.w2(32'hbb2132dc),
	.w3(32'hba79d22a),
	.w4(32'h3b4cdf3e),
	.w5(32'h3b8a3707),
	.w6(32'hbb66e1d4),
	.w7(32'h3aa4fa51),
	.w8(32'h3b234f86),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabec863),
	.w1(32'hb9dc9b55),
	.w2(32'h3c02076c),
	.w3(32'h3a7e34c9),
	.w4(32'h3ba0e9aa),
	.w5(32'hbb64debd),
	.w6(32'h3ae4a048),
	.w7(32'h3b2fc85b),
	.w8(32'h3bb69bbc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7c7f0),
	.w1(32'h3bc8ea82),
	.w2(32'h3c511887),
	.w3(32'h3aff364a),
	.w4(32'hba9e700d),
	.w5(32'hbb8e8c04),
	.w6(32'hbba87b5f),
	.w7(32'hba06a44b),
	.w8(32'h3a00cd3a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf94d06),
	.w1(32'h3bbdc9ce),
	.w2(32'hbac95f76),
	.w3(32'h3a7f3e62),
	.w4(32'h3be5a890),
	.w5(32'h3c088d65),
	.w6(32'hbac7fde9),
	.w7(32'hba55e796),
	.w8(32'hbb6ec90b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7c436),
	.w1(32'hbae41a64),
	.w2(32'hbb068362),
	.w3(32'hbb92c238),
	.w4(32'hba9ac05f),
	.w5(32'hbb3e56d9),
	.w6(32'hbbb71fa4),
	.w7(32'hbaffcb2e),
	.w8(32'h3a4b037c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78806),
	.w1(32'hbb1d5667),
	.w2(32'hbb639873),
	.w3(32'hbb9f5a8a),
	.w4(32'hbbdb884c),
	.w5(32'hbc0051e1),
	.w6(32'hbbe2b866),
	.w7(32'hbb6d36fe),
	.w8(32'hbb954a37),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa72215),
	.w1(32'hbaa6057a),
	.w2(32'h3a6abe2c),
	.w3(32'hbbd3cb2e),
	.w4(32'h39d979ae),
	.w5(32'h3aa1af9b),
	.w6(32'hbaf9f66e),
	.w7(32'hbb5b79d8),
	.w8(32'h3a7d914b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaded88e),
	.w1(32'hbb5ab91e),
	.w2(32'h3a040a14),
	.w3(32'h3bafeead),
	.w4(32'hbbb41950),
	.w5(32'hbb8f8ad1),
	.w6(32'hba22f6e4),
	.w7(32'h3abcf677),
	.w8(32'hbad6e819),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6ff5f),
	.w1(32'hba3ff1e0),
	.w2(32'hba33b3c6),
	.w3(32'hbbbf0720),
	.w4(32'hbb90f1b8),
	.w5(32'hbb8ab60e),
	.w6(32'hbb627add),
	.w7(32'hbad75150),
	.w8(32'h3ac36764),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717ae1),
	.w1(32'hb9561ece),
	.w2(32'h3c1f6362),
	.w3(32'h39fb11ad),
	.w4(32'hbb39dfb4),
	.w5(32'h3aeecd47),
	.w6(32'hba4b5ad6),
	.w7(32'h3a47fccb),
	.w8(32'hbb02a96a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a0fcf),
	.w1(32'hbb5a02b9),
	.w2(32'hba8c4549),
	.w3(32'hbaee7071),
	.w4(32'h3ba44646),
	.w5(32'h3b01361b),
	.w6(32'h3b323f4e),
	.w7(32'h3b89d4f8),
	.w8(32'hb92f1fb3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2aa67e),
	.w1(32'hbb0ac574),
	.w2(32'hbb1d6f3b),
	.w3(32'h3b7cbf22),
	.w4(32'h3a276de1),
	.w5(32'h3b29921c),
	.w6(32'h3b6a1fb2),
	.w7(32'h3c04e7d5),
	.w8(32'h3c189d20),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98e011),
	.w1(32'h3b054532),
	.w2(32'hba2f126d),
	.w3(32'hbace53b4),
	.w4(32'h3a63769c),
	.w5(32'h37a814cd),
	.w6(32'h3badfa10),
	.w7(32'hbb99d39d),
	.w8(32'hba7ab884),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a31f),
	.w1(32'h3bba873f),
	.w2(32'hbb0ffb3b),
	.w3(32'h3a9d4ac3),
	.w4(32'h3ada3bd7),
	.w5(32'hbc110119),
	.w6(32'h3b0c2fce),
	.w7(32'hbb386812),
	.w8(32'hbb417ffb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37101f),
	.w1(32'h3b417d56),
	.w2(32'hbadd4746),
	.w3(32'hbb6334bf),
	.w4(32'hbb4afdd7),
	.w5(32'hbc044e49),
	.w6(32'h39988071),
	.w7(32'hbbc4d5d1),
	.w8(32'hbc00961e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5fd4),
	.w1(32'hbb8bf52c),
	.w2(32'hbbbc8ce6),
	.w3(32'hbba6ebaa),
	.w4(32'h3a1622f7),
	.w5(32'hbb644fff),
	.w6(32'hbb45168b),
	.w7(32'h3ad77e49),
	.w8(32'hbb02e747),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb93e8b),
	.w1(32'h3b43c9d4),
	.w2(32'h3a2a71e4),
	.w3(32'hbb7ea6a6),
	.w4(32'hbb0384d8),
	.w5(32'hbb3e6189),
	.w6(32'hbb55902b),
	.w7(32'h3a68bdba),
	.w8(32'h3af28914),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a0a91),
	.w1(32'h3ad0f1cd),
	.w2(32'h3b17ac2b),
	.w3(32'hbb0fef9a),
	.w4(32'hbbc87584),
	.w5(32'h3b986f07),
	.w6(32'hbae3eeee),
	.w7(32'hbb389835),
	.w8(32'hba3c55d3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf83573),
	.w1(32'hb96993d1),
	.w2(32'hb9a1eec7),
	.w3(32'h3bbecebc),
	.w4(32'hba70017e),
	.w5(32'hbba1f175),
	.w6(32'h3aebe0e5),
	.w7(32'hbb3afd63),
	.w8(32'hbbb0f9b5),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8effde),
	.w1(32'h3a73598d),
	.w2(32'h3b0eac9b),
	.w3(32'hbb16731d),
	.w4(32'h3a7e5bcd),
	.w5(32'hba9158aa),
	.w6(32'hbb575d62),
	.w7(32'hbbb3f6f5),
	.w8(32'hbbbd7b28),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b11d),
	.w1(32'hba2dd2a9),
	.w2(32'h3b08f6b3),
	.w3(32'h3a848ad2),
	.w4(32'hbaaf37f7),
	.w5(32'hbb1e66c0),
	.w6(32'hbafb24f6),
	.w7(32'hbaefef2c),
	.w8(32'hbbc10f9d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7f316),
	.w1(32'h3b4f90eb),
	.w2(32'hbad66e42),
	.w3(32'hbb39302c),
	.w4(32'h3b200652),
	.w5(32'hbc260a5e),
	.w6(32'hbb6614d4),
	.w7(32'h3b62c65b),
	.w8(32'hba4bffc6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecbdd6),
	.w1(32'h3b373c64),
	.w2(32'h3c04d859),
	.w3(32'hbbe6ca44),
	.w4(32'h3ac4adcb),
	.w5(32'hbc3d4d06),
	.w6(32'hbb98a897),
	.w7(32'h394e82f5),
	.w8(32'hbb83d531),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889645),
	.w1(32'hbb8adbf4),
	.w2(32'hb968d297),
	.w3(32'hbb6ede03),
	.w4(32'hbb1dca25),
	.w5(32'h3aa80b83),
	.w6(32'hbbcdbd8c),
	.w7(32'hba5b8c9d),
	.w8(32'hbb1503ae),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdcf16),
	.w1(32'h3b73051c),
	.w2(32'h3919589e),
	.w3(32'hbad76969),
	.w4(32'h39fcf2e2),
	.w5(32'h3a6ddf4a),
	.w6(32'hba8959a6),
	.w7(32'h3b58c22d),
	.w8(32'h3a6c064e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6be67),
	.w1(32'h3b3e6111),
	.w2(32'hbb4d532d),
	.w3(32'h3ae41404),
	.w4(32'h3b11216c),
	.w5(32'hba9e4cd4),
	.w6(32'hb9d9801f),
	.w7(32'hbafeb8f7),
	.w8(32'h3b4810d4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10755c),
	.w1(32'h3abe2a3a),
	.w2(32'h3b807ed8),
	.w3(32'h3b14cbc0),
	.w4(32'h3a76ce92),
	.w5(32'hbb939ce4),
	.w6(32'hb9ed94ae),
	.w7(32'hb9809273),
	.w8(32'hbb193c93),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed9414),
	.w1(32'h3b874b62),
	.w2(32'h3c4cdfed),
	.w3(32'h3b60bd33),
	.w4(32'h3b41eb8c),
	.w5(32'hbc0365b9),
	.w6(32'hbb8979e8),
	.w7(32'h38ad3948),
	.w8(32'hbb73a932),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30453a),
	.w1(32'h3b887ba5),
	.w2(32'h3ac09272),
	.w3(32'h3b9edc34),
	.w4(32'hbb1747f2),
	.w5(32'hba877c07),
	.w6(32'hbaf6ae06),
	.w7(32'h3ace99ee),
	.w8(32'hbb758a08),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bb0e9),
	.w1(32'h3c031952),
	.w2(32'h3c04509f),
	.w3(32'hbbae30d1),
	.w4(32'h3b0cf5ee),
	.w5(32'h3b8dd29b),
	.w6(32'hbc19e1fb),
	.w7(32'h3a5dc09c),
	.w8(32'h38c3735c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998c75e),
	.w1(32'h39169273),
	.w2(32'h3b854d6b),
	.w3(32'hbbdf6c67),
	.w4(32'hbb30fd17),
	.w5(32'h3a17b4a2),
	.w6(32'hbb7cc12d),
	.w7(32'hbbc0fa23),
	.w8(32'hbb5f0f1d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad33bdc),
	.w1(32'hbb863e5d),
	.w2(32'h3c1e8841),
	.w3(32'h3a81c153),
	.w4(32'h3c1e7b96),
	.w5(32'h3c6bf3eb),
	.w6(32'hbb4aab71),
	.w7(32'h3a9bbec3),
	.w8(32'h3b62fdf3),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397dd238),
	.w1(32'hbba83f34),
	.w2(32'hbb315566),
	.w3(32'h3bc00c9a),
	.w4(32'h3b8f9528),
	.w5(32'h3ba20b17),
	.w6(32'h3bb2693b),
	.w7(32'h3bb400a9),
	.w8(32'h3b830c0a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18d54a),
	.w1(32'hb9b58098),
	.w2(32'hbb43253a),
	.w3(32'h3b75cf9b),
	.w4(32'hbb636da7),
	.w5(32'hba940956),
	.w6(32'h3b8ba31c),
	.w7(32'hbb5f7dc4),
	.w8(32'h3a9c72ff),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfedc2),
	.w1(32'h3abcf831),
	.w2(32'h3b182d46),
	.w3(32'hba555ece),
	.w4(32'hbb1f846e),
	.w5(32'hbb77a5da),
	.w6(32'hbb16bf58),
	.w7(32'h3a766f4c),
	.w8(32'hbac982b6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e9f7),
	.w1(32'hbb418a62),
	.w2(32'hbab87d71),
	.w3(32'h3c1bf28e),
	.w4(32'h3b747382),
	.w5(32'h3bde9c1f),
	.w6(32'h3be1bc0f),
	.w7(32'h3bcbf717),
	.w8(32'h3c1b9b10),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b4b06),
	.w1(32'hba4a85a1),
	.w2(32'h3b263295),
	.w3(32'h3ae448f5),
	.w4(32'hbb85fabe),
	.w5(32'hbb9e74c6),
	.w6(32'h3bc49f38),
	.w7(32'hbb8fed77),
	.w8(32'hbc178d9b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5ff24),
	.w1(32'h3b7e6961),
	.w2(32'h38a616d0),
	.w3(32'hbbd58002),
	.w4(32'h3a505dbb),
	.w5(32'hbbddab8f),
	.w6(32'hbc0b1725),
	.w7(32'hbb835f0b),
	.w8(32'hbb3ebecd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6293e1),
	.w1(32'hbb6b3f25),
	.w2(32'hba71ddd1),
	.w3(32'hbb6812a7),
	.w4(32'h3aa481c6),
	.w5(32'h3ad7743a),
	.w6(32'hbb0898d2),
	.w7(32'hbb0a5da5),
	.w8(32'h3ae8b917),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba822566),
	.w1(32'h3a671efa),
	.w2(32'hbbcac88a),
	.w3(32'h3b4884b8),
	.w4(32'hbb572568),
	.w5(32'hbb421886),
	.w6(32'h3ac404c1),
	.w7(32'h388d12f0),
	.w8(32'hbb0332d7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb686fb5),
	.w1(32'h39827a0d),
	.w2(32'hbab5cf4f),
	.w3(32'hbb83b5af),
	.w4(32'hbb9ccd4d),
	.w5(32'hbbb16e2b),
	.w6(32'hbbb53000),
	.w7(32'hbac0cad0),
	.w8(32'h390d3418),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ee3be),
	.w1(32'h3a1978e0),
	.w2(32'hbae2e495),
	.w3(32'hbaf61d41),
	.w4(32'hba9e638e),
	.w5(32'h3b692882),
	.w6(32'h3b272c21),
	.w7(32'hbbbeb2d6),
	.w8(32'hbabf5948),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49dd60),
	.w1(32'h3bc6c490),
	.w2(32'h3c8e3861),
	.w3(32'h3b817869),
	.w4(32'h3a21168f),
	.w5(32'hbbb32243),
	.w6(32'h3b0e9c8f),
	.w7(32'hbab0368d),
	.w8(32'hba518eaa),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e7d74),
	.w1(32'h3c112297),
	.w2(32'h3ccb7b87),
	.w3(32'h3bffbed3),
	.w4(32'h3c05c1e5),
	.w5(32'hbb384b7a),
	.w6(32'h3a8c913b),
	.w7(32'h3ad14ab5),
	.w8(32'hbb80f81f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc12c18),
	.w1(32'hbac0b7e6),
	.w2(32'hbafaa42a),
	.w3(32'hbb66f479),
	.w4(32'hbba3357b),
	.w5(32'h3a515968),
	.w6(32'hbbe21ab7),
	.w7(32'hbb160280),
	.w8(32'h3aa41e08),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2afbcd),
	.w1(32'hbbcd38e0),
	.w2(32'h3aef517f),
	.w3(32'h3a17427b),
	.w4(32'h396e0227),
	.w5(32'hbb5f84b1),
	.w6(32'h392e62cb),
	.w7(32'h3acb2065),
	.w8(32'hba8ed328),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule