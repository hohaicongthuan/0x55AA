module layer_10_featuremap_343(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077e52),
	.w1(32'h3c59aa52),
	.w2(32'h3c3f5380),
	.w3(32'h3bdad071),
	.w4(32'h3be4ac48),
	.w5(32'h3a894a13),
	.w6(32'h3bbaf390),
	.w7(32'h3bd119f5),
	.w8(32'h3a6e17a2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67c82),
	.w1(32'h399a2950),
	.w2(32'hbaa460e4),
	.w3(32'hbbce3beb),
	.w4(32'h3b007a2b),
	.w5(32'hbbb11b18),
	.w6(32'hbb2b2565),
	.w7(32'h3b0b75a8),
	.w8(32'hbc12d3ce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1d9b),
	.w1(32'h3b9fe8ce),
	.w2(32'h3b736a39),
	.w3(32'h3b350483),
	.w4(32'hbb31d98d),
	.w5(32'hbb325545),
	.w6(32'hba4bdfee),
	.w7(32'hba85b8a5),
	.w8(32'hbb04f828),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d4cc5),
	.w1(32'hbaf60790),
	.w2(32'hba844e0a),
	.w3(32'hbac2116b),
	.w4(32'hbae15c9b),
	.w5(32'hbb872da0),
	.w6(32'hbb12faed),
	.w7(32'hbaa73435),
	.w8(32'hbc0d6cab),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec037c),
	.w1(32'hbb86bb36),
	.w2(32'h3a77415f),
	.w3(32'hbb1e8c16),
	.w4(32'h39a9b188),
	.w5(32'hba396e65),
	.w6(32'hbbb1e53e),
	.w7(32'hba78acb1),
	.w8(32'h3b8aabf7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7416f4),
	.w1(32'h3b90d17d),
	.w2(32'h3ba4d2c2),
	.w3(32'hb7d2d2d2),
	.w4(32'h3998cd18),
	.w5(32'h3ab4fb97),
	.w6(32'h3b8e62b8),
	.w7(32'h3ba41f53),
	.w8(32'h3a33e204),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae752f7),
	.w1(32'hbb46e168),
	.w2(32'hb9e59ccd),
	.w3(32'hba87f5bc),
	.w4(32'hbb5a0553),
	.w5(32'h3b59629d),
	.w6(32'h3af670c2),
	.w7(32'h38d8504f),
	.w8(32'h3b590c52),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd96ac1),
	.w1(32'hbb8b009b),
	.w2(32'h3a439feb),
	.w3(32'hbb1f8558),
	.w4(32'hbb915a88),
	.w5(32'h3b5027da),
	.w6(32'hbb90e6d4),
	.w7(32'hbb8bb18e),
	.w8(32'h3bdcb68d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24d138),
	.w1(32'h3c28442d),
	.w2(32'h3c02b249),
	.w3(32'h3ba895fd),
	.w4(32'h3bb7e05c),
	.w5(32'hbb74707a),
	.w6(32'h3baa8dcf),
	.w7(32'h3be8d4bb),
	.w8(32'h3af984d4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d09b2),
	.w1(32'h3b9a5909),
	.w2(32'hbb7c3912),
	.w3(32'hbbe4da73),
	.w4(32'h3ae88498),
	.w5(32'hbbb9ea0a),
	.w6(32'hbb36455e),
	.w7(32'h3bd2fa02),
	.w8(32'hbb89322c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bfa37),
	.w1(32'h3ae0f417),
	.w2(32'h3b0c1c2f),
	.w3(32'hba7e1b39),
	.w4(32'hbad67ded),
	.w5(32'hbb5cdd32),
	.w6(32'h3aa8be04),
	.w7(32'h3b834754),
	.w8(32'hbbd956d6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd69f02),
	.w1(32'h3a870d2d),
	.w2(32'hba537bc1),
	.w3(32'hbb52acec),
	.w4(32'hba9e25c7),
	.w5(32'hbb641f93),
	.w6(32'hbbf0de40),
	.w7(32'hbb6d3b92),
	.w8(32'h3a173792),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9a43e),
	.w1(32'hbba1c7b8),
	.w2(32'hbc331cb2),
	.w3(32'hbc363808),
	.w4(32'hbb6d6793),
	.w5(32'hbbee2972),
	.w6(32'hbc37c850),
	.w7(32'hbbb36fcd),
	.w8(32'hbc0c3603),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc06ce8),
	.w1(32'hbb89db0a),
	.w2(32'hbbfe4cf6),
	.w3(32'hbc00e399),
	.w4(32'hbb934ffb),
	.w5(32'hbbe45c61),
	.w6(32'hbbd984a9),
	.w7(32'hbbd5b26b),
	.w8(32'hbbaef4ce),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46f79),
	.w1(32'hbb65d0cb),
	.w2(32'hbc0ec093),
	.w3(32'hbaee9ec8),
	.w4(32'h3b914685),
	.w5(32'h3afb99f3),
	.w6(32'hbbe33e58),
	.w7(32'hba5b9cad),
	.w8(32'hba16c035),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b965),
	.w1(32'h3ad5e2d4),
	.w2(32'hbb5e11d3),
	.w3(32'hbb8bf8de),
	.w4(32'h3ba964b5),
	.w5(32'hbab3e6c4),
	.w6(32'hbb9e293e),
	.w7(32'h3a63b047),
	.w8(32'hbb83eaea),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93bd99),
	.w1(32'h3aeb2274),
	.w2(32'h3bb774c5),
	.w3(32'h3b09952c),
	.w4(32'h3b1d3dab),
	.w5(32'h3a62d659),
	.w6(32'h3b75ea97),
	.w7(32'h3a5e7df4),
	.w8(32'h3b230a30),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0507c2),
	.w1(32'h3a910121),
	.w2(32'hbb8cc9a0),
	.w3(32'hbb817cc1),
	.w4(32'h3a127137),
	.w5(32'hbc0a3336),
	.w6(32'hbb9e41d9),
	.w7(32'h3b39bc49),
	.w8(32'hbbd4f10b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd071cb),
	.w1(32'hbb2c5508),
	.w2(32'hbbc6b1d3),
	.w3(32'hbb6db7f0),
	.w4(32'hbaada30e),
	.w5(32'hbab468a9),
	.w6(32'hbbec94b6),
	.w7(32'hbac36e58),
	.w8(32'hbaea09c2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a989575),
	.w1(32'h3ab0f865),
	.w2(32'hba4712a3),
	.w3(32'h3b7528c1),
	.w4(32'h3bb1430f),
	.w5(32'h3b2bc76a),
	.w6(32'h3b3791c0),
	.w7(32'hba72ce4e),
	.w8(32'hba6f940e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9eafa),
	.w1(32'h3a861131),
	.w2(32'h3afae2fb),
	.w3(32'hbb61aef3),
	.w4(32'h398c0137),
	.w5(32'hb9bea1ce),
	.w6(32'hbb57ed46),
	.w7(32'hba93bfa3),
	.w8(32'hb94e23de),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd0f4),
	.w1(32'h3a14a5bc),
	.w2(32'hb9e4d15c),
	.w3(32'h3b36fd4a),
	.w4(32'h3bb5449f),
	.w5(32'hbb4e50a3),
	.w6(32'hb96e48f7),
	.w7(32'h3b0ed8fb),
	.w8(32'hbc05b7b3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1706e),
	.w1(32'hbb2bdf54),
	.w2(32'hbc62cb44),
	.w3(32'hbc66a66a),
	.w4(32'h3abfeff0),
	.w5(32'hbc00e025),
	.w6(32'hbc9dfc70),
	.w7(32'hbbf33026),
	.w8(32'hbc6c863b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39545ba8),
	.w1(32'h3bb5a703),
	.w2(32'hbc246ac2),
	.w3(32'hbbc3ac55),
	.w4(32'h3ba1d92a),
	.w5(32'hbbc4216f),
	.w6(32'hbc273adb),
	.w7(32'h3b8f27c7),
	.w8(32'hbbccf7e2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef8679),
	.w1(32'h3b972ff7),
	.w2(32'hbc003fba),
	.w3(32'hbc155e37),
	.w4(32'h3b39e028),
	.w5(32'hbb83e537),
	.w6(32'hbc229505),
	.w7(32'h3a4452ad),
	.w8(32'hbc39ae2b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe3775),
	.w1(32'hbab8d7b9),
	.w2(32'hba71a8f1),
	.w3(32'h3655f6fb),
	.w4(32'h3af9ef7d),
	.w5(32'hba143160),
	.w6(32'h3aa654c3),
	.w7(32'h3ab09298),
	.w8(32'hba4bf533),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af5826),
	.w1(32'hb938eec8),
	.w2(32'h3aad0cd6),
	.w3(32'h3aed2c65),
	.w4(32'h3b23b5d0),
	.w5(32'h3bee7a10),
	.w6(32'hb9d23b78),
	.w7(32'h3a388eb9),
	.w8(32'h3c21c679),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85eece),
	.w1(32'h3c964c29),
	.w2(32'h3c16f7b0),
	.w3(32'h3ba7ebb6),
	.w4(32'h3c0a30e0),
	.w5(32'hbbc372ec),
	.w6(32'h3c3c5d3f),
	.w7(32'h3c6db244),
	.w8(32'hbb938e60),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a8b87),
	.w1(32'h3ae6bd2a),
	.w2(32'h3a9b263f),
	.w3(32'hba7ce7e5),
	.w4(32'hbb564e03),
	.w5(32'hba8cc3ec),
	.w6(32'h3a71bbb9),
	.w7(32'hb9037f47),
	.w8(32'h3b3b63f8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be443d0),
	.w1(32'h3c41f562),
	.w2(32'hb9b6ef17),
	.w3(32'h3bbb7212),
	.w4(32'h3c4b7af2),
	.w5(32'hbab4fc62),
	.w6(32'h39d833a9),
	.w7(32'h3be3ff63),
	.w8(32'hbc16433d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f870e),
	.w1(32'hbbbfa24c),
	.w2(32'hbc2bb773),
	.w3(32'hbb36372d),
	.w4(32'hbb4183fd),
	.w5(32'h3aceb47a),
	.w6(32'h3b619970),
	.w7(32'h3a83e58f),
	.w8(32'h3afbd270),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39583),
	.w1(32'h3b9ae55f),
	.w2(32'h3b2b7cee),
	.w3(32'h3b7e0964),
	.w4(32'hbb930305),
	.w5(32'hbb7c519b),
	.w6(32'hbaa223f4),
	.w7(32'hbb8f193f),
	.w8(32'hbb9a3017),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea9206),
	.w1(32'hbb9ad7b6),
	.w2(32'hbc3aff27),
	.w3(32'hbb95d9d4),
	.w4(32'hbac939c9),
	.w5(32'hbb48d605),
	.w6(32'hbbac5861),
	.w7(32'hbba49abe),
	.w8(32'hbb198b92),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa24d28),
	.w1(32'h3b61eab5),
	.w2(32'hb9d80f59),
	.w3(32'hba9456df),
	.w4(32'h3b84b2ae),
	.w5(32'hba2b2a16),
	.w6(32'h3b098f00),
	.w7(32'h3b0227b3),
	.w8(32'h3b31709d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa30d9),
	.w1(32'h3a60509e),
	.w2(32'h3b919807),
	.w3(32'hbb6f1d90),
	.w4(32'hbad60446),
	.w5(32'h3bae290c),
	.w6(32'h3b43a0df),
	.w7(32'h3affb217),
	.w8(32'h3b00388a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b187fe7),
	.w1(32'h3b1678ec),
	.w2(32'hbac26731),
	.w3(32'hba2ae8f4),
	.w4(32'hbaa53523),
	.w5(32'hbb967215),
	.w6(32'hb967520c),
	.w7(32'h3a025a59),
	.w8(32'hbc1078fb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc873355),
	.w1(32'hbbfd9b23),
	.w2(32'hbc545d0a),
	.w3(32'hbbd6f190),
	.w4(32'h3bbdf800),
	.w5(32'h3b09b797),
	.w6(32'hbb5b7f83),
	.w7(32'h3b3c5db3),
	.w8(32'h3b83f113),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57cc64),
	.w1(32'h3c0803ba),
	.w2(32'h3a36cb51),
	.w3(32'hbb21d2a8),
	.w4(32'h3c76ff8f),
	.w5(32'hbc0db92e),
	.w6(32'hbc3300d5),
	.w7(32'h3c44a989),
	.w8(32'hbc3753ce),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7dfa),
	.w1(32'h3b268d68),
	.w2(32'hbc3eae50),
	.w3(32'hbb6a2d48),
	.w4(32'h3c09435f),
	.w5(32'hbaba2d98),
	.w6(32'hbaa3e88a),
	.w7(32'h3c123549),
	.w8(32'hbc15e064),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d283d3),
	.w1(32'h3a3908cf),
	.w2(32'h39e793f5),
	.w3(32'h3aee48e6),
	.w4(32'h3ba63f0a),
	.w5(32'hb8ce9137),
	.w6(32'hb985a73d),
	.w7(32'h3b014ecd),
	.w8(32'hbb8dd581),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe47fe),
	.w1(32'hbb4a6a51),
	.w2(32'hba88a43b),
	.w3(32'hba60872c),
	.w4(32'hba825430),
	.w5(32'hbab57e1c),
	.w6(32'hbb7cb480),
	.w7(32'hbb25d733),
	.w8(32'hba97f775),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae25fe6),
	.w1(32'hba075ee1),
	.w2(32'h3aaf84f4),
	.w3(32'h3ad9eedd),
	.w4(32'h3ae61607),
	.w5(32'h3a9a2c90),
	.w6(32'h3b471817),
	.w7(32'h3b04fe95),
	.w8(32'h3ba2abce),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82af1ef),
	.w1(32'h3bb0e303),
	.w2(32'hba1251c7),
	.w3(32'h3ad87c62),
	.w4(32'h3b787590),
	.w5(32'hbba27358),
	.w6(32'hba603a2a),
	.w7(32'h3bd96cf9),
	.w8(32'hbb836c6b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42ca67),
	.w1(32'hbb921ff1),
	.w2(32'hbc7f2831),
	.w3(32'hbbf3d8df),
	.w4(32'hbb18010b),
	.w5(32'hbc252aa9),
	.w6(32'hbc52958f),
	.w7(32'hbbb154b4),
	.w8(32'hbc5761df),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b290),
	.w1(32'h3b9b3784),
	.w2(32'hbbe1b091),
	.w3(32'hbaaa37df),
	.w4(32'h3bd2dd0e),
	.w5(32'h3a0844a8),
	.w6(32'hbb71ede7),
	.w7(32'h3b8438c7),
	.w8(32'hbb4952a1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18a16e),
	.w1(32'h3c0e90a7),
	.w2(32'hbb499260),
	.w3(32'h3b7a2454),
	.w4(32'h3c2cafa2),
	.w5(32'hbbaafccc),
	.w6(32'h3b745625),
	.w7(32'h3c1ba515),
	.w8(32'hbc190d26),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde5406),
	.w1(32'hba0b9d5b),
	.w2(32'hbbc3cfcf),
	.w3(32'hbb5220bd),
	.w4(32'h3b4941e0),
	.w5(32'hbb32e1b0),
	.w6(32'hbbc66e15),
	.w7(32'h3a234584),
	.w8(32'hbba29eb2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc086c4f),
	.w1(32'hbb9cda9e),
	.w2(32'hbb21d2d2),
	.w3(32'hbc41c672),
	.w4(32'hbbfce433),
	.w5(32'hbb87e0a1),
	.w6(32'hbc897587),
	.w7(32'hbc023f27),
	.w8(32'hbb0c91e5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95a689),
	.w1(32'h3a78da00),
	.w2(32'hbba85bd1),
	.w3(32'hba806497),
	.w4(32'hbabdefb2),
	.w5(32'h3af02efe),
	.w6(32'hb992fb3e),
	.w7(32'hbabab911),
	.w8(32'h3a4c612d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac47533),
	.w1(32'h3a36d6ed),
	.w2(32'h3b8793f3),
	.w3(32'h3b4e7490),
	.w4(32'h3be3efc0),
	.w5(32'hbb590c81),
	.w6(32'h3b2611c8),
	.w7(32'h3b45bb2d),
	.w8(32'hbbdfc830),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf58dc9),
	.w1(32'h3abd9065),
	.w2(32'hb8e08d1f),
	.w3(32'hbb2ddf6d),
	.w4(32'hbb1038b4),
	.w5(32'hbaa91339),
	.w6(32'hbb02172a),
	.w7(32'hba574cbf),
	.w8(32'hbaa888f1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff7f60),
	.w1(32'hbaf5168a),
	.w2(32'hbbf49160),
	.w3(32'hbb8f0462),
	.w4(32'hbac2d034),
	.w5(32'hbbacee78),
	.w6(32'hbb6355c8),
	.w7(32'hba854381),
	.w8(32'hbc0be91b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bbf4e0),
	.w1(32'h3b94d29c),
	.w2(32'h38fdc7dd),
	.w3(32'h3ae8ed26),
	.w4(32'hb6ead7b1),
	.w5(32'hbb395d88),
	.w6(32'hba93cf47),
	.w7(32'h3b167e94),
	.w8(32'hbbb17b4a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc492609),
	.w1(32'hba217164),
	.w2(32'hbba1e438),
	.w3(32'hbb4086f7),
	.w4(32'hbb40f849),
	.w5(32'hbb56d5e2),
	.w6(32'hba98632f),
	.w7(32'hbab3a769),
	.w8(32'hbb9489d5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888c88),
	.w1(32'h3a35e9e1),
	.w2(32'hbb4a9d9d),
	.w3(32'hba4fcfe6),
	.w4(32'h3a4db45a),
	.w5(32'hbb77c74c),
	.w6(32'hbb7f39f1),
	.w7(32'hbb8b8d02),
	.w8(32'h3b60a294),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ad6c8),
	.w1(32'h3b48a829),
	.w2(32'h3c0b93f0),
	.w3(32'hbaae5ccd),
	.w4(32'hba79fad1),
	.w5(32'h3b58e5f8),
	.w6(32'h3b27e321),
	.w7(32'h3af02749),
	.w8(32'h3b4cb826),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e1a15),
	.w1(32'h3b151e56),
	.w2(32'h3b6da2a3),
	.w3(32'h3ae5a44a),
	.w4(32'h3b10788a),
	.w5(32'hbb390521),
	.w6(32'hba9bcea5),
	.w7(32'h3b2cbd17),
	.w8(32'hba2d0bbf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b1786),
	.w1(32'h3a93df05),
	.w2(32'h3aa50c7e),
	.w3(32'hbaaac577),
	.w4(32'hba399005),
	.w5(32'h3b607705),
	.w6(32'h3b50701a),
	.w7(32'h3847a609),
	.w8(32'h3a55fd0e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825dd7),
	.w1(32'h3b5e1398),
	.w2(32'h3b6f92e2),
	.w3(32'h3b89295b),
	.w4(32'h3bf8d411),
	.w5(32'h3ae39b76),
	.w6(32'h3b374335),
	.w7(32'h3bac031b),
	.w8(32'h3aae47b8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f8fe7),
	.w1(32'h390192bc),
	.w2(32'h3b634a2c),
	.w3(32'h3bbdc087),
	.w4(32'h3c181cac),
	.w5(32'hbbac0e25),
	.w6(32'h3b859994),
	.w7(32'h3bf37320),
	.w8(32'h3afae113),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b817e),
	.w1(32'hbb5c7846),
	.w2(32'hbbb97212),
	.w3(32'hbb9b073e),
	.w4(32'h3b1ead60),
	.w5(32'h3a40bc96),
	.w6(32'h3b9376eb),
	.w7(32'h3ba892bb),
	.w8(32'h3b5d0560),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c09a1),
	.w1(32'h3a986312),
	.w2(32'h39939cf8),
	.w3(32'h3aa1661e),
	.w4(32'h3ba0cefb),
	.w5(32'hbb74035f),
	.w6(32'h3bf0d0d8),
	.w7(32'h3bee8c10),
	.w8(32'hba9b993c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad21fa5),
	.w1(32'hba9f111e),
	.w2(32'h3a14981a),
	.w3(32'hbb72efab),
	.w4(32'hbb3d780b),
	.w5(32'hbb8148da),
	.w6(32'h3b143dee),
	.w7(32'hba5e1cd7),
	.w8(32'hbb3ff915),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99fca8),
	.w1(32'hbb51176a),
	.w2(32'hba164c2a),
	.w3(32'hbb95523d),
	.w4(32'hbaf0081b),
	.w5(32'hbb354563),
	.w6(32'hbb47608b),
	.w7(32'hbb1a5389),
	.w8(32'h3b685b20),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2728a),
	.w1(32'h3b5e4589),
	.w2(32'h3bd1bf65),
	.w3(32'hbb12b1d8),
	.w4(32'h3b369b54),
	.w5(32'h3b26255d),
	.w6(32'h3a01b9a1),
	.w7(32'h3addc48e),
	.w8(32'hbb0b2c72),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91d68a),
	.w1(32'h3bbfdb23),
	.w2(32'h3b873f99),
	.w3(32'h3bed598d),
	.w4(32'h3b7587f2),
	.w5(32'h3ab24620),
	.w6(32'h3b2ad97e),
	.w7(32'hb9af82ea),
	.w8(32'h3a37d838),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc376a5f),
	.w1(32'hbb4577bf),
	.w2(32'hbbece7a2),
	.w3(32'hbaecccd5),
	.w4(32'h3aabbf96),
	.w5(32'hbb24897e),
	.w6(32'hbb55e0a7),
	.w7(32'hbb0373d7),
	.w8(32'hbb0fa6ad),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4521cc),
	.w1(32'hbb0b23c9),
	.w2(32'hbc29c24f),
	.w3(32'hbc4b66a2),
	.w4(32'hbb052b54),
	.w5(32'hbc4e8eb3),
	.w6(32'hbc8c1e10),
	.w7(32'hbb241215),
	.w8(32'hbc4f359b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29cb5e),
	.w1(32'h3b6ff215),
	.w2(32'hbbd1362b),
	.w3(32'hbc210d56),
	.w4(32'h3ba4e18c),
	.w5(32'hbb8fcb43),
	.w6(32'hbc4fbc42),
	.w7(32'h391b8965),
	.w8(32'hbbe98691),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc485c3f),
	.w1(32'h3aef20d2),
	.w2(32'hbc811d60),
	.w3(32'hbb874778),
	.w4(32'h3c35eff9),
	.w5(32'hbb9b2a41),
	.w6(32'hbc825002),
	.w7(32'hba3f55d0),
	.w8(32'hbc85fc04),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30419f),
	.w1(32'hbb6813ff),
	.w2(32'hbb21dda7),
	.w3(32'hba97cc0b),
	.w4(32'h39f0fc6e),
	.w5(32'h38eb02db),
	.w6(32'hbb9987d3),
	.w7(32'hbb028a1b),
	.w8(32'hbb91e613),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68aeacb),
	.w1(32'hbab24e91),
	.w2(32'h3ad0d4c9),
	.w3(32'hbb020632),
	.w4(32'hba8a6d02),
	.w5(32'hb9d3d001),
	.w6(32'hbb6b8235),
	.w7(32'hbb9d60cb),
	.w8(32'hb9c2d0a2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b583a5d),
	.w1(32'h3c265f2c),
	.w2(32'h3c19b2d1),
	.w3(32'h3a617715),
	.w4(32'hbae63f6f),
	.w5(32'hba3c07c6),
	.w6(32'hbb72aeef),
	.w7(32'h3b19124e),
	.w8(32'h3a8a0b0e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ee66),
	.w1(32'hba9bb2c1),
	.w2(32'h39f9cc2a),
	.w3(32'hbb991f4d),
	.w4(32'h3a913f23),
	.w5(32'hb9e955a7),
	.w6(32'h3b035179),
	.w7(32'h3b20c171),
	.w8(32'h3baf9036),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afba31a),
	.w1(32'h3b9f54bd),
	.w2(32'h3b984c04),
	.w3(32'h3b936841),
	.w4(32'h3b29e43c),
	.w5(32'hb81f55c3),
	.w6(32'h3b01cdf9),
	.w7(32'h3aea4f8e),
	.w8(32'h3b4e10b0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e0990),
	.w1(32'hb9af2e7d),
	.w2(32'hbb22f88c),
	.w3(32'hbbfb7f06),
	.w4(32'hbb91b600),
	.w5(32'hb96f495f),
	.w6(32'hbb966805),
	.w7(32'hba979c1c),
	.w8(32'hbbcd7ebb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c5ca1),
	.w1(32'hbb249441),
	.w2(32'hbb6775a6),
	.w3(32'hbb0cf301),
	.w4(32'h37fd4f72),
	.w5(32'hbb4e71b4),
	.w6(32'hbbfe0564),
	.w7(32'h3b216f06),
	.w8(32'hbbae04aa),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebbf06),
	.w1(32'h3a1058d4),
	.w2(32'hbb5effeb),
	.w3(32'hbbac3445),
	.w4(32'h3b0bf5a0),
	.w5(32'h3ab6c7af),
	.w6(32'hbbd1dcd0),
	.w7(32'h3abf7b19),
	.w8(32'hba14f1d9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07cb17),
	.w1(32'h3bd0f182),
	.w2(32'h3ab192fc),
	.w3(32'h3acbf8e9),
	.w4(32'h3b06a342),
	.w5(32'h3b722d51),
	.w6(32'hba4bda78),
	.w7(32'h3b70acdd),
	.w8(32'h3b5ae10b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9f8f),
	.w1(32'h3b4a6d57),
	.w2(32'h39d33582),
	.w3(32'h395deba9),
	.w4(32'h39f220c4),
	.w5(32'hba2bcec0),
	.w6(32'h3b904596),
	.w7(32'h3b20ddf4),
	.w8(32'hba04f4ce),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b237206),
	.w1(32'h3934527c),
	.w2(32'hbaf5c73e),
	.w3(32'h3b0bc255),
	.w4(32'h3ba6f46a),
	.w5(32'h3aff71ea),
	.w6(32'hbbb19a2a),
	.w7(32'hb9a44c6d),
	.w8(32'h3ba719a8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa274e),
	.w1(32'h39d26afe),
	.w2(32'hbb854084),
	.w3(32'hba925be1),
	.w4(32'hba076457),
	.w5(32'hbb8c82bf),
	.w6(32'h3afb334c),
	.w7(32'h3ac1b255),
	.w8(32'hbbd6abc9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6eac6),
	.w1(32'h3af1045d),
	.w2(32'h3a71dac1),
	.w3(32'h3a0fc972),
	.w4(32'h3b2b0555),
	.w5(32'hbba0228f),
	.w6(32'h3aa0f93b),
	.w7(32'h3b96da3a),
	.w8(32'hbbc0189c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7640c),
	.w1(32'hbb873e55),
	.w2(32'hbb8fabe1),
	.w3(32'hbba42df6),
	.w4(32'hbb6c0d2d),
	.w5(32'hbb6897d4),
	.w6(32'hbc1f38ae),
	.w7(32'hbbfbcf54),
	.w8(32'hbbb98024),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae870a8),
	.w1(32'h3a94c4f9),
	.w2(32'h389a85fe),
	.w3(32'hbb5e12a7),
	.w4(32'hbaafa226),
	.w5(32'h3b15c1da),
	.w6(32'hbb5949f2),
	.w7(32'hba89c829),
	.w8(32'h3b9a4783),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ce70e),
	.w1(32'h3be97b94),
	.w2(32'h3b0d6f8d),
	.w3(32'h3bcd24cc),
	.w4(32'hba317704),
	.w5(32'hbb8c21bc),
	.w6(32'h3c3c54d3),
	.w7(32'h3c49fefb),
	.w8(32'hbbcbe2c1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279167),
	.w1(32'hbb29284f),
	.w2(32'hbb5140f8),
	.w3(32'hbb4c8d72),
	.w4(32'h3b3a6ccf),
	.w5(32'h3aa07530),
	.w6(32'hbbf4cdd6),
	.w7(32'hb9a1a235),
	.w8(32'hbad6d049),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399402f3),
	.w1(32'h3ab55df9),
	.w2(32'hbac5c806),
	.w3(32'h3b0231d5),
	.w4(32'h3b6e78ba),
	.w5(32'h3b30cecb),
	.w6(32'h3b97486d),
	.w7(32'h3b3a33fc),
	.w8(32'h3b4927cf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1856a3),
	.w1(32'hb9e060f6),
	.w2(32'hba83951f),
	.w3(32'h3a0b49be),
	.w4(32'h3b99e4ab),
	.w5(32'h3b324c5a),
	.w6(32'h3a13eae3),
	.w7(32'h3b53beb4),
	.w8(32'hb8b1cc15),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2bd2b),
	.w1(32'h3aedfb5c),
	.w2(32'hbbb98b92),
	.w3(32'hbc4b17e8),
	.w4(32'hbb86d64b),
	.w5(32'hbaa6b461),
	.w6(32'hbc9eca1d),
	.w7(32'hbbdeff00),
	.w8(32'hbbdb8062),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc67dfc),
	.w1(32'h3bfc3546),
	.w2(32'hbb535094),
	.w3(32'hbb1ccef8),
	.w4(32'h3b7d1360),
	.w5(32'h3a87c64c),
	.w6(32'hbb8a8a4f),
	.w7(32'h3a016101),
	.w8(32'hbafd886a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d498a),
	.w1(32'hbc171ee4),
	.w2(32'hbb5d87f2),
	.w3(32'hbbba2f2f),
	.w4(32'h3b4214ce),
	.w5(32'hbb8a3c5c),
	.w6(32'hbb7b9f53),
	.w7(32'h3a8e0737),
	.w8(32'hbc3931ee),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e23b7),
	.w1(32'hba2134fd),
	.w2(32'hbbcb6b76),
	.w3(32'hbb96897e),
	.w4(32'hbb35c064),
	.w5(32'hbc257297),
	.w6(32'hbc14b0cc),
	.w7(32'hbbab7671),
	.w8(32'hbc205c57),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54ac6c),
	.w1(32'hbba8f418),
	.w2(32'hbc0b21d1),
	.w3(32'hbc24f176),
	.w4(32'h3a68cb81),
	.w5(32'h3b60ccb0),
	.w6(32'hbc570e4c),
	.w7(32'hbae4aee7),
	.w8(32'h398b7ac7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25d4b6),
	.w1(32'h3bc3fd8b),
	.w2(32'h3baa4498),
	.w3(32'hbafde4c5),
	.w4(32'h3bcbccee),
	.w5(32'hba90ed50),
	.w6(32'hbb6b63a3),
	.w7(32'h3b8d3484),
	.w8(32'hb9a33444),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4686e6),
	.w1(32'h3ba18c4c),
	.w2(32'h39d875cc),
	.w3(32'hba712416),
	.w4(32'h3be7270c),
	.w5(32'hbaf5dead),
	.w6(32'hbb9f9a74),
	.w7(32'h3c01e886),
	.w8(32'hbbad904e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56bf68),
	.w1(32'h3b6aee3c),
	.w2(32'h3afbd458),
	.w3(32'hb9c98bd4),
	.w4(32'hb70c959e),
	.w5(32'hba678554),
	.w6(32'hb9bbd8fc),
	.w7(32'h3a8d8a10),
	.w8(32'hbb93218c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d8a5),
	.w1(32'hbb968b77),
	.w2(32'hbc6caf31),
	.w3(32'hbbfeb60f),
	.w4(32'h3b9b19f7),
	.w5(32'hbc0f54d4),
	.w6(32'hbc17376a),
	.w7(32'h3a251d53),
	.w8(32'hbc3dd510),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc377305),
	.w1(32'hbc09188c),
	.w2(32'hbbe03513),
	.w3(32'hbc42a388),
	.w4(32'hbb71af1f),
	.w5(32'hbbab8ca6),
	.w6(32'hbc57fd91),
	.w7(32'hbbb6a4eb),
	.w8(32'hbb89871e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc481a58),
	.w1(32'hbb859c6d),
	.w2(32'hbb9505c8),
	.w3(32'hbc42dcd6),
	.w4(32'hbb1bf914),
	.w5(32'h3ac42a63),
	.w6(32'hbc412388),
	.w7(32'hbba2aab7),
	.w8(32'hbb978584),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbaaee),
	.w1(32'h3aec582c),
	.w2(32'hbbc840c9),
	.w3(32'hbac6de11),
	.w4(32'h3c2d6b02),
	.w5(32'h3ac63453),
	.w6(32'hbbc3647b),
	.w7(32'h3b8a3173),
	.w8(32'hbbf56237),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34952c),
	.w1(32'h3af7ebd1),
	.w2(32'hbc1a1ab1),
	.w3(32'hb9285a42),
	.w4(32'h3be68de1),
	.w5(32'hbb840d9f),
	.w6(32'hbc219f61),
	.w7(32'hb97ea2fb),
	.w8(32'hbc0181ff),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4141cd),
	.w1(32'hbbfd44a8),
	.w2(32'hbc014ce2),
	.w3(32'hbc08648f),
	.w4(32'hbb86b862),
	.w5(32'hbb744f63),
	.w6(32'hbbce3fc9),
	.w7(32'hbb1d1f79),
	.w8(32'hbb5db193),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a294040),
	.w1(32'hbafbfd5d),
	.w2(32'hbb3820af),
	.w3(32'hbac5864b),
	.w4(32'hbb69ee29),
	.w5(32'hbaac8506),
	.w6(32'hbb88ba91),
	.w7(32'hbb813f5a),
	.w8(32'hbafe6441),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fe5ed),
	.w1(32'hbbeb15d2),
	.w2(32'hbbea7df8),
	.w3(32'hbc380b66),
	.w4(32'hbafa5bfe),
	.w5(32'hbb4a8213),
	.w6(32'hbba78712),
	.w7(32'h3b78f6db),
	.w8(32'hbb87e5ac),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a0f80),
	.w1(32'hba8199c5),
	.w2(32'hbb3bb9a9),
	.w3(32'hbb4e92df),
	.w4(32'hbac4a4fc),
	.w5(32'hbbb64323),
	.w6(32'hbb072ddf),
	.w7(32'hbb17f002),
	.w8(32'hbbaff3c4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964883),
	.w1(32'hba5b2c3f),
	.w2(32'hba216297),
	.w3(32'hbb4ea43f),
	.w4(32'hba9db2e3),
	.w5(32'hb9ae6df4),
	.w6(32'hbb4e20eb),
	.w7(32'hb9513da2),
	.w8(32'hba864897),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506675),
	.w1(32'hbac628d1),
	.w2(32'hba2b6851),
	.w3(32'hba7ea11b),
	.w4(32'h3add8ffa),
	.w5(32'hbbe4e668),
	.w6(32'hba6bb09a),
	.w7(32'h3a606d61),
	.w8(32'hbc220b1c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd941),
	.w1(32'hbc2a4f63),
	.w2(32'hbc51420c),
	.w3(32'hbc3c0df5),
	.w4(32'hbbe50e82),
	.w5(32'hbc110847),
	.w6(32'hbc958d46),
	.w7(32'hbc399b51),
	.w8(32'hbc2fb2d4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12cdf4),
	.w1(32'hb8e8672d),
	.w2(32'hbbf7815a),
	.w3(32'hbb76c1c5),
	.w4(32'h3ab9410f),
	.w5(32'hbbb48cfc),
	.w6(32'hbbd678de),
	.w7(32'hba939695),
	.w8(32'hbbcf8c41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c60c7),
	.w1(32'h3ad10d8c),
	.w2(32'hbb9d417e),
	.w3(32'hbb6155dc),
	.w4(32'h3aaf8447),
	.w5(32'hbb40db66),
	.w6(32'hbb4f8d53),
	.w7(32'h39aaa8f5),
	.w8(32'hbb55102e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ba5d),
	.w1(32'h3a6c76f3),
	.w2(32'hbb3a4503),
	.w3(32'hb9aa41a5),
	.w4(32'h3b138965),
	.w5(32'h3a2df7d9),
	.w6(32'hba033d75),
	.w7(32'h3a9e5646),
	.w8(32'hbb4c257d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9c824),
	.w1(32'hba2c724b),
	.w2(32'hbad35780),
	.w3(32'hbb286bc7),
	.w4(32'h3aa55208),
	.w5(32'hba500493),
	.w6(32'hbb72a204),
	.w7(32'h38932450),
	.w8(32'hbb2968c5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cab56),
	.w1(32'hba2384b7),
	.w2(32'hbb81b466),
	.w3(32'hba93fabb),
	.w4(32'h3b3988aa),
	.w5(32'hba97e83a),
	.w6(32'hbb08e70b),
	.w7(32'h3af7e11d),
	.w8(32'hbb1d638f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06b6b8),
	.w1(32'h3b368e67),
	.w2(32'hbb615190),
	.w3(32'hbaffa74d),
	.w4(32'h3b037749),
	.w5(32'hbb76e7ec),
	.w6(32'hbb376003),
	.w7(32'hb9395c4d),
	.w8(32'hbb90b396),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381930f8),
	.w1(32'hb99614de),
	.w2(32'hba698734),
	.w3(32'hba1d1c4d),
	.w4(32'hb9e9802b),
	.w5(32'hba879b19),
	.w6(32'hba0c5cef),
	.w7(32'hba2e0f6a),
	.w8(32'hbac2ddd9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c687),
	.w1(32'hbb0fafe3),
	.w2(32'hbb291989),
	.w3(32'hbac44669),
	.w4(32'hba849366),
	.w5(32'h3b296356),
	.w6(32'hbadc272f),
	.w7(32'hbacf6ac3),
	.w8(32'hbac5b15b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff5036),
	.w1(32'hbb5519f2),
	.w2(32'h3abee60a),
	.w3(32'h3affd8bd),
	.w4(32'h3b67f29d),
	.w5(32'h3b4584ef),
	.w6(32'hb841969c),
	.w7(32'h3b05466d),
	.w8(32'h3accf69a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b206b80),
	.w1(32'hbadd152f),
	.w2(32'h3af9418d),
	.w3(32'hb810487e),
	.w4(32'h3b3d37c2),
	.w5(32'hbc009e9e),
	.w6(32'hbb2abe7f),
	.w7(32'h3aac88db),
	.w8(32'hbc0d9528),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd815a9),
	.w1(32'hbbe345e2),
	.w2(32'hbc374e10),
	.w3(32'hbc280ef1),
	.w4(32'hbb39ef75),
	.w5(32'hbbb6b79f),
	.w6(32'hbc834807),
	.w7(32'hbbe239fc),
	.w8(32'hbbab8c3b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0342d8),
	.w1(32'hbae2cc32),
	.w2(32'hbb2174f7),
	.w3(32'hbaeec242),
	.w4(32'hbae09073),
	.w5(32'hb9b96db1),
	.w6(32'hba813d26),
	.w7(32'hba73720d),
	.w8(32'hb930dbd4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78f2a2),
	.w1(32'hbb573a30),
	.w2(32'hbb26aa2d),
	.w3(32'hbabec196),
	.w4(32'hbaeb65fc),
	.w5(32'hbb90c0a9),
	.w6(32'hbaadfc4e),
	.w7(32'hb917fa4d),
	.w8(32'hbb9d2dd0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075d04),
	.w1(32'hba82cefe),
	.w2(32'hbc003152),
	.w3(32'hbba92b5f),
	.w4(32'h3a6398f7),
	.w5(32'hbb6e5a6a),
	.w6(32'hbbc14356),
	.w7(32'hba3947f2),
	.w8(32'hbbf9de8f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba646be1),
	.w1(32'hba1e49bf),
	.w2(32'hba4d4d6e),
	.w3(32'h3a9ef7be),
	.w4(32'hb9df43ac),
	.w5(32'hbaa4e0e2),
	.w6(32'h39c395e4),
	.w7(32'hb9df7237),
	.w8(32'hba14a877),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25b0c4),
	.w1(32'h3a445579),
	.w2(32'hba867bf3),
	.w3(32'hbac09531),
	.w4(32'hb953c45c),
	.w5(32'hb9995cb4),
	.w6(32'hba9372e7),
	.w7(32'hb9cd6173),
	.w8(32'hbadd180d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ea434),
	.w1(32'hba10529e),
	.w2(32'h3a2e5206),
	.w3(32'h3a61cb1b),
	.w4(32'h3a4c5fbf),
	.w5(32'h39b84ac7),
	.w6(32'h39a947ba),
	.w7(32'h3a8068fe),
	.w8(32'hb9f25d1d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1b262),
	.w1(32'hba4dac14),
	.w2(32'hb91cc711),
	.w3(32'hbac6d0c9),
	.w4(32'hb96fbc3e),
	.w5(32'h3a85044f),
	.w6(32'hbb4d3b7a),
	.w7(32'hbadccca4),
	.w8(32'hba935fe0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f91c),
	.w1(32'hbb48cb97),
	.w2(32'hbb6418bd),
	.w3(32'hbb3a4d29),
	.w4(32'hbb880567),
	.w5(32'hbb96ac5c),
	.w6(32'hbb8314eb),
	.w7(32'hbba2f0c1),
	.w8(32'hbb075875),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e57fa),
	.w1(32'hbb36367c),
	.w2(32'hbc0592c9),
	.w3(32'hbba0a456),
	.w4(32'hba6309fd),
	.w5(32'hbaf507ec),
	.w6(32'hbbcf3083),
	.w7(32'hbb07a1d9),
	.w8(32'hbb4ec45a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b5663),
	.w1(32'h3a81a0c9),
	.w2(32'h3b36f06c),
	.w3(32'h3aecadd3),
	.w4(32'h3b565448),
	.w5(32'h3ae7fb2a),
	.w6(32'h3b40658b),
	.w7(32'h3b528fcf),
	.w8(32'h3a82bd13),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab81a9e),
	.w1(32'h3aa26764),
	.w2(32'h3a3dddd9),
	.w3(32'hba8d5f4b),
	.w4(32'h3a9b83ab),
	.w5(32'hba88bf20),
	.w6(32'hbb4881ea),
	.w7(32'h3abdfba0),
	.w8(32'hbad0eb6f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aaaab),
	.w1(32'hba1de21a),
	.w2(32'hbacaa93d),
	.w3(32'hbad385c5),
	.w4(32'h3b037240),
	.w5(32'hbb3f43ff),
	.w6(32'hbb15dc76),
	.w7(32'h3aaf34db),
	.w8(32'hbb8e7bc0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e92d2),
	.w1(32'hbac23c04),
	.w2(32'hbb932b2b),
	.w3(32'hbb137367),
	.w4(32'h3b113dd1),
	.w5(32'hbb5f96ca),
	.w6(32'hbb9d95d7),
	.w7(32'h384b72fb),
	.w8(32'hbb857c7d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a1b85),
	.w1(32'hbb53b064),
	.w2(32'hbc07f422),
	.w3(32'hbbcc72f6),
	.w4(32'hba8c4ae0),
	.w5(32'hbaa98de3),
	.w6(32'hbbc7c3bc),
	.w7(32'hbb06b70e),
	.w8(32'hbb544a72),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0ae7d),
	.w1(32'hbb85590d),
	.w2(32'hbbc79beb),
	.w3(32'hbbe9bf79),
	.w4(32'hbac050f7),
	.w5(32'hbb9891d5),
	.w6(32'hbbd0401b),
	.w7(32'hbb21e31e),
	.w8(32'hbbd74494),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5b92d),
	.w1(32'h3aa87b81),
	.w2(32'hbb5623c0),
	.w3(32'hbb4f80bf),
	.w4(32'h3b549e57),
	.w5(32'hbb20eaf8),
	.w6(32'hbb79ec7d),
	.w7(32'h3af244d6),
	.w8(32'hbbd794f3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd54636),
	.w1(32'hbb93f460),
	.w2(32'hbb59cbf3),
	.w3(32'hbb8f96aa),
	.w4(32'h3a11e495),
	.w5(32'hbafcd462),
	.w6(32'hbbd55fd5),
	.w7(32'hbb2bdd75),
	.w8(32'hbba0f2b0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b5085),
	.w1(32'hbbdfa6cd),
	.w2(32'hbc0fb4c6),
	.w3(32'hbc0f4b93),
	.w4(32'hbbba2f6e),
	.w5(32'hbbcc44f4),
	.w6(32'hbbecd524),
	.w7(32'hbb4a5500),
	.w8(32'hbb71674c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb17a3a),
	.w1(32'hba9e1ae3),
	.w2(32'hbb67ac8d),
	.w3(32'hbb6a259a),
	.w4(32'h3a9e806f),
	.w5(32'hba6326e2),
	.w6(32'hbbb89cbc),
	.w7(32'hba1279db),
	.w8(32'hbb86b03d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7c220),
	.w1(32'h3aa16004),
	.w2(32'hbb295d69),
	.w3(32'hba68b0d4),
	.w4(32'h3af719d8),
	.w5(32'hbb964699),
	.w6(32'hbb50423a),
	.w7(32'h3ad0b9f5),
	.w8(32'hbb5c5e7a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad593f9),
	.w1(32'h39c3d0f0),
	.w2(32'hbb906bd7),
	.w3(32'hbad45fc7),
	.w4(32'hbb1ce6f3),
	.w5(32'hbb443c88),
	.w6(32'hba2bc99c),
	.w7(32'hbb0e00ce),
	.w8(32'hbb3c2049),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f57f),
	.w1(32'h3b812112),
	.w2(32'hbb5e9bb5),
	.w3(32'hbb415281),
	.w4(32'h3b6a3a7c),
	.w5(32'hbbcd3839),
	.w6(32'hbb4ab946),
	.w7(32'h3b2bab97),
	.w8(32'hbc003c7c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5138b6),
	.w1(32'h3a1b6122),
	.w2(32'hba9adec5),
	.w3(32'hbba3ff07),
	.w4(32'hba85ab23),
	.w5(32'hba89c23e),
	.w6(32'hbb722a35),
	.w7(32'hb8acdf2c),
	.w8(32'hbb2d7cce),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e6686),
	.w1(32'hba70493d),
	.w2(32'h3a53f87d),
	.w3(32'h38ee079f),
	.w4(32'h3a3840c4),
	.w5(32'h39321487),
	.w6(32'h389aad91),
	.w7(32'h378f6c63),
	.w8(32'hb9caf336),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e7cc6),
	.w1(32'hbae0e44e),
	.w2(32'hbaa7a1ca),
	.w3(32'hba7482db),
	.w4(32'hbacb718b),
	.w5(32'hb9814133),
	.w6(32'hb9834609),
	.w7(32'hbae0482b),
	.w8(32'hb9efa32b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafadcdd),
	.w1(32'h39bab095),
	.w2(32'hba72679e),
	.w3(32'hbb17166e),
	.w4(32'hb88ff9d2),
	.w5(32'hbb09e2b8),
	.w6(32'hbb3da607),
	.w7(32'hba22068f),
	.w8(32'hbb82e26b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4af2),
	.w1(32'hbb9515c3),
	.w2(32'hbbf684ff),
	.w3(32'hbbffcd3e),
	.w4(32'hba8e3b8b),
	.w5(32'hbaba6c0b),
	.w6(32'hbc2639b9),
	.w7(32'hbb658c75),
	.w8(32'hbba55105),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce7a3),
	.w1(32'h3b8cfbd8),
	.w2(32'h3a5278b2),
	.w3(32'hbbda1f71),
	.w4(32'h3a420286),
	.w5(32'hbb2271ae),
	.w6(32'hbb77e57b),
	.w7(32'h3b49984a),
	.w8(32'hbb39b213),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9881055),
	.w1(32'hba8bb4cb),
	.w2(32'hbac02740),
	.w3(32'h3ad1af2b),
	.w4(32'h38be09d3),
	.w5(32'h3a97548c),
	.w6(32'h3a9f888f),
	.w7(32'hba3e1921),
	.w8(32'h3a4921dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5caf82),
	.w1(32'h3a3f4ad6),
	.w2(32'hbbbb3796),
	.w3(32'hbb216608),
	.w4(32'h3b34d2e1),
	.w5(32'hbb62f34c),
	.w6(32'hbbaa4b8c),
	.w7(32'hb99e476b),
	.w8(32'hbb96f304),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba526598),
	.w1(32'h3b012291),
	.w2(32'hbb6d33ee),
	.w3(32'hbb09c014),
	.w4(32'h3a31a65e),
	.w5(32'hbb2bbd27),
	.w6(32'hbb805ae6),
	.w7(32'hba93a6ee),
	.w8(32'hbb707651),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc240a1c),
	.w1(32'hbbcba1a0),
	.w2(32'hbbe2cb64),
	.w3(32'hbbe8317d),
	.w4(32'hbb8bce0b),
	.w5(32'hbb73fb0c),
	.w6(32'hbb7c3383),
	.w7(32'hbb0dcd1a),
	.w8(32'hbbad9a25),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5214),
	.w1(32'h3b3674a0),
	.w2(32'hbbdaad44),
	.w3(32'hbb7c55a3),
	.w4(32'h3b867585),
	.w5(32'hbb0d4ad8),
	.w6(32'hbb9d3de6),
	.w7(32'h3ae41fa3),
	.w8(32'hbbb82163),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c7e9b),
	.w1(32'hbacbcf1c),
	.w2(32'hbb10fefe),
	.w3(32'hbb8abe05),
	.w4(32'hbad43b51),
	.w5(32'hbb406f80),
	.w6(32'hbae88cee),
	.w7(32'hba57c1d0),
	.w8(32'hbb9c7487),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba911ace),
	.w1(32'hbacfdc9c),
	.w2(32'hba960dd3),
	.w3(32'hba6fd9c0),
	.w4(32'hba68bf91),
	.w5(32'hbb06ce42),
	.w6(32'hbacf375b),
	.w7(32'hbafc2c58),
	.w8(32'hbb0fca9a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50531c),
	.w1(32'hb9ae003d),
	.w2(32'hbb6bb251),
	.w3(32'hbad1ba59),
	.w4(32'h3b56e22f),
	.w5(32'h3af06a52),
	.w6(32'hbba44d53),
	.w7(32'h3a29f2fe),
	.w8(32'hbad97bfc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8e48),
	.w1(32'h3a22b6a0),
	.w2(32'hbadd99a2),
	.w3(32'h38cc811e),
	.w4(32'h3bbb054e),
	.w5(32'hba25570b),
	.w6(32'hbb1c580b),
	.w7(32'h3b75a022),
	.w8(32'hbb2b9719),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23d8dc),
	.w1(32'h3b1d1528),
	.w2(32'hbb74cca2),
	.w3(32'h3a81cf96),
	.w4(32'h3b0f989a),
	.w5(32'h39ad23e2),
	.w6(32'hba12e4fb),
	.w7(32'h3af9272d),
	.w8(32'hba83c0b8),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9714e57),
	.w1(32'h39c0946f),
	.w2(32'h3a67e1ed),
	.w3(32'hbb1863bb),
	.w4(32'hb9ab9d0a),
	.w5(32'h39470de1),
	.w6(32'h38d13cda),
	.w7(32'h3b2bb1b1),
	.w8(32'h3afbb5d0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e1136),
	.w1(32'h3ae8370b),
	.w2(32'hba3b1fb2),
	.w3(32'h39788b80),
	.w4(32'hba0b05b7),
	.w5(32'h39c44dea),
	.w6(32'h3a5b436d),
	.w7(32'h3a39514a),
	.w8(32'hba38e0e5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7eaf),
	.w1(32'hbb51232c),
	.w2(32'hbbc1f51f),
	.w3(32'hbba940ba),
	.w4(32'hbb33826f),
	.w5(32'hbac7ab78),
	.w6(32'hbbb06d17),
	.w7(32'hbb6010ff),
	.w8(32'hbb4d92d5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6065fb),
	.w1(32'hba0f6e6b),
	.w2(32'h3a76fa3a),
	.w3(32'h392f4658),
	.w4(32'h39afca3b),
	.w5(32'hbb1694dd),
	.w6(32'h390f07e9),
	.w7(32'h3a1cb768),
	.w8(32'hba86cc2e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4f071),
	.w1(32'h3aa8b5d4),
	.w2(32'hbb19eae6),
	.w3(32'h39a256d8),
	.w4(32'h3b3a7174),
	.w5(32'hba8d29d6),
	.w6(32'h39e60d52),
	.w7(32'h3b44590d),
	.w8(32'hbac728e9),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beca36),
	.w1(32'hbaa8f865),
	.w2(32'hbb181661),
	.w3(32'h3a0a0051),
	.w4(32'hba8b762a),
	.w5(32'h3a7c8fe8),
	.w6(32'hba3b0818),
	.w7(32'hbad118d7),
	.w8(32'hb7b2f0f3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad0a0),
	.w1(32'hbb06b108),
	.w2(32'hbb8894c9),
	.w3(32'hbb1994e0),
	.w4(32'hbaca3d8b),
	.w5(32'hbbbaec68),
	.w6(32'hbacb798c),
	.w7(32'hb982264c),
	.w8(32'hbbd465b3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e94ad),
	.w1(32'hb9fd50e3),
	.w2(32'hba7330f2),
	.w3(32'h3a353e14),
	.w4(32'h3a143987),
	.w5(32'hbabd990f),
	.w6(32'h3a38d486),
	.w7(32'hba34c302),
	.w8(32'hb9e7471c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcc49e),
	.w1(32'hb9aeca15),
	.w2(32'hba419d8b),
	.w3(32'hba34f9ea),
	.w4(32'hbaa52fce),
	.w5(32'h3a44eacf),
	.w6(32'h389c1484),
	.w7(32'hba4d3385),
	.w8(32'hba77d0cf),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ede1),
	.w1(32'hbb346566),
	.w2(32'hbb67bc4b),
	.w3(32'hbab6711f),
	.w4(32'h3b3a62f6),
	.w5(32'hba265548),
	.w6(32'hbc06bf6e),
	.w7(32'hb9a48fc0),
	.w8(32'hbb404bde),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79820a),
	.w1(32'h3b289b36),
	.w2(32'hbbd25c82),
	.w3(32'hbafa0b7d),
	.w4(32'h3b28ae43),
	.w5(32'hbc159c11),
	.w6(32'hbbb10007),
	.w7(32'h3994d99f),
	.w8(32'hbc21bddb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9ceb3),
	.w1(32'h39b5cf51),
	.w2(32'hbb2446bb),
	.w3(32'h3952cbc3),
	.w4(32'h39ca2e22),
	.w5(32'hba2871bc),
	.w6(32'hba80bce3),
	.w7(32'hba45d3b9),
	.w8(32'hbac13536),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7dc9e),
	.w1(32'h3b458f96),
	.w2(32'hbb066dfa),
	.w3(32'h388bab0f),
	.w4(32'h3bc91b0d),
	.w5(32'hbbc4325d),
	.w6(32'hbac9922e),
	.w7(32'h3b99ba2c),
	.w8(32'hbc250c40),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9817ee),
	.w1(32'hb9aa066a),
	.w2(32'h3a67c2e2),
	.w3(32'hbb94aa39),
	.w4(32'hb7a8fdbe),
	.w5(32'hbadf1d9e),
	.w6(32'hbb20d399),
	.w7(32'hb89567a1),
	.w8(32'hbafa241a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0057),
	.w1(32'hba736f21),
	.w2(32'hbbffe9ef),
	.w3(32'hbbfe795c),
	.w4(32'h3af4cf9e),
	.w5(32'h3a90faf6),
	.w6(32'hbc4a018d),
	.w7(32'hbabf70d5),
	.w8(32'hba9bc8d3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe136),
	.w1(32'h3ae8983a),
	.w2(32'hbb4b42b5),
	.w3(32'hbb241a95),
	.w4(32'h3b9515aa),
	.w5(32'hbbafa406),
	.w6(32'hbad02283),
	.w7(32'h3b7872c1),
	.w8(32'hbbda5ace),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52c52f),
	.w1(32'hba1da169),
	.w2(32'hbbe2878d),
	.w3(32'hbb8ffc33),
	.w4(32'h3a3954d2),
	.w5(32'hbb62c798),
	.w6(32'hbbc3756b),
	.w7(32'hba2021ed),
	.w8(32'hbb9a6431),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a944ca5),
	.w1(32'h396d8af0),
	.w2(32'hb60ec3a4),
	.w3(32'h3a9a7b98),
	.w4(32'h3a6c7046),
	.w5(32'hba231422),
	.w6(32'h3a0d7262),
	.w7(32'h396cca84),
	.w8(32'h3a0ac977),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909f8a),
	.w1(32'hba63b0cd),
	.w2(32'hbb918744),
	.w3(32'hbb4606e9),
	.w4(32'hba72d107),
	.w5(32'h3aa64c14),
	.w6(32'hb997d3e7),
	.w7(32'h3a7cccf2),
	.w8(32'h3977b3ac),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ffc90),
	.w1(32'h39ae8634),
	.w2(32'h3ae0f4b0),
	.w3(32'h3aaaae23),
	.w4(32'h3b0c1c6b),
	.w5(32'hbb3cf74a),
	.w6(32'hb916608e),
	.w7(32'h3a7d6c61),
	.w8(32'hbaf86859),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba01dc),
	.w1(32'hbb3fe7e6),
	.w2(32'hba839741),
	.w3(32'hbb880318),
	.w4(32'hba96b083),
	.w5(32'h3b0ea029),
	.w6(32'hbba6a772),
	.w7(32'hbb178f90),
	.w8(32'hbad9390e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba815ebd),
	.w1(32'h39230ee0),
	.w2(32'h3a86efc9),
	.w3(32'h39a66371),
	.w4(32'h3aa2ebda),
	.w5(32'hbb336024),
	.w6(32'h3a0ff4f7),
	.w7(32'h3aebbcca),
	.w8(32'hbab816e2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaa683),
	.w1(32'hbab5467a),
	.w2(32'hbba7067c),
	.w3(32'hbbd66839),
	.w4(32'hbadba19f),
	.w5(32'hbab81e19),
	.w6(32'hbbc238bb),
	.w7(32'hbac6a7ee),
	.w8(32'hbb79b769),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992b2ce),
	.w1(32'h39e79549),
	.w2(32'h3a6f2136),
	.w3(32'hb94f6822),
	.w4(32'hba705b4e),
	.w5(32'hb9f469a8),
	.w6(32'h39218b95),
	.w7(32'h37b2fab2),
	.w8(32'h3a863677),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0512f6),
	.w1(32'h3a8d2a61),
	.w2(32'hb92c779f),
	.w3(32'hba2ff60e),
	.w4(32'hba6e1aa7),
	.w5(32'hbaee371e),
	.w6(32'h39eb8147),
	.w7(32'hb98e13af),
	.w8(32'hbad65620),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7901),
	.w1(32'hba669944),
	.w2(32'hba8571bb),
	.w3(32'hbaa88605),
	.w4(32'h3b004bd9),
	.w5(32'hba44434b),
	.w6(32'h380612db),
	.w7(32'h3aeaaf84),
	.w8(32'hba9cfaeb),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafaf18),
	.w1(32'hbae53947),
	.w2(32'hbb8cfbae),
	.w3(32'hbbb2742a),
	.w4(32'h38c3f523),
	.w5(32'hba26a727),
	.w6(32'hbbb0d337),
	.w7(32'hbb63e1af),
	.w8(32'hbaacc6d7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb259ea4),
	.w1(32'h3a3983a7),
	.w2(32'h379b1de9),
	.w3(32'hb9f1a20f),
	.w4(32'h3aebb910),
	.w5(32'h3b251878),
	.w6(32'h3acb83df),
	.w7(32'h3b7d488d),
	.w8(32'h3a4665a4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0596de),
	.w1(32'h3a02c78f),
	.w2(32'h3a9896cf),
	.w3(32'h3a0ef20f),
	.w4(32'h3b2a6ac3),
	.w5(32'hbb38c56a),
	.w6(32'hba815615),
	.w7(32'h3a3404e5),
	.w8(32'hbb251ef8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99c3c9),
	.w1(32'h3c06d791),
	.w2(32'hbb3becb5),
	.w3(32'hbb25d060),
	.w4(32'h3c00308b),
	.w5(32'hbaf5c6f1),
	.w6(32'hba807db1),
	.w7(32'h3c30d7e2),
	.w8(32'h3a6d50c4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2c5a4),
	.w1(32'h3ad9b5ff),
	.w2(32'hbc186f04),
	.w3(32'hbb636b5c),
	.w4(32'h3c0408df),
	.w5(32'hbb62667c),
	.w6(32'hbb9dbf55),
	.w7(32'h3bc082da),
	.w8(32'hbbb88cad),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83f95f2),
	.w1(32'hb80bda5f),
	.w2(32'hba1dec28),
	.w3(32'hb951f700),
	.w4(32'h387859ea),
	.w5(32'hbb595489),
	.w6(32'h3ac4bc1b),
	.w7(32'h3a7f7a83),
	.w8(32'hbb345b55),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac9676),
	.w1(32'hbad56e13),
	.w2(32'hbab40420),
	.w3(32'hbb123396),
	.w4(32'hbb19af5d),
	.w5(32'hba183380),
	.w6(32'hba8a6d33),
	.w7(32'hba1de915),
	.w8(32'hba375345),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f5f4c),
	.w1(32'h3a397ded),
	.w2(32'h3a362cc0),
	.w3(32'h3a07bb9a),
	.w4(32'h391c7082),
	.w5(32'hb7917857),
	.w6(32'h3a6d6a15),
	.w7(32'hb953da6b),
	.w8(32'h3a9155fd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932cadd),
	.w1(32'hba9a0925),
	.w2(32'hbb25601e),
	.w3(32'hbae18ce3),
	.w4(32'hbb1f5f0a),
	.w5(32'hbb127621),
	.w6(32'hba641131),
	.w7(32'hbb1ebc8e),
	.w8(32'hbaa9dc13),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6ab54),
	.w1(32'hbb0e69b8),
	.w2(32'hbb53378a),
	.w3(32'hbb8b9500),
	.w4(32'hbb7a04c0),
	.w5(32'hbace68a1),
	.w6(32'hbb38b164),
	.w7(32'hbaf91116),
	.w8(32'hbafe2718),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd9287),
	.w1(32'hbb3579e9),
	.w2(32'hbb46f62b),
	.w3(32'hbb51cf80),
	.w4(32'h3ac71e36),
	.w5(32'hbb2bcccf),
	.w6(32'hbb605482),
	.w7(32'hb8810b50),
	.w8(32'hbb4f7fd4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5174b1),
	.w1(32'h3be4c40d),
	.w2(32'h39f0bc32),
	.w3(32'hbb441422),
	.w4(32'h3bc886ce),
	.w5(32'hba330c65),
	.w6(32'hbb6ee4c1),
	.w7(32'h3bba3182),
	.w8(32'hbb65335c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a082e0b),
	.w1(32'h397f71cc),
	.w2(32'hbb185411),
	.w3(32'hba44193b),
	.w4(32'hb937d3a4),
	.w5(32'hb954c821),
	.w6(32'h389a149f),
	.w7(32'hba294f56),
	.w8(32'hbae95367),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8521a),
	.w1(32'h39f322af),
	.w2(32'hbbbceecf),
	.w3(32'hbb8860ee),
	.w4(32'h3b11c17c),
	.w5(32'hbad05204),
	.w6(32'hbb9da8ea),
	.w7(32'h390cd15f),
	.w8(32'hbb962965),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801d1e),
	.w1(32'hb938e252),
	.w2(32'hb9c916d6),
	.w3(32'hba0fb80d),
	.w4(32'h39ba9eb6),
	.w5(32'hbaa2ea08),
	.w6(32'hba274474),
	.w7(32'hb8177f8c),
	.w8(32'hba689e4d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381344fb),
	.w1(32'hb8a84531),
	.w2(32'hb8ced192),
	.w3(32'h3a0c00b8),
	.w4(32'h379c8459),
	.w5(32'h399ff187),
	.w6(32'h38e63cca),
	.w7(32'hb75d24f3),
	.w8(32'hba2549e9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabb0ce),
	.w1(32'hba8849cd),
	.w2(32'hba3635e0),
	.w3(32'hb9ed519a),
	.w4(32'h38f4b00f),
	.w5(32'h3ab80070),
	.w6(32'h3760e93f),
	.w7(32'h39f4ecfb),
	.w8(32'h3afa7904),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a4172),
	.w1(32'h3a883066),
	.w2(32'h3aafe1d7),
	.w3(32'h3a11567e),
	.w4(32'hb9b8def4),
	.w5(32'h3a0c5ac6),
	.w6(32'h3abcbe65),
	.w7(32'h3a151f04),
	.w8(32'h3a88b0f8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12b22d),
	.w1(32'h3a0af03a),
	.w2(32'hbb56ff05),
	.w3(32'hbb0d6f02),
	.w4(32'h3960143a),
	.w5(32'hbb9729cf),
	.w6(32'hbb386048),
	.w7(32'hb81d6b44),
	.w8(32'hbb92420c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094478),
	.w1(32'h3a867e32),
	.w2(32'hbbeecca2),
	.w3(32'hbbaa7ded),
	.w4(32'h3b02792b),
	.w5(32'hbb31da34),
	.w6(32'hbbddd12a),
	.w7(32'h3a5b6628),
	.w8(32'hbbba1b1a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bbc73),
	.w1(32'h3a17b761),
	.w2(32'hbbc3aef4),
	.w3(32'hbb8a51f0),
	.w4(32'h3ae1d482),
	.w5(32'hbb464317),
	.w6(32'hbbc1db88),
	.w7(32'hb9b64edf),
	.w8(32'hbbddb47b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a097d65),
	.w1(32'h3940be48),
	.w2(32'h3a76747c),
	.w3(32'hb9f80e8c),
	.w4(32'h3a2c1e42),
	.w5(32'hbb2ba4a2),
	.w6(32'hbb3876bb),
	.w7(32'hb95b3862),
	.w8(32'hbb1d83e7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba829a4),
	.w1(32'h3a326611),
	.w2(32'hbbca39b7),
	.w3(32'hbbb71d87),
	.w4(32'h3ad49144),
	.w5(32'hbb95556a),
	.w6(32'hbc0b6bda),
	.w7(32'h3884733b),
	.w8(32'hbc1bf95c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833de0),
	.w1(32'hbad08834),
	.w2(32'hbb89a901),
	.w3(32'hbb8acc2a),
	.w4(32'hb9c05690),
	.w5(32'hbae8f8b4),
	.w6(32'hbba765ab),
	.w7(32'hbaae27b7),
	.w8(32'hbafbf84c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f141),
	.w1(32'h3b602141),
	.w2(32'hbb7d9e22),
	.w3(32'hbbdac944),
	.w4(32'h3aac0ffc),
	.w5(32'hbb28d684),
	.w6(32'hbbffb722),
	.w7(32'h3b302d49),
	.w8(32'hbb8d73ba),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb2264),
	.w1(32'h3927d57a),
	.w2(32'h39892338),
	.w3(32'h399e2f53),
	.w4(32'h3a173c51),
	.w5(32'h38a897b3),
	.w6(32'h3a3aa5cd),
	.w7(32'h3a5a3afa),
	.w8(32'h391e9c38),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba304286),
	.w1(32'hbabe20be),
	.w2(32'hbb49903d),
	.w3(32'hbab28ea0),
	.w4(32'hbb26b385),
	.w5(32'h38753ad7),
	.w6(32'hbaf59dce),
	.w7(32'hbb207530),
	.w8(32'h3a0e3e52),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa0f5a),
	.w1(32'h3ab3f537),
	.w2(32'hbb8d0bbd),
	.w3(32'hbb5e1075),
	.w4(32'h3b03ff4b),
	.w5(32'hbb3da672),
	.w6(32'hbbbe6c37),
	.w7(32'hb892a95a),
	.w8(32'hbba160be),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50c705),
	.w1(32'h3b1fe463),
	.w2(32'hbc02e42b),
	.w3(32'hbb61690e),
	.w4(32'h3b16089a),
	.w5(32'hbbe9beca),
	.w6(32'hbbfb3178),
	.w7(32'hb9776b21),
	.w8(32'hbb86f001),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86e57a),
	.w1(32'h3b2e39a0),
	.w2(32'hbba3e931),
	.w3(32'hbb462767),
	.w4(32'h3bb80d9c),
	.w5(32'hbada8cc3),
	.w6(32'hbb9bcd7c),
	.w7(32'h3b4638b0),
	.w8(32'hbba10a2b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad55c26),
	.w1(32'hbb34da3f),
	.w2(32'hb948f7bb),
	.w3(32'hbb417cdb),
	.w4(32'hbb5ecabc),
	.w5(32'hbb2f77b4),
	.w6(32'h3aa3402f),
	.w7(32'h3951d2f2),
	.w8(32'hbb0b7f28),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa93345),
	.w1(32'hbaaa032c),
	.w2(32'hb9315c2e),
	.w3(32'h3a675953),
	.w4(32'h3a1e86d8),
	.w5(32'hba504bb3),
	.w6(32'hb58e4109),
	.w7(32'h39f15339),
	.w8(32'hbaf62045),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8eb7a),
	.w1(32'hbb33012e),
	.w2(32'hbac903aa),
	.w3(32'hbb1aa51c),
	.w4(32'hbaa954dd),
	.w5(32'hb72ee6bb),
	.w6(32'hbb4de03f),
	.w7(32'hbb1e6ea9),
	.w8(32'hba2a400a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba023a5),
	.w1(32'hbaf0bdbc),
	.w2(32'hbb8767c7),
	.w3(32'hbb73a895),
	.w4(32'hba948875),
	.w5(32'hbb838e83),
	.w6(32'hbb79ac55),
	.w7(32'hba3bce7b),
	.w8(32'hbaea3dff),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf76f41),
	.w1(32'h3aed8c5f),
	.w2(32'hbb283e61),
	.w3(32'hbb002dd7),
	.w4(32'h3b0ef302),
	.w5(32'hbb8c029a),
	.w6(32'hba9081c0),
	.w7(32'h3b225ad5),
	.w8(32'hbb3c77ca),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42af9f),
	.w1(32'hbc153113),
	.w2(32'hbbeda2a9),
	.w3(32'hbc1592e9),
	.w4(32'hbbfc5c6e),
	.w5(32'hbbde2499),
	.w6(32'hbc0ffc94),
	.w7(32'hbc008e48),
	.w8(32'hbbe86c87),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb1b4),
	.w1(32'h3b22490f),
	.w2(32'hbb820734),
	.w3(32'hbb91f5c4),
	.w4(32'h3b4784fc),
	.w5(32'h3ab161bf),
	.w6(32'hbbe03042),
	.w7(32'hba0ab984),
	.w8(32'hbb20dd2f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c3e9d),
	.w1(32'h3b97fb83),
	.w2(32'hbb069556),
	.w3(32'h3acd0e8f),
	.w4(32'h3c233631),
	.w5(32'h3ac52631),
	.w6(32'hbb286c6f),
	.w7(32'h3bbc8b4d),
	.w8(32'hbb158caa),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafec37),
	.w1(32'h3ac2c11e),
	.w2(32'h39177df6),
	.w3(32'h3b213cc7),
	.w4(32'h3ad85c26),
	.w5(32'hb7a4cfe1),
	.w6(32'h3b51e960),
	.w7(32'h3acc112b),
	.w8(32'hba356d40),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eac75a),
	.w1(32'hb9823568),
	.w2(32'h3a3f0f4f),
	.w3(32'h38c2eb7b),
	.w4(32'hb8fa933d),
	.w5(32'hbae44a05),
	.w6(32'hb8f23901),
	.w7(32'h3ad40ac6),
	.w8(32'hb9bfd2ee),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f93075),
	.w1(32'hb98482ea),
	.w2(32'h39852d17),
	.w3(32'hbb510759),
	.w4(32'hbb6858c1),
	.w5(32'hb862cffb),
	.w6(32'hbb86cf4b),
	.w7(32'hbb38b12d),
	.w8(32'hb9c13da5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e99e2),
	.w1(32'h3a41a8bf),
	.w2(32'hb8bb920f),
	.w3(32'hba34f27b),
	.w4(32'hba7d04a8),
	.w5(32'hba4f36fa),
	.w6(32'h3a3ffb9e),
	.w7(32'hb896701f),
	.w8(32'hba6db6ce),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d69b6),
	.w1(32'hbad3e24c),
	.w2(32'hbac456d1),
	.w3(32'hba80eb5f),
	.w4(32'hba8c9766),
	.w5(32'hb873e694),
	.w6(32'hba0926aa),
	.w7(32'hbab2c6ff),
	.w8(32'h3a5f88d0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f9f6c),
	.w1(32'h3aab39ac),
	.w2(32'hbb600fd3),
	.w3(32'hbb7719cc),
	.w4(32'hb9d24684),
	.w5(32'hbb1105f8),
	.w6(32'hbb8e11e8),
	.w7(32'h389186dd),
	.w8(32'hbbbb0f21),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacbdd5),
	.w1(32'hbaa4371a),
	.w2(32'hba037b74),
	.w3(32'hb9e7d957),
	.w4(32'h3b14ebd4),
	.w5(32'hbb7ca26e),
	.w6(32'hbb300d1f),
	.w7(32'hb9507785),
	.w8(32'hbbe3f9e4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf4e94),
	.w1(32'hbb49ecad),
	.w2(32'hbb168a80),
	.w3(32'hbb22a3d2),
	.w4(32'hb937aa8f),
	.w5(32'hba9e0416),
	.w6(32'hbb6b0184),
	.w7(32'hbaae85f5),
	.w8(32'h39f23bff),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21cc45),
	.w1(32'hbbfa211d),
	.w2(32'hbc1ca10c),
	.w3(32'hbc4211fe),
	.w4(32'hbbd7c7e5),
	.w5(32'hbc23fedc),
	.w6(32'hbbfc5b39),
	.w7(32'hbbb8c021),
	.w8(32'hbbeb0ab6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58ffd),
	.w1(32'hbb4d4b36),
	.w2(32'hbb84a8e3),
	.w3(32'hbb8731d9),
	.w4(32'hbb713b11),
	.w5(32'hbb19c74e),
	.w6(32'hbb2c81f5),
	.w7(32'hbb5af2fe),
	.w8(32'hbb50810b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb3e8f),
	.w1(32'h38379da4),
	.w2(32'h3939cc0a),
	.w3(32'hbb538cd1),
	.w4(32'hbb25eaa3),
	.w5(32'hbab3457a),
	.w6(32'hbb5bf0f5),
	.w7(32'hbb1b8e76),
	.w8(32'hbb24361c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937182),
	.w1(32'hba0f20a3),
	.w2(32'hbab1db15),
	.w3(32'hbb565f78),
	.w4(32'hbb3b53c1),
	.w5(32'h3b0b91e4),
	.w6(32'hbb52e83a),
	.w7(32'hba0a1ef0),
	.w8(32'h3b0b58bb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a484e73),
	.w1(32'hbab2888f),
	.w2(32'hbad3f737),
	.w3(32'hb9334827),
	.w4(32'hbac99bc6),
	.w5(32'h3a10f493),
	.w6(32'hbb47d3da),
	.w7(32'hbb0fee06),
	.w8(32'h3a95637a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82f9c0),
	.w1(32'hbac99b23),
	.w2(32'hba0b9185),
	.w3(32'hbaa85a46),
	.w4(32'hbac9c67c),
	.w5(32'hbaff7769),
	.w6(32'hba8daae7),
	.w7(32'hba47c156),
	.w8(32'hbb486fe5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e18fe),
	.w1(32'hba8914de),
	.w2(32'hba1667fc),
	.w3(32'hb987392d),
	.w4(32'h3a0db60a),
	.w5(32'hbb9b1734),
	.w6(32'hb9c28cbb),
	.w7(32'hba721632),
	.w8(32'hbbd0178c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc519b7),
	.w1(32'hbb2f4cc1),
	.w2(32'hba7874d7),
	.w3(32'hbb33ceda),
	.w4(32'hbb0076c7),
	.w5(32'h3b004985),
	.w6(32'hbb500b14),
	.w7(32'hbabfe1f1),
	.w8(32'h3b092678),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65b18c),
	.w1(32'h3a92cab7),
	.w2(32'h3aabddef),
	.w3(32'hbb4776a0),
	.w4(32'h3a47cafd),
	.w5(32'hb86e7472),
	.w6(32'hbb53241c),
	.w7(32'h3b1583fb),
	.w8(32'h39ba31b2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29e6f),
	.w1(32'hbb4a834e),
	.w2(32'hbc0cc036),
	.w3(32'hbb68efbf),
	.w4(32'hb9957f9c),
	.w5(32'hbb97ed40),
	.w6(32'hbbb19eb2),
	.w7(32'hba878a42),
	.w8(32'hbbbb5125),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a7f12),
	.w1(32'h3b3ecd9d),
	.w2(32'hbb54aef3),
	.w3(32'hbab8b9f9),
	.w4(32'h3b158df3),
	.w5(32'hbb2d0ce1),
	.w6(32'hbb37eb89),
	.w7(32'h3a6c94f1),
	.w8(32'hbb0c72c2),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc57047),
	.w1(32'h3a4a3d80),
	.w2(32'hbb5a4978),
	.w3(32'hbb80dab0),
	.w4(32'h3a6899f7),
	.w5(32'hbbc1ef35),
	.w6(32'hba9c8559),
	.w7(32'h3a5f3390),
	.w8(32'hbba23bb7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ddcbf),
	.w1(32'h3a8d6f34),
	.w2(32'h3a3259fe),
	.w3(32'hbb05df51),
	.w4(32'h3882a1fc),
	.w5(32'hbad43dae),
	.w6(32'hbb063e67),
	.w7(32'h3987f03b),
	.w8(32'hba72e563),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab35daf),
	.w1(32'hbb820b3b),
	.w2(32'hbabd09e5),
	.w3(32'hba590942),
	.w4(32'hbb2de084),
	.w5(32'h3b8e5c3c),
	.w6(32'hba76d4c9),
	.w7(32'hbb19df75),
	.w8(32'h3ba61d75),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2338fd),
	.w1(32'h3b363fa4),
	.w2(32'h3b41bc1e),
	.w3(32'h3bca962a),
	.w4(32'h3b9621e2),
	.w5(32'hbb58cb98),
	.w6(32'h3bd561ef),
	.w7(32'h3b6d8495),
	.w8(32'hbb8e6c84),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a0261),
	.w1(32'hba908e1f),
	.w2(32'h39ea7c35),
	.w3(32'hbb1f172f),
	.w4(32'h38d08460),
	.w5(32'hba65b7ac),
	.w6(32'hbb988e75),
	.w7(32'hbacbcee0),
	.w8(32'h3a758c0b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc166d01),
	.w1(32'hbb29c93b),
	.w2(32'hbbbd5ca8),
	.w3(32'hbbc3f0c6),
	.w4(32'hb963dc9b),
	.w5(32'hbbde8160),
	.w6(32'hbbd1f4b8),
	.w7(32'h39a91367),
	.w8(32'hbbe7d799),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2e4f),
	.w1(32'hbb8861c0),
	.w2(32'hbb373d29),
	.w3(32'hbb1b8550),
	.w4(32'hb99ff7b1),
	.w5(32'hba84bb3e),
	.w6(32'hbaa6be6c),
	.w7(32'hba916e9a),
	.w8(32'h391be08e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c476e),
	.w1(32'hba905273),
	.w2(32'hbb44fe94),
	.w3(32'hbaa087c0),
	.w4(32'hbb10d6f4),
	.w5(32'hbaa894fc),
	.w6(32'hba2ad416),
	.w7(32'hbaf7016a),
	.w8(32'h380e7d19),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabede24),
	.w1(32'h394b032e),
	.w2(32'h395cfa65),
	.w3(32'hba3df1d8),
	.w4(32'hba0097e0),
	.w5(32'hbb26eabc),
	.w6(32'hb7b652ef),
	.w7(32'h39bb39e2),
	.w8(32'hbb8c74a6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3435ac),
	.w1(32'hbb5b575a),
	.w2(32'hbaad39de),
	.w3(32'hbaab7524),
	.w4(32'hba712461),
	.w5(32'hbb1d1dd5),
	.w6(32'hbbb4ba0a),
	.w7(32'hbb45f042),
	.w8(32'hbab31eaa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87fe14),
	.w1(32'h3a72a2f2),
	.w2(32'h3ac213b7),
	.w3(32'hbb988032),
	.w4(32'hb9f96770),
	.w5(32'h3a5b1af2),
	.w6(32'hbb4be276),
	.w7(32'h3ad54132),
	.w8(32'hbb725350),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29d1bd),
	.w1(32'hbbc17275),
	.w2(32'hbb36c9b4),
	.w3(32'h3a6f0a2c),
	.w4(32'h3ad50162),
	.w5(32'hba335d68),
	.w6(32'hbb95fd4c),
	.w7(32'hba83ec66),
	.w8(32'hbae748c9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61de07),
	.w1(32'hbb5aeea8),
	.w2(32'hbb8aeb55),
	.w3(32'hbb8c29cf),
	.w4(32'h3bb607f6),
	.w5(32'h3881b85b),
	.w6(32'hbba91aaf),
	.w7(32'h3b9805b2),
	.w8(32'hbb04c77f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1f07),
	.w1(32'h3abcba3d),
	.w2(32'h3b71957b),
	.w3(32'hba875107),
	.w4(32'hb9b6a1e2),
	.w5(32'hb9590289),
	.w6(32'h390e1811),
	.w7(32'h3a448729),
	.w8(32'hba95ace6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c9ba),
	.w1(32'h3b1c4a0c),
	.w2(32'h3b174f66),
	.w3(32'hbb5008ee),
	.w4(32'h39e19639),
	.w5(32'hbb6fb830),
	.w6(32'hbb5dfa6b),
	.w7(32'h3ac03487),
	.w8(32'hbb78b900),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule