module layer_8_featuremap_183(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c218600),
	.w1(32'h3ad8c23a),
	.w2(32'hbb88beb0),
	.w3(32'h3b2bbf4e),
	.w4(32'h3bd56df6),
	.w5(32'hbb87b871),
	.w6(32'hba2dc2f8),
	.w7(32'h390f1912),
	.w8(32'h3a917291),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eafa1),
	.w1(32'hbb68a321),
	.w2(32'hbd1a971b),
	.w3(32'h3b874811),
	.w4(32'hbbec4f6c),
	.w5(32'hbd3fd966),
	.w6(32'h3cd4588d),
	.w7(32'h3c921a59),
	.w8(32'h3ce275dd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba5088),
	.w1(32'hbbc004a4),
	.w2(32'h3a82103c),
	.w3(32'hbcee17e2),
	.w4(32'hbb509e72),
	.w5(32'h392d49d4),
	.w6(32'h3b5fd609),
	.w7(32'h3ac4ff34),
	.w8(32'hb915d4fe),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63f78c),
	.w1(32'hbbb39493),
	.w2(32'hbb864988),
	.w3(32'hba8c8b69),
	.w4(32'hbc12ef9a),
	.w5(32'hbc06d42f),
	.w6(32'hba09a504),
	.w7(32'h3b1b5d6c),
	.w8(32'hbb1a7c9b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f0f5f),
	.w1(32'hbca75eb7),
	.w2(32'hbcc22f3a),
	.w3(32'hbba48235),
	.w4(32'h3bf42b3e),
	.w5(32'h3bd6337d),
	.w6(32'hbc63e301),
	.w7(32'hbcbb6fdc),
	.w8(32'hbc1827f1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc604546),
	.w1(32'hba2a6dc6),
	.w2(32'hbc417473),
	.w3(32'h3c035aae),
	.w4(32'h38033a3d),
	.w5(32'hbbab37cd),
	.w6(32'hbb32c5c2),
	.w7(32'hbbcb9af7),
	.w8(32'hbbb971c9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb01720),
	.w1(32'h3bf18810),
	.w2(32'h3d2e0c33),
	.w3(32'h3af3b25f),
	.w4(32'h3cb19b4f),
	.w5(32'h3d6c2628),
	.w6(32'hbceb20c5),
	.w7(32'hbc730a9d),
	.w8(32'hbcc26eb1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc03496),
	.w1(32'hbae72ca5),
	.w2(32'h3a28207f),
	.w3(32'h3d102add),
	.w4(32'hbc28c31d),
	.w5(32'hbc0751bc),
	.w6(32'hbb16baea),
	.w7(32'h3bda69c5),
	.w8(32'hbb24d877),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3280b4),
	.w1(32'hbc12371d),
	.w2(32'h3c4c13a0),
	.w3(32'hbb839f1b),
	.w4(32'h3cddb069),
	.w5(32'h3d548481),
	.w6(32'hbd02a2d5),
	.w7(32'hbcbf22d0),
	.w8(32'hbbd4390c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c869530),
	.w1(32'h3b390256),
	.w2(32'h3b19eb83),
	.w3(32'h3d36b370),
	.w4(32'hbb2fc587),
	.w5(32'h3b830a49),
	.w6(32'h3b95617a),
	.w7(32'hbbb6403e),
	.w8(32'hbb995760),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06be6c),
	.w1(32'hbba809de),
	.w2(32'hbb92bf84),
	.w3(32'h3aeae48f),
	.w4(32'hbaa0518d),
	.w5(32'hbbf07e6f),
	.w6(32'hba3bbb1a),
	.w7(32'hba8719a8),
	.w8(32'hbb9b7a90),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb50c),
	.w1(32'h3b76377d),
	.w2(32'h3b9ad87f),
	.w3(32'hbc09773d),
	.w4(32'h3af1fc86),
	.w5(32'h3b6afda9),
	.w6(32'hba902bcf),
	.w7(32'hba704367),
	.w8(32'h3b53f2a1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abeb3d4),
	.w1(32'hbbbc4e16),
	.w2(32'hbc08bbaf),
	.w3(32'h3b300683),
	.w4(32'h396b2cb3),
	.w5(32'hb86e815c),
	.w6(32'hbb59b093),
	.w7(32'hbb588f36),
	.w8(32'h3910ae57),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cbdd1),
	.w1(32'hbaa1bfaa),
	.w2(32'h3c1601ec),
	.w3(32'h3b5ae340),
	.w4(32'h3a7d9ce9),
	.w5(32'h3b9270fb),
	.w6(32'hbb09b9b4),
	.w7(32'hb9370528),
	.w8(32'hba27efce),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c8bc),
	.w1(32'hbba568f3),
	.w2(32'hbcfe4529),
	.w3(32'hbaadb2af),
	.w4(32'hbd19d67b),
	.w5(32'hbd86a3f6),
	.w6(32'h3ca08c35),
	.w7(32'h3cc70e74),
	.w8(32'h3c59f4bd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb7561),
	.w1(32'h3b721218),
	.w2(32'h3bb231b8),
	.w3(32'hbd5b773c),
	.w4(32'hb9832dc4),
	.w5(32'hbb269766),
	.w6(32'h3b1df2d3),
	.w7(32'hbae3ac64),
	.w8(32'h3b125ea0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4c179),
	.w1(32'hbb46d415),
	.w2(32'hbb44f74a),
	.w3(32'hbb0c93ea),
	.w4(32'hbad1f849),
	.w5(32'hbb2c54d6),
	.w6(32'hbb42ad76),
	.w7(32'h3b271ce9),
	.w8(32'hbb489d75),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a569ee9),
	.w1(32'h3b1e1c07),
	.w2(32'h3ad01938),
	.w3(32'hbb7a087d),
	.w4(32'hb9d40129),
	.w5(32'h39f59716),
	.w6(32'hbb9696bb),
	.w7(32'h3961b310),
	.w8(32'hbad583f8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55dfa9),
	.w1(32'h3c3b18a5),
	.w2(32'h3c76c8ca),
	.w3(32'hb8ba6489),
	.w4(32'hbb9ed53e),
	.w5(32'h3bbc4814),
	.w6(32'hbbe2c8f5),
	.w7(32'h3b5095df),
	.w8(32'h3c106a34),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dc8bb),
	.w1(32'h3bb47882),
	.w2(32'h3d744b93),
	.w3(32'h3a9c3f63),
	.w4(32'h3c507316),
	.w5(32'h3d916021),
	.w6(32'hbd35a1e2),
	.w7(32'hbccfda11),
	.w8(32'hbd1b2bee),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd076d1),
	.w1(32'h3a10d653),
	.w2(32'hbad9db9e),
	.w3(32'h3d12f096),
	.w4(32'hbbf8550b),
	.w5(32'hbbe9bca8),
	.w6(32'hbb5a72b7),
	.w7(32'h3b9b4628),
	.w8(32'h3ab93614),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba921764),
	.w1(32'hbb1cae4b),
	.w2(32'hbb2b4b50),
	.w3(32'h3b220c33),
	.w4(32'h3a908e8b),
	.w5(32'hba2c6a7a),
	.w6(32'h3ba20e44),
	.w7(32'h3b43ab09),
	.w8(32'h3a1e1651),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04b68f),
	.w1(32'h3bb78cf1),
	.w2(32'h3be74486),
	.w3(32'h3b849c21),
	.w4(32'hbb3f1ad6),
	.w5(32'h3c087ebf),
	.w6(32'h3be77c2c),
	.w7(32'h3be57efe),
	.w8(32'hba01ac8d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06527c),
	.w1(32'hb9e309b8),
	.w2(32'hba641b31),
	.w3(32'hba2d2681),
	.w4(32'hbaf2006c),
	.w5(32'h3a97b394),
	.w6(32'hb93f5f7b),
	.w7(32'hbb57ecec),
	.w8(32'hba6c81b1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22881),
	.w1(32'h3b12e50e),
	.w2(32'hbb91c82a),
	.w3(32'h3b2cf09c),
	.w4(32'h3b91b961),
	.w5(32'h3bcbf065),
	.w6(32'hbae04616),
	.w7(32'hbbca5f90),
	.w8(32'h3b68ee0b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8145b2),
	.w1(32'h3c034fd4),
	.w2(32'h3c41cbc7),
	.w3(32'h3c72ee2f),
	.w4(32'h3bc4a9da),
	.w5(32'h3c01ae32),
	.w6(32'h3b31efeb),
	.w7(32'h3ae66f20),
	.w8(32'h3b266ac3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663a84),
	.w1(32'hbc0e7ccb),
	.w2(32'hbc2bc1fd),
	.w3(32'hbafe90d5),
	.w4(32'hbbc8617f),
	.w5(32'hbc14053e),
	.w6(32'h3bcdc945),
	.w7(32'hbb5266c9),
	.w8(32'hbaf8702b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbbfc0),
	.w1(32'hbbf4c75c),
	.w2(32'h3c8a2c90),
	.w3(32'hbcdf51f2),
	.w4(32'hbce81a26),
	.w5(32'hbcb92e9a),
	.w6(32'hbc72bee3),
	.w7(32'h3c2df456),
	.w8(32'h3ccbd20b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab0830),
	.w1(32'hbae9e3dc),
	.w2(32'h3c19930f),
	.w3(32'hbb733a1c),
	.w4(32'hbb94d47d),
	.w5(32'h3b028b2f),
	.w6(32'hbb9f0baf),
	.w7(32'h3c28ff66),
	.w8(32'h37ccc9e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae81235),
	.w1(32'h3c07a451),
	.w2(32'hbb1ad91e),
	.w3(32'hb7603f98),
	.w4(32'h3c91ccf2),
	.w5(32'h3c7482c0),
	.w6(32'h3b9c182a),
	.w7(32'h3c477c14),
	.w8(32'h3bfd93ae),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dff58),
	.w1(32'h3b8171e2),
	.w2(32'hbaecf496),
	.w3(32'h3c630e5f),
	.w4(32'h3a1aa4fd),
	.w5(32'hbaf665b5),
	.w6(32'h3a0072f9),
	.w7(32'hbb31d5de),
	.w8(32'hbbdcae58),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfde2a),
	.w1(32'h3b0d00e1),
	.w2(32'hb9dab255),
	.w3(32'h3b3f0ca1),
	.w4(32'h3bb7f2d2),
	.w5(32'h3aca2d37),
	.w6(32'h3ba329a5),
	.w7(32'h3b64fc28),
	.w8(32'h3b0ba3e3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfb977),
	.w1(32'hb96b550a),
	.w2(32'hb982ca83),
	.w3(32'hb994b9ee),
	.w4(32'h3ad01da1),
	.w5(32'h3b624781),
	.w6(32'h3abf973b),
	.w7(32'h3b75a442),
	.w8(32'hba4b626f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f7308),
	.w1(32'h3b163912),
	.w2(32'h3b49b648),
	.w3(32'h3aaf82ab),
	.w4(32'h3ad6a8cd),
	.w5(32'h3be29852),
	.w6(32'hbaff3b6b),
	.w7(32'hbab8458d),
	.w8(32'h390dca1b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988d350),
	.w1(32'hbb2a03e0),
	.w2(32'h39f9699b),
	.w3(32'h3b7dcd65),
	.w4(32'h3ad8ba8a),
	.w5(32'h3bcfb8b6),
	.w6(32'hbaf5716e),
	.w7(32'h3b3088af),
	.w8(32'h3ab68814),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea8f53),
	.w1(32'hbb61d7d3),
	.w2(32'hba0e9b47),
	.w3(32'h3ab85bb8),
	.w4(32'hba807a15),
	.w5(32'h3af5e7c7),
	.w6(32'hbb5fe86d),
	.w7(32'h39100c1e),
	.w8(32'h39521f53),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4d43f),
	.w1(32'hba919722),
	.w2(32'hb9e92eda),
	.w3(32'hbb876f2a),
	.w4(32'hbac17798),
	.w5(32'h3ada4504),
	.w6(32'h3b53867e),
	.w7(32'h3b7768e5),
	.w8(32'hba74aaba),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5683c6),
	.w1(32'hbc580cbc),
	.w2(32'hbdb662c9),
	.w3(32'h3a1e1014),
	.w4(32'hbd63ff8f),
	.w5(32'hbe0b1326),
	.w6(32'h3d6e441f),
	.w7(32'h3d3b6d4e),
	.w8(32'h3d4bf5b2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd485ae3),
	.w1(32'h3ab83d4e),
	.w2(32'h3a7df16f),
	.w3(32'hbdacdd0a),
	.w4(32'hbb249442),
	.w5(32'hbae5e11f),
	.w6(32'hbb85fb04),
	.w7(32'hbbe3342a),
	.w8(32'hb7eb61d5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1a8b3),
	.w1(32'hbabb7f7f),
	.w2(32'h3b8b362a),
	.w3(32'h3bea4467),
	.w4(32'h3a0ac711),
	.w5(32'h3b732d1c),
	.w6(32'h39ea92be),
	.w7(32'hbbbb6915),
	.w8(32'hb9a8c654),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af90576),
	.w1(32'h3aba94d7),
	.w2(32'h39fe98a5),
	.w3(32'hbbd83a5c),
	.w4(32'hbc5c8ad7),
	.w5(32'hbc11f80b),
	.w6(32'hbb8180eb),
	.w7(32'hbb2446e8),
	.w8(32'hbb446c61),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903a1a),
	.w1(32'h3bb60c30),
	.w2(32'hb9003062),
	.w3(32'hbb82535f),
	.w4(32'h393952ac),
	.w5(32'hba9bd1f2),
	.w6(32'h399113cc),
	.w7(32'hb9605c1d),
	.w8(32'h3b2a1de8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd5f84),
	.w1(32'hbabd6cf6),
	.w2(32'hbbe1422c),
	.w3(32'hbb777f6f),
	.w4(32'hbb4b6e21),
	.w5(32'hbafc4e4d),
	.w6(32'hba890134),
	.w7(32'hbb610c9a),
	.w8(32'h3a1924e6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2e176),
	.w1(32'h3b47bf9a),
	.w2(32'h3b0f4ff2),
	.w3(32'hba9af116),
	.w4(32'hbad7ba6a),
	.w5(32'h3ad96563),
	.w6(32'hbb3b7761),
	.w7(32'hb88bc770),
	.w8(32'hba8130b0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1fa96),
	.w1(32'h3afbdb51),
	.w2(32'h3b953f6b),
	.w3(32'h39f539f7),
	.w4(32'h3b12ff50),
	.w5(32'h3c0d5c9d),
	.w6(32'hbb549a51),
	.w7(32'h3a0f5420),
	.w8(32'h3adfdeb5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09d006),
	.w1(32'h3a83bf88),
	.w2(32'h3ce00000),
	.w3(32'hbb2ded04),
	.w4(32'hbc0b148b),
	.w5(32'h3c72ba6b),
	.w6(32'hbca5f546),
	.w7(32'hbb245e16),
	.w8(32'hbc802f53),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05bab9),
	.w1(32'hbb84ec58),
	.w2(32'hbb3045d0),
	.w3(32'hba810fea),
	.w4(32'hb90fa7ff),
	.w5(32'h3b557bf7),
	.w6(32'hbb8726de),
	.w7(32'hbacc649b),
	.w8(32'hbb8b9888),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4be4c),
	.w1(32'hb9d76121),
	.w2(32'h3ba37fd5),
	.w3(32'h3a84be9b),
	.w4(32'h3b2872f2),
	.w5(32'h3b0ef749),
	.w6(32'hbb9e57d3),
	.w7(32'h3b18623f),
	.w8(32'h3ba55414),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54fdd5),
	.w1(32'hb9900792),
	.w2(32'h38bfe4ca),
	.w3(32'h3bacf3e4),
	.w4(32'h3a8d1d31),
	.w5(32'hbb78ebff),
	.w6(32'hbb74408f),
	.w7(32'h3b997d57),
	.w8(32'hbb2c4d2d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98b80a),
	.w1(32'h3b8f5600),
	.w2(32'hba178792),
	.w3(32'hba98b8b9),
	.w4(32'hbb499e04),
	.w5(32'hbb0fb78d),
	.w6(32'h3b24c7aa),
	.w7(32'hbbd76883),
	.w8(32'hbb967d9f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d604b0),
	.w1(32'hbb94763e),
	.w2(32'hbd15192b),
	.w3(32'hbb58f876),
	.w4(32'hbc80a001),
	.w5(32'hbcf9f4b8),
	.w6(32'h3c8ba578),
	.w7(32'h3c29abc2),
	.w8(32'h3c6e2f30),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc423f18),
	.w1(32'h3bfde480),
	.w2(32'h3c741dea),
	.w3(32'hbcf8ebd5),
	.w4(32'hbc4b8224),
	.w5(32'hbb87808f),
	.w6(32'hbbfff850),
	.w7(32'hbab39883),
	.w8(32'hbbad90e5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15201a),
	.w1(32'hbca72089),
	.w2(32'hbde7ff4a),
	.w3(32'h3b797ffa),
	.w4(32'hbd7790c7),
	.w5(32'hbe271aaa),
	.w6(32'h3d5a22b2),
	.w7(32'h3d0996a0),
	.w8(32'h3d35783e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda18af3),
	.w1(32'h3b50e7ac),
	.w2(32'h3ba5059d),
	.w3(32'hbdea348a),
	.w4(32'hbbc3add6),
	.w5(32'hba947b73),
	.w6(32'hbb9e7cb0),
	.w7(32'hbab11167),
	.w8(32'hbb0e415b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411004),
	.w1(32'hbb08888c),
	.w2(32'hbadfcb80),
	.w3(32'h3af25daa),
	.w4(32'h3b58d7ec),
	.w5(32'h3c116a17),
	.w6(32'h397a3a37),
	.w7(32'hbbe76945),
	.w8(32'h3b2ac250),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047245),
	.w1(32'h3c027440),
	.w2(32'h3c80ae14),
	.w3(32'h3c0524c3),
	.w4(32'h3bbfcb9b),
	.w5(32'h3bb294e1),
	.w6(32'hb9c43bfa),
	.w7(32'h3bd13453),
	.w8(32'h3b822f82),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9071535),
	.w1(32'hbc018317),
	.w2(32'hbb88e269),
	.w3(32'h3b156d95),
	.w4(32'hbbc238b8),
	.w5(32'h39e35636),
	.w6(32'h3a25500a),
	.w7(32'hbb3c7332),
	.w8(32'hbbae7aca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdca667),
	.w1(32'h3aec691b),
	.w2(32'h3bad81af),
	.w3(32'h3ab53481),
	.w4(32'hbb8ea182),
	.w5(32'h3b3161da),
	.w6(32'hbaa093bd),
	.w7(32'h3ae74cae),
	.w8(32'hb850b6e6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5310e3),
	.w1(32'h3bcaab77),
	.w2(32'hbbe47927),
	.w3(32'h3b0325e5),
	.w4(32'hbc22ef48),
	.w5(32'hbcf32487),
	.w6(32'h3ca066ff),
	.w7(32'h3caa5ab5),
	.w8(32'h3c8719b5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf911),
	.w1(32'hbaaec7ab),
	.w2(32'hbb492bcf),
	.w3(32'hbcb9490d),
	.w4(32'hbba16e7b),
	.w5(32'hbbdf9e9d),
	.w6(32'hbbdd32d0),
	.w7(32'hbbea48dc),
	.w8(32'hbb9c6526),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbe6fd),
	.w1(32'hbc420106),
	.w2(32'hbc029651),
	.w3(32'h3bdcdf06),
	.w4(32'hbb56e6c5),
	.w5(32'hbb8ea5bf),
	.w6(32'hbba573ed),
	.w7(32'hbb8b6c53),
	.w8(32'hbb35efc2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9004c6),
	.w1(32'hbc0647c5),
	.w2(32'hbc1033f1),
	.w3(32'hbb0698db),
	.w4(32'hbc820eac),
	.w5(32'hbc90a637),
	.w6(32'h3aa4dd06),
	.w7(32'h3a9bbd37),
	.w8(32'hbb31618d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30e6c3),
	.w1(32'h3bf9745c),
	.w2(32'h3c925db3),
	.w3(32'hbc8af483),
	.w4(32'h3b42cb0e),
	.w5(32'h3b80cd39),
	.w6(32'hbc120c48),
	.w7(32'hbbeb4d34),
	.w8(32'hbc85b454),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba051ff),
	.w1(32'hbb6f2a72),
	.w2(32'h39c5f439),
	.w3(32'hbbb2dbb5),
	.w4(32'hba3e71f0),
	.w5(32'h3b9c90a1),
	.w6(32'hbbeb04a2),
	.w7(32'hbbe181b5),
	.w8(32'hbacb9b4c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a691cda),
	.w1(32'h3c1118a8),
	.w2(32'hbd1f4025),
	.w3(32'h3ba60c9a),
	.w4(32'hbd02d499),
	.w5(32'hbdb22771),
	.w6(32'h3d513c9e),
	.w7(32'h3d45e326),
	.w8(32'h3d3dc2ec),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82148e),
	.w1(32'h3ba66e04),
	.w2(32'h3bdd01c4),
	.w3(32'hbd6145e2),
	.w4(32'hb99b9bad),
	.w5(32'hbabb4084),
	.w6(32'h39b556d3),
	.w7(32'h3bcc4a98),
	.w8(32'h3b025114),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab5d9b),
	.w1(32'h3c45f34c),
	.w2(32'h3bde5fd2),
	.w3(32'hbb817001),
	.w4(32'h3a1f4e5a),
	.w5(32'hbc10945e),
	.w6(32'h3baa816b),
	.w7(32'h3c075148),
	.w8(32'h3bb805d8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb8cc9),
	.w1(32'h3b08670d),
	.w2(32'h3a1f4624),
	.w3(32'h3b05cb36),
	.w4(32'h3b6a2dc9),
	.w5(32'h3be61fc9),
	.w6(32'h3bab506b),
	.w7(32'h3b937846),
	.w8(32'h3be8a9d4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb647409),
	.w1(32'h3b177255),
	.w2(32'h3b578469),
	.w3(32'h3ab6a090),
	.w4(32'hbac3cd89),
	.w5(32'h3b315171),
	.w6(32'hbb43caaa),
	.w7(32'h3b8bdd05),
	.w8(32'hba9e1d0d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb075b2a),
	.w1(32'h3bb1d357),
	.w2(32'h3c4961a1),
	.w3(32'hbbf683e8),
	.w4(32'hbc0239c5),
	.w5(32'h3b693dea),
	.w6(32'hbbe6b6aa),
	.w7(32'hba2024bd),
	.w8(32'h3bea7bd4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f25803),
	.w1(32'h3be78bcd),
	.w2(32'h3b1db55d),
	.w3(32'h3b61fb5c),
	.w4(32'h3c16cdd9),
	.w5(32'hbada8952),
	.w6(32'hbabe5cdf),
	.w7(32'h3aa360ae),
	.w8(32'h3b6d9e3b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b218c2d),
	.w1(32'h3ac7612e),
	.w2(32'h3b7f5633),
	.w3(32'hbb2d3c98),
	.w4(32'h3980e0fe),
	.w5(32'hbbb351b7),
	.w6(32'hb77635a0),
	.w7(32'h3b88cfac),
	.w8(32'hbba12c65),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a90c5),
	.w1(32'h3b9e98dd),
	.w2(32'hba959161),
	.w3(32'hba0ef277),
	.w4(32'h3a7f295e),
	.w5(32'h3b948bc4),
	.w6(32'h3b1a1c20),
	.w7(32'hbb39e099),
	.w8(32'hbabe7008),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba111899),
	.w1(32'h3b743a50),
	.w2(32'h3b653a67),
	.w3(32'hb85e31fa),
	.w4(32'h3b6e8a6b),
	.w5(32'h3954abba),
	.w6(32'hbb088069),
	.w7(32'hbb03ec73),
	.w8(32'hbacce372),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd4e9a),
	.w1(32'hbbca960f),
	.w2(32'hba4c0cf6),
	.w3(32'h398202c1),
	.w4(32'hba1323b5),
	.w5(32'hbb9e6361),
	.w6(32'hbb9cda0f),
	.w7(32'hbbd88c55),
	.w8(32'hbbef1717),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba655c6a),
	.w1(32'h3af5c1c6),
	.w2(32'h3bf5e409),
	.w3(32'h3b157ff7),
	.w4(32'hbbcbf0d6),
	.w5(32'hbb6c5660),
	.w6(32'h3be61b7b),
	.w7(32'hbb28068b),
	.w8(32'hbae461de),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b742dad),
	.w1(32'hbb9f2e7c),
	.w2(32'h3b10c7df),
	.w3(32'h3b974d47),
	.w4(32'h3a97bc5a),
	.w5(32'h3bae0007),
	.w6(32'hbbf56515),
	.w7(32'hbc12fba1),
	.w8(32'hbb692c11),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86ba0e),
	.w1(32'h3a80a893),
	.w2(32'h3be74fae),
	.w3(32'h3bdac794),
	.w4(32'h3a3cc67a),
	.w5(32'h3b9e5410),
	.w6(32'hbb7e570e),
	.w7(32'h38a4201a),
	.w8(32'hbae4ad73),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c070),
	.w1(32'h3c31a64f),
	.w2(32'h3b4f6713),
	.w3(32'h3b5fb63e),
	.w4(32'h3bf7d070),
	.w5(32'h3c3b644e),
	.w6(32'hbb3b75db),
	.w7(32'hbb8d7bdb),
	.w8(32'h3a9a567c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e0fd),
	.w1(32'h3b5f07c4),
	.w2(32'h3b52cb96),
	.w3(32'h3c2d24eb),
	.w4(32'h3b3fcf6f),
	.w5(32'hbb09898e),
	.w6(32'h3bc09ad0),
	.w7(32'h3a92adf4),
	.w8(32'hbba5a46b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e0f9),
	.w1(32'hbbbe15b6),
	.w2(32'hbb852ebb),
	.w3(32'hbb9c0dd2),
	.w4(32'h3b2786fe),
	.w5(32'h3b44fbb6),
	.w6(32'hbb06c747),
	.w7(32'h3ab5a25a),
	.w8(32'hbb1e011e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b563c4),
	.w1(32'h3ba8e741),
	.w2(32'h3ba71952),
	.w3(32'h3b3c5a38),
	.w4(32'hbb888708),
	.w5(32'h3abbfbc2),
	.w6(32'hbb3680b0),
	.w7(32'hbb3a3398),
	.w8(32'h3aba4ece),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bfaf9),
	.w1(32'h3ad7695e),
	.w2(32'h3ad1964c),
	.w3(32'hbb6a8408),
	.w4(32'h3ba52b31),
	.w5(32'hbb992657),
	.w6(32'hbb77559c),
	.w7(32'h3a9e106b),
	.w8(32'hb96eddf0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64d3e4),
	.w1(32'hbab41632),
	.w2(32'hbb7cea7b),
	.w3(32'hbc89d5d6),
	.w4(32'hbc851832),
	.w5(32'hbc6ad0d1),
	.w6(32'hbc254be6),
	.w7(32'hbc494b36),
	.w8(32'hbc69dbae),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a6b24),
	.w1(32'h3bed133a),
	.w2(32'h3bdb3843),
	.w3(32'hbba8cabd),
	.w4(32'hbb23b2e5),
	.w5(32'h3b20915f),
	.w6(32'hbbcf66f1),
	.w7(32'hbba89e98),
	.w8(32'h3b7624bd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8f512),
	.w1(32'h3b062819),
	.w2(32'hbb0bb22d),
	.w3(32'hb9ded21e),
	.w4(32'hbc203b37),
	.w5(32'hbc254c71),
	.w6(32'h3b8b2518),
	.w7(32'hbacebf79),
	.w8(32'hb995d85f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61276c),
	.w1(32'h3c2d1991),
	.w2(32'h3c294601),
	.w3(32'hbaa81a93),
	.w4(32'h3c421ec9),
	.w5(32'h3c59b56e),
	.w6(32'h3bced523),
	.w7(32'h3bd3f549),
	.w8(32'h3b217e09),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3ea4),
	.w1(32'h3a4ef755),
	.w2(32'h3bfe7715),
	.w3(32'h3c299020),
	.w4(32'h39846298),
	.w5(32'hbb6d76ee),
	.w6(32'h3ba1b3e9),
	.w7(32'h3c3c91f7),
	.w8(32'h3c0ab7cb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd48bb),
	.w1(32'h3bb781ea),
	.w2(32'h3b66cf7a),
	.w3(32'h3b4ea1e8),
	.w4(32'h3c088387),
	.w5(32'h3c4a07bf),
	.w6(32'h3b66482c),
	.w7(32'hb889341c),
	.w8(32'hbb13e42c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938060d),
	.w1(32'hbaab65d7),
	.w2(32'h3ac4174f),
	.w3(32'h3c4ec3df),
	.w4(32'h3b20912d),
	.w5(32'hbac30b58),
	.w6(32'h3addac44),
	.w7(32'hbb2934c8),
	.w8(32'hb9e440b7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05099c),
	.w1(32'hbb3ee9f9),
	.w2(32'hbaeba132),
	.w3(32'h3b7f0454),
	.w4(32'h3a8a2e33),
	.w5(32'hbb3d8a38),
	.w6(32'hba888284),
	.w7(32'h3a1976a4),
	.w8(32'hba81b6e9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f57f3),
	.w1(32'hbb185ab7),
	.w2(32'h3b093e3d),
	.w3(32'hbb4efd4f),
	.w4(32'h3bba390f),
	.w5(32'h3bb60a3d),
	.w6(32'hbb32800d),
	.w7(32'hba85db74),
	.w8(32'h3b038089),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e31c),
	.w1(32'h3bc4868a),
	.w2(32'h3cb5fff4),
	.w3(32'h3a2c344b),
	.w4(32'h3c7edd43),
	.w5(32'h3d2546f0),
	.w6(32'hbc83135d),
	.w7(32'hbc4e89db),
	.w8(32'hbc5432d1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e9d20),
	.w1(32'hba9e7c44),
	.w2(32'hba09c0f0),
	.w3(32'h3ce83c45),
	.w4(32'h3a056fd5),
	.w5(32'h3b0be7d5),
	.w6(32'h3a937a0a),
	.w7(32'h3b74e4a9),
	.w8(32'h3bf3bafe),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a881681),
	.w1(32'hba9b007e),
	.w2(32'hbaae5896),
	.w3(32'h3c09f098),
	.w4(32'h3bd5fecd),
	.w5(32'h3a8f9125),
	.w6(32'h3a5622dd),
	.w7(32'hbad0c74d),
	.w8(32'hbb1efc62),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f902),
	.w1(32'h3bf7f9e5),
	.w2(32'h3c62c059),
	.w3(32'h3b4ee7f2),
	.w4(32'h3b73066a),
	.w5(32'h3c2e1f5c),
	.w6(32'h3b36dbdc),
	.w7(32'h3bf146e5),
	.w8(32'h3aebee1e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33b091),
	.w1(32'h3bfb85a9),
	.w2(32'h3c2cf6f5),
	.w3(32'h3ba624ff),
	.w4(32'h3a39f110),
	.w5(32'h3b973378),
	.w6(32'h3abf7aea),
	.w7(32'h3bb0d181),
	.w8(32'h3bb528cc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b53e6),
	.w1(32'h39db2366),
	.w2(32'hba71b878),
	.w3(32'h3bd00cb7),
	.w4(32'h3b205448),
	.w5(32'hbac678e7),
	.w6(32'hbb38a239),
	.w7(32'hbb203408),
	.w8(32'hbb343d02),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb27a3),
	.w1(32'hbb51104a),
	.w2(32'hbb3676f7),
	.w3(32'h3ba20bb7),
	.w4(32'hba9ef763),
	.w5(32'hba3da8ea),
	.w6(32'hbac40546),
	.w7(32'hba36199b),
	.w8(32'hbb9cd7a9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce14c),
	.w1(32'h3b1961cd),
	.w2(32'hbb29aa0d),
	.w3(32'hbbdc0014),
	.w4(32'h3bad25fd),
	.w5(32'h3bdbfe8c),
	.w6(32'hbb09ced4),
	.w7(32'h3b6e3289),
	.w8(32'h3ac24503),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe157),
	.w1(32'hbb2857d2),
	.w2(32'h3aca7a9f),
	.w3(32'hbb946f66),
	.w4(32'h3b3f4efc),
	.w5(32'h3ae73725),
	.w6(32'hbb5aa582),
	.w7(32'h3b10e226),
	.w8(32'hbb3bab5e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3eeb1),
	.w1(32'hbb9369cd),
	.w2(32'h3b80e8ff),
	.w3(32'hbb4dfc6c),
	.w4(32'hba8f4fb1),
	.w5(32'h3bd86e08),
	.w6(32'hbc1c7a24),
	.w7(32'hbb13bc5c),
	.w8(32'h3aaa9a1c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacba7f8),
	.w1(32'h3b10ed31),
	.w2(32'hbb8216c9),
	.w3(32'h3a531c1a),
	.w4(32'h3aaa93b9),
	.w5(32'h3ad0d1b1),
	.w6(32'h3ae5b02e),
	.w7(32'hbb0b0051),
	.w8(32'h3b03a85b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec9176),
	.w1(32'h3b25c54a),
	.w2(32'hbae0b7f3),
	.w3(32'hbb52beab),
	.w4(32'h3a661652),
	.w5(32'hba2538e7),
	.w6(32'hbb1b2920),
	.w7(32'hbc0541df),
	.w8(32'h3aac7501),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b136974),
	.w1(32'hbaa5008a),
	.w2(32'hba1b3fa1),
	.w3(32'hbb556ad5),
	.w4(32'hba82a76c),
	.w5(32'hbc09f717),
	.w6(32'hbb04b21e),
	.w7(32'hbb822951),
	.w8(32'hbaed00f8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ce081),
	.w1(32'h3cd09d99),
	.w2(32'h3c1d53b6),
	.w3(32'hbc0f4e42),
	.w4(32'hbcd5d59e),
	.w5(32'hbd773754),
	.w6(32'h3d29685c),
	.w7(32'h3d731e53),
	.w8(32'h3d34f850),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f154fd),
	.w1(32'h3b994b7d),
	.w2(32'h3b9c385d),
	.w3(32'hbd459cf0),
	.w4(32'h3bc82a2b),
	.w5(32'h3c29cf22),
	.w6(32'h3b1d3d3e),
	.w7(32'hbac429e8),
	.w8(32'hbb78202a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affa374),
	.w1(32'h3af6fb2c),
	.w2(32'hbaa31590),
	.w3(32'h3c0a2a9f),
	.w4(32'h3b297454),
	.w5(32'h3bafae85),
	.w6(32'hb935d352),
	.w7(32'hbb654e84),
	.w8(32'hb9e6669b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3037),
	.w1(32'h3a4f46d9),
	.w2(32'h3a8eddfc),
	.w3(32'h3c101ac0),
	.w4(32'hbb69f05b),
	.w5(32'hba4226ae),
	.w6(32'h3b44bed3),
	.w7(32'h3a725b5b),
	.w8(32'h3b9ef41d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b554e90),
	.w1(32'hbb93eccd),
	.w2(32'hbd26a0dd),
	.w3(32'h3b7154bb),
	.w4(32'hbc775c10),
	.w5(32'hbd644066),
	.w6(32'h3cd57417),
	.w7(32'h3c9591a2),
	.w8(32'h3cd13832),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdd906),
	.w1(32'h3b83fb03),
	.w2(32'h3b9198e3),
	.w3(32'hbd0b3925),
	.w4(32'h3b2be1e9),
	.w5(32'h3c0d256a),
	.w6(32'hba18f272),
	.w7(32'h3baa5a3c),
	.w8(32'hb9160ad8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba56dd1),
	.w1(32'h3c33af94),
	.w2(32'h3d00ad9b),
	.w3(32'hbb0e9d88),
	.w4(32'h3c88b70c),
	.w5(32'h3d260d4f),
	.w6(32'hbba19091),
	.w7(32'hbab942c6),
	.w8(32'hbbb7f555),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1977b),
	.w1(32'h3ac6445c),
	.w2(32'hbc1c8ce2),
	.w3(32'h3cf5f947),
	.w4(32'h39f9c219),
	.w5(32'hbae7b617),
	.w6(32'h3c083625),
	.w7(32'h3b3f5a53),
	.w8(32'h3b8d60ab),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab34dc2),
	.w1(32'h3b4126c7),
	.w2(32'hbb767591),
	.w3(32'h3a2b3c24),
	.w4(32'hba36ce1b),
	.w5(32'hbba0d59c),
	.w6(32'h3be798af),
	.w7(32'h3b6b8581),
	.w8(32'h3bf12ad9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c3e2),
	.w1(32'hb70cee6f),
	.w2(32'hbb369821),
	.w3(32'hbaf41ec9),
	.w4(32'h3b58dac2),
	.w5(32'h3b1bf3ce),
	.w6(32'h3af36e6f),
	.w7(32'hbb087e9c),
	.w8(32'h3ab1db1c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb668398),
	.w1(32'hbc79adc3),
	.w2(32'hbd81d515),
	.w3(32'h3badd66a),
	.w4(32'hbd170255),
	.w5(32'hbdbd4f10),
	.w6(32'h3cf0d0bd),
	.w7(32'h3ca5b3e1),
	.w8(32'h3cc79625),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e9acb),
	.w1(32'h3af126e6),
	.w2(32'hb9cd8f3c),
	.w3(32'hbd80c090),
	.w4(32'h3c235d5c),
	.w5(32'h3c1f41f7),
	.w6(32'hb9baf5b1),
	.w7(32'hba8ac0f8),
	.w8(32'hb9ddbaf4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3418),
	.w1(32'h3ba42c97),
	.w2(32'h3c0c27d1),
	.w3(32'h3b9d1514),
	.w4(32'hbbb50d74),
	.w5(32'hbb29cdc9),
	.w6(32'h3b353581),
	.w7(32'h3b32a98c),
	.w8(32'h3b59d5c9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f7ad9),
	.w1(32'hbb9f16b2),
	.w2(32'hbbc5ff87),
	.w3(32'hbb591809),
	.w4(32'hba0f674d),
	.w5(32'h39a54926),
	.w6(32'h3b822ace),
	.w7(32'h3b2bdc9a),
	.w8(32'h3bdea53d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26dbd3),
	.w1(32'h3a0072c2),
	.w2(32'hbb1a79cb),
	.w3(32'hbb61226a),
	.w4(32'h3ba33c97),
	.w5(32'h3ac5a161),
	.w6(32'hb9e88df1),
	.w7(32'hbba48373),
	.w8(32'hbb9fb007),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57fe48),
	.w1(32'h3b81c7cf),
	.w2(32'h3b132fbc),
	.w3(32'hbb299d95),
	.w4(32'hbb9a5d73),
	.w5(32'hbba12488),
	.w6(32'h3b6b6ef6),
	.w7(32'hbb0c4d8e),
	.w8(32'h392479ef),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6e933),
	.w1(32'h3b2f36b9),
	.w2(32'h3a74661e),
	.w3(32'hbb95504c),
	.w4(32'h3b75d91c),
	.w5(32'h3b1960e4),
	.w6(32'hba8cf72f),
	.w7(32'h39af84f5),
	.w8(32'hbb3802a3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ab9ba),
	.w1(32'h3b2f8e14),
	.w2(32'h3c8479f2),
	.w3(32'hbaeb503a),
	.w4(32'h3c890daf),
	.w5(32'h3cf63e13),
	.w6(32'hbc03df06),
	.w7(32'hbbafc813),
	.w8(32'hba111157),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a56e3),
	.w1(32'h3b38fe8a),
	.w2(32'hba0711c9),
	.w3(32'h3cd57c6c),
	.w4(32'hbac70938),
	.w5(32'hba90e756),
	.w6(32'h3a6a75f2),
	.w7(32'h3aa53389),
	.w8(32'h3baced0d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491149),
	.w1(32'hbb92fa1d),
	.w2(32'hbaae40b3),
	.w3(32'hbb8af387),
	.w4(32'hbaafe168),
	.w5(32'h3bcaf781),
	.w6(32'h3b1832e1),
	.w7(32'h3a94fe11),
	.w8(32'h3ae643f3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7fdd7),
	.w1(32'hb9d3e272),
	.w2(32'h3b092e19),
	.w3(32'hba84cd7a),
	.w4(32'hbb1e12a2),
	.w5(32'hb9f36b36),
	.w6(32'hbb6fb638),
	.w7(32'h3a851851),
	.w8(32'hbae92b39),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c13e),
	.w1(32'hba43f543),
	.w2(32'h3a2ac2dd),
	.w3(32'hbae06f0e),
	.w4(32'hba4dbe7d),
	.w5(32'h3abf438f),
	.w6(32'hba896326),
	.w7(32'h3a7e12f5),
	.w8(32'hb8e803db),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb8664),
	.w1(32'h3ad1b523),
	.w2(32'h3c153216),
	.w3(32'hbb19a7cd),
	.w4(32'hbbbf95bf),
	.w5(32'h3b36f8b5),
	.w6(32'hba7e6d05),
	.w7(32'h3b0dc80f),
	.w8(32'h3bf33fc0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule