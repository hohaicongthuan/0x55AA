module layer_8_featuremap_159(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1296dd),
	.w1(32'h3a084cae),
	.w2(32'h3c0a1622),
	.w3(32'hbaa1df0d),
	.w4(32'h3b4d9e93),
	.w5(32'h3b0d08fe),
	.w6(32'hb9d3e2f5),
	.w7(32'h3b98019f),
	.w8(32'h3b8ea4e5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc2ca0),
	.w1(32'hbb1faacc),
	.w2(32'hbb8b6fe4),
	.w3(32'h3a3d11e1),
	.w4(32'hb9de2d55),
	.w5(32'hbaf6162e),
	.w6(32'hbad86167),
	.w7(32'hbb274f9d),
	.w8(32'hb983e1fb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1713),
	.w1(32'hba7e8a96),
	.w2(32'h3b0ca71f),
	.w3(32'hba4208c3),
	.w4(32'hba8739d6),
	.w5(32'h3a114402),
	.w6(32'h3af576ae),
	.w7(32'hba109afa),
	.w8(32'h3b203c1d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae95f3),
	.w1(32'hb9885c4d),
	.w2(32'hbb2e3e25),
	.w3(32'h3b03c31e),
	.w4(32'h3a606b48),
	.w5(32'h3b8e9d93),
	.w6(32'h3b1570e5),
	.w7(32'h3b20474f),
	.w8(32'h3bc69734),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dafee),
	.w1(32'hbba4c306),
	.w2(32'hbc0111c6),
	.w3(32'h3b15d998),
	.w4(32'hbb40f1a4),
	.w5(32'hbbbb67f1),
	.w6(32'hbb8ea3cd),
	.w7(32'hbb8b6a0f),
	.w8(32'hbb7a5016),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17c07a),
	.w1(32'hbad4c5a5),
	.w2(32'h38edfb5e),
	.w3(32'hbbd92117),
	.w4(32'hbb810eeb),
	.w5(32'h3b33758e),
	.w6(32'h3a9f877b),
	.w7(32'hba384e2b),
	.w8(32'hbb45fb31),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33d000),
	.w1(32'h3b4f9941),
	.w2(32'h3b4a3269),
	.w3(32'hba601e80),
	.w4(32'h3a54fd24),
	.w5(32'h3b02e640),
	.w6(32'h3b016c80),
	.w7(32'h3b62047d),
	.w8(32'h3a9b07b8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56454b),
	.w1(32'h3c00dcf5),
	.w2(32'h3bfa0e63),
	.w3(32'h3b0cf4b4),
	.w4(32'h3bd7a112),
	.w5(32'hba6c6712),
	.w6(32'h3bb89b80),
	.w7(32'h3b4f86ab),
	.w8(32'h3b2665cf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9540b80),
	.w1(32'h3b89b99c),
	.w2(32'hb6cbb375),
	.w3(32'hbb001ee2),
	.w4(32'h3bc8ebc0),
	.w5(32'h3b8653b9),
	.w6(32'h3badba67),
	.w7(32'h3b711ecb),
	.w8(32'h3b608c84),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996a9a),
	.w1(32'h3a2af26c),
	.w2(32'hb9fd549f),
	.w3(32'h3b0b2dc3),
	.w4(32'h3b2a3474),
	.w5(32'h3abd1792),
	.w6(32'h3b0a899c),
	.w7(32'h3b9b2544),
	.w8(32'h3ae3cdde),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c3c5e),
	.w1(32'h3b5654ba),
	.w2(32'hba07fffd),
	.w3(32'hbb349746),
	.w4(32'h3b087fc6),
	.w5(32'h3aa6a6a3),
	.w6(32'hbb754cce),
	.w7(32'hbab23be5),
	.w8(32'h39a5ca87),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2f6ac),
	.w1(32'h3b1ceec8),
	.w2(32'h3b336f55),
	.w3(32'h3b428dc8),
	.w4(32'h3af5d958),
	.w5(32'h3ae62b7d),
	.w6(32'h3a90e330),
	.w7(32'h3b327ec7),
	.w8(32'h3af00a7b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a361c3b),
	.w1(32'hba4f7f60),
	.w2(32'h3aa94ba6),
	.w3(32'h3b32bb2a),
	.w4(32'h3a81b6b4),
	.w5(32'h3b01fc07),
	.w6(32'hbb217710),
	.w7(32'hbb291962),
	.w8(32'hbb5aff58),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a44a),
	.w1(32'hbac67f6c),
	.w2(32'h3b7121cc),
	.w3(32'hba123f59),
	.w4(32'h39826cea),
	.w5(32'hb8ce8a85),
	.w6(32'h3ab853df),
	.w7(32'h3aa27682),
	.w8(32'h3b26e2b9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f32d),
	.w1(32'h3c00f4d0),
	.w2(32'h3c31a3b8),
	.w3(32'hb908c40b),
	.w4(32'h3bbdcc19),
	.w5(32'h3c196bdf),
	.w6(32'h3bd8503c),
	.w7(32'h3c10acd2),
	.w8(32'h3bc0777f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d82c4),
	.w1(32'h3abcb2a1),
	.w2(32'h3b712f97),
	.w3(32'h3be087ad),
	.w4(32'hbb1d8ae0),
	.w5(32'h3b049119),
	.w6(32'h3abb5b90),
	.w7(32'h3a337eed),
	.w8(32'hba99bdb6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78b7ef),
	.w1(32'h3b203de8),
	.w2(32'h3b333154),
	.w3(32'hbb1fb13d),
	.w4(32'h3b216a73),
	.w5(32'h3b76e856),
	.w6(32'hb95c55aa),
	.w7(32'h3a86474d),
	.w8(32'h3be8f3c7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3421f),
	.w1(32'h3926e306),
	.w2(32'h3aaaaf8f),
	.w3(32'h3b8e3344),
	.w4(32'h3b7a2fc6),
	.w5(32'h3b117360),
	.w6(32'h3a869a93),
	.w7(32'hbad949d1),
	.w8(32'h3b963a98),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1765e6),
	.w1(32'h3afa040b),
	.w2(32'hbafcbaed),
	.w3(32'h3b28bd15),
	.w4(32'h3b378881),
	.w5(32'h3b9853c6),
	.w6(32'h39ad6ee8),
	.w7(32'h3aeb870d),
	.w8(32'h39f22dbb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd6a4a),
	.w1(32'h3b32abc8),
	.w2(32'h3c09920d),
	.w3(32'hbb3b76ec),
	.w4(32'h3a6074ee),
	.w5(32'h3bb2ae4a),
	.w6(32'h39cd87ee),
	.w7(32'h3b3998e9),
	.w8(32'h39afbb3a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b100a9f),
	.w1(32'hbc003fe0),
	.w2(32'hbc319348),
	.w3(32'hba35b5d5),
	.w4(32'hbba6bf5b),
	.w5(32'hbb881b57),
	.w6(32'hbb6132c8),
	.w7(32'hbb765caf),
	.w8(32'hba2edda3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7e9d),
	.w1(32'h3b2696a0),
	.w2(32'h3b56fb6b),
	.w3(32'h3b083fa3),
	.w4(32'hb9023a34),
	.w5(32'h39c1bebb),
	.w6(32'hbac63dcc),
	.w7(32'h3aa4e0e4),
	.w8(32'hbb053033),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf6493),
	.w1(32'h3acf81d0),
	.w2(32'hb9b70e6b),
	.w3(32'h3ad39f43),
	.w4(32'hb968dbf7),
	.w5(32'h39ecc0ab),
	.w6(32'hbb210c3c),
	.w7(32'h3ac7dcff),
	.w8(32'h3aa0d9f9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb083722),
	.w1(32'h3ad7efd2),
	.w2(32'h3af454a7),
	.w3(32'hba8b402d),
	.w4(32'h3a6d3f17),
	.w5(32'hb88464a8),
	.w6(32'h3b865d7a),
	.w7(32'h3ad143d9),
	.w8(32'hba50b0bc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ff971),
	.w1(32'h39be686b),
	.w2(32'h3b149723),
	.w3(32'h3ab47540),
	.w4(32'hba101fd2),
	.w5(32'h3b30d78e),
	.w6(32'h3bc0f1c7),
	.w7(32'h3b1fc715),
	.w8(32'h3b688236),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0e17),
	.w1(32'hbacba1d3),
	.w2(32'h38825a26),
	.w3(32'h3b187d96),
	.w4(32'hbb0526d0),
	.w5(32'hbb8a71d1),
	.w6(32'hbbe2eb4b),
	.w7(32'hbaa1e4c2),
	.w8(32'hbb8968d2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902dfc8),
	.w1(32'h3ac09d74),
	.w2(32'h3b411164),
	.w3(32'hbafa1c4a),
	.w4(32'hba1ad6a1),
	.w5(32'h3baaf3ad),
	.w6(32'h3a135616),
	.w7(32'h3b20815f),
	.w8(32'h3b307e5f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b136318),
	.w1(32'hbba9de5d),
	.w2(32'hbc3442ca),
	.w3(32'h3b31972c),
	.w4(32'h3bf9fb12),
	.w5(32'h3c608677),
	.w6(32'hbc2f9a98),
	.w7(32'h3b92b0de),
	.w8(32'h3bd6050d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc09f7),
	.w1(32'hbbf9dd48),
	.w2(32'h3b17c301),
	.w3(32'h3afdce53),
	.w4(32'hbb3667d2),
	.w5(32'h3bbb8720),
	.w6(32'hbc2e4c34),
	.w7(32'hba7f5d46),
	.w8(32'h3c07be93),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45c3e6),
	.w1(32'h3acaa323),
	.w2(32'h3b2cbb51),
	.w3(32'h3c6d9824),
	.w4(32'h3bc03ff6),
	.w5(32'h3be87d75),
	.w6(32'h3ab83b80),
	.w7(32'h3b05f444),
	.w8(32'h3b17bc6a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a889d23),
	.w1(32'h3b182503),
	.w2(32'h3b79d305),
	.w3(32'h3bcf89bd),
	.w4(32'h3c12a400),
	.w5(32'h3c15a649),
	.w6(32'hbaabe43f),
	.w7(32'hb91e84d8),
	.w8(32'hba36e684),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaa633),
	.w1(32'hbabde95c),
	.w2(32'hbb335fa2),
	.w3(32'h3c0d7810),
	.w4(32'hba1d3181),
	.w5(32'hbb9578a1),
	.w6(32'hbaefa099),
	.w7(32'hbb486061),
	.w8(32'hbb003052),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b09f8),
	.w1(32'hbb01495e),
	.w2(32'h3b4be9cc),
	.w3(32'hbb4a9c7d),
	.w4(32'hba61c4b5),
	.w5(32'h3b3085e5),
	.w6(32'hbb498049),
	.w7(32'h3a483a9a),
	.w8(32'h3a2be82a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a012185),
	.w1(32'hbaff2a7b),
	.w2(32'hbb6eb7ba),
	.w3(32'hbabb251a),
	.w4(32'hba41617e),
	.w5(32'hba23704d),
	.w6(32'h3a14a0dc),
	.w7(32'hbb95e09b),
	.w8(32'hbb604e67),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22349e),
	.w1(32'h3a9974fd),
	.w2(32'h3935b343),
	.w3(32'hbb4408dc),
	.w4(32'h3a1c6a17),
	.w5(32'hbace08ed),
	.w6(32'h3a6aa402),
	.w7(32'hba997ee7),
	.w8(32'hba2ac038),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa975a6),
	.w1(32'h3a45c633),
	.w2(32'h3b8d07c7),
	.w3(32'hba23f34d),
	.w4(32'hbaa1042d),
	.w5(32'h3a292ab0),
	.w6(32'hb9f1767e),
	.w7(32'h3b57598c),
	.w8(32'h3b08162a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ecf81),
	.w1(32'hbb2cbbbf),
	.w2(32'hbb26435d),
	.w3(32'h3abbef1d),
	.w4(32'hbaf7b7f4),
	.w5(32'hbb318597),
	.w6(32'hb87f9e28),
	.w7(32'h39e83808),
	.w8(32'h3ac6b0bb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d7386),
	.w1(32'h3adecb99),
	.w2(32'h3b1f9401),
	.w3(32'hba8841be),
	.w4(32'h3b21f5c8),
	.w5(32'h3b8178c7),
	.w6(32'h3b103bf1),
	.w7(32'h3b401003),
	.w8(32'h3b2299d8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7f898),
	.w1(32'h3a75c031),
	.w2(32'h394f4b26),
	.w3(32'h3b0945d1),
	.w4(32'hb9d53d09),
	.w5(32'hb98a660f),
	.w6(32'h3a8b12e4),
	.w7(32'hbb0b4712),
	.w8(32'hb85a5413),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0841df),
	.w1(32'hbb389c6e),
	.w2(32'hbaffba3d),
	.w3(32'h3aa68f63),
	.w4(32'h3b247859),
	.w5(32'hbb5cf1a1),
	.w6(32'hba8d9742),
	.w7(32'hbb523eb1),
	.w8(32'hbaab8d7e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafee42e),
	.w1(32'hba68cebd),
	.w2(32'hbb902c5c),
	.w3(32'h3a3eb025),
	.w4(32'hbaeb2622),
	.w5(32'hbb8bf358),
	.w6(32'hbb767dc0),
	.w7(32'hbb113a54),
	.w8(32'hbb64a207),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bc889),
	.w1(32'h3bfbfe09),
	.w2(32'hba89052d),
	.w3(32'hbb1f37a2),
	.w4(32'h3be98e7f),
	.w5(32'h3a2eea65),
	.w6(32'h3c3204f3),
	.w7(32'hba131535),
	.w8(32'hbbf2abed),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db643),
	.w1(32'hbb214331),
	.w2(32'h3a61a409),
	.w3(32'hbbe55598),
	.w4(32'hbaa9d6a3),
	.w5(32'h3adb4cce),
	.w6(32'hbb270e00),
	.w7(32'h3b30feb0),
	.w8(32'h3bbd6308),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2938c6),
	.w1(32'h3ab54131),
	.w2(32'h3a802736),
	.w3(32'h3b181d51),
	.w4(32'h3af13c6a),
	.w5(32'h3b0ce8be),
	.w6(32'hb9c6fcc1),
	.w7(32'h3b02fa1c),
	.w8(32'h3b5f9ce2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c3e8f),
	.w1(32'h3a1d34a7),
	.w2(32'h3b40ef3a),
	.w3(32'h3b30804b),
	.w4(32'h3a0c21b0),
	.w5(32'h3b213715),
	.w6(32'hbaedc219),
	.w7(32'hbb06c10b),
	.w8(32'hbb521fc0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab367d8),
	.w1(32'h3b9ee9cf),
	.w2(32'h3be67efb),
	.w3(32'hb9d6a93f),
	.w4(32'h3b3f498f),
	.w5(32'h3bd0346a),
	.w6(32'h3b9a2e69),
	.w7(32'h3bb1f898),
	.w8(32'h3b28f893),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f774d),
	.w1(32'h3bc784e7),
	.w2(32'h3c0b56bd),
	.w3(32'h3ac150dc),
	.w4(32'h3bcfe7cb),
	.w5(32'h3bd84f4d),
	.w6(32'h3b9fffad),
	.w7(32'h3bda3db1),
	.w8(32'h3b8d3b7d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba05e3f),
	.w1(32'h3b0b3b4b),
	.w2(32'h3b29413e),
	.w3(32'h3b54755e),
	.w4(32'h3b36f129),
	.w5(32'h3aee8323),
	.w6(32'h39bee6ea),
	.w7(32'h3aa42671),
	.w8(32'h3b448776),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857d5c),
	.w1(32'h3bae23ba),
	.w2(32'h3b44fcf6),
	.w3(32'hb8fc45f7),
	.w4(32'hba9888dd),
	.w5(32'h374aa87c),
	.w6(32'hbad74f04),
	.w7(32'h3ac299db),
	.w8(32'h3b0a9a8f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5a56e),
	.w1(32'hb6120d07),
	.w2(32'h3b982a15),
	.w3(32'h3a898bcc),
	.w4(32'h3bb92fa2),
	.w5(32'h3b8ea1c7),
	.w6(32'h3a131fd0),
	.w7(32'h3b347e11),
	.w8(32'hb9c5c702),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8fd41),
	.w1(32'hba19c85a),
	.w2(32'hbb17e5f9),
	.w3(32'h3ae6aaf5),
	.w4(32'h3a3ec29f),
	.w5(32'hbada34fd),
	.w6(32'h3898df3b),
	.w7(32'hba85bd7e),
	.w8(32'h3a0d633a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f9621),
	.w1(32'hba07503b),
	.w2(32'hbb67eab5),
	.w3(32'h3a0cf89c),
	.w4(32'h3b621691),
	.w5(32'h3a605efd),
	.w6(32'h3b6b7822),
	.w7(32'h39d17c7e),
	.w8(32'h3a727c24),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3da30),
	.w1(32'hbb2be612),
	.w2(32'hbb6642e8),
	.w3(32'h3a244b1a),
	.w4(32'h3a706bc4),
	.w5(32'hba1a109a),
	.w6(32'hba921149),
	.w7(32'hbadbbd01),
	.w8(32'h39fd4051),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dd473),
	.w1(32'h3b23913a),
	.w2(32'h3b23c759),
	.w3(32'h3a133d0f),
	.w4(32'h3b146c24),
	.w5(32'hbb48cab9),
	.w6(32'h3a76ebd7),
	.w7(32'h3a44fe18),
	.w8(32'h3a92f86a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f80e95),
	.w1(32'hbac90034),
	.w2(32'h3b524baf),
	.w3(32'h39af8f18),
	.w4(32'h3b4f5372),
	.w5(32'h3ba9bb28),
	.w6(32'h39cbe1c5),
	.w7(32'h3ba70609),
	.w8(32'h3af5fddf),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae60455),
	.w1(32'hbb21374b),
	.w2(32'h3b10ed60),
	.w3(32'h3b08630f),
	.w4(32'h3b855d68),
	.w5(32'h3b9990d4),
	.w6(32'hba3d0f8d),
	.w7(32'h38d2e0db),
	.w8(32'h3b3ef680),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b508aaf),
	.w1(32'h3ac7543f),
	.w2(32'hbabd6480),
	.w3(32'h39a95c29),
	.w4(32'hbaa9f8aa),
	.w5(32'h3b25c028),
	.w6(32'hba5a497a),
	.w7(32'h3a46394f),
	.w8(32'hb9cd8ad2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110ffc),
	.w1(32'hbbdce86a),
	.w2(32'hb9955269),
	.w3(32'h3b95c3e5),
	.w4(32'hbb78ebd1),
	.w5(32'h3abd5f02),
	.w6(32'hbbce429d),
	.w7(32'hb9a2e052),
	.w8(32'h3b7e0909),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa188ae),
	.w1(32'h3a90aa5d),
	.w2(32'h3a5dc8d6),
	.w3(32'h3b59e4a8),
	.w4(32'h3a120ae4),
	.w5(32'h3af02f19),
	.w6(32'hba772796),
	.w7(32'h38f0f207),
	.w8(32'h3a62810d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08d084),
	.w1(32'hba85cfe0),
	.w2(32'hbacadb9b),
	.w3(32'h3b2cdd45),
	.w4(32'hbaf6f3bc),
	.w5(32'h3aea8b1a),
	.w6(32'h3afd912e),
	.w7(32'hbae6789d),
	.w8(32'h3ad66fde),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915c191),
	.w1(32'h3b2db35a),
	.w2(32'hb95695c3),
	.w3(32'h39ad5851),
	.w4(32'h3ab694b7),
	.w5(32'h3a99a6d4),
	.w6(32'h3b9fa73c),
	.w7(32'h3b51f46a),
	.w8(32'h3b367d21),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae95124),
	.w1(32'h3b2a9df2),
	.w2(32'h3a537880),
	.w3(32'hba124551),
	.w4(32'hb7726625),
	.w5(32'h3ae34b90),
	.w6(32'h3b814d48),
	.w7(32'h3b8e251a),
	.w8(32'h3b9bd4a3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1d650),
	.w1(32'hbb5a9e98),
	.w2(32'hbbe26cf7),
	.w3(32'hba841b09),
	.w4(32'hbb6e6a7c),
	.w5(32'hbba670af),
	.w6(32'hbb93e1fb),
	.w7(32'hbb75c221),
	.w8(32'hbb0aabb3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eb0ee),
	.w1(32'h3a5e4f2a),
	.w2(32'h3ac9f1dd),
	.w3(32'hbb62042b),
	.w4(32'hb765b2fd),
	.w5(32'h398a6ffe),
	.w6(32'h3a62c21f),
	.w7(32'h3a8d86eb),
	.w8(32'h398550ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46a5cd),
	.w1(32'h3aabfeda),
	.w2(32'h3b400008),
	.w3(32'hb9517b27),
	.w4(32'h3aa20e4d),
	.w5(32'h3b0f36dc),
	.w6(32'h3a2255c2),
	.w7(32'h3a373419),
	.w8(32'hb95787f6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29bb59),
	.w1(32'h3a826e59),
	.w2(32'h3afd6ef3),
	.w3(32'h3b31588e),
	.w4(32'hbaff69de),
	.w5(32'hb9169b84),
	.w6(32'hba4c7252),
	.w7(32'h3aaf3b3e),
	.w8(32'h3875e344),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3439aa),
	.w1(32'hbb713c01),
	.w2(32'h3b19c93a),
	.w3(32'hba25678f),
	.w4(32'hbb804adf),
	.w5(32'h3b29b474),
	.w6(32'hbb2bad9c),
	.w7(32'h39f11d48),
	.w8(32'hbb346fb8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c410),
	.w1(32'h3a0f111d),
	.w2(32'h3aeee987),
	.w3(32'hbb643ebf),
	.w4(32'h3b818cdf),
	.w5(32'h3b0bd7b0),
	.w6(32'hb9c84c92),
	.w7(32'h3aa07103),
	.w8(32'h3b0363a8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b177063),
	.w1(32'h3b6220af),
	.w2(32'h3b518336),
	.w3(32'h3b09319f),
	.w4(32'h388e6077),
	.w5(32'h39b478e3),
	.w6(32'hb9e11c49),
	.w7(32'h3a49d7cc),
	.w8(32'h3b629d46),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47be05),
	.w1(32'h3bdc9f43),
	.w2(32'h3a1c6f47),
	.w3(32'h39ba1b22),
	.w4(32'h3b119d9b),
	.w5(32'h3b62a74f),
	.w6(32'h3b224bf0),
	.w7(32'h3c01085a),
	.w8(32'h3ba2b04b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237c43),
	.w1(32'h3b186308),
	.w2(32'h397494cd),
	.w3(32'h3b8fc931),
	.w4(32'h3a1d9598),
	.w5(32'h3a98fd57),
	.w6(32'h3bb66fc5),
	.w7(32'h3b5f867e),
	.w8(32'h3b647471),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a916c63),
	.w1(32'h3a1a45f9),
	.w2(32'hbb2df246),
	.w3(32'hb9bf8e7d),
	.w4(32'hba223dc6),
	.w5(32'h3b13e53d),
	.w6(32'hb9d6e18d),
	.w7(32'h3b0c1c68),
	.w8(32'h3a7b35a1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994cee7),
	.w1(32'h39c708a5),
	.w2(32'h3b651437),
	.w3(32'hba85af80),
	.w4(32'h3abbc463),
	.w5(32'hb929a2f2),
	.w6(32'hb9bdb812),
	.w7(32'hba91d626),
	.w8(32'h3a78fb2d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1888a),
	.w1(32'hbb5e4af9),
	.w2(32'h3a784008),
	.w3(32'h3b3a7684),
	.w4(32'hbafbced3),
	.w5(32'h3ae22990),
	.w6(32'hbaf11fec),
	.w7(32'h3aab87d3),
	.w8(32'hbaa62cec),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad069dd),
	.w1(32'hba304c76),
	.w2(32'hbb3e0718),
	.w3(32'h3a9310d4),
	.w4(32'hbb012e58),
	.w5(32'hba855886),
	.w6(32'h3b0dfe8b),
	.w7(32'hbaf80d32),
	.w8(32'hba3c0da0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb171a08),
	.w1(32'h3b152698),
	.w2(32'hba5d1d8a),
	.w3(32'hbadfd808),
	.w4(32'h3aa933be),
	.w5(32'hba76d749),
	.w6(32'h3b6a2fae),
	.w7(32'h3a87a7fe),
	.w8(32'h3ad67fe5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb97a),
	.w1(32'h3ab16857),
	.w2(32'h3b8ac8fb),
	.w3(32'h3bb60d8a),
	.w4(32'h3af6b5d8),
	.w5(32'h3b9be72b),
	.w6(32'h3b22138e),
	.w7(32'h3bafaf4c),
	.w8(32'h3b36088c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35bd09),
	.w1(32'h3b3d39ec),
	.w2(32'h3b5be13e),
	.w3(32'h3bbf325d),
	.w4(32'h3b4ee197),
	.w5(32'h3bc5ee70),
	.w6(32'h3ab740a7),
	.w7(32'h3b8a26cb),
	.w8(32'h3b64469e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0ef6),
	.w1(32'h3a16500c),
	.w2(32'h3b6bede3),
	.w3(32'h3b8d6174),
	.w4(32'h3ac6ba6e),
	.w5(32'h3b41c6a6),
	.w6(32'h3b12c08c),
	.w7(32'h3bb29905),
	.w8(32'h3b9885c8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ded9),
	.w1(32'h3b150b6e),
	.w2(32'h3b1358d2),
	.w3(32'h3b8483b8),
	.w4(32'h3b393607),
	.w5(32'h3b1a7bf6),
	.w6(32'h3ae3acaf),
	.w7(32'h3a9171ee),
	.w8(32'h3b76c622),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ed236),
	.w1(32'h3b06b4ba),
	.w2(32'h38f30fe2),
	.w3(32'h3b3bea7e),
	.w4(32'hb929fd39),
	.w5(32'h38778c59),
	.w6(32'hbb1a4002),
	.w7(32'hba4b94b7),
	.w8(32'h3a130d11),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393315c6),
	.w1(32'h3b3051f5),
	.w2(32'h3b120cef),
	.w3(32'h38161146),
	.w4(32'h3b90d551),
	.w5(32'h3a08bc77),
	.w6(32'h3ae7e4b0),
	.w7(32'h3b189a26),
	.w8(32'h3af8d737),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b70cf),
	.w1(32'h3b2aefb2),
	.w2(32'hbb13fb9c),
	.w3(32'hbacfb3ee),
	.w4(32'h3b92bca3),
	.w5(32'h3b70b820),
	.w6(32'h3b798ad3),
	.w7(32'h3a862960),
	.w8(32'hbb02aaab),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a287819),
	.w1(32'h3ad5ea3b),
	.w2(32'hbb508151),
	.w3(32'hba798a8c),
	.w4(32'h3b739298),
	.w5(32'h3ac0a3c6),
	.w6(32'h3b9e7419),
	.w7(32'h3a8975e0),
	.w8(32'hbae31997),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35c2dc),
	.w1(32'h3a2fe129),
	.w2(32'h3b167510),
	.w3(32'hba34bba9),
	.w4(32'h3bd6fc50),
	.w5(32'h3bdd8646),
	.w6(32'hbadb5d18),
	.w7(32'h3b497bc8),
	.w8(32'h3b3516a5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41027b),
	.w1(32'h3aa3b018),
	.w2(32'h3b204155),
	.w3(32'h3b2fc35c),
	.w4(32'h3b65f272),
	.w5(32'h3b994352),
	.w6(32'hba036151),
	.w7(32'h39c32bf3),
	.w8(32'h3b151e22),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3efc60),
	.w1(32'hbb189b36),
	.w2(32'hbb1e23fa),
	.w3(32'h3b3f1c50),
	.w4(32'h39b40c93),
	.w5(32'h3a81fefe),
	.w6(32'hbb4f6824),
	.w7(32'hbb56d196),
	.w8(32'hbb25c8c2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9da87a),
	.w1(32'h39a27b45),
	.w2(32'hbab7a4f1),
	.w3(32'h3abe2072),
	.w4(32'hbc080b1d),
	.w5(32'hbc1c67a6),
	.w6(32'h3bc15d7b),
	.w7(32'h3ba8bbf1),
	.w8(32'h3b768fd3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c6e08),
	.w1(32'hbae14f25),
	.w2(32'hb99ded75),
	.w3(32'hbc09bb49),
	.w4(32'h3ab2cc69),
	.w5(32'h3b6265a4),
	.w6(32'hbb503249),
	.w7(32'hbb666433),
	.w8(32'hbb167f81),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6bd72),
	.w1(32'h3a467491),
	.w2(32'h3af17bcf),
	.w3(32'h3b8fed17),
	.w4(32'h3b57c577),
	.w5(32'h3b0e763a),
	.w6(32'h3b1dd4ab),
	.w7(32'h3b7f1ffc),
	.w8(32'h3b19e6ab),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7ca0a),
	.w1(32'hbb7c68fe),
	.w2(32'hbaf87d8c),
	.w3(32'h3a44624c),
	.w4(32'h39c01487),
	.w5(32'h3b2a00ff),
	.w6(32'hba3c154d),
	.w7(32'h3a6a24f5),
	.w8(32'h3b5b4769),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e79c51),
	.w1(32'hba4829b1),
	.w2(32'hbaacbc4f),
	.w3(32'h3a1cda4f),
	.w4(32'hb8b706c4),
	.w5(32'hba89d4fc),
	.w6(32'h38bec8be),
	.w7(32'h3b68e472),
	.w8(32'h3b13a70f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f92dc2),
	.w1(32'h39ab7b7c),
	.w2(32'hb74e9b72),
	.w3(32'h3ac2c2c3),
	.w4(32'h3a40affc),
	.w5(32'h398b6481),
	.w6(32'h3a049411),
	.w7(32'h3a112ced),
	.w8(32'hb976898c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40da1f),
	.w1(32'hb96d31f2),
	.w2(32'h38bffa25),
	.w3(32'hba86fdde),
	.w4(32'h3ab43fb0),
	.w5(32'h3ad5f734),
	.w6(32'hba4e3ae8),
	.w7(32'hb8cbbab5),
	.w8(32'h3a6d763a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a72d4),
	.w1(32'hbb019636),
	.w2(32'h3be1c9a2),
	.w3(32'h3a8c3833),
	.w4(32'h3af9a319),
	.w5(32'h3b9e75da),
	.w6(32'hba36ba14),
	.w7(32'h3bdf7a6f),
	.w8(32'h3b4f777e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39316117),
	.w1(32'hbb6a8cce),
	.w2(32'hb9952639),
	.w3(32'h3b34d968),
	.w4(32'hb9e6c7eb),
	.w5(32'h3b5f1559),
	.w6(32'hbb983740),
	.w7(32'hbb0fe64e),
	.w8(32'h39b8c0d8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a918ab2),
	.w1(32'h3b4f38b1),
	.w2(32'h3a0f153a),
	.w3(32'h3b264ce2),
	.w4(32'h3adcda62),
	.w5(32'h3bbe7ead),
	.w6(32'h3b909bfd),
	.w7(32'h3b8709e8),
	.w8(32'h3a43e47c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc351c7),
	.w1(32'hbb7d15a2),
	.w2(32'hbb226fc8),
	.w3(32'h3c0ca975),
	.w4(32'hbab5f65a),
	.w5(32'h3a1ea9e4),
	.w6(32'hbacf4e81),
	.w7(32'hbab830ff),
	.w8(32'h3ac81b6b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e63c2),
	.w1(32'hba054b23),
	.w2(32'h3ad4495a),
	.w3(32'h3b12c28b),
	.w4(32'h3adf9d86),
	.w5(32'h3a9e9600),
	.w6(32'h3ac42f42),
	.w7(32'h3aa7f471),
	.w8(32'hba8f1de8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8dfd2),
	.w1(32'hbba6d744),
	.w2(32'hbb8a9242),
	.w3(32'h3aaf313d),
	.w4(32'h3a6b0a5b),
	.w5(32'hbb936395),
	.w6(32'hbbc5cf35),
	.w7(32'hbb3a3bf5),
	.w8(32'h3a29c271),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824dfb),
	.w1(32'hba8967fa),
	.w2(32'hbad56e95),
	.w3(32'hbb6338d4),
	.w4(32'h39be96ff),
	.w5(32'hbb077c4f),
	.w6(32'h3a3dbf84),
	.w7(32'hbb99caa6),
	.w8(32'h3ad41a53),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba21213),
	.w1(32'hbc13b178),
	.w2(32'hbc0e677b),
	.w3(32'h3aeebd48),
	.w4(32'hbc127727),
	.w5(32'hbc05b011),
	.w6(32'hbb96973f),
	.w7(32'hbb22d378),
	.w8(32'hbb571cb7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ae2a),
	.w1(32'hb96a840a),
	.w2(32'hba5afadf),
	.w3(32'hbc0e9c9f),
	.w4(32'hbab97616),
	.w5(32'h3b1ef9d7),
	.w6(32'h3b71095b),
	.w7(32'h39a698c2),
	.w8(32'h3a5f42e4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e01ad),
	.w1(32'h3b68ba81),
	.w2(32'hbb0c3695),
	.w3(32'h3a833052),
	.w4(32'hbb148704),
	.w5(32'h3a82d2fc),
	.w6(32'h3b9e96ed),
	.w7(32'h3bda887d),
	.w8(32'h3a456cf6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ed1a8),
	.w1(32'hb9ca117b),
	.w2(32'hbb3779ee),
	.w3(32'h3b8e4252),
	.w4(32'hbb9a2ce4),
	.w5(32'hbb58baf1),
	.w6(32'hba8b4eec),
	.w7(32'hba841874),
	.w8(32'h3b4bfc23),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb39811),
	.w1(32'h3ba1e087),
	.w2(32'h3be412a1),
	.w3(32'h3b94b078),
	.w4(32'h3b8ab8f3),
	.w5(32'h3bd400c4),
	.w6(32'h3b6ede7c),
	.w7(32'h3b912ba6),
	.w8(32'h3b781e36),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba61e29),
	.w1(32'h3935270a),
	.w2(32'h3aa59e37),
	.w3(32'h3b8f4965),
	.w4(32'hba409ea0),
	.w5(32'h3a94d643),
	.w6(32'h3b80ec53),
	.w7(32'h3b69c40d),
	.w8(32'h3b14c547),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55e64d),
	.w1(32'hbb8e5657),
	.w2(32'h396aa702),
	.w3(32'h3b624836),
	.w4(32'hbb2dcde6),
	.w5(32'hb94f4721),
	.w6(32'hbb46a137),
	.w7(32'h3ad8f4ae),
	.w8(32'h399e3c51),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90b2de),
	.w1(32'h3b18e536),
	.w2(32'h3a872b7f),
	.w3(32'hb9ff4209),
	.w4(32'h3a35625d),
	.w5(32'hb9e01a41),
	.w6(32'h3b7c8b8a),
	.w7(32'h3b67ced5),
	.w8(32'h3adb9deb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a026f93),
	.w1(32'hbade79c5),
	.w2(32'hbb817c8f),
	.w3(32'h39110029),
	.w4(32'h39de79f3),
	.w5(32'hbaf0f8bc),
	.w6(32'hb906ef0e),
	.w7(32'hbaf421bd),
	.w8(32'h3ad0e4ab),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac75ef5),
	.w1(32'hbb04bb99),
	.w2(32'hbb225c46),
	.w3(32'h3a5b1915),
	.w4(32'hba89562f),
	.w5(32'hbacd6f3d),
	.w6(32'hbab55b04),
	.w7(32'hbb33f801),
	.w8(32'hbaf3a1ba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba371a26),
	.w1(32'hbb7c9d7a),
	.w2(32'hbb7a03fd),
	.w3(32'h3af44fe6),
	.w4(32'hbb790ec7),
	.w5(32'hbb84ac0c),
	.w6(32'hbb59f24a),
	.w7(32'hbb889e9f),
	.w8(32'hbbbca4d2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2e4dd),
	.w1(32'h3a9d87b2),
	.w2(32'hb9e9aa27),
	.w3(32'hbbc998b2),
	.w4(32'h3b0541d2),
	.w5(32'h3b3bf9a0),
	.w6(32'h3b25738c),
	.w7(32'h390b72ff),
	.w8(32'h3940dbe9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a691b62),
	.w1(32'h3a104de0),
	.w2(32'h3ae603b8),
	.w3(32'h3b2aeff6),
	.w4(32'h3a244339),
	.w5(32'h38dabb74),
	.w6(32'h3ac8c008),
	.w7(32'hb996a2e0),
	.w8(32'hbb219837),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b571),
	.w1(32'h3abbfc56),
	.w2(32'hba8e4098),
	.w3(32'h39addfa7),
	.w4(32'h3b941935),
	.w5(32'h3af07ab5),
	.w6(32'h3a0fb75d),
	.w7(32'hba080885),
	.w8(32'hbb3b9e38),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bd7e7),
	.w1(32'hbab1c47d),
	.w2(32'hbb0847f3),
	.w3(32'hb9df75b6),
	.w4(32'h398edaf5),
	.w5(32'hb9ef2ae2),
	.w6(32'hba238724),
	.w7(32'hbab3152e),
	.w8(32'h3a80e3dc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd57bd),
	.w1(32'hbb23d9fc),
	.w2(32'hbb415a43),
	.w3(32'h3b003aab),
	.w4(32'h3aa89d86),
	.w5(32'h3a657518),
	.w6(32'hba6bf652),
	.w7(32'hbb2ea460),
	.w8(32'h3982e72c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55685c),
	.w1(32'h3990aa77),
	.w2(32'h3ac42c20),
	.w3(32'hbae8e512),
	.w4(32'h3b061f58),
	.w5(32'h3a26881b),
	.w6(32'hbaa0f53a),
	.w7(32'h3b52ad5e),
	.w8(32'h3b067cc6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39944d44),
	.w1(32'h3abb4c0a),
	.w2(32'h3b584b94),
	.w3(32'h3ae7979e),
	.w4(32'h3b0c7fec),
	.w5(32'h3a9784de),
	.w6(32'hbb30b6fb),
	.w7(32'hba82d0a3),
	.w8(32'hbbddc161),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7814aa),
	.w1(32'hb98f81b9),
	.w2(32'hbb012437),
	.w3(32'hbb2338b6),
	.w4(32'h3a0354a0),
	.w5(32'hbad10236),
	.w6(32'h3aa9f5db),
	.w7(32'hbb477133),
	.w8(32'hbb3ee91a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa78ee0),
	.w1(32'h3ae6e746),
	.w2(32'hbac4bb1b),
	.w3(32'hba7856a4),
	.w4(32'h3b2d6855),
	.w5(32'h3b8eedfc),
	.w6(32'h3b0adb27),
	.w7(32'h3b87b6ae),
	.w8(32'h3a681b9c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af175ff),
	.w1(32'h3b5780fa),
	.w2(32'h3b0ede1a),
	.w3(32'h3b02129b),
	.w4(32'h3af517fc),
	.w5(32'hb88124a6),
	.w6(32'hba8126bd),
	.w7(32'h3b353f0d),
	.w8(32'h3a4e6f1d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8da40),
	.w1(32'h3b8eeceb),
	.w2(32'h3b665841),
	.w3(32'hbadd38f6),
	.w4(32'h3b9619ab),
	.w5(32'h3b6247d8),
	.w6(32'h3b9faf2b),
	.w7(32'h3b90fdda),
	.w8(32'h3b860a66),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219f0f),
	.w1(32'h3b545986),
	.w2(32'h39ec2d60),
	.w3(32'h3b39a99d),
	.w4(32'h3b95b00b),
	.w5(32'hb9b30c92),
	.w6(32'h3b2ec1a2),
	.w7(32'h3b91e9f5),
	.w8(32'h3a8be031),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c44b27),
	.w1(32'hb920fd1f),
	.w2(32'h3b6de6d0),
	.w3(32'h3b390161),
	.w4(32'h3bd0048e),
	.w5(32'h3b214dce),
	.w6(32'hbad2df0a),
	.w7(32'hba21b515),
	.w8(32'hb9d01267),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2ad4f),
	.w1(32'h3b012b9a),
	.w2(32'h3a40f967),
	.w3(32'hbb0daac5),
	.w4(32'h3a0db678),
	.w5(32'hbac911e3),
	.w6(32'h3a994d8a),
	.w7(32'h3ac9aa29),
	.w8(32'h3b107b60),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390087ed),
	.w1(32'hba974518),
	.w2(32'h3b298b1f),
	.w3(32'h3b3fa5e1),
	.w4(32'h39c758c6),
	.w5(32'h3a5e5ece),
	.w6(32'h3a212ab7),
	.w7(32'h3a6dc754),
	.w8(32'h3a208a79),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb333d31),
	.w1(32'hbc30a47f),
	.w2(32'hbbf64cef),
	.w3(32'hbac902eb),
	.w4(32'h3ad2e5ca),
	.w5(32'h3bbfa8aa),
	.w6(32'h3ada5a32),
	.w7(32'h3bd42500),
	.w8(32'hba93da3d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule