module layer_10_featuremap_174(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fc6c0),
	.w1(32'hb99c9c15),
	.w2(32'h3a155607),
	.w3(32'hb89c10b8),
	.w4(32'hb9a90875),
	.w5(32'h38c66015),
	.w6(32'hb8bd7dc3),
	.w7(32'hb99cf86d),
	.w8(32'hb8f05e6c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8865478),
	.w1(32'h39bb0bff),
	.w2(32'h394c44db),
	.w3(32'h399ddfee),
	.w4(32'h39e171b8),
	.w5(32'h38957987),
	.w6(32'h3a4d1932),
	.w7(32'h393dd7f3),
	.w8(32'hb8923976),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38973221),
	.w1(32'h37764da1),
	.w2(32'h39a72bb0),
	.w3(32'h394f5d79),
	.w4(32'h37509611),
	.w5(32'h391732ff),
	.w6(32'h39252eed),
	.w7(32'h397eacb2),
	.w8(32'h38b345c7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95975b9),
	.w1(32'hb9cbd39e),
	.w2(32'hba0cbb7e),
	.w3(32'hb93d1282),
	.w4(32'h37c08a13),
	.w5(32'hb95b20d1),
	.w6(32'h3983a8b1),
	.w7(32'h38582ae5),
	.w8(32'hb87e5e60),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab2f37),
	.w1(32'hb9bdb51f),
	.w2(32'hba758b14),
	.w3(32'hb8189635),
	.w4(32'h39e2f1e1),
	.w5(32'hba3ad857),
	.w6(32'hb92b0c26),
	.w7(32'hb7eb9279),
	.w8(32'h39ba5749),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e8a2c),
	.w1(32'hb8c401c9),
	.w2(32'hb98d18a5),
	.w3(32'hba22abef),
	.w4(32'h39b1c2e2),
	.w5(32'hb825e13d),
	.w6(32'hb92bab36),
	.w7(32'hb9856fe9),
	.w8(32'hb9bfd1cf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba763165),
	.w1(32'hb9360e01),
	.w2(32'h38ec154f),
	.w3(32'hb99aa45c),
	.w4(32'h3983eb21),
	.w5(32'h3a2b19b1),
	.w6(32'h39f37eb1),
	.w7(32'h3a5307e8),
	.w8(32'h3a3ba031),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ceb22),
	.w1(32'hbaecb158),
	.w2(32'hbabfe497),
	.w3(32'hbae7acc3),
	.w4(32'hba9116cc),
	.w5(32'hb9e776e3),
	.w6(32'hb861d148),
	.w7(32'hba578126),
	.w8(32'hba890bd7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d6f17),
	.w1(32'hba308af4),
	.w2(32'hba6e1b32),
	.w3(32'h392f50ce),
	.w4(32'hb87b6c41),
	.w5(32'hba07d322),
	.w6(32'h3a01cd62),
	.w7(32'h39ba12c7),
	.w8(32'hba161c5e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af269),
	.w1(32'hbb0d9953),
	.w2(32'hbaf55f61),
	.w3(32'hbb826252),
	.w4(32'hbabb61ff),
	.w5(32'hba934f21),
	.w6(32'hbb296951),
	.w7(32'hba1e5d4e),
	.w8(32'hb9e71e6b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81caa39),
	.w1(32'hb9c99c97),
	.w2(32'hba21b9ba),
	.w3(32'hb9616507),
	.w4(32'hba8d3762),
	.w5(32'hbae36dfa),
	.w6(32'hb8f5ca7d),
	.w7(32'hba6bf91b),
	.w8(32'hba78b60b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86aadc),
	.w1(32'h3a4d15cd),
	.w2(32'h3a596fe5),
	.w3(32'h3a8837b8),
	.w4(32'h3a810e7f),
	.w5(32'h3aa401b3),
	.w6(32'h3b09dea1),
	.w7(32'h3aa865c1),
	.w8(32'h3ab5213e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb537d52),
	.w1(32'hbb179673),
	.w2(32'hbb294a5f),
	.w3(32'hbb6c39e3),
	.w4(32'hbb045282),
	.w5(32'hbb2eacab),
	.w6(32'hbb13f74e),
	.w7(32'hbaa59325),
	.w8(32'hbb07d91f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dab7c),
	.w1(32'h3a35deee),
	.w2(32'h3a1e5854),
	.w3(32'hba80fd90),
	.w4(32'hba66a4a3),
	.w5(32'hba1fb5de),
	.w6(32'hba3136d5),
	.w7(32'hba07b2b4),
	.w8(32'hba27a29b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036b5e),
	.w1(32'hbb07cf00),
	.w2(32'hbab9c75c),
	.w3(32'h3a6aea10),
	.w4(32'h3aa73fe9),
	.w5(32'h3aa311a6),
	.w6(32'hbae806bf),
	.w7(32'h3a5c30e6),
	.w8(32'h3b1a6ecb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0540b6),
	.w1(32'h38c9e4a4),
	.w2(32'hba07da54),
	.w3(32'hbb03ad2e),
	.w4(32'h39d8d9ba),
	.w5(32'hb9657987),
	.w6(32'hbb100c82),
	.w7(32'hb96b7902),
	.w8(32'hbaeb074c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13a1ce),
	.w1(32'h3a47f80e),
	.w2(32'h39f42524),
	.w3(32'h39916e17),
	.w4(32'hba2cf8e7),
	.w5(32'hba24e6e2),
	.w6(32'hba027ebf),
	.w7(32'hba87cc31),
	.w8(32'hb6a7b6b8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c9e5),
	.w1(32'hbab03b60),
	.w2(32'hbb601013),
	.w3(32'hba9efb94),
	.w4(32'hba818b37),
	.w5(32'hbb82297e),
	.w6(32'h395d1c98),
	.w7(32'hba8413db),
	.w8(32'hbb2b4c2f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd666f),
	.w1(32'hbabc7135),
	.w2(32'hbad026cb),
	.w3(32'hbaa006c2),
	.w4(32'hbb0db085),
	.w5(32'hbb213be2),
	.w6(32'hba28f397),
	.w7(32'hba553da1),
	.w8(32'hbae98338),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7351c5a),
	.w1(32'hb99671ca),
	.w2(32'hb95cf19a),
	.w3(32'h376f3f75),
	.w4(32'hb94ba72a),
	.w5(32'hb9588722),
	.w6(32'hb9821f64),
	.w7(32'hb9b19621),
	.w8(32'hb8a27eb8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92acca7),
	.w1(32'h380ad46b),
	.w2(32'hb8ea1a56),
	.w3(32'hb84cb718),
	.w4(32'h399abc18),
	.w5(32'h3894354e),
	.w6(32'h38463a85),
	.w7(32'hb90a7b5e),
	.w8(32'h38a712f1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09fc03),
	.w1(32'h39dc6d2b),
	.w2(32'h39484c52),
	.w3(32'h3adc3607),
	.w4(32'hb6a892e3),
	.w5(32'h399b18a3),
	.w6(32'h3a9de73a),
	.w7(32'h3a665d4c),
	.w8(32'h39dc7881),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05113f),
	.w1(32'hbadd778d),
	.w2(32'hb991a259),
	.w3(32'hbb57cc9f),
	.w4(32'h3b4e50a2),
	.w5(32'h3b62fd5b),
	.w6(32'hbb449ddf),
	.w7(32'h3b55645a),
	.w8(32'h3aec80d2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcd814),
	.w1(32'hbaaae526),
	.w2(32'hbaee4cd5),
	.w3(32'hba88c54d),
	.w4(32'h3a373af3),
	.w5(32'hb9330f6d),
	.w6(32'hbafd65f4),
	.w7(32'h3947ed1d),
	.w8(32'h39c70d07),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae1119),
	.w1(32'hb9f74139),
	.w2(32'hbac0706e),
	.w3(32'h39c82a76),
	.w4(32'h39f82b83),
	.w5(32'hb97d56cb),
	.w6(32'hba0b0866),
	.w7(32'hb9470e3f),
	.w8(32'hba4dfe06),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb47cb),
	.w1(32'h3a892866),
	.w2(32'h3ad5f106),
	.w3(32'h3a08808f),
	.w4(32'h39938c4f),
	.w5(32'h3a2a9524),
	.w6(32'hb6513664),
	.w7(32'h3a1d8f4a),
	.w8(32'h3a84918e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d3abd),
	.w1(32'hb915e018),
	.w2(32'hb87bc569),
	.w3(32'h39817e45),
	.w4(32'hb811d137),
	.w5(32'hb9049f97),
	.w6(32'hb8b857bb),
	.w7(32'hb949e4d8),
	.w8(32'hb7590c2e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c32c),
	.w1(32'h3a4f4268),
	.w2(32'h39fcb94f),
	.w3(32'h3af457e5),
	.w4(32'hb7f6d3ee),
	.w5(32'hb9b39405),
	.w6(32'h3aebd402),
	.w7(32'h3a3737fc),
	.w8(32'hb8b77ea3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ee3d9),
	.w1(32'h39fe331f),
	.w2(32'hb981e2bc),
	.w3(32'h3a797bec),
	.w4(32'h39e395e1),
	.w5(32'hb9943a1b),
	.w6(32'h3a2df70e),
	.w7(32'hb91b59e8),
	.w8(32'h3a7f1aa0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30e8cb),
	.w1(32'hb9fede5c),
	.w2(32'h3972619e),
	.w3(32'hbacc6106),
	.w4(32'h3a28a5e1),
	.w5(32'h3aa21ca6),
	.w6(32'hbb1772ed),
	.w7(32'h399272b3),
	.w8(32'h3a94b42c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92af5f0),
	.w1(32'hb7df4b8b),
	.w2(32'h37869c4f),
	.w3(32'hb77780ce),
	.w4(32'h38e35e81),
	.w5(32'h3807156c),
	.w6(32'hb8cba691),
	.w7(32'hb8fad8af),
	.w8(32'h385525c8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889f211),
	.w1(32'hb999d5c7),
	.w2(32'h398e8a10),
	.w3(32'hb946b9c7),
	.w4(32'hb8c86c50),
	.w5(32'h3939ba9e),
	.w6(32'hb919efd3),
	.w7(32'hb8807247),
	.w8(32'h393d19a8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc3296),
	.w1(32'hba3bdb47),
	.w2(32'hba4f4024),
	.w3(32'hb9564986),
	.w4(32'hb9a79338),
	.w5(32'hba0748ef),
	.w6(32'hba431be9),
	.w7(32'h39b823ea),
	.w8(32'h3a5d40e8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad623b8),
	.w1(32'hba5c507d),
	.w2(32'h396aa96f),
	.w3(32'hba9617f8),
	.w4(32'h390fa853),
	.w5(32'h3a14e83d),
	.w6(32'hba940933),
	.w7(32'hb9b85995),
	.w8(32'hb9ce7b69),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9a790),
	.w1(32'h3964772c),
	.w2(32'h39cea42b),
	.w3(32'hb9fe5c9a),
	.w4(32'h3990029d),
	.w5(32'h398f3853),
	.w6(32'h393a2872),
	.w7(32'h39938724),
	.w8(32'hb91c47d4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98da536),
	.w1(32'hb7f718c6),
	.w2(32'h3901dc41),
	.w3(32'hb96d01c2),
	.w4(32'h38faf5fd),
	.w5(32'h395d0b18),
	.w6(32'h3908294f),
	.w7(32'h39cfb3a3),
	.w8(32'h3a178abd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb629c94),
	.w1(32'hbade9347),
	.w2(32'h3b6c134d),
	.w3(32'hbb09039c),
	.w4(32'hbad1e830),
	.w5(32'h3b5373b8),
	.w6(32'hbb2d9e29),
	.w7(32'h394885fb),
	.w8(32'h3b154d08),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb369d19),
	.w1(32'hbb0e3c11),
	.w2(32'h3a462003),
	.w3(32'h3a47f85f),
	.w4(32'h3b2ddd86),
	.w5(32'h3b782b80),
	.w6(32'h3ac1658e),
	.w7(32'h3b247239),
	.w8(32'h3b81e0a2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bf455),
	.w1(32'h3b367466),
	.w2(32'h3b29c1f6),
	.w3(32'h3bad4f2e),
	.w4(32'h3b7acfcc),
	.w5(32'h3b6bf7bc),
	.w6(32'h3bb12fe2),
	.w7(32'h3b24d860),
	.w8(32'h3b33872f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39361142),
	.w1(32'h39a83552),
	.w2(32'h39a8425f),
	.w3(32'h39e1cc13),
	.w4(32'h3a07ed47),
	.w5(32'h3a13798a),
	.w6(32'h3a077f79),
	.w7(32'h3a366156),
	.w8(32'h39f90eff),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e6e30a),
	.w1(32'hba49bab2),
	.w2(32'hba1dd187),
	.w3(32'hb93f02b2),
	.w4(32'hba6fd250),
	.w5(32'hb9f6c6ce),
	.w6(32'hba4bcc7a),
	.w7(32'hba810371),
	.w8(32'hba302ab1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e53b6e),
	.w1(32'h38e32695),
	.w2(32'h398a8213),
	.w3(32'hb9bc5d3a),
	.w4(32'h39b05ec7),
	.w5(32'h3a066508),
	.w6(32'h392aa017),
	.w7(32'h38b2f60a),
	.w8(32'hb9837458),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b534fd),
	.w1(32'h395d7211),
	.w2(32'h3acb0a70),
	.w3(32'h3a03d88c),
	.w4(32'h3a88bb56),
	.w5(32'h3aba2872),
	.w6(32'h39b3ca38),
	.w7(32'h3a093f17),
	.w8(32'h3a114584),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7569fc),
	.w1(32'hb99e8723),
	.w2(32'hbb223880),
	.w3(32'hbb6d8355),
	.w4(32'h3a83c52b),
	.w5(32'hba3d2be0),
	.w6(32'hbab8ef9b),
	.w7(32'h3af6a816),
	.w8(32'h3b250997),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1378d4),
	.w1(32'hba3c03ec),
	.w2(32'hb8297572),
	.w3(32'hb99e56ea),
	.w4(32'h3a9d7e99),
	.w5(32'h3ac2b7f4),
	.w6(32'hba361adb),
	.w7(32'h3aecedd1),
	.w8(32'h3b1bba6c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aa9e5),
	.w1(32'hba6dbc46),
	.w2(32'hba39c3f9),
	.w3(32'hba51a7eb),
	.w4(32'h3aa574b0),
	.w5(32'h3a9a311f),
	.w6(32'hba9ea169),
	.w7(32'h3af97146),
	.w8(32'h3af30f3b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46ae4a),
	.w1(32'hbaab46da),
	.w2(32'hbab6fc72),
	.w3(32'hbaf980db),
	.w4(32'h394e935b),
	.w5(32'hba156142),
	.w6(32'hbb31ca67),
	.w7(32'h39f34e0e),
	.w8(32'h3a053695),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3768df),
	.w1(32'hbb4cfccb),
	.w2(32'hbbb6a1ca),
	.w3(32'hbb2c47c3),
	.w4(32'hbb4b43e7),
	.w5(32'hbba5d3e1),
	.w6(32'h38fced66),
	.w7(32'hbae6fb62),
	.w8(32'hbb6a2045),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba052baa),
	.w1(32'h39c52c9e),
	.w2(32'h39da0eeb),
	.w3(32'hba0dcf24),
	.w4(32'h39ffb164),
	.w5(32'h3a0da9f3),
	.w6(32'hb98ae0f9),
	.w7(32'h39bea607),
	.w8(32'h3a317591),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad282b8),
	.w1(32'h3a037020),
	.w2(32'h389399c0),
	.w3(32'hba1ae0b9),
	.w4(32'h3a098a0d),
	.w5(32'h37ab1edf),
	.w6(32'hba29e352),
	.w7(32'h38c3193c),
	.w8(32'hb8e26abb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f43cc),
	.w1(32'h3ac0cd24),
	.w2(32'h3aa3a2fc),
	.w3(32'h39faf1f7),
	.w4(32'h3ae19817),
	.w5(32'h3aa9a33e),
	.w6(32'h3aacb22f),
	.w7(32'h3b02f4f1),
	.w8(32'h3ad7f1bb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367b847a),
	.w1(32'hb87507d2),
	.w2(32'h382caaf6),
	.w3(32'h3983d208),
	.w4(32'hba3ced88),
	.w5(32'hb9edeb00),
	.w6(32'h3990b478),
	.w7(32'hb952c0b9),
	.w8(32'hba3343e7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba781910),
	.w1(32'hba2383f8),
	.w2(32'hba11d27f),
	.w3(32'hb935f97d),
	.w4(32'h39d713d2),
	.w5(32'hb802a64d),
	.w6(32'hb9617bf4),
	.w7(32'h38214bd0),
	.w8(32'h38449256),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf22c4),
	.w1(32'hbb75d5dd),
	.w2(32'hbb698130),
	.w3(32'hbbae973a),
	.w4(32'hbb2d584c),
	.w5(32'hbb187034),
	.w6(32'hb954c867),
	.w7(32'h3ab933ec),
	.w8(32'h39e02bcf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39760f0b),
	.w1(32'h372dd5d0),
	.w2(32'h399b51d7),
	.w3(32'h393d1c35),
	.w4(32'h39b48f7d),
	.w5(32'h39c3ef07),
	.w6(32'h3a4b2c68),
	.w7(32'h39d08bbd),
	.w8(32'h39722171),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d9dfb),
	.w1(32'hb9876c3a),
	.w2(32'hba414c6e),
	.w3(32'h39900e33),
	.w4(32'hb689eb40),
	.w5(32'hba0aed51),
	.w6(32'hb9b2477e),
	.w7(32'hba601d47),
	.w8(32'hba02345b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9993a32),
	.w1(32'h39e6018f),
	.w2(32'h3a4bfd3b),
	.w3(32'hb98653a6),
	.w4(32'h39bf3065),
	.w5(32'h3a332631),
	.w6(32'h39ce4349),
	.w7(32'h3a06cfe1),
	.w8(32'h39abaa07),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecbdae),
	.w1(32'hb9c65776),
	.w2(32'hb9a081fa),
	.w3(32'h3a222dea),
	.w4(32'h381ec020),
	.w5(32'hb99bf2c5),
	.w6(32'hba46bd23),
	.w7(32'hb9e693cf),
	.w8(32'h384dbd2c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f76bc),
	.w1(32'h3a8b9043),
	.w2(32'h3ab68792),
	.w3(32'h3a0f9c68),
	.w4(32'h3a77868e),
	.w5(32'h3a91360a),
	.w6(32'h3a90e6da),
	.w7(32'h3a7391e9),
	.w8(32'h3a34d2aa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4127ae),
	.w1(32'h39b9372f),
	.w2(32'hb8f35974),
	.w3(32'h3a6084a0),
	.w4(32'h39041b99),
	.w5(32'hb9740463),
	.w6(32'h399afbe6),
	.w7(32'hb9aa7036),
	.w8(32'hba09e674),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a505),
	.w1(32'hb9fc68ba),
	.w2(32'hba93473b),
	.w3(32'hbab8d4d7),
	.w4(32'hba0e4bbf),
	.w5(32'hba81ddde),
	.w6(32'hb9ab0ddd),
	.w7(32'h39c8db13),
	.w8(32'hba2fd834),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e9348b),
	.w1(32'hba0a02e8),
	.w2(32'hb9b6bbf6),
	.w3(32'hb96302af),
	.w4(32'hb99d5d7b),
	.w5(32'hb995fe5d),
	.w6(32'hb88c49fe),
	.w7(32'hb8b12fb5),
	.w8(32'hba009d38),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996d099),
	.w1(32'hba220b8d),
	.w2(32'h3a0fb291),
	.w3(32'hb9176918),
	.w4(32'hba707db5),
	.w5(32'h3731bc00),
	.w6(32'hb9e32e70),
	.w7(32'hba0cd535),
	.w8(32'h37a6dbdf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a6867),
	.w1(32'h3a3fffeb),
	.w2(32'h39bbb8ff),
	.w3(32'hb8dea065),
	.w4(32'h3a589615),
	.w5(32'h3a176ff1),
	.w6(32'h3a84d966),
	.w7(32'h3a225602),
	.w8(32'h3a345197),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53e3a5),
	.w1(32'h38a5b1f1),
	.w2(32'h392e7181),
	.w3(32'h3a830c91),
	.w4(32'hb74b2ca9),
	.w5(32'h38a624a7),
	.w6(32'h39de4edd),
	.w7(32'h3926b402),
	.w8(32'h390961b9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38364ab8),
	.w1(32'hb978a941),
	.w2(32'hb822b7ac),
	.w3(32'h3824ab17),
	.w4(32'hb90ee652),
	.w5(32'h3955c2af),
	.w6(32'hb95f7a69),
	.w7(32'hb85dd8e8),
	.w8(32'hb86e1be9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9662bb),
	.w1(32'hba3283d0),
	.w2(32'hbac8d16a),
	.w3(32'hb9aa43f5),
	.w4(32'hbaf77af5),
	.w5(32'hbb3785cb),
	.w6(32'hba52a345),
	.w7(32'hbacde53f),
	.w8(32'hbb4dc40c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b65e),
	.w1(32'hbab13e0a),
	.w2(32'hbacd33ee),
	.w3(32'hbae377b6),
	.w4(32'h3974c5ab),
	.w5(32'h398beb35),
	.w6(32'hb9bc5a3f),
	.w7(32'h39409033),
	.w8(32'hb9cdd9cc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb1999),
	.w1(32'hb83fc3d8),
	.w2(32'hb9da9817),
	.w3(32'h3a1855b4),
	.w4(32'h3add7a7d),
	.w5(32'h3a98c764),
	.w6(32'h3ab91211),
	.w7(32'h3a7e0e5b),
	.w8(32'h391964bf),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f74ed),
	.w1(32'hbb14ed0f),
	.w2(32'hbaef03ba),
	.w3(32'hba182041),
	.w4(32'h39522753),
	.w5(32'h3a0e6ab6),
	.w6(32'hba538984),
	.w7(32'h39977492),
	.w8(32'h3a9a3b18),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1e77e),
	.w1(32'h395dc71a),
	.w2(32'h39f5c33d),
	.w3(32'h39be9347),
	.w4(32'h39aa7e8c),
	.w5(32'h39ff717d),
	.w6(32'h3994d7a9),
	.w7(32'h39af3dcd),
	.w8(32'h391e3bdd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dc416),
	.w1(32'hb8f8a8aa),
	.w2(32'hb8ec3e4b),
	.w3(32'h39aacd54),
	.w4(32'h3908cf18),
	.w5(32'hb834a033),
	.w6(32'hb910fa87),
	.w7(32'hb946b655),
	.w8(32'hb8d6f1d1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92498cd),
	.w1(32'hb93714a7),
	.w2(32'hb978352f),
	.w3(32'hb8da5e6a),
	.w4(32'h3821b2a6),
	.w5(32'hb91bc739),
	.w6(32'hb8d2d299),
	.w7(32'hb999578b),
	.w8(32'hb98a8b64),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9890e72),
	.w1(32'hba06bdda),
	.w2(32'hba030a2a),
	.w3(32'h3879f612),
	.w4(32'h392bd930),
	.w5(32'hba02ca67),
	.w6(32'h3a29f2fd),
	.w7(32'hb8bd38c6),
	.w8(32'hba7a92bd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e92d98),
	.w1(32'h395940ba),
	.w2(32'h39c77976),
	.w3(32'h395ce126),
	.w4(32'h39884937),
	.w5(32'h39edbbb8),
	.w6(32'h399e08b9),
	.w7(32'h39a6928d),
	.w8(32'h391c66e7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b04898),
	.w1(32'h39454421),
	.w2(32'hba928f5f),
	.w3(32'hb61e2873),
	.w4(32'hb9c6caf8),
	.w5(32'hba2778fc),
	.w6(32'h3a126c23),
	.w7(32'h39df1c02),
	.w8(32'h3987ede7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d0cda),
	.w1(32'hba9bb4d9),
	.w2(32'hbb36f7e2),
	.w3(32'hb8de93ff),
	.w4(32'hb9c853c3),
	.w5(32'hbaa8880c),
	.w6(32'hb9ee0be2),
	.w7(32'hba3aa388),
	.w8(32'h38ac16f6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81583),
	.w1(32'hba4d0ffc),
	.w2(32'hb99e4acd),
	.w3(32'hba8910ba),
	.w4(32'hba16238d),
	.w5(32'hba36c81c),
	.w6(32'hba9f4aaf),
	.w7(32'hba298f35),
	.w8(32'hba50abc8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab9bf9),
	.w1(32'hba8115e3),
	.w2(32'hba42ebc1),
	.w3(32'hb9c985fc),
	.w4(32'hb9e86ed1),
	.w5(32'hba17ba18),
	.w6(32'h39049b07),
	.w7(32'h38fa6b03),
	.w8(32'hbace62f2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb750ee59),
	.w1(32'hba07530f),
	.w2(32'hb9bad628),
	.w3(32'h39e8503e),
	.w4(32'hb9b72bd4),
	.w5(32'hba370b5e),
	.w6(32'hb9a56777),
	.w7(32'hb9b3f6a4),
	.w8(32'hba22f5b6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba769305),
	.w1(32'hba95332d),
	.w2(32'hba90a4b4),
	.w3(32'hb9d0bfea),
	.w4(32'h3910caec),
	.w5(32'hb97b3c73),
	.w6(32'hbab4e455),
	.w7(32'hba58e189),
	.w8(32'hba0a795c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e090f),
	.w1(32'h39835ae6),
	.w2(32'h376d3acb),
	.w3(32'hb98a588d),
	.w4(32'hb8a85fb9),
	.w5(32'hba065a04),
	.w6(32'h3a24d7a4),
	.w7(32'h394dc582),
	.w8(32'hb9f3faa4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a3660),
	.w1(32'hb94ca6ce),
	.w2(32'hb90ac7a1),
	.w3(32'h3928596e),
	.w4(32'hb810bdb4),
	.w5(32'hb89091f0),
	.w6(32'hb984d412),
	.w7(32'hb9b9d6d4),
	.w8(32'hb8b154c5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3832eeaf),
	.w1(32'h3974d70c),
	.w2(32'h39e4251f),
	.w3(32'h3967b1a1),
	.w4(32'h38d7106b),
	.w5(32'h39915c11),
	.w6(32'h39c93e33),
	.w7(32'h399ca389),
	.w8(32'h3945cdd3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f10153),
	.w1(32'hb9cac0e0),
	.w2(32'h3936a821),
	.w3(32'h396228ae),
	.w4(32'hb9b8e777),
	.w5(32'hb81550f2),
	.w6(32'hb9c99b78),
	.w7(32'hb8e38747),
	.w8(32'hb9c04fad),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91069d5),
	.w1(32'hb8300349),
	.w2(32'h3909ede2),
	.w3(32'hba2fd31a),
	.w4(32'h381ef2f2),
	.w5(32'h3971da81),
	.w6(32'hb8e63031),
	.w7(32'hb87c138a),
	.w8(32'hb8ec7f6e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99b786),
	.w1(32'hb7ef0bc1),
	.w2(32'h38dce527),
	.w3(32'h3a51bd71),
	.w4(32'h3aeae199),
	.w5(32'h3b115f14),
	.w6(32'h3afe811d),
	.w7(32'h3a9e4466),
	.w8(32'h3acda33a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ed715),
	.w1(32'h39b7fa26),
	.w2(32'h3a104f35),
	.w3(32'h3a00e48f),
	.w4(32'h39b2d822),
	.w5(32'h398de005),
	.w6(32'hba091473),
	.w7(32'hb93f0018),
	.w8(32'h3953e215),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace3f02),
	.w1(32'hbab646b4),
	.w2(32'hbaa1301f),
	.w3(32'hba445e1e),
	.w4(32'h38979af1),
	.w5(32'hba1b1fdd),
	.w6(32'h39ffc766),
	.w7(32'h3a70a741),
	.w8(32'hb9411da3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875b82),
	.w1(32'hba831422),
	.w2(32'hba63655a),
	.w3(32'hba75b632),
	.w4(32'hba018bb7),
	.w5(32'hba82dc6e),
	.w6(32'hba30a3d0),
	.w7(32'hba07c2aa),
	.w8(32'hba8efb3e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a004f33),
	.w1(32'h3a3bf207),
	.w2(32'h3aadd304),
	.w3(32'h3a4c6c3f),
	.w4(32'h3a960f75),
	.w5(32'h3b06ee03),
	.w6(32'h39ef0551),
	.w7(32'h39d34b7f),
	.w8(32'h3adacea9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aca04),
	.w1(32'hbafec9d0),
	.w2(32'hbb0d1e5b),
	.w3(32'hb8d53a74),
	.w4(32'hba10bded),
	.w5(32'hba3cef2f),
	.w6(32'h3b05cf97),
	.w7(32'h3b3fd23f),
	.w8(32'h3a6ea06e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accae71),
	.w1(32'h3a3243de),
	.w2(32'hb86db1e4),
	.w3(32'h3b113016),
	.w4(32'h3aa92a8c),
	.w5(32'h37e64680),
	.w6(32'h3ac36c23),
	.w7(32'h3a76ac3e),
	.w8(32'h388ca6ce),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdeb29),
	.w1(32'hbbd0f56b),
	.w2(32'hbbaf9e54),
	.w3(32'hbb6f18cc),
	.w4(32'hbaee4e78),
	.w5(32'hbafb81aa),
	.w6(32'hbae32c41),
	.w7(32'hbb11ed28),
	.w8(32'hbb472e10),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8baeb4),
	.w1(32'h3a667e29),
	.w2(32'h3a97c403),
	.w3(32'h3a8b91a6),
	.w4(32'h3ad8113c),
	.w5(32'h3b3045c8),
	.w6(32'h3a8f0d30),
	.w7(32'h3b2b8181),
	.w8(32'h3ad19afd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa66d94),
	.w1(32'hba4de5aa),
	.w2(32'hba93b3be),
	.w3(32'hba1e8b27),
	.w4(32'h382d7a19),
	.w5(32'h3a04068c),
	.w6(32'hb95f7417),
	.w7(32'h37a130ed),
	.w8(32'h3a800cb8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf9f3d),
	.w1(32'h3ac838ed),
	.w2(32'h3a26e12a),
	.w3(32'h3aee4fa2),
	.w4(32'h3abec3de),
	.w5(32'h39f70988),
	.w6(32'h3a8fa31c),
	.w7(32'h3a9ebc81),
	.w8(32'hb942b94c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1c3b),
	.w1(32'hbaaeb497),
	.w2(32'hba8e064e),
	.w3(32'hbac1c120),
	.w4(32'h3a4c4812),
	.w5(32'hb75369e0),
	.w6(32'hbb09d2aa),
	.w7(32'h3a975b1f),
	.w8(32'h3a2dd34f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba952777),
	.w1(32'h39bd064a),
	.w2(32'h3b4b5950),
	.w3(32'h3ab6f6c8),
	.w4(32'h3b17546f),
	.w5(32'h3b55415f),
	.w6(32'h3b3c2221),
	.w7(32'h3ae7edcb),
	.w8(32'h39eeeb8e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67a4bc),
	.w1(32'hb973610e),
	.w2(32'hb9b100b7),
	.w3(32'hba9d97ce),
	.w4(32'hbb14e2e1),
	.w5(32'hbaaec71d),
	.w6(32'hba9a5323),
	.w7(32'hb9c31546),
	.w8(32'hb9c32c2a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc289793),
	.w1(32'hbbddb2c8),
	.w2(32'hbb37fe13),
	.w3(32'hbabcac5a),
	.w4(32'h3b4aaec4),
	.w5(32'h3bcf6be5),
	.w6(32'h3a9ee499),
	.w7(32'h3b8c0471),
	.w8(32'h3c0de64e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a7f2c),
	.w1(32'hbb298de5),
	.w2(32'hbb0b407b),
	.w3(32'hbabd016b),
	.w4(32'h3928f490),
	.w5(32'hba99536e),
	.w6(32'hbb3e2d5f),
	.w7(32'h3930cd25),
	.w8(32'h3a4ff072),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a1b9),
	.w1(32'hbaef01df),
	.w2(32'hbaaeadec),
	.w3(32'h3a072a37),
	.w4(32'h3a4cceac),
	.w5(32'hbaa8a342),
	.w6(32'hb8bd912e),
	.w7(32'hb92fc1ec),
	.w8(32'hb9d4541b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25b517),
	.w1(32'h3a8b9eea),
	.w2(32'h3a26a90c),
	.w3(32'hba428c5a),
	.w4(32'h3a85c9ca),
	.w5(32'h3abcc53f),
	.w6(32'hb9969ebf),
	.w7(32'h3aac59e6),
	.w8(32'h3b2070dc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fd467),
	.w1(32'hbb0db9ff),
	.w2(32'hbaae7a1b),
	.w3(32'hbb16d0a1),
	.w4(32'hbb18ceea),
	.w5(32'hba526484),
	.w6(32'hb9cd7316),
	.w7(32'hba9ae85a),
	.w8(32'hb84c60c9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac91e8b),
	.w1(32'hb9ab5d22),
	.w2(32'hba9281a2),
	.w3(32'h3a102c11),
	.w4(32'hb9d72159),
	.w5(32'hb84da4f2),
	.w6(32'h3941950a),
	.w7(32'hba29da39),
	.w8(32'h39df5f89),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8b7f8),
	.w1(32'h3954f763),
	.w2(32'h39897c8b),
	.w3(32'h39939a9a),
	.w4(32'h37225502),
	.w5(32'h3841bc4a),
	.w6(32'h3a6541e7),
	.w7(32'h39b7d8e3),
	.w8(32'hb936f28a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9fd9d),
	.w1(32'hb9ab102a),
	.w2(32'hb8c22914),
	.w3(32'h378c51ef),
	.w4(32'h3965436c),
	.w5(32'h394b2077),
	.w6(32'hb79b6ed3),
	.w7(32'hb8b0a138),
	.w8(32'hb95226b8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba718839),
	.w1(32'hb9e1d153),
	.w2(32'hb9f1a5e4),
	.w3(32'hba3b8db6),
	.w4(32'h380d6f3e),
	.w5(32'hba844f0a),
	.w6(32'hbb085a1d),
	.w7(32'hb9b37ada),
	.w8(32'h38b80bf5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002109),
	.w1(32'h3af65209),
	.w2(32'h3b037ec5),
	.w3(32'hb9cec2d9),
	.w4(32'h3b33bc31),
	.w5(32'h3b286485),
	.w6(32'hba3a21b1),
	.w7(32'h3b30f7aa),
	.w8(32'h3b3a0cf4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e71d16),
	.w1(32'hbab855fa),
	.w2(32'hb9c5b1bd),
	.w3(32'h3a22faad),
	.w4(32'h3a383a5e),
	.w5(32'h3a5a81c5),
	.w6(32'h37a80367),
	.w7(32'h3a30c010),
	.w8(32'h3b2152f7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb685081),
	.w1(32'hbb66a48b),
	.w2(32'hba7f4d80),
	.w3(32'hbb0d6e97),
	.w4(32'hbb28623c),
	.w5(32'hba64a281),
	.w6(32'hbac4436b),
	.w7(32'hbb28aac9),
	.w8(32'hba786839),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2c698),
	.w1(32'hba8ccca9),
	.w2(32'h3886e288),
	.w3(32'hba135163),
	.w4(32'h37b90ac3),
	.w5(32'h3a685908),
	.w6(32'h381c03a4),
	.w7(32'h39b645f7),
	.w8(32'h3a910b77),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba28d3),
	.w1(32'h3a0c27b7),
	.w2(32'h3a2f10bb),
	.w3(32'hba715c05),
	.w4(32'h39d6a70f),
	.w5(32'hb8170d61),
	.w6(32'hba76584e),
	.w7(32'hba67bb74),
	.w8(32'hba9ff514),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5201a3),
	.w1(32'hb9ab4c52),
	.w2(32'hb9041484),
	.w3(32'hb9d4ebc0),
	.w4(32'h399e71b6),
	.w5(32'hb8bbe555),
	.w6(32'hba135eef),
	.w7(32'h392f01d4),
	.w8(32'h389d1270),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba239d08),
	.w1(32'hb951bafa),
	.w2(32'hba346c92),
	.w3(32'hb9eb26b8),
	.w4(32'h391697c9),
	.w5(32'hb9206e01),
	.w6(32'hb983131e),
	.w7(32'hb9f5b1d8),
	.w8(32'hb8c9a353),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce950d),
	.w1(32'hb93d16e8),
	.w2(32'hb9720147),
	.w3(32'hb7f53b3e),
	.w4(32'h38d3cb16),
	.w5(32'hb77f5517),
	.w6(32'hb9022419),
	.w7(32'hb9ac6365),
	.w8(32'hb9900b16),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b34f9),
	.w1(32'hb955d930),
	.w2(32'hb9da6d45),
	.w3(32'hb8778fdb),
	.w4(32'h39141a9c),
	.w5(32'hb90b56b1),
	.w6(32'hb8dd247e),
	.w7(32'hb99633ba),
	.w8(32'hb94a6788),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba0a2d),
	.w1(32'h3a2ead39),
	.w2(32'h3a3ab8fb),
	.w3(32'h3a0fc758),
	.w4(32'h3a156bf5),
	.w5(32'h3a60dbba),
	.w6(32'h3a4abf59),
	.w7(32'h3a964867),
	.w8(32'h3932f935),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08cc27),
	.w1(32'hba02d278),
	.w2(32'hb93a5aa7),
	.w3(32'hb93315d7),
	.w4(32'h3b28dc58),
	.w5(32'h3aea1e8e),
	.w6(32'hb9d553bf),
	.w7(32'h3ab48a3c),
	.w8(32'h3acd086a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393dd1a7),
	.w1(32'hba8596a9),
	.w2(32'hbaa6fa0b),
	.w3(32'hb853c174),
	.w4(32'hb988eeca),
	.w5(32'hba4db5e2),
	.w6(32'h39b5fb5a),
	.w7(32'h39a62046),
	.w8(32'hb9e84020),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c986),
	.w1(32'hbab5668c),
	.w2(32'hbaa53274),
	.w3(32'hbaae3ace),
	.w4(32'hba2e8e3f),
	.w5(32'hba3d79fc),
	.w6(32'hbab7140c),
	.w7(32'hba5adabc),
	.w8(32'hb9c315e3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04ff85),
	.w1(32'hba83f1f0),
	.w2(32'hba15edd5),
	.w3(32'hb99af1d4),
	.w4(32'hb9ae397f),
	.w5(32'hb998e6ab),
	.w6(32'hba6ad42c),
	.w7(32'hbaa46264),
	.w8(32'hb9d3ef24),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9815bc2),
	.w1(32'hb8d9a56d),
	.w2(32'hba2b2e83),
	.w3(32'hb7fbe569),
	.w4(32'hb99d6c94),
	.w5(32'hb8d6c8c7),
	.w6(32'h393b5940),
	.w7(32'h395e6b4f),
	.w8(32'hb8e2c564),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e6703),
	.w1(32'hb8c5fd9e),
	.w2(32'hba214ec8),
	.w3(32'hb96319a1),
	.w4(32'h39b01019),
	.w5(32'hb92aead8),
	.w6(32'hb892662f),
	.w7(32'hba0c9ccc),
	.w8(32'hb99b07f5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a31e6),
	.w1(32'hb971039a),
	.w2(32'hb96b9410),
	.w3(32'h38c3912e),
	.w4(32'h37dace1c),
	.w5(32'hb8e3799e),
	.w6(32'hb91d75e5),
	.w7(32'hb9ad01a0),
	.w8(32'h3650c813),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c6a64),
	.w1(32'h3ab4e10c),
	.w2(32'hbb03a9a0),
	.w3(32'h39bf6ca7),
	.w4(32'h3b1909d8),
	.w5(32'hbaaf0252),
	.w6(32'h3b25cdbf),
	.w7(32'hba5788e0),
	.w8(32'h39d477e6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cfc12),
	.w1(32'hbba354b5),
	.w2(32'hbbf26171),
	.w3(32'hba91d153),
	.w4(32'hbb8223b4),
	.w5(32'hbbb87186),
	.w6(32'hbb8a561c),
	.w7(32'hbba4306d),
	.w8(32'hbb5fbd1a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd04b00),
	.w1(32'h3bf57eb9),
	.w2(32'hbb00f0aa),
	.w3(32'hbbb709f9),
	.w4(32'h3c87d38d),
	.w5(32'h3c04ae24),
	.w6(32'h3a47b869),
	.w7(32'hbbd219e0),
	.w8(32'hbc5c6eca),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf69b27),
	.w1(32'h3b15b562),
	.w2(32'h3c08b9ab),
	.w3(32'hbb58dabf),
	.w4(32'hb99feba7),
	.w5(32'h3bb5c241),
	.w6(32'hbb0c96cb),
	.w7(32'h3b54fc95),
	.w8(32'hba4a8412),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cbe31),
	.w1(32'h3b2e670e),
	.w2(32'h3bb857c8),
	.w3(32'h3826ed93),
	.w4(32'hb823635f),
	.w5(32'h3ad6c757),
	.w6(32'h3ac06298),
	.w7(32'h3b794543),
	.w8(32'h3b1d629d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4480c0),
	.w1(32'h3bc96d89),
	.w2(32'h3bf8eeaf),
	.w3(32'hba501d83),
	.w4(32'h3b3ce454),
	.w5(32'h3b4835a8),
	.w6(32'h3c3eed96),
	.w7(32'h3c40d864),
	.w8(32'h3c147c91),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a25bd),
	.w1(32'hbbd2968c),
	.w2(32'h394a2f4e),
	.w3(32'h3b196d04),
	.w4(32'hbbb92c4e),
	.w5(32'hba4ff0fe),
	.w6(32'hbb9ba80a),
	.w7(32'h39f83f7c),
	.w8(32'h3bc6f3c8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8139c),
	.w1(32'hbb740274),
	.w2(32'hbad6a212),
	.w3(32'h3bb5c3cc),
	.w4(32'hbb04f444),
	.w5(32'hba305f75),
	.w6(32'hbb4e3f6c),
	.w7(32'hbad704b1),
	.w8(32'hba74f607),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8983eb6),
	.w1(32'hbb12ba6d),
	.w2(32'h3b9707db),
	.w3(32'h3a01075b),
	.w4(32'hbb1f57d0),
	.w5(32'h3b780cee),
	.w6(32'hbbe6ea98),
	.w7(32'h394f1169),
	.w8(32'hba81a07e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f656),
	.w1(32'hbc0cbeae),
	.w2(32'hbc453698),
	.w3(32'h3b1a52c6),
	.w4(32'hbbd33e20),
	.w5(32'hbc2d3913),
	.w6(32'hbbf5f9b1),
	.w7(32'hbc251f71),
	.w8(32'hbc0167ec),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d13a2),
	.w1(32'hb972d3e1),
	.w2(32'hbb18bb87),
	.w3(32'hbc18b3a9),
	.w4(32'h3aa8460c),
	.w5(32'hba86758b),
	.w6(32'hb8a181e5),
	.w7(32'hbb268aec),
	.w8(32'hbaeb37db),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb309821),
	.w1(32'h3b85e20c),
	.w2(32'h3c458841),
	.w3(32'hbb096584),
	.w4(32'h3a64d743),
	.w5(32'h3c0a39ea),
	.w6(32'h3a334087),
	.w7(32'h3c07eba8),
	.w8(32'h3b6e3590),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf77131),
	.w1(32'h3b34fac2),
	.w2(32'h3b0c2b9a),
	.w3(32'h3ba76c77),
	.w4(32'h3b501b6e),
	.w5(32'h3b709752),
	.w6(32'h3b44fc3b),
	.w7(32'h3aec6fc3),
	.w8(32'h3add9d98),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab55b9e),
	.w1(32'hbb6ec286),
	.w2(32'hbb53729e),
	.w3(32'h3b0650cb),
	.w4(32'hbac09836),
	.w5(32'hbb416acc),
	.w6(32'hba9a31e4),
	.w7(32'hbaa6cc5a),
	.w8(32'hbaecd6bb),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4954),
	.w1(32'h38eed078),
	.w2(32'hbaa6ccc0),
	.w3(32'hbb66fe51),
	.w4(32'h3a76120f),
	.w5(32'hba18c8c7),
	.w6(32'h38ebffe1),
	.w7(32'hba674124),
	.w8(32'hb66c5efd),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee7d52),
	.w1(32'hbc6ef9ca),
	.w2(32'hbc918f38),
	.w3(32'h3a8e7992),
	.w4(32'hbc2c0127),
	.w5(32'hbc844998),
	.w6(32'hbc2dfe30),
	.w7(32'hbc6aa369),
	.w8(32'hbc55c9d5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79a50b),
	.w1(32'hbb349348),
	.w2(32'hb9c91b3a),
	.w3(32'hbc5d3f65),
	.w4(32'hbb27c1fa),
	.w5(32'hbadd155a),
	.w6(32'h39e11115),
	.w7(32'hb9ed05b5),
	.w8(32'h3a10ed5e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade465b),
	.w1(32'hb9a89cf9),
	.w2(32'hbad034a6),
	.w3(32'hbb1116bc),
	.w4(32'hba26acaa),
	.w5(32'hbb1ebb76),
	.w6(32'hba3b0ee6),
	.w7(32'hbac569d9),
	.w8(32'hbb0ed497),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb162fa7),
	.w1(32'hbb1d243c),
	.w2(32'hbb1e69f9),
	.w3(32'hbb444b2d),
	.w4(32'hba464a31),
	.w5(32'hba923872),
	.w6(32'hbb1125a9),
	.w7(32'hbb2733a2),
	.w8(32'hba4e220a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39f2d),
	.w1(32'h3a93536b),
	.w2(32'h3be8ed9e),
	.w3(32'h37f74674),
	.w4(32'hbacd1c1e),
	.w5(32'h3b903634),
	.w6(32'hbb45dd12),
	.w7(32'h3ae7f775),
	.w8(32'hba8bc19e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a8e5),
	.w1(32'hba45e248),
	.w2(32'h3b2aaa89),
	.w3(32'h3a4f06fc),
	.w4(32'hbaa5c9e2),
	.w5(32'h3aeec050),
	.w6(32'hbb527f3c),
	.w7(32'hb9ccdaa9),
	.w8(32'hbaf90670),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f6bf),
	.w1(32'hba807a10),
	.w2(32'hbb0616a7),
	.w3(32'hbba0fc8f),
	.w4(32'hbaa5d4ba),
	.w5(32'hbb2e7ae4),
	.w6(32'h3a1eca9a),
	.w7(32'hbacf1322),
	.w8(32'hbb2dbb9c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc75f4),
	.w1(32'h3aac555b),
	.w2(32'hbb16c64d),
	.w3(32'h38cb9402),
	.w4(32'h3afdc475),
	.w5(32'hbb0ad3ba),
	.w6(32'h3b47427a),
	.w7(32'hba4a9fec),
	.w8(32'h39bfc5df),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78d37f),
	.w1(32'hbb5410ed),
	.w2(32'hbb04c6e7),
	.w3(32'hbaf1a725),
	.w4(32'hba9bb6ae),
	.w5(32'hbbb883b6),
	.w6(32'hbb4400d0),
	.w7(32'h37c45d7a),
	.w8(32'hba2bd2a1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11a43),
	.w1(32'hb9baf343),
	.w2(32'hbb4ae331),
	.w3(32'hbb92df62),
	.w4(32'hb9e6415f),
	.w5(32'hbb4020e4),
	.w6(32'hbac39cb8),
	.w7(32'hbaa8b2d3),
	.w8(32'hbb3f2e38),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94a26e),
	.w1(32'hbc084ff2),
	.w2(32'hbc401545),
	.w3(32'hbb244190),
	.w4(32'hbbeb38e3),
	.w5(32'hbc346739),
	.w6(32'hbc0e0be5),
	.w7(32'hbc38d848),
	.w8(32'hbc254004),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e71fc),
	.w1(32'h3baa5780),
	.w2(32'h3b98af94),
	.w3(32'hbc08bd0d),
	.w4(32'h3aa1e389),
	.w5(32'hba5b9e57),
	.w6(32'h3be60a0f),
	.w7(32'h3be3d051),
	.w8(32'h3a796bc8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb065d0e),
	.w1(32'hba6583b9),
	.w2(32'h3abbd28e),
	.w3(32'hbc00dcf6),
	.w4(32'hbaf6b426),
	.w5(32'hbb5dd742),
	.w6(32'hb6ce8e4c),
	.w7(32'h3b41a8d1),
	.w8(32'h3b104686),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60966a),
	.w1(32'h3ab5c41b),
	.w2(32'h39cb7d48),
	.w3(32'hbb0b3262),
	.w4(32'h3b2a58e1),
	.w5(32'h3b03a4c8),
	.w6(32'h3b0958d7),
	.w7(32'h3a4f7d54),
	.w8(32'h3a977d72),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02adf4),
	.w1(32'h3bb57b04),
	.w2(32'h3bb3ed7b),
	.w3(32'hbaae7738),
	.w4(32'h3b256522),
	.w5(32'h3b39eae0),
	.w6(32'h3ae6930c),
	.w7(32'h3b9854d1),
	.w8(32'hb99ef4c5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ec934),
	.w1(32'h3ba1c94a),
	.w2(32'hb949a477),
	.w3(32'hbbd89d42),
	.w4(32'h3bb7f5d7),
	.w5(32'hba016cf6),
	.w6(32'h3c08cf05),
	.w7(32'hb99443b2),
	.w8(32'hb953a11b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39039c97),
	.w1(32'h39e0d2a0),
	.w2(32'hbac9806a),
	.w3(32'h396f4537),
	.w4(32'h39db8147),
	.w5(32'hbac2671e),
	.w6(32'h3b056ae0),
	.w7(32'hb94edd56),
	.w8(32'hb9a7ea95),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e1012),
	.w1(32'h3a51e721),
	.w2(32'hba9e344c),
	.w3(32'hbb51ac12),
	.w4(32'h3aa34e05),
	.w5(32'hba80d905),
	.w6(32'h3adb1ddf),
	.w7(32'hb9e56c58),
	.w8(32'h3a027677),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa0240),
	.w1(32'h3ab61c91),
	.w2(32'h3921a4ad),
	.w3(32'hb95a207f),
	.w4(32'h3b0e8909),
	.w5(32'h3a33ade8),
	.w6(32'h3ae34243),
	.w7(32'h398adbb3),
	.w8(32'h3a8e7607),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32637),
	.w1(32'h3aec731a),
	.w2(32'h3ba713d9),
	.w3(32'hb9b79f0e),
	.w4(32'h3b3fc247),
	.w5(32'h3bc8c881),
	.w6(32'hb8bd15a0),
	.w7(32'h3b5c177a),
	.w8(32'hb8bd00fa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3596a1),
	.w1(32'hbadfa0c8),
	.w2(32'h3b13c1f4),
	.w3(32'hba9846bf),
	.w4(32'hbb138478),
	.w5(32'h3a97eea6),
	.w6(32'hba824f7c),
	.w7(32'h3ad2099a),
	.w8(32'h3b2c8b77),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e91f),
	.w1(32'h3b3d0560),
	.w2(32'h3c3930a1),
	.w3(32'h3b2f7d24),
	.w4(32'hba890bf2),
	.w5(32'h3bffe01a),
	.w6(32'hbb365d4b),
	.w7(32'h3bb5f804),
	.w8(32'h3b3d1fcf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012dc6),
	.w1(32'h3b20f916),
	.w2(32'h3ab8f47b),
	.w3(32'h3b8583a2),
	.w4(32'h3b21a067),
	.w5(32'h3a85a098),
	.w6(32'h3b35d7fb),
	.w7(32'h3add2578),
	.w8(32'h3b161c84),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb87440),
	.w1(32'h3aca7f9d),
	.w2(32'h3c185fc9),
	.w3(32'h3bb45100),
	.w4(32'hbb05c5ae),
	.w5(32'h3bbfdd75),
	.w6(32'h3ab1c78d),
	.w7(32'h3bc38029),
	.w8(32'h3b620ed3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5b5d3),
	.w1(32'h3a48b747),
	.w2(32'h3bcd66bb),
	.w3(32'h3b7f6176),
	.w4(32'hbabbf978),
	.w5(32'h3b80777f),
	.w6(32'hbb2d5854),
	.w7(32'h3b1a629a),
	.w8(32'hb96c3830),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f96b9),
	.w1(32'hbbb0a6a6),
	.w2(32'hbc0d94b2),
	.w3(32'h3ae69473),
	.w4(32'hbb8af301),
	.w5(32'hbbf9f799),
	.w6(32'hbb842f1b),
	.w7(32'hbbfe457c),
	.w8(32'hbbe1cb68),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e9bf2),
	.w1(32'hbbcc8bd3),
	.w2(32'h389abcb5),
	.w3(32'hbbd0662f),
	.w4(32'hbbc40b83),
	.w5(32'h39e6d5ba),
	.w6(32'hbc088de7),
	.w7(32'hbab2ea9d),
	.w8(32'hb9b30bcf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf665f),
	.w1(32'hbb333ef5),
	.w2(32'hbba7ec88),
	.w3(32'hbb87142b),
	.w4(32'hb9d1601a),
	.w5(32'hbb57826d),
	.w6(32'hbb8de99e),
	.w7(32'hbacc585a),
	.w8(32'hbabb9a89),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37ff84),
	.w1(32'h3b3d2a12),
	.w2(32'h3bc16190),
	.w3(32'hbb2d451f),
	.w4(32'hba9d3899),
	.w5(32'h3ad7d6d9),
	.w6(32'h3a6da191),
	.w7(32'h3b81a2de),
	.w8(32'h3afff6c6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c053f4),
	.w1(32'hbac0158d),
	.w2(32'hbac738ce),
	.w3(32'hbab55875),
	.w4(32'h393b7b0c),
	.w5(32'hba936a85),
	.w6(32'h3aac7c8c),
	.w7(32'h39c76a40),
	.w8(32'hb8115b60),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7506d0),
	.w1(32'h3ae57177),
	.w2(32'h3c2b51d0),
	.w3(32'h3ab0852e),
	.w4(32'hba5d729c),
	.w5(32'h3c009283),
	.w6(32'hbb7e2c42),
	.w7(32'h3b8a0c31),
	.w8(32'h3b229535),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee53bc),
	.w1(32'h3925e85d),
	.w2(32'h3b0d4efa),
	.w3(32'h3bd27b8d),
	.w4(32'h3a5dd827),
	.w5(32'h3b029034),
	.w6(32'h3b130f2f),
	.w7(32'h3b2e3738),
	.w8(32'h3a04a317),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9344f),
	.w1(32'hbb2aeb31),
	.w2(32'h3a833d4e),
	.w3(32'h3a274ae7),
	.w4(32'hbadc7cf9),
	.w5(32'h3af0b201),
	.w6(32'hbb824ddd),
	.w7(32'hbb06287e),
	.w8(32'hbb319108),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955dcc),
	.w1(32'hba861345),
	.w2(32'hbaba15a0),
	.w3(32'hbb0e169b),
	.w4(32'hb8c1ec6e),
	.w5(32'hbab32de5),
	.w6(32'h3ac34730),
	.w7(32'h3b5a7192),
	.w8(32'h3af1f341),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60d441),
	.w1(32'h3b6ea28d),
	.w2(32'hba8607f4),
	.w3(32'hbb5509bc),
	.w4(32'h3b6b8fe3),
	.w5(32'h395d0b1b),
	.w6(32'h3b245ab5),
	.w7(32'h39bd8215),
	.w8(32'h3ab78d0d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21748b),
	.w1(32'h3a091e74),
	.w2(32'h3a21d4bb),
	.w3(32'hba347f7b),
	.w4(32'h3ab115c7),
	.w5(32'h3a830ecd),
	.w6(32'h3a17d136),
	.w7(32'h39559178),
	.w8(32'h3a3c8338),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96cba0),
	.w1(32'hbbd812a3),
	.w2(32'hbc1bccbb),
	.w3(32'h3abfa484),
	.w4(32'hbbb0e2da),
	.w5(32'hbc11648e),
	.w6(32'hbbb47671),
	.w7(32'hbc0a7f93),
	.w8(32'hbbf8cc00),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a69e),
	.w1(32'h3b890583),
	.w2(32'h3bba8a5c),
	.w3(32'hbc04eef5),
	.w4(32'h3b150f12),
	.w5(32'h3b60c789),
	.w6(32'h3b01a229),
	.w7(32'h3b4ca7e0),
	.w8(32'h3a175e21),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0efb31),
	.w1(32'h3c3609d4),
	.w2(32'h3b75dacd),
	.w3(32'h39e8875b),
	.w4(32'h3bf0c6f6),
	.w5(32'h39eaf05a),
	.w6(32'h3c2ca632),
	.w7(32'h3b7b5a07),
	.w8(32'hbbdb6352),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2ec0),
	.w1(32'h3a85e157),
	.w2(32'h3b4567ca),
	.w3(32'hbc4e09fc),
	.w4(32'hb9960915),
	.w5(32'h3a7759c3),
	.w6(32'hb9a45d23),
	.w7(32'h3a4ddd72),
	.w8(32'hba9eb2a9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19cfad),
	.w1(32'hbc7e3d29),
	.w2(32'hba845d80),
	.w3(32'h39322d7e),
	.w4(32'hbc68d1c7),
	.w5(32'hbb38005c),
	.w6(32'hbc7a85c2),
	.w7(32'hbb924de2),
	.w8(32'h3b291ab4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7aabc),
	.w1(32'h3ac4c915),
	.w2(32'h3c101865),
	.w3(32'h3babd7a1),
	.w4(32'hbade2e13),
	.w5(32'h3b955171),
	.w6(32'h3a0c12c3),
	.w7(32'h3ba9b51c),
	.w8(32'h3b2bf4ac),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88a94f),
	.w1(32'hbb46def2),
	.w2(32'hbbbf4e6f),
	.w3(32'h3aaa5a12),
	.w4(32'hbad8ae1c),
	.w5(32'hbb9b3356),
	.w6(32'hba6f24a8),
	.w7(32'hbb728206),
	.w8(32'hbb57508b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd31127),
	.w1(32'h3c1a6722),
	.w2(32'h3c59bfc9),
	.w3(32'hbb6ae444),
	.w4(32'h3c0a6597),
	.w5(32'h3c3616ed),
	.w6(32'h3c32155d),
	.w7(32'h3c3ed0fe),
	.w8(32'h3c096098),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c138cee),
	.w1(32'hba75cba3),
	.w2(32'hba97f982),
	.w3(32'h3bb43b19),
	.w4(32'hba5c9463),
	.w5(32'hba75d21a),
	.w6(32'hbb1d61b0),
	.w7(32'hbb74c6d5),
	.w8(32'hbb0eafb0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8db9aa),
	.w1(32'h39128c16),
	.w2(32'h3ba3db5c),
	.w3(32'hbb299461),
	.w4(32'hbb433557),
	.w5(32'h3ace590a),
	.w6(32'hbb0f5409),
	.w7(32'h3a9c0eb8),
	.w8(32'hbb9592d4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eb9fe),
	.w1(32'hbc092106),
	.w2(32'hbc73caac),
	.w3(32'hbbb53b51),
	.w4(32'hbbb2c648),
	.w5(32'hbc470ef5),
	.w6(32'hbbf4924c),
	.w7(32'hbc0b9e7d),
	.w8(32'hbc251b91),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185b9f),
	.w1(32'hbc0d31f7),
	.w2(32'hbacd8dcc),
	.w3(32'hbbca4f0c),
	.w4(32'hbbdbf93f),
	.w5(32'hbac7d16e),
	.w6(32'hbc3cdcc4),
	.w7(32'hbb8c2bef),
	.w8(32'hbbf337e7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc33d),
	.w1(32'hbb743d64),
	.w2(32'hbbb60a51),
	.w3(32'hbbed2735),
	.w4(32'hbb0ea2db),
	.w5(32'hbb990cdb),
	.w6(32'hbb70a7f0),
	.w7(32'hbbaf6a7a),
	.w8(32'hbb8142c7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2acdf),
	.w1(32'hbb30debf),
	.w2(32'hbaee6d60),
	.w3(32'hbb963f60),
	.w4(32'hbb77e04b),
	.w5(32'hbb02248f),
	.w6(32'hbac4a678),
	.w7(32'hbace67b6),
	.w8(32'h3ad46723),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3af499),
	.w1(32'h3aec94ed),
	.w2(32'h3c0fd753),
	.w3(32'h3a9a1161),
	.w4(32'hb68bf789),
	.w5(32'h3bde9620),
	.w6(32'hbb24ff01),
	.w7(32'h3b86fa02),
	.w8(32'h3b32b969),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be566d1),
	.w1(32'h3bab5e75),
	.w2(32'h3be2a7c8),
	.w3(32'h3b9d4833),
	.w4(32'h3b10cb97),
	.w5(32'h3ba6d3e4),
	.w6(32'h3b34ad46),
	.w7(32'h3b597ce3),
	.w8(32'hba9a1eeb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c07ea6),
	.w1(32'hba0324b4),
	.w2(32'hbae8e938),
	.w3(32'hba87c7bd),
	.w4(32'hba4057be),
	.w5(32'hbb1bad21),
	.w6(32'hba19e1a3),
	.w7(32'hbb443971),
	.w8(32'hba874a95),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce4ec),
	.w1(32'hbb907468),
	.w2(32'hbbb5076a),
	.w3(32'hbb2899e8),
	.w4(32'hbb55fa91),
	.w5(32'hbb99c3b2),
	.w6(32'hbb0112e1),
	.w7(32'hbb75b0ec),
	.w8(32'hbb819a35),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1593d0),
	.w1(32'hbaddfcb1),
	.w2(32'hbb803864),
	.w3(32'hbbf0dbf4),
	.w4(32'hb9ec06d6),
	.w5(32'hbb20e02e),
	.w6(32'hbac072b6),
	.w7(32'hbb1189e0),
	.w8(32'hbab30135),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c04d),
	.w1(32'hbaf98eac),
	.w2(32'hbb27806b),
	.w3(32'hb7424c3c),
	.w4(32'hbab753c7),
	.w5(32'hbb2f5bdb),
	.w6(32'hba802b30),
	.w7(32'hbac5d190),
	.w8(32'hbae0ba2c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00ef3),
	.w1(32'hbb11bc02),
	.w2(32'hbb7be49b),
	.w3(32'hbb928ed0),
	.w4(32'hbb8cf4e8),
	.w5(32'hbbba269c),
	.w6(32'hbb878eb4),
	.w7(32'hbb921307),
	.w8(32'hbbd16f63),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcb9fb),
	.w1(32'h3a45bc55),
	.w2(32'h3bc505a2),
	.w3(32'hbbdf17e7),
	.w4(32'hbab738ff),
	.w5(32'h3b6d4926),
	.w6(32'hbb396d92),
	.w7(32'h3a51ceda),
	.w8(32'hba8141da),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b665ac2),
	.w1(32'hbb5777fd),
	.w2(32'hbbacd2ed),
	.w3(32'h3abb6ffa),
	.w4(32'hbb0b0b03),
	.w5(32'hbb9a171f),
	.w6(32'hbb4f3764),
	.w7(32'hbba7cb65),
	.w8(32'hbb6119d2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73695c),
	.w1(32'hbb97fc4a),
	.w2(32'hbbd7b585),
	.w3(32'hbb5a9137),
	.w4(32'hbb6e02c6),
	.w5(32'hbbcebf58),
	.w6(32'hbb8626af),
	.w7(32'hbbe08e8f),
	.w8(32'hbbb9aa16),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd88fa3),
	.w1(32'h3b0bc3eb),
	.w2(32'h3a40ef9b),
	.w3(32'hbbba6cf2),
	.w4(32'h3b3dd9af),
	.w5(32'h3a8150e7),
	.w6(32'h3b484f63),
	.w7(32'h3a9df736),
	.w8(32'h3afa53f6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39273e88),
	.w1(32'h3ab21adb),
	.w2(32'h3bb58542),
	.w3(32'h3a9f5140),
	.w4(32'hbac51807),
	.w5(32'h3b3fce81),
	.w6(32'hba6f5c63),
	.w7(32'h3b43fb62),
	.w8(32'hbb55979f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a918ff6),
	.w1(32'hbbce045c),
	.w2(32'hbb8be90e),
	.w3(32'hba1e05dd),
	.w4(32'hbb70356c),
	.w5(32'hbaa6f975),
	.w6(32'hbbb9370f),
	.w7(32'hbb9434f9),
	.w8(32'hbba62b2d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9858d6),
	.w1(32'hbb8e8e17),
	.w2(32'hbc375c8a),
	.w3(32'hbb0217ca),
	.w4(32'hbabb97fb),
	.w5(32'hbc1529cd),
	.w6(32'hba2afcd2),
	.w7(32'hbbc74a34),
	.w8(32'hbb8f13b9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccd391),
	.w1(32'hba961949),
	.w2(32'hb94e1048),
	.w3(32'hbb9a9923),
	.w4(32'hbb33fe3e),
	.w5(32'hba61178c),
	.w6(32'hbb86316d),
	.w7(32'hbb1f82d4),
	.w8(32'hbbc1ca1e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55e994),
	.w1(32'h3a86553b),
	.w2(32'h3bb80247),
	.w3(32'hbb90ff68),
	.w4(32'h3a547841),
	.w5(32'h3b1fabd6),
	.w6(32'hba8830fa),
	.w7(32'h3b634c08),
	.w8(32'h3a88359f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393dca64),
	.w1(32'h39b832db),
	.w2(32'hbb640627),
	.w3(32'hb999ebd7),
	.w4(32'h3ab79425),
	.w5(32'hbb408a53),
	.w6(32'h3a2a0339),
	.w7(32'hbadfeabf),
	.w8(32'h397ed169),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7533),
	.w1(32'hbb5460d2),
	.w2(32'hbbb40ac0),
	.w3(32'hbb9ed91c),
	.w4(32'hbb37f438),
	.w5(32'hbb943e21),
	.w6(32'hbb4d6b6c),
	.w7(32'hbb8681d6),
	.w8(32'hbb864c47),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb523280),
	.w1(32'hbb3b6c75),
	.w2(32'h3b856240),
	.w3(32'hbaff1e3e),
	.w4(32'hbb8fe913),
	.w5(32'h3b2119d1),
	.w6(32'hbbd5fe64),
	.w7(32'h3a5b4b2e),
	.w8(32'hb9733968),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a11b8),
	.w1(32'h3b838feb),
	.w2(32'h3b443873),
	.w3(32'h3ab852c6),
	.w4(32'h3ae3c13c),
	.w5(32'h38f89b96),
	.w6(32'h3b8af9dc),
	.w7(32'h3b7657dc),
	.w8(32'h3a4390c9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0a0a5),
	.w1(32'hbb94bdb0),
	.w2(32'h3a036750),
	.w3(32'hbb500e68),
	.w4(32'hbb718137),
	.w5(32'h3b152b36),
	.w6(32'hbc0b8d00),
	.w7(32'hbb479fcc),
	.w8(32'hbbdd509b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5e895),
	.w1(32'hba89defa),
	.w2(32'hbb70e736),
	.w3(32'hbb87f549),
	.w4(32'h3b884870),
	.w5(32'h3ab4a468),
	.w6(32'h3a2f9353),
	.w7(32'h3ab69194),
	.w8(32'h3b2360de),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1d64d),
	.w1(32'hb97cbcf4),
	.w2(32'h3a42420d),
	.w3(32'h3a3f82e6),
	.w4(32'h39a03996),
	.w5(32'h3ab5026f),
	.w6(32'hbaa966f2),
	.w7(32'h3ad14bfd),
	.w8(32'h3af4f159),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03e62f),
	.w1(32'h3ae82163),
	.w2(32'h3b8e1cc2),
	.w3(32'h3ab8e435),
	.w4(32'h3aa412b0),
	.w5(32'h3b406416),
	.w6(32'h3a8cbc57),
	.w7(32'h3b0158d7),
	.w8(32'h3b12d2f6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd9d9),
	.w1(32'h3a0c6abc),
	.w2(32'hbabd2d26),
	.w3(32'h3b7e7660),
	.w4(32'h3a72ca93),
	.w5(32'hbaae666f),
	.w6(32'h3abe821f),
	.w7(32'hba1ec97b),
	.w8(32'h393cf441),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa177),
	.w1(32'h3a6da63b),
	.w2(32'h3c212a5d),
	.w3(32'hbb02472a),
	.w4(32'hbb4a2a0f),
	.w5(32'h3b91a9ec),
	.w6(32'hba5e05d1),
	.w7(32'h3ba96898),
	.w8(32'h3b6924fd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6f1de),
	.w1(32'h38b4e33d),
	.w2(32'hbb01dcf4),
	.w3(32'h3af676a2),
	.w4(32'h3a174172),
	.w5(32'hba964f79),
	.w6(32'h3a6b5f11),
	.w7(32'hbad3ea4d),
	.w8(32'h3a61e4ae),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89205f),
	.w1(32'hbb48e9a0),
	.w2(32'hbb93dda2),
	.w3(32'hbb9cb390),
	.w4(32'hbac796a1),
	.w5(32'hbb622152),
	.w6(32'h3a87c793),
	.w7(32'hba6ee554),
	.w8(32'hbb1117a0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33fbc9),
	.w1(32'h3b0b5443),
	.w2(32'h3c03d43b),
	.w3(32'h3a560c92),
	.w4(32'h3a912d56),
	.w5(32'h3bd899ac),
	.w6(32'hba15acf1),
	.w7(32'h3b938250),
	.w8(32'h3b1262e7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be322e0),
	.w1(32'h3bb8e33e),
	.w2(32'h3c3fc102),
	.w3(32'h3bd81f52),
	.w4(32'h3b6e9e61),
	.w5(32'h3c218181),
	.w6(32'h3b23aa92),
	.w7(32'h3bdc2888),
	.w8(32'h3b84ac0f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9295e4),
	.w1(32'hbb7008dc),
	.w2(32'hbbb31413),
	.w3(32'h3b675ffb),
	.w4(32'hbac4dfa8),
	.w5(32'hbb5d083f),
	.w6(32'hbb3c06c8),
	.w7(32'hbb8ce445),
	.w8(32'hbb00624a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51255b),
	.w1(32'hb98be7f2),
	.w2(32'h3b116ed2),
	.w3(32'hbaffd80f),
	.w4(32'hbb30ab15),
	.w5(32'hba9a70bc),
	.w6(32'hbaf481c4),
	.w7(32'h386fb650),
	.w8(32'hba8ca612),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c1394),
	.w1(32'hbc1a8891),
	.w2(32'hbb84d591),
	.w3(32'hbb2e61bb),
	.w4(32'hbb61b0f7),
	.w5(32'h3affd6e8),
	.w6(32'hbc7e8bdf),
	.w7(32'hbc51b755),
	.w8(32'hbc1e5370),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0834a8),
	.w1(32'hb8cd4db0),
	.w2(32'hbb2017dc),
	.w3(32'h3b7a2e07),
	.w4(32'hb8fa22db),
	.w5(32'hbb1e2f32),
	.w6(32'hb9b0cfa7),
	.w7(32'hbb0172cd),
	.w8(32'hbaff78f1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05f5b0),
	.w1(32'h3c2ea147),
	.w2(32'h3bd10eac),
	.w3(32'hbaffe969),
	.w4(32'h3c39a1e8),
	.w5(32'h3be98df4),
	.w6(32'h3c098285),
	.w7(32'h3b8eccf2),
	.w8(32'hbb06fc37),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba853),
	.w1(32'hbb078b67),
	.w2(32'h3bf3372a),
	.w3(32'hbb2553f5),
	.w4(32'hbb181352),
	.w5(32'h3bfede17),
	.w6(32'hbbd795d2),
	.w7(32'h3a29401a),
	.w8(32'hbac77201),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8c7c1),
	.w1(32'h3b96c00c),
	.w2(32'h3c107050),
	.w3(32'h3bba1051),
	.w4(32'h3b45ed44),
	.w5(32'h3baea5f5),
	.w6(32'h3ba84ffd),
	.w7(32'h3c0939ff),
	.w8(32'h3b81fb38),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0612e),
	.w1(32'h3afab229),
	.w2(32'h3b6730ce),
	.w3(32'h3a3274d8),
	.w4(32'h3b4b0f11),
	.w5(32'h3b1a2c3a),
	.w6(32'h38e21fdf),
	.w7(32'hbb359c9c),
	.w8(32'hbb30e39f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966593),
	.w1(32'hbbcf9ad4),
	.w2(32'hba4cd449),
	.w3(32'hbb6f8d1d),
	.w4(32'hbb977584),
	.w5(32'hbacf7d36),
	.w6(32'hbbff0e93),
	.w7(32'hbbac53cb),
	.w8(32'hbb4d4a40),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65ce24),
	.w1(32'hbbf06fe0),
	.w2(32'hbc7cf96e),
	.w3(32'hba2898bc),
	.w4(32'hbb86355b),
	.w5(32'hbc66bd06),
	.w6(32'hbb0bde93),
	.w7(32'hbc1ba7b1),
	.w8(32'hbbc4953f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55b860),
	.w1(32'hbb52d558),
	.w2(32'hbbabca0a),
	.w3(32'hbc0d0411),
	.w4(32'hba9ef3c6),
	.w5(32'hbb87024d),
	.w6(32'hbb07b664),
	.w7(32'hbb6c19e4),
	.w8(32'hbafd74af),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4daa20),
	.w1(32'hbb3a49b2),
	.w2(32'hbbf32e1d),
	.w3(32'hbb1d71fa),
	.w4(32'hbaaadb2e),
	.w5(32'hbbcea1b9),
	.w6(32'hba53c702),
	.w7(32'hbba517a3),
	.w8(32'hbb49c6b0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc71b3b),
	.w1(32'hb99a97af),
	.w2(32'hba92f47d),
	.w3(32'hbb993b8a),
	.w4(32'h37813399),
	.w5(32'hbab29b0d),
	.w6(32'h39554acd),
	.w7(32'hba125937),
	.w8(32'hbaaac450),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd8fc6),
	.w1(32'h3b0f85b4),
	.w2(32'h3bdd2d03),
	.w3(32'hb9a13c5b),
	.w4(32'hbac62fe1),
	.w5(32'h3b6767d5),
	.w6(32'h39d149d2),
	.w7(32'h3b7bb3bd),
	.w8(32'h3b1da148),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba441d0),
	.w1(32'h3ab08ffa),
	.w2(32'hbab912c4),
	.w3(32'h3b3372f1),
	.w4(32'h3aeb2679),
	.w5(32'hba8310da),
	.w6(32'h3b23ac25),
	.w7(32'h3a682ec8),
	.w8(32'h3aa6c124),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94a09),
	.w1(32'hbb53c1fe),
	.w2(32'hbc045caa),
	.w3(32'hba2612a3),
	.w4(32'hbae11e5f),
	.w5(32'hbbe78cfe),
	.w6(32'hba4478ad),
	.w7(32'hbbab3e61),
	.w8(32'hbb564e36),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc9d5),
	.w1(32'h3ae90a00),
	.w2(32'h3b98757b),
	.w3(32'hbb8e56a2),
	.w4(32'hb9ab0c51),
	.w5(32'h3b329b80),
	.w6(32'h3968d90d),
	.w7(32'h3b13f1fa),
	.w8(32'h3a8de21a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4525e9),
	.w1(32'h39e29b1d),
	.w2(32'hbb20d6e1),
	.w3(32'h381b9d39),
	.w4(32'hb8d538c9),
	.w5(32'hbb489f29),
	.w6(32'hb88601a5),
	.w7(32'hbb35b48b),
	.w8(32'hbb56eb83),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb3648),
	.w1(32'hbb7cb801),
	.w2(32'hbb5f06d4),
	.w3(32'hbbc7f567),
	.w4(32'hbb250abe),
	.w5(32'hbb946b20),
	.w6(32'hbbb6cfe6),
	.w7(32'hbb83043a),
	.w8(32'hbab2ac27),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2e8c5),
	.w1(32'hbb85f0e1),
	.w2(32'hbbc5eb01),
	.w3(32'hbbb95abe),
	.w4(32'hbb2d76cc),
	.w5(32'hbbb58264),
	.w6(32'hbb1b305a),
	.w7(32'hbb29f634),
	.w8(32'hbb88d4e9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1b424),
	.w1(32'hba9ea522),
	.w2(32'h3aa17805),
	.w3(32'hbc097332),
	.w4(32'hbb833f07),
	.w5(32'hbb028025),
	.w6(32'hbb1082e4),
	.w7(32'hb9fd4ac7),
	.w8(32'hbb174706),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a716335),
	.w1(32'hbb427a6c),
	.w2(32'hbb5c5e47),
	.w3(32'hbaebeeed),
	.w4(32'hbb445dd4),
	.w5(32'hbb7f3db2),
	.w6(32'hbb44de37),
	.w7(32'hbb79a68a),
	.w8(32'hbb651f66),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dc46d),
	.w1(32'hbb93a406),
	.w2(32'hbc38f7b7),
	.w3(32'hbb7d5578),
	.w4(32'hbb192d39),
	.w5(32'hbc20f767),
	.w6(32'hba8c9431),
	.w7(32'hbbf36189),
	.w8(32'hbb9723c1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c0c0),
	.w1(32'hbb8079f7),
	.w2(32'hbbe69d55),
	.w3(32'hbbc68bf7),
	.w4(32'hbb0da0ba),
	.w5(32'hbbaaf2a4),
	.w6(32'hbb604306),
	.w7(32'hbbd755bf),
	.w8(32'hbb8dbdd5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba68461),
	.w1(32'hbb08ddf4),
	.w2(32'hbbaa6b53),
	.w3(32'hbb55ce7d),
	.w4(32'hb999de2b),
	.w5(32'hbb5e7688),
	.w6(32'hba916a9c),
	.w7(32'hbb8a8dba),
	.w8(32'hbaf26d7d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb779691),
	.w1(32'hbb32c50f),
	.w2(32'hbb21962a),
	.w3(32'hbab71272),
	.w4(32'hb9d3e27b),
	.w5(32'hbb3a4185),
	.w6(32'hbb16983a),
	.w7(32'hba61da05),
	.w8(32'hba8caf3b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2975c6),
	.w1(32'hba5bfed1),
	.w2(32'h3ae40bba),
	.w3(32'hbb522e17),
	.w4(32'hbaadc7b6),
	.w5(32'hb8d68bd1),
	.w6(32'hbb1cb316),
	.w7(32'hbace50cf),
	.w8(32'hbb91904e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9bb6),
	.w1(32'h3b32672e),
	.w2(32'h3b8736d0),
	.w3(32'hbb79ec17),
	.w4(32'h3b0ad2ee),
	.w5(32'h3b2f815c),
	.w6(32'h3b377119),
	.w7(32'h3b7173de),
	.w8(32'h3b8e3e7e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7f4c9),
	.w1(32'h3b014753),
	.w2(32'h3af5413d),
	.w3(32'h3b9c93bf),
	.w4(32'h3ae54fb2),
	.w5(32'h3ad90773),
	.w6(32'h3a230d34),
	.w7(32'hb9bc3c97),
	.w8(32'hbb057c8c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9749870),
	.w1(32'hbbf4137f),
	.w2(32'hbc2fbe73),
	.w3(32'hb9b10273),
	.w4(32'hbbc2ef8f),
	.w5(32'hbc1e8a02),
	.w6(32'hbbd9f49a),
	.w7(32'hbc207d8e),
	.w8(32'hbc0d450b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2303e6),
	.w1(32'hbb8400f6),
	.w2(32'hba2ce9e0),
	.w3(32'hbc115c33),
	.w4(32'h3959102d),
	.w5(32'h3a6c097e),
	.w6(32'hbc00baa0),
	.w7(32'hbbd4d553),
	.w8(32'hbbe01194),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbb90a),
	.w1(32'hbadfa7ab),
	.w2(32'h3b5ed6b4),
	.w3(32'h3adb9d9c),
	.w4(32'hbacb2c5d),
	.w5(32'h3b691573),
	.w6(32'hbb8c2767),
	.w7(32'hba56e35f),
	.w8(32'h39f1f6fe),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9bb8),
	.w1(32'h3aa355e6),
	.w2(32'hbb2d068c),
	.w3(32'h3b8b9ae5),
	.w4(32'h3b0098b4),
	.w5(32'hbb143277),
	.w6(32'h3b8adbd2),
	.w7(32'hb956c725),
	.w8(32'hb99fda80),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f9573),
	.w1(32'h389cb356),
	.w2(32'h37fb1749),
	.w3(32'h3ab4af94),
	.w4(32'h3877e0a8),
	.w5(32'h38b585db),
	.w6(32'h37dceaae),
	.w7(32'h3787d4a4),
	.w8(32'h3892ca48),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b4cbb),
	.w1(32'hbb53a426),
	.w2(32'hbb304dd8),
	.w3(32'hbb2ce73e),
	.w4(32'hbaa6f263),
	.w5(32'h364fb5c6),
	.w6(32'h3abed865),
	.w7(32'h3aa8edd3),
	.w8(32'h3a2e7612),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule