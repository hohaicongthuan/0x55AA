module layer_10_featuremap_396(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bdc52),
	.w1(32'h3aa9fc19),
	.w2(32'h3ab6d827),
	.w3(32'hbbfd499c),
	.w4(32'hbb2725a9),
	.w5(32'hbbac3ea6),
	.w6(32'hbbda1c5c),
	.w7(32'h3bcf6e59),
	.w8(32'hb9584174),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0305b),
	.w1(32'h3b02519e),
	.w2(32'h3c1c0680),
	.w3(32'h39ec7ff7),
	.w4(32'h3bc130b6),
	.w5(32'h3b6e0c2c),
	.w6(32'h3b3d2b41),
	.w7(32'h3a876d3b),
	.w8(32'h3bf45508),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393722a8),
	.w1(32'hbbbb4d6b),
	.w2(32'hbb521897),
	.w3(32'h3b6262b6),
	.w4(32'hbb876a59),
	.w5(32'h3b95fca2),
	.w6(32'hb99e9228),
	.w7(32'h3befe33a),
	.w8(32'h3af0c37e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd2b38),
	.w1(32'hbc01a4f9),
	.w2(32'hbb27c29b),
	.w3(32'hbba4f2e2),
	.w4(32'hbbbb8005),
	.w5(32'h3a4d0fe0),
	.w6(32'hbaf2bcbe),
	.w7(32'hbbd45fc5),
	.w8(32'hbb858ffe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c61e),
	.w1(32'h3b841073),
	.w2(32'hbb6dc836),
	.w3(32'hbb5b77d9),
	.w4(32'h3b8232a5),
	.w5(32'h3c108c1b),
	.w6(32'hba961207),
	.w7(32'h38cbb7ab),
	.w8(32'hbad6762a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e98cb),
	.w1(32'h3bdfea46),
	.w2(32'h3c5532e7),
	.w3(32'hba6c8e85),
	.w4(32'h3b191e99),
	.w5(32'h3c8471f7),
	.w6(32'h3a698741),
	.w7(32'h3ad976b6),
	.w8(32'hbb354b32),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc44334),
	.w1(32'h3a1a7c34),
	.w2(32'h3b45f657),
	.w3(32'h3c26cab9),
	.w4(32'h3c1eb87a),
	.w5(32'h3c09b00c),
	.w6(32'h3bbc44a0),
	.w7(32'hbc1abb0e),
	.w8(32'hbbc4317d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9c01),
	.w1(32'hbbc5ad46),
	.w2(32'hbc11eeb1),
	.w3(32'hbc2232ad),
	.w4(32'hbc50012b),
	.w5(32'hbb797aac),
	.w6(32'hbc92a8e8),
	.w7(32'hbc0882ce),
	.w8(32'hbb32f157),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0be426),
	.w1(32'h3b0d0579),
	.w2(32'hba11ef7f),
	.w3(32'hbaef6288),
	.w4(32'h3a013d54),
	.w5(32'hbb7106fa),
	.w6(32'hba8a460c),
	.w7(32'h3b32efe1),
	.w8(32'hbba01c60),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5e0e8),
	.w1(32'h3b3068a7),
	.w2(32'h3c240a1b),
	.w3(32'h3b39657b),
	.w4(32'h3b3161be),
	.w5(32'h3beb6a1e),
	.w6(32'hbbac9ec4),
	.w7(32'hbbed8131),
	.w8(32'hbba31d7b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ffd7a),
	.w1(32'hb8c682d5),
	.w2(32'h3ba62367),
	.w3(32'hbb6a5e99),
	.w4(32'h3a8f1f3e),
	.w5(32'h3b8b1ef6),
	.w6(32'h3b69224a),
	.w7(32'h3b754547),
	.w8(32'h3ba53ecd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a866f40),
	.w1(32'hbc068313),
	.w2(32'hbc1bbcad),
	.w3(32'h3c244de8),
	.w4(32'hbb58d3b8),
	.w5(32'hbadeeeb0),
	.w6(32'h3c183cc3),
	.w7(32'hbb873e21),
	.w8(32'h399615cf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847b52),
	.w1(32'hbb6e17f3),
	.w2(32'h3a9cbc51),
	.w3(32'h3b8c7852),
	.w4(32'hba673800),
	.w5(32'hbbc31c6a),
	.w6(32'h3b207bc8),
	.w7(32'hbb37367e),
	.w8(32'h3ad22e7f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb646ff5),
	.w1(32'h3b0295cc),
	.w2(32'h3a642217),
	.w3(32'h3b9159af),
	.w4(32'h3aed6463),
	.w5(32'h3becf363),
	.w6(32'h3b1f40fc),
	.w7(32'hba903796),
	.w8(32'hb94f9b5f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86024c),
	.w1(32'h3b876531),
	.w2(32'h3c1fdd3f),
	.w3(32'h3c08c76e),
	.w4(32'hbafa2b9c),
	.w5(32'h3c5954a7),
	.w6(32'h3ab1d294),
	.w7(32'h3abfe58b),
	.w8(32'h3ba857f6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52bd68),
	.w1(32'hbc013f68),
	.w2(32'h3b2cbbc0),
	.w3(32'h3c339f76),
	.w4(32'hbbb8a8db),
	.w5(32'hbb2159fb),
	.w6(32'h3bd62278),
	.w7(32'hbbc8de69),
	.w8(32'hbbb1ccf8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fed13),
	.w1(32'hbba77f7d),
	.w2(32'hbb09da3b),
	.w3(32'h3c13737d),
	.w4(32'hbb340f1a),
	.w5(32'hbc2a5546),
	.w6(32'h3abab6f3),
	.w7(32'hb890b344),
	.w8(32'hbabbd914),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119a8c),
	.w1(32'hbc722858),
	.w2(32'hbc964e76),
	.w3(32'hbcbbc4ac),
	.w4(32'hbcbc35a0),
	.w5(32'hbc9e4312),
	.w6(32'hbcaf6d7f),
	.w7(32'hbc9f93a4),
	.w8(32'hbca11245),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff8023),
	.w1(32'hbbb274b2),
	.w2(32'hbbbc0f87),
	.w3(32'hbc6d9715),
	.w4(32'hbb96cfe9),
	.w5(32'h3a3f5782),
	.w6(32'hbc921118),
	.w7(32'hbbcd78c2),
	.w8(32'hbb24d3ec),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac98785),
	.w1(32'h3c4a7ab1),
	.w2(32'h3bf1f60d),
	.w3(32'h3b606fbf),
	.w4(32'h3b20d21d),
	.w5(32'hbc1ccaa4),
	.w6(32'h3b66965f),
	.w7(32'h3c4f7cc1),
	.w8(32'hbb318a04),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21fb29),
	.w1(32'hbbcebbdf),
	.w2(32'hbbbca484),
	.w3(32'h3c261886),
	.w4(32'hbb61c95c),
	.w5(32'h3a44083a),
	.w6(32'hbb320408),
	.w7(32'hb9a439c4),
	.w8(32'h37e65335),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bd77c),
	.w1(32'hbb79e23b),
	.w2(32'h39a559c9),
	.w3(32'h3aa31bd0),
	.w4(32'hbb5a0836),
	.w5(32'hbbe9fea9),
	.w6(32'h3bc87e15),
	.w7(32'h3b026c7c),
	.w8(32'h3a7e4a49),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2517),
	.w1(32'hbcbd0170),
	.w2(32'hbcfb7a31),
	.w3(32'hbcfd33cf),
	.w4(32'hbc78c2be),
	.w5(32'hbc2d1dd3),
	.w6(32'hbd02247b),
	.w7(32'hbc90b37a),
	.w8(32'hbc6e5fb4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41a4d1),
	.w1(32'h3ba16f6c),
	.w2(32'h3b7238a7),
	.w3(32'h3b9bfe80),
	.w4(32'h3b970d7f),
	.w5(32'h3bac338d),
	.w6(32'h3bc25730),
	.w7(32'hbb9be3e9),
	.w8(32'hbc15d223),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acba8),
	.w1(32'h3c10ac67),
	.w2(32'h3ad0a4c7),
	.w3(32'hbb1c37c2),
	.w4(32'h3c24d4dc),
	.w5(32'hbb263faf),
	.w6(32'hbbf1cd78),
	.w7(32'h3b802874),
	.w8(32'hbbcf524b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5189a),
	.w1(32'hbb80f232),
	.w2(32'h3bbbc7b2),
	.w3(32'hbbd2e0a7),
	.w4(32'hbbb108f8),
	.w5(32'h3b1eeeb6),
	.w6(32'hbc0ca6e6),
	.w7(32'hbab33815),
	.w8(32'h3b85e83d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d2900),
	.w1(32'hbba57992),
	.w2(32'hb9334ea4),
	.w3(32'hbb4926f4),
	.w4(32'h3a95d9bf),
	.w5(32'hb9e2e72d),
	.w6(32'h3a858746),
	.w7(32'hbabd3964),
	.w8(32'hb986ecb5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b6c33),
	.w1(32'h3b9857c6),
	.w2(32'h3baf4aca),
	.w3(32'h3b7cfc0d),
	.w4(32'h3b11e00f),
	.w5(32'hbb41c5cd),
	.w6(32'h3bfb0215),
	.w7(32'h394e3145),
	.w8(32'hbb578de6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf687c3),
	.w1(32'hbc3ddb28),
	.w2(32'hbba1e76a),
	.w3(32'hbbf20ac0),
	.w4(32'h3b63d3d7),
	.w5(32'hbb42dde7),
	.w6(32'hbbfcfdd4),
	.w7(32'hba576686),
	.w8(32'h396fff6a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b714e5a),
	.w1(32'hba3f49ab),
	.w2(32'hbb5ff39e),
	.w3(32'h3b2196e6),
	.w4(32'h3bbebd0c),
	.w5(32'h3c20f86b),
	.w6(32'h3c24e4de),
	.w7(32'hba421291),
	.w8(32'h3be8657c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe007d),
	.w1(32'h3bedee67),
	.w2(32'h3cb69303),
	.w3(32'h3a075981),
	.w4(32'hbab7b828),
	.w5(32'hbc00b107),
	.w6(32'h3b2ba96f),
	.w7(32'h3ab8035c),
	.w8(32'hbacb0192),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf37c0),
	.w1(32'hbbafe9e4),
	.w2(32'hbb3277b5),
	.w3(32'hbbcb186c),
	.w4(32'hbb0a003a),
	.w5(32'h3af8a5f6),
	.w6(32'hba61e434),
	.w7(32'hbb4d8d97),
	.w8(32'h3bb54c98),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad38925),
	.w1(32'hba9a21b3),
	.w2(32'h3b2faca5),
	.w3(32'h3b66a0bf),
	.w4(32'h3b6fdaf6),
	.w5(32'hba966ac5),
	.w6(32'h37a9ffdb),
	.w7(32'h3c342c20),
	.w8(32'h3c288e0b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074d38),
	.w1(32'h3b7d1619),
	.w2(32'h3b189617),
	.w3(32'hbaf66bf4),
	.w4(32'h3b2b80be),
	.w5(32'h3b4622ab),
	.w6(32'h3bcee8d3),
	.w7(32'hbb293b22),
	.w8(32'h3ac0736f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b0d57),
	.w1(32'hba53ae13),
	.w2(32'hbb2973cd),
	.w3(32'h3b26bca1),
	.w4(32'hbbb4008b),
	.w5(32'hbc368f69),
	.w6(32'h3bc5ef9f),
	.w7(32'hbb8f40ca),
	.w8(32'hb9ce150b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cf45e),
	.w1(32'h3c0cd968),
	.w2(32'h3b47751a),
	.w3(32'hbb6a907c),
	.w4(32'h3b4ea7b8),
	.w5(32'hba0190c5),
	.w6(32'hbbc3b251),
	.w7(32'hbb111511),
	.w8(32'h38c67ad6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91d058),
	.w1(32'hbb5e35ad),
	.w2(32'h39d5b6dd),
	.w3(32'hbbc23cab),
	.w4(32'hbb0ac3d4),
	.w5(32'h3c04290d),
	.w6(32'hbc1f346d),
	.w7(32'hbb9d638c),
	.w8(32'hbbb8e460),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3d24),
	.w1(32'h3c0eebfd),
	.w2(32'h3c751b56),
	.w3(32'h3ca60ee9),
	.w4(32'h3c370ad6),
	.w5(32'h3b07f2d2),
	.w6(32'h3c792426),
	.w7(32'h3b80b031),
	.w8(32'h3bc1c070),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fab0e5),
	.w1(32'h3c57a8a8),
	.w2(32'h3c08077d),
	.w3(32'h3c8ad188),
	.w4(32'h3c0ae4ce),
	.w5(32'hba1d689a),
	.w6(32'h3c33b8a2),
	.w7(32'h3c4a8cc2),
	.w8(32'hba0f9d3a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952e51),
	.w1(32'hba6214fc),
	.w2(32'h3aeb8ca9),
	.w3(32'h3a936bd9),
	.w4(32'hba917bf7),
	.w5(32'h3a0ff109),
	.w6(32'hbb79c412),
	.w7(32'h3ab2338f),
	.w8(32'h3a75bf1e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998b877),
	.w1(32'h3b87ed99),
	.w2(32'h3ba1b2aa),
	.w3(32'hbbb6f589),
	.w4(32'h3b383625),
	.w5(32'h3c1b12c8),
	.w6(32'hbb7d224a),
	.w7(32'h3b37f056),
	.w8(32'h3b893379),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b764a76),
	.w1(32'hbaf87ffd),
	.w2(32'h3b811d50),
	.w3(32'h3c1fc6ff),
	.w4(32'hbba9470d),
	.w5(32'h3b6437ff),
	.w6(32'h3b42ed9c),
	.w7(32'hba1d342b),
	.w8(32'hbb5103db),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae472c5),
	.w1(32'hbb26433e),
	.w2(32'hbb1c24d0),
	.w3(32'h3b50db26),
	.w4(32'h3bc36ab4),
	.w5(32'hbb865b58),
	.w6(32'hbb604397),
	.w7(32'h399077a6),
	.w8(32'h3b5073c0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98ca9e),
	.w1(32'hb8e41015),
	.w2(32'hbb47b676),
	.w3(32'hbbbc35a1),
	.w4(32'hba6c4080),
	.w5(32'hbbe06ef3),
	.w6(32'hbc086ee7),
	.w7(32'hba27f713),
	.w8(32'hbb7161b0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d839),
	.w1(32'h3b93fec5),
	.w2(32'h3b6b7ec5),
	.w3(32'hbb959398),
	.w4(32'hba79e07f),
	.w5(32'hbb6b1566),
	.w6(32'hbb61a0c2),
	.w7(32'hba8cdde5),
	.w8(32'hbbaef8d6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974a9e),
	.w1(32'hbaf44e25),
	.w2(32'h3b23b44a),
	.w3(32'hbb636dfa),
	.w4(32'hb8ae1210),
	.w5(32'h3a52a9a7),
	.w6(32'hbba9fd9b),
	.w7(32'hbaeae5a3),
	.w8(32'h3ad47c0a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42f2d5),
	.w1(32'hbb935a6b),
	.w2(32'hba1d9a33),
	.w3(32'h39c167b0),
	.w4(32'hbb334136),
	.w5(32'h3b322c39),
	.w6(32'hbb1ec292),
	.w7(32'hbba652f1),
	.w8(32'h398aa1e3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272dfd),
	.w1(32'hbca108eb),
	.w2(32'hbce2937a),
	.w3(32'hbca3bdf0),
	.w4(32'hbc8c7c96),
	.w5(32'hbc3c81bd),
	.w6(32'hbcb40122),
	.w7(32'hbc34e8e9),
	.w8(32'hbbe6241b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8326d),
	.w1(32'hbb4150fa),
	.w2(32'hbb4f59b8),
	.w3(32'h3a035407),
	.w4(32'hb8a5c304),
	.w5(32'h392e3549),
	.w6(32'hba392e39),
	.w7(32'h37835958),
	.w8(32'hb8c4ba04),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fa2c0),
	.w1(32'hbafcaaca),
	.w2(32'hbb264b33),
	.w3(32'h3af34a94),
	.w4(32'hbbe468b2),
	.w5(32'hbb89c790),
	.w6(32'h3addf5a9),
	.w7(32'hbbe89f60),
	.w8(32'hbb31efaa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b741554),
	.w1(32'h3a9f50a2),
	.w2(32'h3b010dc6),
	.w3(32'h3a979eec),
	.w4(32'hbb07db63),
	.w5(32'hbb265015),
	.w6(32'hbab1b453),
	.w7(32'h3c2a6426),
	.w8(32'hbb8471c1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a4efe),
	.w1(32'h3b506004),
	.w2(32'h3bb1df7a),
	.w3(32'hbb695319),
	.w4(32'h3c3d8a28),
	.w5(32'h3af3058a),
	.w6(32'hbb844f20),
	.w7(32'hb92ca3af),
	.w8(32'h3c2d59de),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480fc6),
	.w1(32'h3b2ccba4),
	.w2(32'h3ba1cd9b),
	.w3(32'h3b994f5e),
	.w4(32'h3ac8d93e),
	.w5(32'h3ba16550),
	.w6(32'hb98c15e8),
	.w7(32'hba83ee3b),
	.w8(32'h3a309157),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb553c44),
	.w1(32'hbc876ecf),
	.w2(32'hbcade457),
	.w3(32'hbc2f9b3a),
	.w4(32'hbc69cd16),
	.w5(32'hbc2e70e6),
	.w6(32'hbc0c4c7b),
	.w7(32'hbc061a87),
	.w8(32'hba0dd966),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167b69),
	.w1(32'hbb8db581),
	.w2(32'hbb5ae86a),
	.w3(32'hbb5bc122),
	.w4(32'h3a942c4c),
	.w5(32'hbbf65eec),
	.w6(32'hb90ad181),
	.w7(32'h3baba20a),
	.w8(32'h3b099b97),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba914d85),
	.w1(32'hbbccd3c7),
	.w2(32'h3ab8865b),
	.w3(32'hbb7a97a0),
	.w4(32'hbc09e1d6),
	.w5(32'hbb2c88cf),
	.w6(32'hbb97cce6),
	.w7(32'hbb2bb935),
	.w8(32'hb9aca29d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982d7a),
	.w1(32'h3a662519),
	.w2(32'hbb32177f),
	.w3(32'h3bbb7f88),
	.w4(32'h3bd525aa),
	.w5(32'h3c01fc64),
	.w6(32'hbb904bb0),
	.w7(32'hb9946e1b),
	.w8(32'h3b80e1f3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a346d),
	.w1(32'h39247a0b),
	.w2(32'h3b67c4d5),
	.w3(32'h3bced164),
	.w4(32'hbbb82216),
	.w5(32'h3c968612),
	.w6(32'h3b34abb3),
	.w7(32'hbb1449ad),
	.w8(32'h3bac5bf1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9002),
	.w1(32'h3b393108),
	.w2(32'hbaf7e03e),
	.w3(32'h3ac5c48e),
	.w4(32'h3b8cf204),
	.w5(32'hbc0852e3),
	.w6(32'h3c53a2e5),
	.w7(32'h3c56e9e3),
	.w8(32'hbb1211e4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb2b6),
	.w1(32'h3bfcc4a6),
	.w2(32'hbbb70131),
	.w3(32'h39c2ce79),
	.w4(32'h3c1f9726),
	.w5(32'h3b97c227),
	.w6(32'hbb92e677),
	.w7(32'h3ba46eb6),
	.w8(32'h3a679801),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6123a),
	.w1(32'hbbd4ed31),
	.w2(32'hbc27cf8c),
	.w3(32'hbb2d48b9),
	.w4(32'hbbd1136e),
	.w5(32'hbb8b1557),
	.w6(32'hba80277a),
	.w7(32'h3ab9512e),
	.w8(32'hba90e80e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0935a2),
	.w1(32'hbc1f8508),
	.w2(32'hbc1d9233),
	.w3(32'hbc499f6b),
	.w4(32'hbc37984d),
	.w5(32'hbb9e888c),
	.w6(32'hbc406128),
	.w7(32'hbb702608),
	.w8(32'hbb0fb504),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355ed465),
	.w1(32'h3a639c34),
	.w2(32'hbad82c07),
	.w3(32'hbbdc1453),
	.w4(32'h3b00dc0f),
	.w5(32'hbb792ef6),
	.w6(32'h3a8f3677),
	.w7(32'hbb9b24f6),
	.w8(32'hbbbe2636),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db0db),
	.w1(32'h3a819f9d),
	.w2(32'hbb52f40f),
	.w3(32'hbbcdde43),
	.w4(32'hbb3e5218),
	.w5(32'hbb72a15e),
	.w6(32'hbbc27813),
	.w7(32'h3b840d63),
	.w8(32'h396afd48),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb39f),
	.w1(32'h3b16937d),
	.w2(32'hb9e8c207),
	.w3(32'h392d6708),
	.w4(32'h3959c997),
	.w5(32'hb92c782f),
	.w6(32'h3a1e45e6),
	.w7(32'h3966b2f2),
	.w8(32'h3aff0622),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8e0e),
	.w1(32'h3ab45fc2),
	.w2(32'h3b67b86e),
	.w3(32'h3b813424),
	.w4(32'hba9cb306),
	.w5(32'hbb600d1f),
	.w6(32'h3af519f2),
	.w7(32'hba699979),
	.w8(32'hbbbd97ad),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2414),
	.w1(32'hbb977ebd),
	.w2(32'hbb9cad04),
	.w3(32'h3a86136c),
	.w4(32'hbb0d0f0b),
	.w5(32'hbaa493d5),
	.w6(32'hbbe4c50c),
	.w7(32'h3afdc8f8),
	.w8(32'h3ad3111d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98c984),
	.w1(32'h3bd44aa9),
	.w2(32'h3c4eceab),
	.w3(32'hbb704b54),
	.w4(32'h3c063bfd),
	.w5(32'h3c5a5257),
	.w6(32'hb90f0775),
	.w7(32'h3b3eb316),
	.w8(32'h3c8c7932),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5046e3),
	.w1(32'hbc87ddb9),
	.w2(32'hbc33722a),
	.w3(32'hbc467c25),
	.w4(32'hbba68d45),
	.w5(32'hbb5f73ae),
	.w6(32'hbc053997),
	.w7(32'h3adf6e6b),
	.w8(32'hbc221b97),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fa2ff),
	.w1(32'h3c09e8f7),
	.w2(32'h3c403161),
	.w3(32'h3c1be359),
	.w4(32'h3bcdf416),
	.w5(32'h3af2543c),
	.w6(32'h3c1492a0),
	.w7(32'hbaaf1354),
	.w8(32'h3ad09f85),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a43e2),
	.w1(32'h3b563afd),
	.w2(32'hbba8a27d),
	.w3(32'hbb4a1070),
	.w4(32'hb81d236d),
	.w5(32'h3bb0a06e),
	.w6(32'h3aab68a8),
	.w7(32'h3907401a),
	.w8(32'h3bf49900),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dd546),
	.w1(32'hbb2b7a3b),
	.w2(32'h3b6aee7a),
	.w3(32'h3b1b7bd2),
	.w4(32'h3c0d4f24),
	.w5(32'h3caa32ad),
	.w6(32'h3bed3eea),
	.w7(32'hbbbb7dbe),
	.w8(32'hbbc1fa90),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad520a7),
	.w1(32'h3b72e8f9),
	.w2(32'h3b8136cf),
	.w3(32'h3b0fe2fe),
	.w4(32'hbb5f2e31),
	.w5(32'hba978ff5),
	.w6(32'hbc5e1fb9),
	.w7(32'hbc2b4f06),
	.w8(32'hbc05e7e3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ced37),
	.w1(32'hbb212c7d),
	.w2(32'hbc0dce00),
	.w3(32'h37e22805),
	.w4(32'hbc16e47c),
	.w5(32'hbbc65b76),
	.w6(32'hbba4e127),
	.w7(32'hbbd98e89),
	.w8(32'hbbf99a80),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebd400),
	.w1(32'hbba0133c),
	.w2(32'hbc21d25c),
	.w3(32'hbbf8fb4d),
	.w4(32'hbbd14a7e),
	.w5(32'hbcb19337),
	.w6(32'hbba2c8c8),
	.w7(32'hbc33ff7d),
	.w8(32'hbc87d9fc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88b7ce),
	.w1(32'hbc5afc30),
	.w2(32'hbc5ca405),
	.w3(32'hbccc1433),
	.w4(32'hbc8142ff),
	.w5(32'hbc09df94),
	.w6(32'hbc822bd1),
	.w7(32'hbc4f8499),
	.w8(32'hbc1b019d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a1118),
	.w1(32'hbc1cdf7f),
	.w2(32'hbbca8d9a),
	.w3(32'hbc6ecdc6),
	.w4(32'hbc90fb4b),
	.w5(32'hbc26b57a),
	.w6(32'hbcc9ed3a),
	.w7(32'hbc75e34b),
	.w8(32'hbc28a72e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa10a8a),
	.w1(32'h3b1b3e9e),
	.w2(32'h3ba05c3c),
	.w3(32'h3b2c0e0e),
	.w4(32'h3ab7e05e),
	.w5(32'h3b619dff),
	.w6(32'h3b37752d),
	.w7(32'h3c24689a),
	.w8(32'h3c3271dc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a740a),
	.w1(32'hb90ffdcb),
	.w2(32'hbb5621ca),
	.w3(32'hbb7a768a),
	.w4(32'hbb5d026c),
	.w5(32'hbbaa0547),
	.w6(32'h3ae28d7b),
	.w7(32'hbaa1673b),
	.w8(32'hbba66fcc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68aece),
	.w1(32'hbaa9118a),
	.w2(32'h3be1967b),
	.w3(32'hbaf4bbb6),
	.w4(32'hbb0f087e),
	.w5(32'h3b85a402),
	.w6(32'h39d32efb),
	.w7(32'hbab09fd5),
	.w8(32'h3b2ff1da),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a7392),
	.w1(32'h3c3a1e5b),
	.w2(32'h3c37714a),
	.w3(32'h3aba31d1),
	.w4(32'h3b984b15),
	.w5(32'h399c8d2c),
	.w6(32'hbb563e03),
	.w7(32'hbb2bbb45),
	.w8(32'hbc42674c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0682ad),
	.w1(32'hbc3b6eb3),
	.w2(32'hbc2d4762),
	.w3(32'hbbb926ef),
	.w4(32'hbc194ac0),
	.w5(32'hbbc8aa58),
	.w6(32'hbc5dcbd3),
	.w7(32'hbc28b5ac),
	.w8(32'hbb45cadc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b2cb),
	.w1(32'h3baaec78),
	.w2(32'h3ba4592f),
	.w3(32'hbb285405),
	.w4(32'h3c321bfb),
	.w5(32'h3c8ec945),
	.w6(32'hb9eb8bc8),
	.w7(32'h3b8c3640),
	.w8(32'h3b940863),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e31c6),
	.w1(32'h3b665ee6),
	.w2(32'hba88b49c),
	.w3(32'h3b769841),
	.w4(32'hbb20b898),
	.w5(32'h38bacee9),
	.w6(32'hb7d2a24d),
	.w7(32'hb9941790),
	.w8(32'hbbdaac76),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29db67),
	.w1(32'h3b4f621e),
	.w2(32'hbc274d65),
	.w3(32'hbbf3bac3),
	.w4(32'h3bcb6a2d),
	.w5(32'hbb631446),
	.w6(32'hbb5b4f03),
	.w7(32'hbb9cddb6),
	.w8(32'hbc00792d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0cd8a),
	.w1(32'hba8ac0c6),
	.w2(32'hbb21ca98),
	.w3(32'h3b3b0537),
	.w4(32'hbbc7e6af),
	.w5(32'h3b2a2f18),
	.w6(32'hbba6bed4),
	.w7(32'h3c0e84a6),
	.w8(32'h3b301ff4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba973152),
	.w1(32'h39aa63d7),
	.w2(32'hba3dda52),
	.w3(32'h3ba991f3),
	.w4(32'hba87ab01),
	.w5(32'hbba7861d),
	.w6(32'h3c34fea8),
	.w7(32'h3bcec669),
	.w8(32'hbb632f5a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e82b4),
	.w1(32'h3b8714be),
	.w2(32'hbaa5a447),
	.w3(32'h3ad06fcc),
	.w4(32'h3b9e56f4),
	.w5(32'h3bd61c2d),
	.w6(32'hbb7870ec),
	.w7(32'h3b2b33a1),
	.w8(32'hbbc66576),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99971e0),
	.w1(32'h398e07ec),
	.w2(32'h3881d73d),
	.w3(32'h392ca4f4),
	.w4(32'h3aa7cf41),
	.w5(32'hbb2b6292),
	.w6(32'hbbaf7be6),
	.w7(32'hbbd7b429),
	.w8(32'hbb383ccb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77c60d),
	.w1(32'hbca231fd),
	.w2(32'hbca0aba6),
	.w3(32'hbcc1d632),
	.w4(32'hbc4e92ca),
	.w5(32'hbbb11df7),
	.w6(32'hbcd8ee5b),
	.w7(32'hbbf59926),
	.w8(32'hbc18f597),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b25898),
	.w1(32'h3ba1250c),
	.w2(32'hb9d2a41e),
	.w3(32'h3bcdffc8),
	.w4(32'h3b326eec),
	.w5(32'h397705f4),
	.w6(32'h3afa35fd),
	.w7(32'h3a8f3cc6),
	.w8(32'h3af4b8d4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41064f),
	.w1(32'hbb65edc2),
	.w2(32'hbc3f84df),
	.w3(32'hbaf876e3),
	.w4(32'h3b4a9280),
	.w5(32'hbbf2277b),
	.w6(32'h3ba38921),
	.w7(32'hba951de4),
	.w8(32'hbbd8f288),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a508258),
	.w1(32'h3c81e13b),
	.w2(32'h3c0702a6),
	.w3(32'h3a063d09),
	.w4(32'h3c51d419),
	.w5(32'h3c294570),
	.w6(32'h3baa389d),
	.w7(32'h3b815171),
	.w8(32'hb9121cfe),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9822f),
	.w1(32'hbbc0faf5),
	.w2(32'hbc8a6690),
	.w3(32'h3b02e939),
	.w4(32'hbc89e2da),
	.w5(32'hbcbab4e8),
	.w6(32'hbb78761a),
	.w7(32'hbc6e4465),
	.w8(32'hbc8852ed),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc487ed7),
	.w1(32'hb960d894),
	.w2(32'hba65e2bb),
	.w3(32'hbc7c2698),
	.w4(32'h3b9a875b),
	.w5(32'h3b3fd266),
	.w6(32'hbb98817c),
	.w7(32'hbb4961e7),
	.w8(32'hbc2f4525),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990f2cc),
	.w1(32'h3a77b992),
	.w2(32'hbba22df6),
	.w3(32'h3b6a5766),
	.w4(32'h3a4c5552),
	.w5(32'h3b07f36a),
	.w6(32'hbb6c8da0),
	.w7(32'h3ad41d7c),
	.w8(32'h3c2277ad),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa63704),
	.w1(32'h3bacb2a0),
	.w2(32'hbb7c4ae0),
	.w3(32'h3b763e4f),
	.w4(32'hbabdfac6),
	.w5(32'hbb27a323),
	.w6(32'h3c051adb),
	.w7(32'hbbb195d2),
	.w8(32'hbc04108e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d381c),
	.w1(32'h3ada3ef0),
	.w2(32'h3b96210e),
	.w3(32'hbc050df5),
	.w4(32'h3b51738a),
	.w5(32'h3b1799c5),
	.w6(32'hbc4c706b),
	.w7(32'hba8081f7),
	.w8(32'hbc0c5170),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b606968),
	.w1(32'hbb915cb3),
	.w2(32'hba337408),
	.w3(32'hbb6df8cc),
	.w4(32'h3b95ee69),
	.w5(32'hbb7a8037),
	.w6(32'hbc732463),
	.w7(32'h3c1cf9ba),
	.w8(32'h3a3cee14),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc017b8c),
	.w1(32'hbc51b2ce),
	.w2(32'hbc4c1ae4),
	.w3(32'hbca2b235),
	.w4(32'hbc5cf584),
	.w5(32'hbc0cf70f),
	.w6(32'hbc5a1f0f),
	.w7(32'hbc8468fa),
	.w8(32'hbbe36e35),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2af2f),
	.w1(32'h3bf78fb7),
	.w2(32'hbbac9a4e),
	.w3(32'h3c831c64),
	.w4(32'h3b9c8b05),
	.w5(32'h3ae907c9),
	.w6(32'h3c80eeb9),
	.w7(32'h3b800810),
	.w8(32'hbc0f0e06),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8a660),
	.w1(32'h3b7cdc5a),
	.w2(32'h3bb6bce0),
	.w3(32'hbb392f84),
	.w4(32'h3b86bcab),
	.w5(32'h39d88076),
	.w6(32'hbb8826d1),
	.w7(32'hbb02e6d8),
	.w8(32'hb9895a90),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba552ee8),
	.w1(32'hbc2e9098),
	.w2(32'hbc8bb9c0),
	.w3(32'hbb0b68ab),
	.w4(32'hbb74d4c5),
	.w5(32'h3cb0d86c),
	.w6(32'hbbb0e6a2),
	.w7(32'hbb8e8217),
	.w8(32'hbc055dd3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103667),
	.w1(32'hbbb83c0a),
	.w2(32'hbca31a9c),
	.w3(32'h3c378edc),
	.w4(32'h3a438374),
	.w5(32'hbc1d5c4d),
	.w6(32'hbb2936b2),
	.w7(32'hbb852927),
	.w8(32'hbc636458),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2eabc),
	.w1(32'hbc8f30c4),
	.w2(32'hbcf495e1),
	.w3(32'hbcb4bece),
	.w4(32'hbc9be826),
	.w5(32'hbbe221fa),
	.w6(32'hbcc3d853),
	.w7(32'hbccd8217),
	.w8(32'hbcb1f41c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38280d5f),
	.w1(32'h3b93b068),
	.w2(32'h3b32a305),
	.w3(32'h3b41f41d),
	.w4(32'h396d9244),
	.w5(32'hbbd62acb),
	.w6(32'h3b6de180),
	.w7(32'h3b3c8c57),
	.w8(32'hb93096b7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6367b0),
	.w1(32'h3b4d1f73),
	.w2(32'h3ba4043b),
	.w3(32'h3aaec279),
	.w4(32'hbaadad50),
	.w5(32'hbb759233),
	.w6(32'hbadb6359),
	.w7(32'h3b3c5af5),
	.w8(32'h3b4bff47),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b3be7),
	.w1(32'h3b698515),
	.w2(32'hbb58e390),
	.w3(32'hbb616dac),
	.w4(32'h3b09dc7e),
	.w5(32'h3b77cbe7),
	.w6(32'h3bd02cce),
	.w7(32'hbc152156),
	.w8(32'h3b2224c0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a7ae2),
	.w1(32'h3b9b1476),
	.w2(32'h39892e37),
	.w3(32'hba7dbea6),
	.w4(32'h3bb0e556),
	.w5(32'h3ba313ed),
	.w6(32'hbb11e983),
	.w7(32'hbb90505a),
	.w8(32'hbb8293af),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ce5fe),
	.w1(32'h3a9db2ed),
	.w2(32'hb9878f05),
	.w3(32'h3b460879),
	.w4(32'hba40edd0),
	.w5(32'hba532820),
	.w6(32'h37116247),
	.w7(32'hbae89a89),
	.w8(32'hbabed020),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f74f),
	.w1(32'hbbb415a8),
	.w2(32'hbc0fb0a2),
	.w3(32'hba3072e7),
	.w4(32'h3b04c2de),
	.w5(32'hbbcfcbc9),
	.w6(32'hbb62882e),
	.w7(32'hbb962315),
	.w8(32'hbc51816d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bcac1),
	.w1(32'h3bf01a72),
	.w2(32'h3ba40e03),
	.w3(32'h3a65f887),
	.w4(32'h3b1db5e8),
	.w5(32'h3b933b22),
	.w6(32'hbbfd29d4),
	.w7(32'h3ba587b4),
	.w8(32'hbb843270),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89cd9f),
	.w1(32'h3b032110),
	.w2(32'hba84daac),
	.w3(32'hba501761),
	.w4(32'h3aa00527),
	.w5(32'h3b1d98ff),
	.w6(32'hbbca93e7),
	.w7(32'hbabea6e0),
	.w8(32'hbb06bd42),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80ab6),
	.w1(32'h3c02853b),
	.w2(32'h3bb58a14),
	.w3(32'hbae82678),
	.w4(32'h38b3fccf),
	.w5(32'hbc463fdf),
	.w6(32'hbbac368b),
	.w7(32'hbc14c534),
	.w8(32'hbc8074d5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cf125),
	.w1(32'hbbbe9473),
	.w2(32'h3baf719a),
	.w3(32'hbc09e5cf),
	.w4(32'h3bc645dc),
	.w5(32'h3be6bc23),
	.w6(32'hbbf1b1f4),
	.w7(32'h3be9c34b),
	.w8(32'hba83baf5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b36a4),
	.w1(32'h3b49808f),
	.w2(32'hbb51b576),
	.w3(32'h3ba17430),
	.w4(32'h3ae809c1),
	.w5(32'h3aca444b),
	.w6(32'hbae50139),
	.w7(32'hbb620fbe),
	.w8(32'h3c0387f8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad16d72),
	.w1(32'hb9e8500c),
	.w2(32'h3ad5274a),
	.w3(32'hb985a41c),
	.w4(32'h3a054281),
	.w5(32'hbb727895),
	.w6(32'h39c1b7b9),
	.w7(32'hbace18f3),
	.w8(32'hba3cbbcd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb056161),
	.w1(32'h3b5105d7),
	.w2(32'hbaff41ae),
	.w3(32'h3a79f7d1),
	.w4(32'hbb497332),
	.w5(32'hbbff054e),
	.w6(32'h3a8644bf),
	.w7(32'hbba72d50),
	.w8(32'hbb9aee0c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954629),
	.w1(32'hbab62312),
	.w2(32'hbb11cfd3),
	.w3(32'hbc1b86a2),
	.w4(32'hbb6a2e10),
	.w5(32'h3a4bd8f6),
	.w6(32'hbc16ec83),
	.w7(32'hbb2c528b),
	.w8(32'hbaab1f14),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb496d6e),
	.w1(32'hbc3c6d70),
	.w2(32'hb99e49f2),
	.w3(32'hbb040325),
	.w4(32'h3af7df29),
	.w5(32'h3ca1f810),
	.w6(32'h3af2c2e0),
	.w7(32'h3b730449),
	.w8(32'h3b187dd3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c152298),
	.w1(32'h3b702c7b),
	.w2(32'h3ad5561f),
	.w3(32'h3bdb664b),
	.w4(32'h3b49d296),
	.w5(32'hba34a3c3),
	.w6(32'hbbddd2a7),
	.w7(32'h3bc33012),
	.w8(32'h3ab471d5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6388b),
	.w1(32'hbc0300ea),
	.w2(32'hbc18998c),
	.w3(32'hbb61e672),
	.w4(32'hba92fbb5),
	.w5(32'hbb14df7b),
	.w6(32'hbb97a76b),
	.w7(32'hbc11d742),
	.w8(32'h3a9e5521),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293aa6),
	.w1(32'h3c62985c),
	.w2(32'h3c0978fe),
	.w3(32'h3bd07aba),
	.w4(32'h3c0ca3e8),
	.w5(32'h3c532a6a),
	.w6(32'h3c084391),
	.w7(32'h3b006fa7),
	.w8(32'h3bcf693f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7de46),
	.w1(32'h3bc974c1),
	.w2(32'h3b1f0f9f),
	.w3(32'h3baab058),
	.w4(32'h3aa0beaa),
	.w5(32'hbac9625d),
	.w6(32'h3c0efa6f),
	.w7(32'hbb2f1dc5),
	.w8(32'hbb154742),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b515849),
	.w1(32'h3bedad39),
	.w2(32'hbad50f46),
	.w3(32'hba027859),
	.w4(32'h3b3466cb),
	.w5(32'h3b81f52d),
	.w6(32'h3b861179),
	.w7(32'hbc0dfeb5),
	.w8(32'hbb3183e1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c5903),
	.w1(32'hb8d06cde),
	.w2(32'hbb43f78e),
	.w3(32'hbbcda1a1),
	.w4(32'hb9883968),
	.w5(32'h3bd6af48),
	.w6(32'hbba5b648),
	.w7(32'hbb963e3a),
	.w8(32'hbb9d32f8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e22e1),
	.w1(32'hbc45c950),
	.w2(32'hbb7f4776),
	.w3(32'hbaea6ed5),
	.w4(32'hbaec30f6),
	.w5(32'hbbd0dbaa),
	.w6(32'hbb17c451),
	.w7(32'h3ace135c),
	.w8(32'h3a5d2fa9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf92159),
	.w1(32'hbc2ad01d),
	.w2(32'hbc1f75d5),
	.w3(32'hbc16a054),
	.w4(32'hbc533375),
	.w5(32'hbc2246f7),
	.w6(32'hbbe261d2),
	.w7(32'hbc8049bb),
	.w8(32'hbc216751),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41fd76),
	.w1(32'h3b12acf7),
	.w2(32'h3bdd2be1),
	.w3(32'hbc0cb479),
	.w4(32'h3b9c4270),
	.w5(32'h3bfe8313),
	.w6(32'hbb0f222f),
	.w7(32'h3b02d39b),
	.w8(32'hb9fe6d4b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b116207),
	.w1(32'hbb9782d8),
	.w2(32'h3a5f20a3),
	.w3(32'h3b108809),
	.w4(32'h3b1b2e34),
	.w5(32'h39e11c2f),
	.w6(32'hba9a1105),
	.w7(32'h3bbd45d0),
	.w8(32'hba6db1ca),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba976b1),
	.w1(32'hbbf12f9a),
	.w2(32'h3a4f5289),
	.w3(32'hbb48cae0),
	.w4(32'hbc13bacc),
	.w5(32'hbc2f0a88),
	.w6(32'hbbbb137e),
	.w7(32'hbbba8d3e),
	.w8(32'hbc4ccb8c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c915e),
	.w1(32'h3abc5d2f),
	.w2(32'hbb0bcc7a),
	.w3(32'hbbf129e7),
	.w4(32'hbb0eb7d5),
	.w5(32'h395c4ef3),
	.w6(32'hbc4a4b25),
	.w7(32'hbbd7cb06),
	.w8(32'hbaf7f1fd),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd73c1d),
	.w1(32'h3ba3f864),
	.w2(32'h3bbf9943),
	.w3(32'hbbc2302b),
	.w4(32'h3b252767),
	.w5(32'hbb0add63),
	.w6(32'hbb5e073e),
	.w7(32'h38771ccd),
	.w8(32'hbb4721e4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f597b),
	.w1(32'h3a20c029),
	.w2(32'h3bf5ad89),
	.w3(32'hbaf241fb),
	.w4(32'h3b9c751e),
	.w5(32'h3c22540c),
	.w6(32'hbb0ab02c),
	.w7(32'h39a6bced),
	.w8(32'h3a6d04d8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc053cfa),
	.w1(32'hbbf5e4be),
	.w2(32'hbc1eeb3e),
	.w3(32'hbbf41ac2),
	.w4(32'hbc7a3035),
	.w5(32'hbba01419),
	.w6(32'hbc283f14),
	.w7(32'hbc5715ef),
	.w8(32'hbc3723fb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a84a0),
	.w1(32'hba241ac4),
	.w2(32'hbba76b00),
	.w3(32'hb9a340c2),
	.w4(32'hbc4ce651),
	.w5(32'hbca69d89),
	.w6(32'h3a90b3ac),
	.w7(32'hbb0b4f80),
	.w8(32'hbbbd9e78),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a1cd4),
	.w1(32'hbbe1d21e),
	.w2(32'hbc93c608),
	.w3(32'hbc8682f0),
	.w4(32'hbbc44b01),
	.w5(32'hbbab642a),
	.w6(32'hbb8f6f5a),
	.w7(32'hbbfc9486),
	.w8(32'hbc1dbe67),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89c6de),
	.w1(32'h3bcf6845),
	.w2(32'hba7f6963),
	.w3(32'hbc6d062a),
	.w4(32'hbb7a18d9),
	.w5(32'h3bb67262),
	.w6(32'hbc65382a),
	.w7(32'h3b309fc2),
	.w8(32'hbb5e51ac),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8d199),
	.w1(32'h3c002d0e),
	.w2(32'h3c0832e0),
	.w3(32'hbb8ea104),
	.w4(32'h3c151f25),
	.w5(32'h3bfa0ea9),
	.w6(32'h3b555a4c),
	.w7(32'h3aa1781e),
	.w8(32'hbb432523),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6a07f),
	.w1(32'h3b0e8cf3),
	.w2(32'hba73645b),
	.w3(32'h3b1033e4),
	.w4(32'h3a9b2189),
	.w5(32'hbbed67d1),
	.w6(32'hbb8ba0b7),
	.w7(32'hbaaad5d6),
	.w8(32'hbba9df1f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf6d69),
	.w1(32'hbb65f860),
	.w2(32'hbbb3bfd8),
	.w3(32'hbb4c7a25),
	.w4(32'hbb235f97),
	.w5(32'hbaaf9de4),
	.w6(32'hbb96e77c),
	.w7(32'hbc0054aa),
	.w8(32'h3a94f4e1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3cbae),
	.w1(32'h3bcc9148),
	.w2(32'hba682ddd),
	.w3(32'hba497516),
	.w4(32'h3c5587b8),
	.w5(32'h3bdc6ab6),
	.w6(32'h3bae83aa),
	.w7(32'h3b804766),
	.w8(32'hbc03f20b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2fda),
	.w1(32'hba571c5e),
	.w2(32'hbb899b21),
	.w3(32'hb9614f7d),
	.w4(32'hbb52da77),
	.w5(32'hbb766117),
	.w6(32'hbc080f92),
	.w7(32'hbbda40f9),
	.w8(32'h3b08e6c5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4f0ab),
	.w1(32'hba208417),
	.w2(32'hbb84bbf3),
	.w3(32'hbb46b957),
	.w4(32'h3ad1008f),
	.w5(32'hba18e955),
	.w6(32'hbb19791f),
	.w7(32'hbb71abdc),
	.w8(32'h3ba7368a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bd4e8),
	.w1(32'hba75cceb),
	.w2(32'hbbd5b602),
	.w3(32'hbb4e6e8c),
	.w4(32'hbb8a2054),
	.w5(32'hb9bcd7fd),
	.w6(32'hbb2a9d35),
	.w7(32'hbc1345af),
	.w8(32'hbae90d2c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46768),
	.w1(32'h3ae1ae89),
	.w2(32'h3c20894b),
	.w3(32'hbb87e076),
	.w4(32'h3ade8109),
	.w5(32'h3c0e120e),
	.w6(32'hbba3f4a2),
	.w7(32'h3bc90f94),
	.w8(32'h3a13aaa9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1163d1),
	.w1(32'h3c12d6ad),
	.w2(32'hbb4bfd76),
	.w3(32'hba5a9035),
	.w4(32'hbb85ee43),
	.w5(32'hbbe0b033),
	.w6(32'hbbb24591),
	.w7(32'hbc0d51df),
	.w8(32'hbc315389),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bab41),
	.w1(32'h3b64ca5e),
	.w2(32'hbab2c817),
	.w3(32'hbb2126ad),
	.w4(32'h3bc466a2),
	.w5(32'hbaee208b),
	.w6(32'hbb923522),
	.w7(32'h3ac76d61),
	.w8(32'h3818e1f4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7908dc),
	.w1(32'h3b847258),
	.w2(32'hbaaded9b),
	.w3(32'hbad55654),
	.w4(32'hbb4b0c08),
	.w5(32'hbc497c99),
	.w6(32'hbbe006eb),
	.w7(32'hbb602979),
	.w8(32'hbbdcafff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cfdbd),
	.w1(32'h3ad92eb4),
	.w2(32'h3bc94d50),
	.w3(32'hbbee8a2a),
	.w4(32'hb8f652a3),
	.w5(32'h3acf0bd0),
	.w6(32'hb8870275),
	.w7(32'hbbe6972e),
	.w8(32'hba2d576d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e68a32),
	.w1(32'hba251e6f),
	.w2(32'h3bb19770),
	.w3(32'hbb4117e2),
	.w4(32'h3a592466),
	.w5(32'hba93418d),
	.w6(32'h3afff748),
	.w7(32'h3a778e9d),
	.w8(32'h39b74b54),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38e1ef),
	.w1(32'hbb55a7e0),
	.w2(32'hbc65df86),
	.w3(32'hbb895c85),
	.w4(32'hbc4cbf51),
	.w5(32'hbc24dc37),
	.w6(32'hb96a97db),
	.w7(32'hbc0438fc),
	.w8(32'hbc28cd54),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae69588),
	.w1(32'hba4191fe),
	.w2(32'hbc0eab43),
	.w3(32'hbaab2e5e),
	.w4(32'h3bff9c51),
	.w5(32'hbbc99966),
	.w6(32'h3bd38011),
	.w7(32'h3c02a04a),
	.w8(32'hbb02c756),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf2ad0),
	.w1(32'h3b9b3ae9),
	.w2(32'h3b620efb),
	.w3(32'hbb963be1),
	.w4(32'h3aeeeb41),
	.w5(32'hbbf803e7),
	.w6(32'hb9ef0bd4),
	.w7(32'hbb33cced),
	.w8(32'hbb9625c2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968108d),
	.w1(32'h3bd43435),
	.w2(32'h3ca22f02),
	.w3(32'h3b0db79d),
	.w4(32'h3ca4ac63),
	.w5(32'h3ca22784),
	.w6(32'h3b86d1e1),
	.w7(32'h3b41713b),
	.w8(32'hbb941030),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4e67e),
	.w1(32'h3b637e7b),
	.w2(32'hbb15043c),
	.w3(32'hba5eacdd),
	.w4(32'h3b476c91),
	.w5(32'hb9f973b5),
	.w6(32'hbc2f20e0),
	.w7(32'h39f24857),
	.w8(32'h3a463b48),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29e0b8),
	.w1(32'hba0bafe1),
	.w2(32'h3b89d111),
	.w3(32'h3a884ab3),
	.w4(32'h3b4e5196),
	.w5(32'h38ad8188),
	.w6(32'h3a81ac47),
	.w7(32'hbb449d4e),
	.w8(32'hbb8d5743),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc02ebf),
	.w1(32'h3b89873a),
	.w2(32'h3a520660),
	.w3(32'h39d1ca42),
	.w4(32'h3c052884),
	.w5(32'hba8c1d20),
	.w6(32'h3ac01669),
	.w7(32'h3bb3e14e),
	.w8(32'hba874c1b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38529f18),
	.w1(32'hbb9aba69),
	.w2(32'hbb031695),
	.w3(32'hba328df5),
	.w4(32'hbb77f049),
	.w5(32'h3bfff737),
	.w6(32'hbb620f02),
	.w7(32'h3a0ac3e6),
	.w8(32'h3b9c03cb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57c2ec),
	.w1(32'hbc17bf86),
	.w2(32'h3b0e179c),
	.w3(32'h3bbb970b),
	.w4(32'h3a2a9828),
	.w5(32'h3a3f0c87),
	.w6(32'h3b8cad5b),
	.w7(32'h3bd89c08),
	.w8(32'hbb3641ab),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e38b0),
	.w1(32'h3a873d14),
	.w2(32'h3a974b8a),
	.w3(32'hbbf4f45a),
	.w4(32'hbc149f8c),
	.w5(32'hbb56518c),
	.w6(32'hbc5379ae),
	.w7(32'hbb3cc03c),
	.w8(32'hbc5947f3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ffde),
	.w1(32'h3a2ffaca),
	.w2(32'h3aa27d20),
	.w3(32'hbba0e5a8),
	.w4(32'h3a625d9e),
	.w5(32'hb8c4566c),
	.w6(32'hbbee37cc),
	.w7(32'h3baa7a31),
	.w8(32'h39fba1b0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a001b41),
	.w1(32'h3c3a0ada),
	.w2(32'h3c90f1c0),
	.w3(32'hb92aff3a),
	.w4(32'h3cb1e2d4),
	.w5(32'h3ca3a36d),
	.w6(32'h3bdeabae),
	.w7(32'h3c114b1f),
	.w8(32'h3b101b9e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f52d3),
	.w1(32'hbb803622),
	.w2(32'hba58984e),
	.w3(32'h3c0cb0dd),
	.w4(32'h3a0d527c),
	.w5(32'h3affcb83),
	.w6(32'hbbe40dd6),
	.w7(32'h3a961583),
	.w8(32'h39a9e570),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b1f5f),
	.w1(32'hba9aafad),
	.w2(32'hbbde4971),
	.w3(32'h3b27d435),
	.w4(32'hbb5febaf),
	.w5(32'hbb04e0c1),
	.w6(32'h3aa11fd8),
	.w7(32'hbc05cbdf),
	.w8(32'hbbe3f2cf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f656),
	.w1(32'hbb060e09),
	.w2(32'h3b927be8),
	.w3(32'h3abaf757),
	.w4(32'hbb745aff),
	.w5(32'hbb621320),
	.w6(32'hbba42c31),
	.w7(32'hbb851022),
	.w8(32'hbbc734b7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae8c6),
	.w1(32'hbb5a9734),
	.w2(32'hbb582b05),
	.w3(32'hbb445369),
	.w4(32'hbc023428),
	.w5(32'hbb9b0c63),
	.w6(32'hbba7086c),
	.w7(32'hbaeb65dd),
	.w8(32'h3b0e96c2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05809b),
	.w1(32'h3ae5064e),
	.w2(32'hbb62df66),
	.w3(32'h3b528935),
	.w4(32'h3b19af70),
	.w5(32'hbb1ea8c0),
	.w6(32'hbad71d10),
	.w7(32'hbb36699b),
	.w8(32'hbae7bc24),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd342),
	.w1(32'hbc8b884e),
	.w2(32'hbcce4d9e),
	.w3(32'hbbc2855c),
	.w4(32'hbc3c4d81),
	.w5(32'hb9fc6449),
	.w6(32'hbc679d00),
	.w7(32'hbc1a8b44),
	.w8(32'h3a531936),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9426),
	.w1(32'hbb3ccf54),
	.w2(32'h39d147f6),
	.w3(32'h3b814af9),
	.w4(32'hbad951f8),
	.w5(32'h3b6868df),
	.w6(32'hbb50044a),
	.w7(32'h3a208ea4),
	.w8(32'h3bdce34f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b216b17),
	.w1(32'hbb284188),
	.w2(32'h3a78725b),
	.w3(32'h3bdd700b),
	.w4(32'h3b2b7b92),
	.w5(32'h3bcc0dbb),
	.w6(32'h3b9ba322),
	.w7(32'h389659d1),
	.w8(32'hbaf9a3ce),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd57a3),
	.w1(32'h3ac91577),
	.w2(32'h3a7c4e4a),
	.w3(32'h3a6b65e1),
	.w4(32'h3b8b68b8),
	.w5(32'hbbc00869),
	.w6(32'hbb8dfa42),
	.w7(32'hbaf10bad),
	.w8(32'h3ac04a73),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85bb6a),
	.w1(32'h3b2a5133),
	.w2(32'hbb26f47b),
	.w3(32'h39b99ae3),
	.w4(32'hba938425),
	.w5(32'hba13c6bd),
	.w6(32'hbaaf755e),
	.w7(32'hbb5f3b38),
	.w8(32'hbb62c87a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a26f),
	.w1(32'hbbece56a),
	.w2(32'hbc0c51c6),
	.w3(32'hbb85ee8c),
	.w4(32'hbb01aa41),
	.w5(32'hba907a47),
	.w6(32'hbb47abb3),
	.w7(32'hb9c3fa2b),
	.w8(32'h3afe4393),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca857),
	.w1(32'hbb9bc04f),
	.w2(32'hbbbb3406),
	.w3(32'hbc161def),
	.w4(32'hbbf7a05c),
	.w5(32'h3b63e879),
	.w6(32'hbc12d013),
	.w7(32'hbb197fcb),
	.w8(32'h3b2e4dec),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386257f0),
	.w1(32'hbc330ea5),
	.w2(32'hbb97f749),
	.w3(32'h3b032682),
	.w4(32'hbbba9d70),
	.w5(32'h3b33484a),
	.w6(32'h3c246733),
	.w7(32'h3ae65ce6),
	.w8(32'h3bcc0d4f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae007fa),
	.w1(32'hb917cf38),
	.w2(32'hbc5d3fd4),
	.w3(32'h3b141efa),
	.w4(32'hbbd3b9ba),
	.w5(32'hbc85e705),
	.w6(32'hbb5d6ecc),
	.w7(32'hba61b1ef),
	.w8(32'hbc19e98b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b288),
	.w1(32'hbab19214),
	.w2(32'h3c13122a),
	.w3(32'hbc068a38),
	.w4(32'h3c356fa0),
	.w5(32'h3c2c7347),
	.w6(32'h3a8fa492),
	.w7(32'h3c9c9789),
	.w8(32'h3bb9cab5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c524d96),
	.w1(32'h3b4f83c2),
	.w2(32'h3b209b90),
	.w3(32'h3bce5462),
	.w4(32'hbbaaaa2c),
	.w5(32'hba82a01b),
	.w6(32'h3989a1c4),
	.w7(32'h3ae38aee),
	.w8(32'hbabdd2f0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b584311),
	.w1(32'h3b0110e9),
	.w2(32'hbb48ba2c),
	.w3(32'hba212784),
	.w4(32'hbba4939e),
	.w5(32'hbbbe5312),
	.w6(32'hbab8cc07),
	.w7(32'hbaeb6ef2),
	.w8(32'hbb1894aa),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902abe3),
	.w1(32'hbad850b0),
	.w2(32'h3b021823),
	.w3(32'hbb9ff699),
	.w4(32'h3a857673),
	.w5(32'h3ba3002f),
	.w6(32'hbbeb5d44),
	.w7(32'h3ae87ac9),
	.w8(32'hbb7a2044),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3a0a4),
	.w1(32'h3beab5ff),
	.w2(32'h3c015f1d),
	.w3(32'h3b79230b),
	.w4(32'h3a62d413),
	.w5(32'hbae79f07),
	.w6(32'h3a58bea4),
	.w7(32'h3be6581f),
	.w8(32'hbbcf3dbc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baca44b),
	.w1(32'h3a4741df),
	.w2(32'hb5dee552),
	.w3(32'h389d5a39),
	.w4(32'h3a9bbe5b),
	.w5(32'hbb00ec44),
	.w6(32'hbaf6b1ab),
	.w7(32'hbbc51da5),
	.w8(32'hbb89d3a8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79c622),
	.w1(32'h3b1532c8),
	.w2(32'h3b3edb2c),
	.w3(32'hbac4857b),
	.w4(32'hb9935aba),
	.w5(32'hbbbfce62),
	.w6(32'hbb8c65b6),
	.w7(32'h3b09994e),
	.w8(32'hbbf63c96),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c78a),
	.w1(32'h3924d211),
	.w2(32'h3b76b135),
	.w3(32'hb8dab586),
	.w4(32'h3b21abf7),
	.w5(32'h3b8b9534),
	.w6(32'hbb3c19f2),
	.w7(32'hbb097b26),
	.w8(32'hbb9d6611),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214bc4),
	.w1(32'hbb701009),
	.w2(32'hbb3ea157),
	.w3(32'h3b111afd),
	.w4(32'h3afde4a9),
	.w5(32'hbb37c885),
	.w6(32'hbb8f531c),
	.w7(32'hbb62867c),
	.w8(32'hbb60dae0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1639d3),
	.w1(32'h3a304642),
	.w2(32'h396e65d1),
	.w3(32'hbbc07d2c),
	.w4(32'h3a891baa),
	.w5(32'hbb648628),
	.w6(32'hbb6ee996),
	.w7(32'hbb92600b),
	.w8(32'hbaf5bc37),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc468ab7),
	.w1(32'hbc2b0f9a),
	.w2(32'hbbed0c07),
	.w3(32'hbc1c6bed),
	.w4(32'hbb2b9f0b),
	.w5(32'hbba4af72),
	.w6(32'hbb8361fa),
	.w7(32'hbbccdd36),
	.w8(32'h3b6b41d9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bbc80),
	.w1(32'h3bfcdc0a),
	.w2(32'h3c55dde2),
	.w3(32'h3bc73e7c),
	.w4(32'h3c0469c3),
	.w5(32'hb950e0d6),
	.w6(32'h3b9f8f25),
	.w7(32'h3baddab5),
	.w8(32'hbbe33530),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b602b66),
	.w1(32'h3b4b7a89),
	.w2(32'h3b130f41),
	.w3(32'hbbb8e468),
	.w4(32'hb9fd504c),
	.w5(32'hbb9976ef),
	.w6(32'hbc0e4b44),
	.w7(32'hbb807bd4),
	.w8(32'hbbdbebce),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab90ba6),
	.w1(32'hbc24eb72),
	.w2(32'hbbec9759),
	.w3(32'hbb14a98f),
	.w4(32'hb9a04383),
	.w5(32'h3ad0deef),
	.w6(32'hbbcfffc3),
	.w7(32'h3a90de16),
	.w8(32'hbb721788),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907ec6),
	.w1(32'h3ba59422),
	.w2(32'h3b9941b4),
	.w3(32'hbb867865),
	.w4(32'h39c847d2),
	.w5(32'hbba9f61a),
	.w6(32'hbb38777b),
	.w7(32'h3ac267e5),
	.w8(32'h3ac873b3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94cf27),
	.w1(32'h3c07f75a),
	.w2(32'h3bc8da28),
	.w3(32'hba19d80e),
	.w4(32'hbac39744),
	.w5(32'hbb9628e8),
	.w6(32'hbb03c71d),
	.w7(32'hbb20bf36),
	.w8(32'hbbbd10be),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658b20),
	.w1(32'h3a74723c),
	.w2(32'hbb5af013),
	.w3(32'hbb3a28f8),
	.w4(32'h3adacb12),
	.w5(32'hbb9bf5c7),
	.w6(32'hbb439240),
	.w7(32'hbba3925b),
	.w8(32'hbc1760ab),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10a03),
	.w1(32'hbba5fc96),
	.w2(32'hbbaf8b02),
	.w3(32'h3b6f9d94),
	.w4(32'h392d13d4),
	.w5(32'hbb820036),
	.w6(32'hbbc9f7d7),
	.w7(32'hbb31dd9c),
	.w8(32'hbb915198),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8c0d6),
	.w1(32'hbc042fa4),
	.w2(32'hbae95873),
	.w3(32'h3b1f08f4),
	.w4(32'h3a5acb42),
	.w5(32'h390c4264),
	.w6(32'h3b50278e),
	.w7(32'h3c00bb53),
	.w8(32'h3bea4ded),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c1729),
	.w1(32'hbbc1ed46),
	.w2(32'h3ae4d505),
	.w3(32'hbba86cbc),
	.w4(32'h3b1cfe9f),
	.w5(32'h3baa0f32),
	.w6(32'h3a23420b),
	.w7(32'h3c47ac7f),
	.w8(32'h3b929fdb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b687424),
	.w1(32'h3c0f6234),
	.w2(32'hbb94a230),
	.w3(32'h3a9d3535),
	.w4(32'h3b16b658),
	.w5(32'hbbf20328),
	.w6(32'hbbbd4e11),
	.w7(32'hbc6643eb),
	.w8(32'hbbf4a7a3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab10f),
	.w1(32'hbbfa5554),
	.w2(32'hbad77643),
	.w3(32'hbc26c008),
	.w4(32'hbc3e3cfe),
	.w5(32'hbca6d2ab),
	.w6(32'hbc011a48),
	.w7(32'hbc3207c9),
	.w8(32'hbaff8c28),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc535d20),
	.w1(32'hbc3d8da9),
	.w2(32'hbc9411cf),
	.w3(32'hbc21925c),
	.w4(32'h3b02133c),
	.w5(32'h3ca7e2f1),
	.w6(32'hb954c84a),
	.w7(32'hbbde329f),
	.w8(32'hbc8967ea),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bb9e3),
	.w1(32'hbb02b081),
	.w2(32'hbc33a135),
	.w3(32'hbc55d5d9),
	.w4(32'h3a40bb8b),
	.w5(32'h3b0d133e),
	.w6(32'hbc881d8c),
	.w7(32'hbb09234a),
	.w8(32'hb8eeea1f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba041ddd),
	.w1(32'h3c082204),
	.w2(32'h3a90ea1e),
	.w3(32'hbbb1f429),
	.w4(32'h3c221a02),
	.w5(32'h3ba9d186),
	.w6(32'hbbe22b48),
	.w7(32'h3ac779b0),
	.w8(32'h39f24638),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf6f58),
	.w1(32'h3b8a13b4),
	.w2(32'hba50321a),
	.w3(32'hbab9994b),
	.w4(32'h3c2c221f),
	.w5(32'h3d026c64),
	.w6(32'h3b06aca0),
	.w7(32'h3b1d1fe6),
	.w8(32'hbc18bc64),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b31007),
	.w1(32'hba888334),
	.w2(32'h3ba8c05c),
	.w3(32'h3c863bdb),
	.w4(32'h3c2588b0),
	.w5(32'h3cdf612c),
	.w6(32'h3c1038c4),
	.w7(32'h3bc2ccef),
	.w8(32'hba07a993),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1da14),
	.w1(32'h3b94642b),
	.w2(32'h3c1e7d2f),
	.w3(32'h3c2567f6),
	.w4(32'h3b81397c),
	.w5(32'h3b010f27),
	.w6(32'h3c09d44e),
	.w7(32'h3b3b4092),
	.w8(32'hbb340204),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a3f94),
	.w1(32'h3cfc33d1),
	.w2(32'h3c42b14a),
	.w3(32'h3a27ad21),
	.w4(32'h3cc9051b),
	.w5(32'h3c7d1817),
	.w6(32'h38f17334),
	.w7(32'h3c4bd647),
	.w8(32'h3c2b7c92),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18a035),
	.w1(32'h3bf20675),
	.w2(32'h3bc050c4),
	.w3(32'h3ce0e5b1),
	.w4(32'h3bfcc82b),
	.w5(32'hba5179dc),
	.w6(32'h3ccba718),
	.w7(32'h3bcdc77d),
	.w8(32'h3b9879e5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1ac1d),
	.w1(32'hbb9c4b06),
	.w2(32'hbbbd976e),
	.w3(32'h3bd38213),
	.w4(32'hbc45e0b5),
	.w5(32'hbc567049),
	.w6(32'h3b2b444e),
	.w7(32'hbbe1b66c),
	.w8(32'hbc106f84),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1631b4),
	.w1(32'h3a2aba29),
	.w2(32'h3b5ed080),
	.w3(32'hba463a33),
	.w4(32'h3bc25531),
	.w5(32'h3b9cf711),
	.w6(32'hbbaa7f74),
	.w7(32'h3b0470c1),
	.w8(32'hbb027593),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364b7d),
	.w1(32'hbb2d4ddc),
	.w2(32'hbb43cb02),
	.w3(32'h3b1d0993),
	.w4(32'hbb582e9a),
	.w5(32'hbbb394a4),
	.w6(32'h39251230),
	.w7(32'hbc0a63e4),
	.w8(32'hbba08f0e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadfa5f),
	.w1(32'hbae42125),
	.w2(32'h3c043848),
	.w3(32'h3b075d15),
	.w4(32'h3bda9c91),
	.w5(32'h3b89743f),
	.w6(32'h3a7b2182),
	.w7(32'h3abd4daf),
	.w8(32'hbb1d82b5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcc960),
	.w1(32'hbb5922e9),
	.w2(32'hbb593b9c),
	.w3(32'h3b9ff49f),
	.w4(32'h3b8ccc65),
	.w5(32'hbc471238),
	.w6(32'h3aee6de4),
	.w7(32'hbb3b86c0),
	.w8(32'h39109d2d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ddd90),
	.w1(32'hbc789cb1),
	.w2(32'hbc8aa87d),
	.w3(32'hbc1b091e),
	.w4(32'hbc1d5459),
	.w5(32'hbb3340c7),
	.w6(32'hbc1f8602),
	.w7(32'hbc9687af),
	.w8(32'hbc7d8dd5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451c3e),
	.w1(32'hba9e7ae6),
	.w2(32'h3aaa13c5),
	.w3(32'hb9e2f86f),
	.w4(32'h3a4e04e0),
	.w5(32'hbc1b2bbc),
	.w6(32'hbb920fa5),
	.w7(32'hbb84a237),
	.w8(32'h3a5e5912),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb202d71),
	.w1(32'hbc690e8d),
	.w2(32'hbc174bbe),
	.w3(32'hbb4c926d),
	.w4(32'hbc29dc55),
	.w5(32'hbc3b7db4),
	.w6(32'hbc543e99),
	.w7(32'hbcb4c90f),
	.w8(32'hbcab9c6a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7127c5),
	.w1(32'h3a2acdf5),
	.w2(32'h3b4a738b),
	.w3(32'hbc27e5ab),
	.w4(32'h3aaebd60),
	.w5(32'h3ca46e47),
	.w6(32'hbc86b19f),
	.w7(32'hbc1f511a),
	.w8(32'hbc4dde83),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad56c96),
	.w1(32'hba671f9f),
	.w2(32'h3b98adb8),
	.w3(32'hbb0d5078),
	.w4(32'h3a17d028),
	.w5(32'hbb442021),
	.w6(32'hbc59f574),
	.w7(32'h3b949a17),
	.w8(32'hbbab0689),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80afc),
	.w1(32'h3b7a0da6),
	.w2(32'hbb44732f),
	.w3(32'h3b7f0bf7),
	.w4(32'hb9a69f6e),
	.w5(32'h3c165006),
	.w6(32'h3b049ffc),
	.w7(32'h3b0be99e),
	.w8(32'h3c9bc67c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d8c44),
	.w1(32'hbc239371),
	.w2(32'hbc117e6f),
	.w3(32'hbc0cfb34),
	.w4(32'hbc6102e9),
	.w5(32'hbb9c3b32),
	.w6(32'h3ac614e9),
	.w7(32'hbc88fa6e),
	.w8(32'hba82d226),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ffb8),
	.w1(32'hbb6405ae),
	.w2(32'hbbb21419),
	.w3(32'hbc107ce2),
	.w4(32'hbc2c44bf),
	.w5(32'hbb5abc18),
	.w6(32'hbc282752),
	.w7(32'hbc64f50b),
	.w8(32'hbb86449d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab76e35),
	.w1(32'h3b472c2b),
	.w2(32'h3c1e93bc),
	.w3(32'h3b2de04a),
	.w4(32'h3bcde009),
	.w5(32'hbc54f94b),
	.w6(32'hbb0d0a5b),
	.w7(32'h3c0a7a24),
	.w8(32'h3c980963),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b299287),
	.w1(32'h3b024487),
	.w2(32'h3c0fc4e1),
	.w3(32'h3bc486f7),
	.w4(32'h3b8c71f6),
	.w5(32'hbbbc1fec),
	.w6(32'h3c0c5a45),
	.w7(32'hb9cebd76),
	.w8(32'hba5d5f3c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae14daf),
	.w1(32'h3ab541fa),
	.w2(32'h3b453243),
	.w3(32'hbaef5117),
	.w4(32'h3b73a691),
	.w5(32'h3bb80871),
	.w6(32'hbb532229),
	.w7(32'h3b0cf6d1),
	.w8(32'hbaac4035),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe933f9),
	.w1(32'h3c83bf99),
	.w2(32'h3c3dc997),
	.w3(32'hb9ed6136),
	.w4(32'h3c6ad026),
	.w5(32'h3cce8619),
	.w6(32'hbabf3da4),
	.w7(32'h3c9aa7c5),
	.w8(32'h3c9701bf),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb093f9),
	.w1(32'h3946e47f),
	.w2(32'hbb48aa43),
	.w3(32'h3c29f3bd),
	.w4(32'h3b91b731),
	.w5(32'h3c09f0b7),
	.w6(32'h3bb90a31),
	.w7(32'hbc1e48f1),
	.w8(32'hbc39ef4b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4798a5),
	.w1(32'hbbca59ff),
	.w2(32'hbc04e150),
	.w3(32'hbb4deaf4),
	.w4(32'hbc10839d),
	.w5(32'h3aac88af),
	.w6(32'hbc797aa8),
	.w7(32'hbc571ded),
	.w8(32'hbb4b414d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23da71),
	.w1(32'h3b27502a),
	.w2(32'hbb0b8b5f),
	.w3(32'hbbcb9558),
	.w4(32'hbb654a4d),
	.w5(32'hbac4fdd8),
	.w6(32'hbb5efd1f),
	.w7(32'h3a923eb6),
	.w8(32'h3c3a119f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c1449),
	.w1(32'hbc1c0bb3),
	.w2(32'hbc4e92c0),
	.w3(32'hbad00c16),
	.w4(32'hba869e93),
	.w5(32'h3b2c2714),
	.w6(32'hb9a6915e),
	.w7(32'hbb1e9c0a),
	.w8(32'hbace75d7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05ee60),
	.w1(32'hbacd8b25),
	.w2(32'hbb2cbd25),
	.w3(32'h39c7cd71),
	.w4(32'h3b7eccc5),
	.w5(32'h3c001043),
	.w6(32'h3b947365),
	.w7(32'hba269992),
	.w8(32'hbaa04d0c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be9fd),
	.w1(32'hbafb41f1),
	.w2(32'hbbbf8fd9),
	.w3(32'h3a51d240),
	.w4(32'hbbfcd3ef),
	.w5(32'hbbbe0e8e),
	.w6(32'hbad4cabf),
	.w7(32'hbb54923e),
	.w8(32'hbb35d37c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94f570),
	.w1(32'h3b86a8ae),
	.w2(32'hbbdaf821),
	.w3(32'hbcbb1810),
	.w4(32'h3c59401d),
	.w5(32'h3c8593ba),
	.w6(32'hbcb00c9d),
	.w7(32'h3ba32032),
	.w8(32'h3bb9203d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8975655),
	.w1(32'hbb899087),
	.w2(32'hbc4a9182),
	.w3(32'hbad6b52a),
	.w4(32'hbc04608c),
	.w5(32'h3b67bf90),
	.w6(32'h3ad379fb),
	.w7(32'hbc2a6284),
	.w8(32'hb9f64114),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29d643),
	.w1(32'h3c0b9d98),
	.w2(32'h3caaaccd),
	.w3(32'hbb36180e),
	.w4(32'hbbbd5b04),
	.w5(32'hbce5a5e1),
	.w6(32'h3b331144),
	.w7(32'h369c9f41),
	.w8(32'h3c27a382),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be81c8f),
	.w1(32'hbb70a030),
	.w2(32'hbbdcbd49),
	.w3(32'hbc3b7862),
	.w4(32'hbc233f9b),
	.w5(32'hbc188191),
	.w6(32'h3bf2e6d3),
	.w7(32'hbc3cf207),
	.w8(32'hbb380c88),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2565d3),
	.w1(32'h3c0fa4d4),
	.w2(32'h3c416b19),
	.w3(32'hbb5c8545),
	.w4(32'h3be0ca44),
	.w5(32'hba2bbcb6),
	.w6(32'hba9c0cea),
	.w7(32'h39a02b53),
	.w8(32'hbb09baae),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e510),
	.w1(32'hbb81516d),
	.w2(32'hbba5b61e),
	.w3(32'hb9ed24cd),
	.w4(32'h3ba0460f),
	.w5(32'h391b98b8),
	.w6(32'hbb7b3cba),
	.w7(32'hbc159ef3),
	.w8(32'hb8ffc0c6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf67df2),
	.w1(32'h3bc2e341),
	.w2(32'h3c0601be),
	.w3(32'hbc19e636),
	.w4(32'h3b0b1606),
	.w5(32'h3bd5ae68),
	.w6(32'h3ac11420),
	.w7(32'hbba00353),
	.w8(32'hbc1d7e66),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8abab5),
	.w1(32'h3c2da2af),
	.w2(32'h3c7b36b0),
	.w3(32'h3ac36a55),
	.w4(32'hbba37a8f),
	.w5(32'hbcf769a5),
	.w6(32'hba9eecd2),
	.w7(32'h3c94b193),
	.w8(32'h3cb9274c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f889d),
	.w1(32'hbc18c102),
	.w2(32'hbb9ca4c2),
	.w3(32'h3a5d08b3),
	.w4(32'hbc0f5441),
	.w5(32'hbab20e2c),
	.w6(32'h3c2cd9b5),
	.w7(32'h3bf5407f),
	.w8(32'h3c24e6e7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39890035),
	.w1(32'hbb4d5f12),
	.w2(32'hbb58bbbf),
	.w3(32'hbbbfaf00),
	.w4(32'hbb0c6036),
	.w5(32'hbb0496d2),
	.w6(32'hbb7764ba),
	.w7(32'hbb494876),
	.w8(32'h39285c44),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83522e),
	.w1(32'hba71e567),
	.w2(32'hbb567e41),
	.w3(32'hbbda7daa),
	.w4(32'hbb930ef1),
	.w5(32'hbaa46f82),
	.w6(32'hbbba55db),
	.w7(32'hbac5690a),
	.w8(32'h3b896013),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabe6b9),
	.w1(32'hbab85d5c),
	.w2(32'hb7656db1),
	.w3(32'hb4c33ad8),
	.w4(32'h3a5210ef),
	.w5(32'h3b839155),
	.w6(32'h3af1b913),
	.w7(32'h3be63a84),
	.w8(32'h3c2f39f9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6221b),
	.w1(32'hbb9f6cb1),
	.w2(32'h3ab18676),
	.w3(32'h3bce2988),
	.w4(32'h3c126902),
	.w5(32'hbc08a40a),
	.w6(32'h3b00d1b2),
	.w7(32'h3bd59a02),
	.w8(32'h3a36f3b0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb059d96),
	.w1(32'hbb0fa39d),
	.w2(32'hbba3c9f2),
	.w3(32'hbbbc6eac),
	.w4(32'hbc141306),
	.w5(32'hbc0a7995),
	.w6(32'h3a92bb9d),
	.w7(32'hbc1d6953),
	.w8(32'hba3e7836),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5e0e3),
	.w1(32'h3b19cce3),
	.w2(32'h3bb5e53e),
	.w3(32'hbb284bbd),
	.w4(32'hba8c8a8f),
	.w5(32'h3aafde32),
	.w6(32'h3ba8aeed),
	.w7(32'h3ab2ac91),
	.w8(32'h3b909244),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babccd2),
	.w1(32'h3b2619e6),
	.w2(32'h3c302a3c),
	.w3(32'h3c0cd5fd),
	.w4(32'h3af9a74a),
	.w5(32'hbbb94084),
	.w6(32'h3b336c85),
	.w7(32'h3b61972e),
	.w8(32'h3bff7b5c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa50ceb),
	.w1(32'h3bdb282d),
	.w2(32'hbc556f76),
	.w3(32'hba9642a5),
	.w4(32'h3ba98bd3),
	.w5(32'h3c4c24d6),
	.w6(32'h3ba36972),
	.w7(32'h3bdf040a),
	.w8(32'hbbdf7e07),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebde09),
	.w1(32'hbbbbc6cc),
	.w2(32'hbbf8963e),
	.w3(32'h3b9f7991),
	.w4(32'hbb730d57),
	.w5(32'hbc33bb3b),
	.w6(32'h3c42192b),
	.w7(32'hbb90cc18),
	.w8(32'hbc07fd09),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10b694),
	.w1(32'h3bcbc212),
	.w2(32'h3b9a004d),
	.w3(32'hbc3b5bba),
	.w4(32'hbb74dde6),
	.w5(32'hbc0d3d36),
	.w6(32'hbc3ecd91),
	.w7(32'hba7389d7),
	.w8(32'hbaa0f79b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb126576),
	.w1(32'h3b53c107),
	.w2(32'h3afd3a2b),
	.w3(32'h3b2b1c7d),
	.w4(32'hba6fdb1a),
	.w5(32'h3b8e1ab5),
	.w6(32'h3bdd3046),
	.w7(32'h3c5a3afa),
	.w8(32'h3c952a4d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395bf5),
	.w1(32'hbbed017c),
	.w2(32'h3a86047c),
	.w3(32'h3be91ab4),
	.w4(32'hbc38b0d8),
	.w5(32'hbc6710f8),
	.w6(32'h3b896ebc),
	.w7(32'hbc704a6f),
	.w8(32'hbc77c090),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cb353),
	.w1(32'hbb7a1880),
	.w2(32'hbc321ae2),
	.w3(32'hbc3b11a9),
	.w4(32'h3a89e0dc),
	.w5(32'h3ae142e5),
	.w6(32'hbc220fbc),
	.w7(32'hbba79bc8),
	.w8(32'h386bcfe9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe14a0f),
	.w1(32'hbc10e67f),
	.w2(32'hbc6268f0),
	.w3(32'hbb8130bc),
	.w4(32'h3af4086d),
	.w5(32'h3c7f69bd),
	.w6(32'h3b85336e),
	.w7(32'hbc185bbb),
	.w8(32'hbc4aab19),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc2153),
	.w1(32'hbb601b90),
	.w2(32'hba2f004c),
	.w3(32'hbba7be21),
	.w4(32'hbc253dfe),
	.w5(32'hbc930a2b),
	.w6(32'hbc80db8f),
	.w7(32'hbb173929),
	.w8(32'h3c7453d7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1487a3),
	.w1(32'hbb100fd0),
	.w2(32'h3a90b2ea),
	.w3(32'hbbe9b406),
	.w4(32'h3bc83a82),
	.w5(32'h3b8b2c26),
	.w6(32'h3b19ca22),
	.w7(32'h3c08bac4),
	.w8(32'h3c4f2d0d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf50fce),
	.w1(32'hbc02b31d),
	.w2(32'hbb9edee3),
	.w3(32'hbb26feda),
	.w4(32'hbb5a37fb),
	.w5(32'h3c36a873),
	.w6(32'h3980cb62),
	.w7(32'h39b3f047),
	.w8(32'hbc0d25be),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule