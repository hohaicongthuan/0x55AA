module layer_10_featuremap_249(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2227b9),
	.w1(32'h3c4abea1),
	.w2(32'h3b9c2b83),
	.w3(32'h3c171814),
	.w4(32'h3c042d12),
	.w5(32'h3bda7754),
	.w6(32'h3c1d4181),
	.w7(32'h3bae8c2e),
	.w8(32'h3bf032c0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3fa94),
	.w1(32'h3b07c9f9),
	.w2(32'h3c012629),
	.w3(32'hba87dc57),
	.w4(32'hbb2881e8),
	.w5(32'hbc0c5a54),
	.w6(32'hbbd9c69c),
	.w7(32'h3b27391f),
	.w8(32'hbb345f8e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a3ed4),
	.w1(32'hbb709e97),
	.w2(32'hbb28a46f),
	.w3(32'hbb80ba55),
	.w4(32'hbb82098b),
	.w5(32'h3bae9585),
	.w6(32'hbb42b7ec),
	.w7(32'hbbe99819),
	.w8(32'h3c1e030b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bf946),
	.w1(32'h3bfc7977),
	.w2(32'h3bae239f),
	.w3(32'h3b7b3f0e),
	.w4(32'h3bc0f6ff),
	.w5(32'h3ad8ca97),
	.w6(32'h3c9b0f74),
	.w7(32'h3c07621a),
	.w8(32'hbbb270bf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb247ee0),
	.w1(32'hbb03deec),
	.w2(32'hbb2d165e),
	.w3(32'h39e1e51f),
	.w4(32'h3b42a3fd),
	.w5(32'hbb03b1c2),
	.w6(32'hbc167660),
	.w7(32'hbbbc4cc0),
	.w8(32'h3a9eba45),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dfee8),
	.w1(32'hb9d58a57),
	.w2(32'hbb4a8d28),
	.w3(32'hb9e19667),
	.w4(32'hbb35258e),
	.w5(32'hba9ba50a),
	.w6(32'h3b955b42),
	.w7(32'hba0ba8ae),
	.w8(32'h38582b5a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11d35e),
	.w1(32'hba711ff1),
	.w2(32'h3ab5c477),
	.w3(32'hbc12c287),
	.w4(32'hbb6dc8eb),
	.w5(32'h3bb8b503),
	.w6(32'h38b2c180),
	.w7(32'hba99f11e),
	.w8(32'h3c3a0a89),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc7265),
	.w1(32'h3c9d54d4),
	.w2(32'h3bce4bc6),
	.w3(32'h3cae2d6f),
	.w4(32'h3cd2ab28),
	.w5(32'h3bad46e9),
	.w6(32'h3d003bf9),
	.w7(32'h3cd3c160),
	.w8(32'h3c3751db),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4160e),
	.w1(32'h3c133e60),
	.w2(32'h3bcff07c),
	.w3(32'h3ba32fbe),
	.w4(32'h3b22258f),
	.w5(32'h3a9206cb),
	.w6(32'h3bbb1ca1),
	.w7(32'h3bb4d5d1),
	.w8(32'h3b6735d3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02a2f5),
	.w1(32'h3ade5a10),
	.w2(32'hbbe1435a),
	.w3(32'h38a3067a),
	.w4(32'hbba2ad86),
	.w5(32'hbbdc9a16),
	.w6(32'h3be17c4b),
	.w7(32'hbb0654f7),
	.w8(32'hbb0766a0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16b41d),
	.w1(32'h3ab36467),
	.w2(32'hbb47c833),
	.w3(32'hbac82eb8),
	.w4(32'h3ad3d6ef),
	.w5(32'h3918aaad),
	.w6(32'h3b9094ef),
	.w7(32'hb94ceec4),
	.w8(32'h3a46a3be),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8dc4a),
	.w1(32'hbc006f2d),
	.w2(32'hbb4cbc9d),
	.w3(32'hbbfdc3b2),
	.w4(32'h3ba4b1c5),
	.w5(32'h3bc31354),
	.w6(32'hbb89b31e),
	.w7(32'hbc0dffbc),
	.w8(32'h3b4b5578),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1daec8),
	.w1(32'h3b944b3e),
	.w2(32'h3a6c75e5),
	.w3(32'h3ac9cf29),
	.w4(32'hbab92eef),
	.w5(32'hbb74e2f1),
	.w6(32'hba208fcf),
	.w7(32'hbb59bfb7),
	.w8(32'hbb245c32),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c35b0),
	.w1(32'h3b15a9df),
	.w2(32'h3b884627),
	.w3(32'hbb841b13),
	.w4(32'hbaf60ada),
	.w5(32'hbb646219),
	.w6(32'hbb5298f2),
	.w7(32'h3b7f1625),
	.w8(32'h3b3ea872),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a6ab8),
	.w1(32'h3be87b8b),
	.w2(32'h3aacefc3),
	.w3(32'hbbab0cf3),
	.w4(32'hbb8434d9),
	.w5(32'h3bd1e37e),
	.w6(32'h3c34112a),
	.w7(32'h3b00b1ca),
	.w8(32'h3c1a1a6f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a0508),
	.w1(32'h3bdb1eb9),
	.w2(32'hba119132),
	.w3(32'h3bff06c6),
	.w4(32'h3a7f4637),
	.w5(32'hbbc32104),
	.w6(32'h3c40eee5),
	.w7(32'h3b8e5bc4),
	.w8(32'h3b33d969),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545c53),
	.w1(32'h3b05b09a),
	.w2(32'hbb4ddba6),
	.w3(32'h3a92a1ba),
	.w4(32'hbbc8065d),
	.w5(32'hbb4deb22),
	.w6(32'h3a6e0706),
	.w7(32'h39dae92e),
	.w8(32'hbb36d430),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10512f),
	.w1(32'h3b142068),
	.w2(32'hb9560ff3),
	.w3(32'h3bcb26dd),
	.w4(32'h3b96763f),
	.w5(32'hbbdcd62d),
	.w6(32'h3c41b46b),
	.w7(32'h3bc656c0),
	.w8(32'h3be38f39),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b2e74),
	.w1(32'hbb489417),
	.w2(32'hbb5761e2),
	.w3(32'hbadbc4f1),
	.w4(32'h38c1b45d),
	.w5(32'hbb2243ba),
	.w6(32'h3bf53d51),
	.w7(32'h3b5ed9e2),
	.w8(32'h3b60a67a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ffbca),
	.w1(32'h3a8f39a3),
	.w2(32'h3bb573ca),
	.w3(32'hb93a1f25),
	.w4(32'hb9c1c7f8),
	.w5(32'h3bac1198),
	.w6(32'h3aeebf0c),
	.w7(32'h3aacce00),
	.w8(32'h3c3cd924),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e9756),
	.w1(32'h3b328227),
	.w2(32'h3b7edcc1),
	.w3(32'h3b8821d9),
	.w4(32'hb9d66ed0),
	.w5(32'h3a92257e),
	.w6(32'h3bd6224d),
	.w7(32'h3b82fd38),
	.w8(32'h3aeb67f2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c93aa),
	.w1(32'h3b627f73),
	.w2(32'h3b1368c5),
	.w3(32'h3b89342c),
	.w4(32'h39a53c11),
	.w5(32'h3b5d2936),
	.w6(32'h3bfebb8b),
	.w7(32'h3b124075),
	.w8(32'h39715711),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083336),
	.w1(32'h3bdad5b6),
	.w2(32'hba93d468),
	.w3(32'h3c3a962f),
	.w4(32'h3c740c17),
	.w5(32'h39e74a1c),
	.w6(32'h3c36487e),
	.w7(32'h3b8f4e4b),
	.w8(32'h3c673417),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb48c34),
	.w1(32'h3a2e1cc9),
	.w2(32'hbb67654c),
	.w3(32'hbb17e5e1),
	.w4(32'h3ba25b9b),
	.w5(32'h3a30a906),
	.w6(32'h3bb4838a),
	.w7(32'h3bc32e2f),
	.w8(32'hbad04d4b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0487b),
	.w1(32'h3be15c90),
	.w2(32'h3c13ef5e),
	.w3(32'h3b64bc56),
	.w4(32'h386b1d52),
	.w5(32'hbb66bbd5),
	.w6(32'hbaa588f2),
	.w7(32'h3b539c68),
	.w8(32'h3ac8e540),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63e7d3),
	.w1(32'h3b413364),
	.w2(32'hbba30f34),
	.w3(32'hbb58be52),
	.w4(32'hbbac5e09),
	.w5(32'hbb3ffad1),
	.w6(32'h3be23241),
	.w7(32'h39636809),
	.w8(32'h3b644bb5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14b944),
	.w1(32'hba405c05),
	.w2(32'h38b970a8),
	.w3(32'hbacec1b2),
	.w4(32'h36889d2b),
	.w5(32'h3bf2cebd),
	.w6(32'h3bb27c15),
	.w7(32'h3bc4d4a5),
	.w8(32'h3c1467c6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61ba05),
	.w1(32'h3c421d45),
	.w2(32'h3bbecdfc),
	.w3(32'h3c2f54dd),
	.w4(32'hbbd7d729),
	.w5(32'h3bc90c6a),
	.w6(32'h3a2d0ee4),
	.w7(32'hbb6b55a7),
	.w8(32'hbb1bc3c8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fce82c),
	.w1(32'hbb01aea9),
	.w2(32'h3aba37aa),
	.w3(32'hbab1909b),
	.w4(32'hb9ae326c),
	.w5(32'h3aa23b60),
	.w6(32'h3a70fa2e),
	.w7(32'hbabbd410),
	.w8(32'h3b9267f7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf828a),
	.w1(32'h3bde81db),
	.w2(32'h3c45850e),
	.w3(32'hbb38fad6),
	.w4(32'h3ad702ae),
	.w5(32'hb9218cbd),
	.w6(32'hbb531195),
	.w7(32'h3a4232f0),
	.w8(32'hbbb49a5b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be85515),
	.w1(32'hb9fe04e4),
	.w2(32'hbacc06e0),
	.w3(32'hbb850b4c),
	.w4(32'hbb54f5af),
	.w5(32'h3b7b87d6),
	.w6(32'hbc0163eb),
	.w7(32'hba6e4150),
	.w8(32'h3ab065da),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d8f0),
	.w1(32'hbaa32227),
	.w2(32'h3b1a575c),
	.w3(32'h3ab8b21c),
	.w4(32'h3c181be8),
	.w5(32'hbbada16a),
	.w6(32'hbb8c8e2a),
	.w7(32'hba9186d8),
	.w8(32'hbbbc3dcc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2561d1),
	.w1(32'h3aa4d8b2),
	.w2(32'hbb50f926),
	.w3(32'hbc015cd1),
	.w4(32'hbb4f5397),
	.w5(32'hbb429352),
	.w6(32'h3b069490),
	.w7(32'hba166abc),
	.w8(32'hbb1e301d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecd3a7),
	.w1(32'h3b26edc9),
	.w2(32'h3b494a41),
	.w3(32'hbbb64d21),
	.w4(32'hbb03ea71),
	.w5(32'h3a92d4d9),
	.w6(32'hbb166dd2),
	.w7(32'hba8d4ef6),
	.w8(32'hbb5c5a98),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab032e1),
	.w1(32'hbb1925e6),
	.w2(32'hbaea798f),
	.w3(32'hba1cd6fc),
	.w4(32'hbb1af3cd),
	.w5(32'hbbaac716),
	.w6(32'h3a81de7d),
	.w7(32'h39d5deca),
	.w8(32'hb9042413),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb657b7),
	.w1(32'hbb3e6e36),
	.w2(32'hbbdf8639),
	.w3(32'hbb6f6119),
	.w4(32'hbba278e6),
	.w5(32'hbb3f57b4),
	.w6(32'hbc09d2c1),
	.w7(32'hba3854ce),
	.w8(32'hbb419240),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c24eb),
	.w1(32'h3c61560b),
	.w2(32'h3b0f37c9),
	.w3(32'hbc32bc21),
	.w4(32'h3b433ed9),
	.w5(32'hbc40a1e3),
	.w6(32'hbc0458dd),
	.w7(32'h3a8aa7a2),
	.w8(32'h3b04cbb7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b332e41),
	.w1(32'h3bd42b8f),
	.w2(32'h3bcd2e81),
	.w3(32'h39166a97),
	.w4(32'hbc0b2fd3),
	.w5(32'h3bd6748b),
	.w6(32'h3bcf4207),
	.w7(32'h3aad5f94),
	.w8(32'h3a5212c4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb914350),
	.w1(32'hba90b660),
	.w2(32'h3c31a1f5),
	.w3(32'hbb5c9c3b),
	.w4(32'hbbe36710),
	.w5(32'h3be510ec),
	.w6(32'hbca4eb47),
	.w7(32'hbc165903),
	.w8(32'hbb922126),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3a67b),
	.w1(32'hbbf213e6),
	.w2(32'hbad85be5),
	.w3(32'hbac98219),
	.w4(32'hbb5b177e),
	.w5(32'h3b48ce86),
	.w6(32'hbbc61444),
	.w7(32'hbbc5c834),
	.w8(32'h3a6a4b3a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7a965),
	.w1(32'h3b6712eb),
	.w2(32'h3c05ea7f),
	.w3(32'h3a3a25eb),
	.w4(32'h3b9fc524),
	.w5(32'hbb6fb98e),
	.w6(32'h3bbc002c),
	.w7(32'h3ba0c6dc),
	.w8(32'hbb632bed),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6afb8a),
	.w1(32'hba8b2023),
	.w2(32'hbb85c461),
	.w3(32'hbb02f269),
	.w4(32'hbb92d39d),
	.w5(32'hb9dc0ef4),
	.w6(32'h3b4814b4),
	.w7(32'hbb3ad1a7),
	.w8(32'h3a69cec8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc30fa),
	.w1(32'h39083e5b),
	.w2(32'hbba22850),
	.w3(32'h3b5e4292),
	.w4(32'h3abc7062),
	.w5(32'hbc3147c4),
	.w6(32'h3c1d2fdf),
	.w7(32'hb9be07e9),
	.w8(32'h3b16107d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1b71),
	.w1(32'h3a7e2831),
	.w2(32'hbc3f271c),
	.w3(32'hba32f1f0),
	.w4(32'hbc75d6b5),
	.w5(32'hba843d2a),
	.w6(32'hba4953aa),
	.w7(32'h37d8e430),
	.w8(32'hbc0aa945),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a825b1b),
	.w1(32'hbb676c7c),
	.w2(32'h3b182380),
	.w3(32'hba7e16d8),
	.w4(32'h398193f9),
	.w5(32'hba95b50e),
	.w6(32'h3ac7fecc),
	.w7(32'hba87ea72),
	.w8(32'hbb670abd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfa75e),
	.w1(32'h3b0ce6d9),
	.w2(32'hbbd794a7),
	.w3(32'hb9b064bd),
	.w4(32'hbb727289),
	.w5(32'h39f53e5c),
	.w6(32'hbc2aad21),
	.w7(32'hbc107875),
	.w8(32'h3bcd57d3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46b135),
	.w1(32'h3b20175f),
	.w2(32'hbb6e8478),
	.w3(32'h3b73449f),
	.w4(32'hbb76a777),
	.w5(32'h3b83fdf8),
	.w6(32'h3c186516),
	.w7(32'hbb133967),
	.w8(32'h3bdec9fc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc7868),
	.w1(32'h3c3a819f),
	.w2(32'h3b945453),
	.w3(32'h3c857ed4),
	.w4(32'h3c342871),
	.w5(32'h3aa95841),
	.w6(32'h3cb0d85e),
	.w7(32'h3c8aacc3),
	.w8(32'h3c0bca50),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9e0c8),
	.w1(32'h3b8274c8),
	.w2(32'h3ba2ea8b),
	.w3(32'h3ba280c1),
	.w4(32'h3b94df0b),
	.w5(32'h3b27c046),
	.w6(32'h3b73745c),
	.w7(32'h3b6addb4),
	.w8(32'h3af2b251),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca3bab),
	.w1(32'h3bd0391d),
	.w2(32'h3b2ff072),
	.w3(32'h3c145f7e),
	.w4(32'h3b1773f9),
	.w5(32'hba1d8d1f),
	.w6(32'h3c4a5359),
	.w7(32'h3bb18d29),
	.w8(32'hbbea63fc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08ade6),
	.w1(32'hb97b7340),
	.w2(32'h3a1fd9d8),
	.w3(32'hbbf35999),
	.w4(32'hbbee24bd),
	.w5(32'hbc24c25a),
	.w6(32'hbbcd9bd5),
	.w7(32'h38980733),
	.w8(32'hbba98f64),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d60de),
	.w1(32'hbbbc980c),
	.w2(32'hbc0e1679),
	.w3(32'hbbd5aa7f),
	.w4(32'hbb891860),
	.w5(32'hba430d8d),
	.w6(32'hbb365eda),
	.w7(32'hbb121a43),
	.w8(32'h39cb84ad),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa79dcf),
	.w1(32'hb98deda5),
	.w2(32'hbb86c9c3),
	.w3(32'hbb42ac2c),
	.w4(32'h3a4738b5),
	.w5(32'hbab0774c),
	.w6(32'hbaedb5d4),
	.w7(32'hbaff37fb),
	.w8(32'h39642971),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ce0d7),
	.w1(32'h3b3c1a89),
	.w2(32'h3bb3100c),
	.w3(32'h3a64e82e),
	.w4(32'h3b82de1c),
	.w5(32'hbb2529cd),
	.w6(32'h3c3600ab),
	.w7(32'h3b2be05e),
	.w8(32'h39cc93e8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21824f),
	.w1(32'h3a0ed615),
	.w2(32'h3b7be046),
	.w3(32'h3ab265f0),
	.w4(32'hbb155725),
	.w5(32'h3ba81555),
	.w6(32'hbab3ca0c),
	.w7(32'h3a2ba025),
	.w8(32'h3b3629af),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b312b45),
	.w1(32'h3a0a1092),
	.w2(32'hbb0fc434),
	.w3(32'h3a6c571e),
	.w4(32'h3b611f40),
	.w5(32'h3bcf04e4),
	.w6(32'hba9c49c3),
	.w7(32'hba507636),
	.w8(32'h3b8b73ab),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9e581),
	.w1(32'h3b4d9028),
	.w2(32'h3bd8fa3c),
	.w3(32'h3ba6e904),
	.w4(32'h3bcd4ec6),
	.w5(32'h3b095a57),
	.w6(32'h3ba76177),
	.w7(32'h3bad515a),
	.w8(32'h3ad6370f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeda0f),
	.w1(32'h3b533a42),
	.w2(32'h3c08f759),
	.w3(32'h3a956c60),
	.w4(32'h3b84f08a),
	.w5(32'hba90f424),
	.w6(32'h3bb1700e),
	.w7(32'h38a0046d),
	.w8(32'hb9a0863f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b365ead),
	.w1(32'h3bc462b2),
	.w2(32'h3b3d89c1),
	.w3(32'h3b8e9ef0),
	.w4(32'h39e90544),
	.w5(32'h3b99f335),
	.w6(32'h3c10a88f),
	.w7(32'h3b2fa568),
	.w8(32'hb9d21b3e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128c1c),
	.w1(32'hbb0d4211),
	.w2(32'hbb70fb8c),
	.w3(32'h3be8fcff),
	.w4(32'h3b9f65c5),
	.w5(32'h3af93a56),
	.w6(32'hbc40a45d),
	.w7(32'hbbb3a7bc),
	.w8(32'h3aaaed8a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92ef62),
	.w1(32'h3c05cfdb),
	.w2(32'h3ba2e4b2),
	.w3(32'h3bd929b8),
	.w4(32'h3b3922e1),
	.w5(32'h3afbdddd),
	.w6(32'h3bc9fe44),
	.w7(32'h3becf4b3),
	.w8(32'h3bc4a553),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49bdd0),
	.w1(32'h3c12fb5d),
	.w2(32'h3b662a12),
	.w3(32'h3bfdd0a3),
	.w4(32'h3a87a010),
	.w5(32'h3b56511e),
	.w6(32'h3bc9a6aa),
	.w7(32'h3a00c68d),
	.w8(32'hbba5c281),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13181f),
	.w1(32'h39699cef),
	.w2(32'hbb3ae31d),
	.w3(32'hb6d383be),
	.w4(32'hba9d692f),
	.w5(32'h3b688260),
	.w6(32'hbc186f98),
	.w7(32'hbb93be30),
	.w8(32'h374b5c5f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba391b6d),
	.w1(32'hba9fea78),
	.w2(32'h397a4ed9),
	.w3(32'hb9c5c8b2),
	.w4(32'hbac31e7f),
	.w5(32'h3ba38639),
	.w6(32'h3b4731f2),
	.w7(32'h3aa11de9),
	.w8(32'h3adf6485),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38532917),
	.w1(32'hbb273ff5),
	.w2(32'h3be3c7e4),
	.w3(32'h39a10649),
	.w4(32'h3b408c87),
	.w5(32'h3b8f27b6),
	.w6(32'h3b603743),
	.w7(32'h3b9c8a62),
	.w8(32'hba1c4e23),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83a562),
	.w1(32'h3ab64d63),
	.w2(32'hba092153),
	.w3(32'h3b378748),
	.w4(32'h3b55bf82),
	.w5(32'h389869dc),
	.w6(32'hbbaa892d),
	.w7(32'hbb3de077),
	.w8(32'h3b31c3c6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40046d),
	.w1(32'h3bcbac2e),
	.w2(32'hbbaa6824),
	.w3(32'h3c161545),
	.w4(32'h3a1cf282),
	.w5(32'hba9b32df),
	.w6(32'h3c8c73de),
	.w7(32'h3a747d7b),
	.w8(32'hbb1050ee),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072335),
	.w1(32'h3c1ddde8),
	.w2(32'h3b0aeaa0),
	.w3(32'h3c0f285b),
	.w4(32'h3b0ec139),
	.w5(32'h3a6853b0),
	.w6(32'h3c266967),
	.w7(32'h3c3c03af),
	.w8(32'h3b960bd8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba65107),
	.w1(32'h3b8cc9a8),
	.w2(32'h3a722cbc),
	.w3(32'h3bb3c522),
	.w4(32'h3adc9585),
	.w5(32'hbb01ae73),
	.w6(32'h3c1ec489),
	.w7(32'h3bded0af),
	.w8(32'h3bb2be34),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0da12),
	.w1(32'h3b7aaf82),
	.w2(32'h3ad88d17),
	.w3(32'h38fe7d64),
	.w4(32'hbb970226),
	.w5(32'hb993b799),
	.w6(32'hba288e35),
	.w7(32'h3aefe460),
	.w8(32'h3b119d4b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f3e5),
	.w1(32'h3b98ac71),
	.w2(32'hb912f941),
	.w3(32'h3b3f8a47),
	.w4(32'hba2a59fb),
	.w5(32'h3a14f2f3),
	.w6(32'h3c5a7f02),
	.w7(32'h3b9b96cd),
	.w8(32'h3bd9658b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b47aa),
	.w1(32'h3baad49d),
	.w2(32'hbb6c83c3),
	.w3(32'hba127323),
	.w4(32'h3b60f181),
	.w5(32'hbb95695e),
	.w6(32'hbb1faa9a),
	.w7(32'h3b5b2031),
	.w8(32'hbaa38b06),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b670c),
	.w1(32'hbae7668d),
	.w2(32'hbba9d4ee),
	.w3(32'hbb3a7672),
	.w4(32'hbaf0e12e),
	.w5(32'h3a5aff14),
	.w6(32'hbc315208),
	.w7(32'hbae226ca),
	.w8(32'hbb854840),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb82be0),
	.w1(32'hba3dedc8),
	.w2(32'h3b895b6e),
	.w3(32'hbaa02f39),
	.w4(32'hbb8c8227),
	.w5(32'hbafc29ed),
	.w6(32'hbb6ebcf9),
	.w7(32'hbb1d8ead),
	.w8(32'h3a979ece),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbca96),
	.w1(32'h3b9bcba3),
	.w2(32'hb969f675),
	.w3(32'h3a9a32ae),
	.w4(32'h3a5b8fa3),
	.w5(32'h3b67143f),
	.w6(32'h3b6963c0),
	.w7(32'hba852229),
	.w8(32'hba80dc04),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada7902),
	.w1(32'h3b83bfea),
	.w2(32'h3ba5b43e),
	.w3(32'h3baf7698),
	.w4(32'h3c02f3f9),
	.w5(32'h3a9a33c0),
	.w6(32'h3a04772c),
	.w7(32'h3b7dc0dd),
	.w8(32'h3aabd951),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f2ff3),
	.w1(32'h3c18f2d7),
	.w2(32'h3b1f0038),
	.w3(32'h3c13bd8a),
	.w4(32'h3c526dfd),
	.w5(32'hbb19f396),
	.w6(32'h3bffbc16),
	.w7(32'h3c3d0842),
	.w8(32'hbbab0b4f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf5f8f),
	.w1(32'hbc0b39e3),
	.w2(32'hbbaa5a8b),
	.w3(32'hbba7cca4),
	.w4(32'hbb9484f6),
	.w5(32'hbae615a0),
	.w6(32'hbbd2d64d),
	.w7(32'hbbbbad5b),
	.w8(32'hba59de16),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0852),
	.w1(32'h3a89e30c),
	.w2(32'hbb6f1802),
	.w3(32'hb954148f),
	.w4(32'h3b86703c),
	.w5(32'hbb5410f7),
	.w6(32'h3b2f85e1),
	.w7(32'h3b7a31d2),
	.w8(32'h3b5a14fd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80db59),
	.w1(32'h3c24cb80),
	.w2(32'h3a0c073e),
	.w3(32'h3afa96c7),
	.w4(32'hbb5c5c79),
	.w5(32'h3bb960b5),
	.w6(32'h3b71a57f),
	.w7(32'h39814564),
	.w8(32'h3b95ef63),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d2578),
	.w1(32'h3c342a00),
	.w2(32'h3c2cc9fb),
	.w3(32'h3c411c1a),
	.w4(32'h3c31b24d),
	.w5(32'hbaee8aaf),
	.w6(32'h3c6fe4bb),
	.w7(32'h3bed42f2),
	.w8(32'hbbfbd981),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae80cd),
	.w1(32'hbb5c60db),
	.w2(32'hbb626de1),
	.w3(32'h39c2f8ec),
	.w4(32'hba2a0102),
	.w5(32'hbb3c0b48),
	.w6(32'h38919979),
	.w7(32'hba8a500c),
	.w8(32'hb9e88c28),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b441e02),
	.w1(32'hbab27ed7),
	.w2(32'h3909f8c8),
	.w3(32'hbb2bbe3c),
	.w4(32'h3baa4e6b),
	.w5(32'hbb29d4b0),
	.w6(32'h39234f23),
	.w7(32'h3b5ab137),
	.w8(32'hbae0c545),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a6017),
	.w1(32'hbbe96c6b),
	.w2(32'hbb910ae1),
	.w3(32'hbbfa3ccc),
	.w4(32'hba8b4ef2),
	.w5(32'h3b5756ad),
	.w6(32'hbc05e914),
	.w7(32'hbaf9379d),
	.w8(32'hb8dec28a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb0c8e),
	.w1(32'hb99905d6),
	.w2(32'h3a3ccb0d),
	.w3(32'h3ba4d701),
	.w4(32'h3b90c3a7),
	.w5(32'hb8e92e49),
	.w6(32'hb9f7d259),
	.w7(32'h39e90764),
	.w8(32'hb9c3bda5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee9ffc),
	.w1(32'h3bac04f6),
	.w2(32'h3b1ff70f),
	.w3(32'hbb62e93a),
	.w4(32'h3b823fcc),
	.w5(32'hbbdf8ac8),
	.w6(32'hbc269fe0),
	.w7(32'hbadb8a12),
	.w8(32'hbb7429b7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8373e74),
	.w1(32'hbb87cb9a),
	.w2(32'hb94487bf),
	.w3(32'hbbc668ff),
	.w4(32'hbbca00c4),
	.w5(32'h3b28ee15),
	.w6(32'h39cfd6c3),
	.w7(32'hbb96fef5),
	.w8(32'hbb4980e9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8940),
	.w1(32'h3b1fdef8),
	.w2(32'h3b820691),
	.w3(32'h3b490ac5),
	.w4(32'h3b25b2ef),
	.w5(32'h3a99158c),
	.w6(32'hbbffceb1),
	.w7(32'hbb236ba0),
	.w8(32'h3b569dc3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babfc1e),
	.w1(32'h3c0fabab),
	.w2(32'h3b7f631f),
	.w3(32'h3be0ae39),
	.w4(32'hbabbbd5e),
	.w5(32'h3b2def4b),
	.w6(32'h3bc6adc9),
	.w7(32'h3ae38d59),
	.w8(32'h3b6854e6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba17dc5),
	.w1(32'h3ac63f7e),
	.w2(32'hba66f2b0),
	.w3(32'h3c104276),
	.w4(32'h3b953c82),
	.w5(32'hb9714709),
	.w6(32'h3c76bdc2),
	.w7(32'h3c3dcbe5),
	.w8(32'h3bf98faa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0623d1),
	.w1(32'h3b1cff14),
	.w2(32'h3c189057),
	.w3(32'hbbc540d5),
	.w4(32'h397d1dc8),
	.w5(32'h3ba0c2ee),
	.w6(32'hbbca2874),
	.w7(32'h3b3c4b2e),
	.w8(32'h3ab5d72f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88e37d),
	.w1(32'hbb27ce5a),
	.w2(32'hbb9ce24f),
	.w3(32'hbb43989b),
	.w4(32'h3b150ca5),
	.w5(32'hb84240e1),
	.w6(32'h3a9616e5),
	.w7(32'hba49884d),
	.w8(32'hbb75ac4f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb9765),
	.w1(32'hbb2f0bb6),
	.w2(32'h3b6add3e),
	.w3(32'hba1637b7),
	.w4(32'h3b2e78f4),
	.w5(32'h3852ec77),
	.w6(32'hb7f73c62),
	.w7(32'h3bb999d9),
	.w8(32'h3be03d55),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032023),
	.w1(32'h3c6e6ee1),
	.w2(32'h3bb25062),
	.w3(32'h3c6bb1a4),
	.w4(32'h3b247dc8),
	.w5(32'hba98d82d),
	.w6(32'h3caba59a),
	.w7(32'h3c4fb0ec),
	.w8(32'h3bb70fec),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b442f89),
	.w1(32'h3b29703f),
	.w2(32'hbb43562d),
	.w3(32'h3ad4188a),
	.w4(32'hbb7171c6),
	.w5(32'hbb1c7714),
	.w6(32'h3bb77d3e),
	.w7(32'hba3a093c),
	.w8(32'hba9e17ea),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ccc30),
	.w1(32'h3b8c16bd),
	.w2(32'hbabdc175),
	.w3(32'h3ad2ad3d),
	.w4(32'hba8c3f12),
	.w5(32'h3c33ddc5),
	.w6(32'h3a86887d),
	.w7(32'hbc4b4eb6),
	.w8(32'hbb1ec673),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38bf07),
	.w1(32'hbb662ca0),
	.w2(32'h3bb2ecbd),
	.w3(32'hb901bfe3),
	.w4(32'h3b681744),
	.w5(32'hbb961016),
	.w6(32'hbbab99d0),
	.w7(32'h3a422cc9),
	.w8(32'hbb9b3f27),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dac97),
	.w1(32'hb980cb2e),
	.w2(32'hbbf884ed),
	.w3(32'hbbac32b4),
	.w4(32'hbba6eada),
	.w5(32'hbba18ce2),
	.w6(32'h3b19672a),
	.w7(32'hb954ca5e),
	.w8(32'hb9c411fb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9bccd),
	.w1(32'h3a94f55d),
	.w2(32'hbb41a1f8),
	.w3(32'h3a9d0809),
	.w4(32'hbb8c9e82),
	.w5(32'h3b7f95ad),
	.w6(32'hba7742c5),
	.w7(32'hbba1ec4a),
	.w8(32'h3b235a10),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0bd29),
	.w1(32'h3c853049),
	.w2(32'h3ba35c97),
	.w3(32'h3c34a016),
	.w4(32'h3c860dc9),
	.w5(32'hbb12a0c9),
	.w6(32'h3c711c40),
	.w7(32'h3bf0b134),
	.w8(32'hbb2f31ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd991ad),
	.w1(32'h3c056597),
	.w2(32'h3bcffbd0),
	.w3(32'hbba7bac1),
	.w4(32'hbae4bb37),
	.w5(32'h3bb9d415),
	.w6(32'hbbc05f9a),
	.w7(32'hbbdd741e),
	.w8(32'hbb1a0c4f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4e781),
	.w1(32'h3a78fba3),
	.w2(32'h3a81c25c),
	.w3(32'hbb5f3bdf),
	.w4(32'hbbaf1330),
	.w5(32'hba972f06),
	.w6(32'hbbdb4c32),
	.w7(32'hbb1a9742),
	.w8(32'hbb76c90e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46beb2),
	.w1(32'h3b914b5f),
	.w2(32'h393874b3),
	.w3(32'hbc0bb38c),
	.w4(32'h3b88ab1a),
	.w5(32'hbb2916e1),
	.w6(32'hb9e97b33),
	.w7(32'hba938405),
	.w8(32'h3a952f53),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbacaf1),
	.w1(32'h3babecfc),
	.w2(32'hba5fd4ae),
	.w3(32'h3b2eaf13),
	.w4(32'h390ca304),
	.w5(32'hbb06deb0),
	.w6(32'h3ac8ea02),
	.w7(32'h369eeec8),
	.w8(32'h3b8f4077),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8763e2),
	.w1(32'h3c984add),
	.w2(32'h3cad8d4e),
	.w3(32'h3bdfbc70),
	.w4(32'h3c5794a7),
	.w5(32'h3b018f2c),
	.w6(32'h3bba754d),
	.w7(32'h3c3d0db9),
	.w8(32'h3b9940d9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1996a),
	.w1(32'h391ac05a),
	.w2(32'h3b194460),
	.w3(32'hbb8ec54b),
	.w4(32'hbaca60de),
	.w5(32'hbadf7b4b),
	.w6(32'h3a444eae),
	.w7(32'hbb9cc163),
	.w8(32'h3aaa912d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ae470),
	.w1(32'hb9b49b1c),
	.w2(32'hb9ef0e0f),
	.w3(32'h3b88eb80),
	.w4(32'hbbc08c4d),
	.w5(32'hba734ab1),
	.w6(32'h3c3facdf),
	.w7(32'hbbd46a79),
	.w8(32'hbabf6cc0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7d00),
	.w1(32'h3ad9a655),
	.w2(32'h3afd2b11),
	.w3(32'h3a19ebda),
	.w4(32'hba297264),
	.w5(32'hbac757e1),
	.w6(32'h3bcf933e),
	.w7(32'h3a0d3ab6),
	.w8(32'hbb3b62c3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80fcdb),
	.w1(32'hbb12b762),
	.w2(32'hbb905069),
	.w3(32'h39f1114c),
	.w4(32'hbbcd20d3),
	.w5(32'hbb382ed2),
	.w6(32'hbb09e263),
	.w7(32'hbb4845bb),
	.w8(32'hba4d8ae1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c44a),
	.w1(32'hb9b832aa),
	.w2(32'h3a698d8c),
	.w3(32'hbb5cd193),
	.w4(32'hbb47ead8),
	.w5(32'h3b301929),
	.w6(32'hbb7769c1),
	.w7(32'hbb30250a),
	.w8(32'h3b940af0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba9767),
	.w1(32'h3b42dc86),
	.w2(32'h3c171063),
	.w3(32'h3c06bfb1),
	.w4(32'hb8a2d19f),
	.w5(32'h3a372066),
	.w6(32'h3c02c7a1),
	.w7(32'h3b29e6b1),
	.w8(32'h3a2e78af),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad99456),
	.w1(32'h3a95bb2d),
	.w2(32'h3b1ff3b8),
	.w3(32'hbb022264),
	.w4(32'hbb8e2ff7),
	.w5(32'h3ad6dc23),
	.w6(32'hbab3fb9c),
	.w7(32'hbb12608c),
	.w8(32'h3b247338),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1974c),
	.w1(32'hbb519082),
	.w2(32'hb9f4e89e),
	.w3(32'h3bafe308),
	.w4(32'h3bc28179),
	.w5(32'hba023125),
	.w6(32'h3ab87461),
	.w7(32'hba8613b5),
	.w8(32'hbb80f97c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06340e),
	.w1(32'h3ba09139),
	.w2(32'h3947f6d8),
	.w3(32'h3b317b95),
	.w4(32'h3bcac989),
	.w5(32'hb985c400),
	.w6(32'h3aa91959),
	.w7(32'h3b30acbb),
	.w8(32'hbb6d0654),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b573d),
	.w1(32'hba486751),
	.w2(32'h3a232fa0),
	.w3(32'h383941a9),
	.w4(32'h3a4c6191),
	.w5(32'h3a5a9873),
	.w6(32'hbab0ff9e),
	.w7(32'hb9ab943b),
	.w8(32'h3aef1533),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0c5c4),
	.w1(32'h3b34f5bc),
	.w2(32'h3af875b5),
	.w3(32'h3ae2172b),
	.w4(32'h3709ccb4),
	.w5(32'h3b3c9118),
	.w6(32'h3aa1ddb5),
	.w7(32'hba158394),
	.w8(32'h3aa3a5c2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b040ac1),
	.w1(32'h3b03fb26),
	.w2(32'h3abed9d7),
	.w3(32'h3a88a772),
	.w4(32'h3aa1c851),
	.w5(32'hbadbff3a),
	.w6(32'hba169e1d),
	.w7(32'h3a708c28),
	.w8(32'h3a923bb2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b508c28),
	.w1(32'h3ad5eeba),
	.w2(32'h399bf6a2),
	.w3(32'hbb17e361),
	.w4(32'hbb05ee7d),
	.w5(32'hbb49e162),
	.w6(32'hb782f7e9),
	.w7(32'hbb333702),
	.w8(32'h3a1d7df4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96e012),
	.w1(32'hbac7510e),
	.w2(32'hbae3740a),
	.w3(32'hbb0ba24d),
	.w4(32'hb9dd5b6f),
	.w5(32'h3a61462d),
	.w6(32'h3a403ed9),
	.w7(32'hbb06a51d),
	.w8(32'hba944d66),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a7ff1),
	.w1(32'h3b4f1968),
	.w2(32'h3970e850),
	.w3(32'h3ae136f6),
	.w4(32'hb929f189),
	.w5(32'hbad754e2),
	.w6(32'hbb294eec),
	.w7(32'hb92dd1fc),
	.w8(32'hbaab69e5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb930),
	.w1(32'hbaba1f15),
	.w2(32'hbb3bb3ba),
	.w3(32'h39193f9e),
	.w4(32'hba897a52),
	.w5(32'hba99a45f),
	.w6(32'h394da1b5),
	.w7(32'h39a44fd0),
	.w8(32'hbae8b2dd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2afc65),
	.w1(32'h3a48e94b),
	.w2(32'hbab9ee11),
	.w3(32'hbaffa68e),
	.w4(32'h3b2ef208),
	.w5(32'hba7f9190),
	.w6(32'h3bbcea2e),
	.w7(32'h3b5fbdc9),
	.w8(32'hbad2dd41),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39854828),
	.w1(32'hbacfff3e),
	.w2(32'h3bcb60da),
	.w3(32'hbba2015c),
	.w4(32'hbbc0c90d),
	.w5(32'hba651e54),
	.w6(32'hbc0d0f04),
	.w7(32'hbbade986),
	.w8(32'hba8565e1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a280066),
	.w1(32'hbb463993),
	.w2(32'hba6614a8),
	.w3(32'hbb2885bb),
	.w4(32'h3b6ffc0d),
	.w5(32'hba8b5591),
	.w6(32'hbabfee0e),
	.w7(32'h3b264df3),
	.w8(32'hbb282ec6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71ad1a),
	.w1(32'hba61d553),
	.w2(32'h390975a7),
	.w3(32'hbacbb452),
	.w4(32'hb9ce0ea8),
	.w5(32'hba355497),
	.w6(32'hbb51e05e),
	.w7(32'hbb54c475),
	.w8(32'hbb2cf567),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40776f),
	.w1(32'hbaa9d432),
	.w2(32'hba407061),
	.w3(32'hb8b06a69),
	.w4(32'hba6a617d),
	.w5(32'h3aad7f74),
	.w6(32'hbac89f13),
	.w7(32'hb98de698),
	.w8(32'h3a9e9266),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c70ed),
	.w1(32'h380f2a7d),
	.w2(32'h3a6fe266),
	.w3(32'h39b01a05),
	.w4(32'h3a74ad8f),
	.w5(32'hbb2ac970),
	.w6(32'h39aaccc4),
	.w7(32'h3a6b6103),
	.w8(32'hbb90ebda),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe22d8e),
	.w1(32'hbbc1d852),
	.w2(32'hbad4025a),
	.w3(32'hbadbf2fb),
	.w4(32'h3b779346),
	.w5(32'h3b2a4718),
	.w6(32'h3a6d4b8c),
	.w7(32'hbb97796f),
	.w8(32'h3b68cf69),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932710e),
	.w1(32'hbab3c689),
	.w2(32'hbb9f218c),
	.w3(32'h397f674c),
	.w4(32'hbb47cb87),
	.w5(32'hbbabebe7),
	.w6(32'h3bc49e9a),
	.w7(32'hba1cb2b8),
	.w8(32'hbafed803),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989c385),
	.w1(32'hba9e1649),
	.w2(32'hb9dc1ccb),
	.w3(32'h398c98a7),
	.w4(32'h3a93c527),
	.w5(32'hbabc4253),
	.w6(32'h3aa45b5f),
	.w7(32'h3a562318),
	.w8(32'h3a4982a3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52cb2c),
	.w1(32'h3b8e108e),
	.w2(32'h3b825395),
	.w3(32'h3b56a214),
	.w4(32'h3b4d5c9c),
	.w5(32'h3af04d2c),
	.w6(32'h3c35180b),
	.w7(32'h3b7c0815),
	.w8(32'h3bab45c6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a59b),
	.w1(32'h3b2540d3),
	.w2(32'h3b103078),
	.w3(32'h3a5e42c0),
	.w4(32'hba230cd7),
	.w5(32'hba887ad7),
	.w6(32'hba617beb),
	.w7(32'hb93700f2),
	.w8(32'hba847134),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7efb3),
	.w1(32'hba9d184c),
	.w2(32'hbb2390cf),
	.w3(32'h390839cb),
	.w4(32'hba03bab5),
	.w5(32'hba0fba32),
	.w6(32'hbafa7149),
	.w7(32'hbb2dae72),
	.w8(32'h3a97a282),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835244),
	.w1(32'h3acc9cea),
	.w2(32'hb9687be2),
	.w3(32'h3ae1fd25),
	.w4(32'hbb192894),
	.w5(32'h3926be8c),
	.w6(32'h3abec2d6),
	.w7(32'hb9c35cd7),
	.w8(32'hbb1a0759),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c9c5),
	.w1(32'h3b04ee3f),
	.w2(32'hba775d73),
	.w3(32'h3bea2748),
	.w4(32'h3bbab2b5),
	.w5(32'h39e6e0c8),
	.w6(32'h3c1d896d),
	.w7(32'h3b8e10c9),
	.w8(32'h3bc3d382),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b430140),
	.w1(32'h3b8d9121),
	.w2(32'h3b9bc10b),
	.w3(32'hbadbd390),
	.w4(32'hbb240a9e),
	.w5(32'h3a914e84),
	.w6(32'hbb055967),
	.w7(32'hba393382),
	.w8(32'h39a488e9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892a2e),
	.w1(32'h3ad3e924),
	.w2(32'hbb07b028),
	.w3(32'h39eb789d),
	.w4(32'hb9354540),
	.w5(32'h39d68824),
	.w6(32'h3b34838e),
	.w7(32'h39d1874c),
	.w8(32'h3a72d93f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85015e),
	.w1(32'h3b43e23d),
	.w2(32'hbaef1b0c),
	.w3(32'h3b880af4),
	.w4(32'h3b7b32e5),
	.w5(32'hba3c1c4e),
	.w6(32'h3bba0461),
	.w7(32'h3b7dc308),
	.w8(32'h3b880a83),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bb952),
	.w1(32'h3b580def),
	.w2(32'h3b46029f),
	.w3(32'h3b6ffe23),
	.w4(32'h3b29720c),
	.w5(32'hbb4f8a47),
	.w6(32'h3b312dfd),
	.w7(32'h3b2ea755),
	.w8(32'hbbaad055),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c578fa),
	.w1(32'hba5abab0),
	.w2(32'hbb70c471),
	.w3(32'hbb1ebdf3),
	.w4(32'hbb1371a0),
	.w5(32'hbb3050f2),
	.w6(32'h3c31dd77),
	.w7(32'hbba8fc03),
	.w8(32'hb6cc85f7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace63f1),
	.w1(32'h3b0bb9d3),
	.w2(32'h3ade944c),
	.w3(32'h3b48499b),
	.w4(32'h3a85bc37),
	.w5(32'h3ab794fd),
	.w6(32'h3b6d9473),
	.w7(32'h3b601e02),
	.w8(32'h3ad5e664),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd36a38),
	.w1(32'h3ba099e2),
	.w2(32'h3b967af8),
	.w3(32'hbb024ed3),
	.w4(32'hbb2e369d),
	.w5(32'h3bc56240),
	.w6(32'hbc0163fd),
	.w7(32'hbc2dbeee),
	.w8(32'h3b52dc7f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a808d),
	.w1(32'h3bbf6658),
	.w2(32'h3ba6452e),
	.w3(32'h3bcb7adf),
	.w4(32'h3b96bd36),
	.w5(32'h382311f9),
	.w6(32'h3bb9fc31),
	.w7(32'h3b72b03d),
	.w8(32'h39988cf5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ff86b),
	.w1(32'hbb5edc11),
	.w2(32'hbb5ed3bd),
	.w3(32'hba96fa7e),
	.w4(32'hbabac602),
	.w5(32'hbaa3df08),
	.w6(32'h3a66eb49),
	.w7(32'hbb40d07d),
	.w8(32'hbb114c52),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2cfa),
	.w1(32'hbaa504cb),
	.w2(32'hb7e73cff),
	.w3(32'hba5a0496),
	.w4(32'h39181b5b),
	.w5(32'hba552985),
	.w6(32'h3aeb16ae),
	.w7(32'h39945406),
	.w8(32'h3aa09d8a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c6065),
	.w1(32'h3a08838a),
	.w2(32'hbb08b978),
	.w3(32'h3a2e8d74),
	.w4(32'hba4e641c),
	.w5(32'h3ba28022),
	.w6(32'h3b13c8aa),
	.w7(32'hbafb3852),
	.w8(32'h3c2df5b2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe842b),
	.w1(32'h3b5b4bbb),
	.w2(32'h3b9920a8),
	.w3(32'h3bb62800),
	.w4(32'h3b6748a5),
	.w5(32'hb8c0bf9d),
	.w6(32'h3ab307e6),
	.w7(32'h3b512963),
	.w8(32'hb69a1e70),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91de9b),
	.w1(32'hba32c287),
	.w2(32'hbb6d4ecd),
	.w3(32'hba21cc84),
	.w4(32'hba76379f),
	.w5(32'hbb73d1e6),
	.w6(32'h3a5e94ee),
	.w7(32'hbab5545f),
	.w8(32'hbb6ab2b5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804d7e),
	.w1(32'h3a16d892),
	.w2(32'hb9915d7d),
	.w3(32'h3903e2af),
	.w4(32'hba93ded8),
	.w5(32'h3b19c336),
	.w6(32'h3a7e7900),
	.w7(32'h3acd7c28),
	.w8(32'h3aaf2801),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b774b6c),
	.w1(32'h3a88369a),
	.w2(32'hbb54965f),
	.w3(32'h3a90a815),
	.w4(32'hbaeca243),
	.w5(32'hbb2a9c33),
	.w6(32'h390366ef),
	.w7(32'hb7d20e1f),
	.w8(32'hbae18d06),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bce0c4),
	.w1(32'hbafe3737),
	.w2(32'hbb5849e4),
	.w3(32'hbb18f870),
	.w4(32'hb948b35b),
	.w5(32'h392281a7),
	.w6(32'h384efd70),
	.w7(32'hba614c1e),
	.w8(32'h3b22f696),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d9648),
	.w1(32'h3a912ef8),
	.w2(32'hbb53b8dc),
	.w3(32'h3a7c4af9),
	.w4(32'hba92e72b),
	.w5(32'hbbef34fe),
	.w6(32'h3bcfb885),
	.w7(32'hb6e12be8),
	.w8(32'h38b0d3be),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f4e2),
	.w1(32'h3b592657),
	.w2(32'h3b4022cf),
	.w3(32'h3afe0494),
	.w4(32'hbc02c18e),
	.w5(32'h39fbc92b),
	.w6(32'hbb812636),
	.w7(32'hb94215f6),
	.w8(32'hbac0ffa6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9618f49),
	.w1(32'h3b8e2f5e),
	.w2(32'h3b9524e7),
	.w3(32'hb9cf8915),
	.w4(32'h3aa22e5e),
	.w5(32'h3b1fa238),
	.w6(32'h3a2b49ae),
	.w7(32'hb8c09147),
	.w8(32'h38135002),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc687b),
	.w1(32'h3a732865),
	.w2(32'hba85f6bd),
	.w3(32'h3a85da60),
	.w4(32'hbaa62184),
	.w5(32'hb9128757),
	.w6(32'h3b198fed),
	.w7(32'hbad664cb),
	.w8(32'hb9c4d15f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af66b8),
	.w1(32'hbb122582),
	.w2(32'hbb02c7c5),
	.w3(32'hbb5ed512),
	.w4(32'hbb462c52),
	.w5(32'hb912fb73),
	.w6(32'hbb208341),
	.w7(32'hbb32a293),
	.w8(32'hbb19ce10),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82308e),
	.w1(32'hb9d21e91),
	.w2(32'hb945eb47),
	.w3(32'h39e8c1ba),
	.w4(32'h3953070b),
	.w5(32'hbb3a3c62),
	.w6(32'hbb0091a7),
	.w7(32'hbb04f70b),
	.w8(32'hbb59db28),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f3d65),
	.w1(32'hba8ad4a2),
	.w2(32'h3b23136b),
	.w3(32'hbbaf242d),
	.w4(32'h39277771),
	.w5(32'h3b0ca90f),
	.w6(32'h3a107adc),
	.w7(32'h39de70b0),
	.w8(32'hba80a908),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9d6d9),
	.w1(32'h3b115af5),
	.w2(32'h3a8d8bba),
	.w3(32'h3ae7c1e1),
	.w4(32'h3b056c5d),
	.w5(32'hbb42ca0c),
	.w6(32'hbae71765),
	.w7(32'hba9450b2),
	.w8(32'hbb900458),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8765e),
	.w1(32'hbb9144e1),
	.w2(32'hb8ad8cd6),
	.w3(32'hbb33b623),
	.w4(32'hbb52ffac),
	.w5(32'h3bb7d26a),
	.w6(32'hbb6abd33),
	.w7(32'h3ad8b52b),
	.w8(32'h3bbbd1d8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43eaff),
	.w1(32'h3ab761e0),
	.w2(32'hbb51a429),
	.w3(32'h3b28fe72),
	.w4(32'h3b831d89),
	.w5(32'hbb813c6f),
	.w6(32'hbaa17199),
	.w7(32'h3b415f20),
	.w8(32'hbb039f3d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aac1bf),
	.w1(32'h3895d9d2),
	.w2(32'hbb421826),
	.w3(32'hb920533e),
	.w4(32'hbb856798),
	.w5(32'hbb1d2a9c),
	.w6(32'h3b886db0),
	.w7(32'hbbdcfca8),
	.w8(32'h3a30f78b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c013133),
	.w1(32'h3b44b070),
	.w2(32'h3aa8a548),
	.w3(32'h3a539bfd),
	.w4(32'hbb01c6ae),
	.w5(32'hbb1455b4),
	.w6(32'hba8c3b9e),
	.w7(32'hb97f4916),
	.w8(32'hb9d504ae),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48e285),
	.w1(32'h3ae368b7),
	.w2(32'hbb211a2b),
	.w3(32'h3b0d32a9),
	.w4(32'h3a95ea12),
	.w5(32'hba63be9d),
	.w6(32'h3babab5d),
	.w7(32'hba796dc9),
	.w8(32'h3a8b2241),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a389c),
	.w1(32'hbaaa8761),
	.w2(32'hbbd8def7),
	.w3(32'hbbc950c6),
	.w4(32'hbac57ad0),
	.w5(32'h3b1dbc21),
	.w6(32'hbba4906b),
	.w7(32'h3ac547b7),
	.w8(32'h3ba52d8c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d61ba8),
	.w1(32'h3acfc493),
	.w2(32'h39e36a5a),
	.w3(32'hb8c0446f),
	.w4(32'h39bdb1a8),
	.w5(32'hbad5a072),
	.w6(32'h393ca349),
	.w7(32'hba359087),
	.w8(32'hba5981b1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f89b41),
	.w1(32'hba02d0fc),
	.w2(32'hba8e81dd),
	.w3(32'hba589795),
	.w4(32'hb972bb65),
	.w5(32'hbb8b584e),
	.w6(32'hbb3ce25e),
	.w7(32'hba5d559a),
	.w8(32'hba061de2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0338ad),
	.w1(32'h39dff8e1),
	.w2(32'hbbbc2c13),
	.w3(32'hbb88e15e),
	.w4(32'hbc214045),
	.w5(32'h3b09152c),
	.w6(32'hbb450af3),
	.w7(32'hbbe28e69),
	.w8(32'hb8bfeee2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b308e),
	.w1(32'h3a0e930d),
	.w2(32'h39a87892),
	.w3(32'h3abd4dbb),
	.w4(32'h3b4bb4c8),
	.w5(32'hbb38b6f0),
	.w6(32'h3bf71fe0),
	.w7(32'h3b95932a),
	.w8(32'h3b1a7e43),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dfa1d2),
	.w1(32'h3aa975e6),
	.w2(32'hb9a934f6),
	.w3(32'h39850e08),
	.w4(32'h3982a0a9),
	.w5(32'hb9d85a7d),
	.w6(32'h3b0a72ff),
	.w7(32'h3a22017a),
	.w8(32'h3a408bd2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d9e45),
	.w1(32'hbb808774),
	.w2(32'h3a6df0a0),
	.w3(32'hbb98d269),
	.w4(32'hbacedd17),
	.w5(32'hba9048d0),
	.w6(32'hbb8644fa),
	.w7(32'hbbe7fe46),
	.w8(32'hbb8ee336),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4449),
	.w1(32'hbbc91224),
	.w2(32'h3b18049c),
	.w3(32'h39b73443),
	.w4(32'h3a9be6af),
	.w5(32'h3b2b4445),
	.w6(32'hbb413b4e),
	.w7(32'hbb80f7b0),
	.w8(32'hb9f6c868),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d9d8),
	.w1(32'hba087524),
	.w2(32'hbbcbab86),
	.w3(32'h3b9245af),
	.w4(32'hbb215cc1),
	.w5(32'h3ba68697),
	.w6(32'hbb15aa92),
	.w7(32'hbb2ab312),
	.w8(32'h3b23a38d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf66042),
	.w1(32'h3b9cf38c),
	.w2(32'h3b4a2127),
	.w3(32'h3ba8fc0f),
	.w4(32'h3b4c2d44),
	.w5(32'h3b816a2c),
	.w6(32'h3c01e127),
	.w7(32'h3a971cfc),
	.w8(32'h3ba1f4cc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c573),
	.w1(32'h3bcfcdfe),
	.w2(32'hb92d9403),
	.w3(32'h3c07abf2),
	.w4(32'h3b5f682f),
	.w5(32'hbaf5dba8),
	.w6(32'h3c7cb089),
	.w7(32'h3baf5ace),
	.w8(32'h3a2b32de),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2e43c),
	.w1(32'h3a0bb101),
	.w2(32'hb97f7ce6),
	.w3(32'hb95daefb),
	.w4(32'h3a93b448),
	.w5(32'hba7a25d6),
	.w6(32'hbaedeb0b),
	.w7(32'hb92b7514),
	.w8(32'hba3bb561),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2f380),
	.w1(32'h39c2b9af),
	.w2(32'h3ab1cbdf),
	.w3(32'h3ad68019),
	.w4(32'h3ad991db),
	.w5(32'h3b077c82),
	.w6(32'h3ad35f4b),
	.w7(32'h3ae35c35),
	.w8(32'hba7c9060),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985487),
	.w1(32'h3a143a05),
	.w2(32'hba5b4fe6),
	.w3(32'hba24ca85),
	.w4(32'hb9f6b815),
	.w5(32'h3b1a6978),
	.w6(32'hbb0cc460),
	.w7(32'hba43fb8a),
	.w8(32'h3b864a0a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dcc99),
	.w1(32'hbabc7f9b),
	.w2(32'hbb052085),
	.w3(32'h3b4cd33f),
	.w4(32'hbadb5446),
	.w5(32'hb974bb22),
	.w6(32'hba41f202),
	.w7(32'hbb5c9bdf),
	.w8(32'hba9a500c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba0e5a),
	.w1(32'h39e3e4c7),
	.w2(32'h3b71f262),
	.w3(32'hbae67e12),
	.w4(32'h3ab48029),
	.w5(32'h3aa2e970),
	.w6(32'hbaf98928),
	.w7(32'hba5d862b),
	.w8(32'h3b8ddc94),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8266ab),
	.w1(32'hba794f88),
	.w2(32'hbb36c431),
	.w3(32'h3bc26b50),
	.w4(32'hbb485097),
	.w5(32'h3948b39d),
	.w6(32'h3b9fb9b5),
	.w7(32'hbb38681a),
	.w8(32'h390baec5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c32f2),
	.w1(32'h3b7a26b9),
	.w2(32'hba50c884),
	.w3(32'hbaf0c441),
	.w4(32'h39939be0),
	.w5(32'hb9babe0b),
	.w6(32'h3ba8264e),
	.w7(32'hbaedf363),
	.w8(32'hb9d2a1a9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b31c2c),
	.w1(32'h3a017667),
	.w2(32'hba51cb4f),
	.w3(32'hba3fe9fa),
	.w4(32'h3af57b11),
	.w5(32'hba9e8c86),
	.w6(32'hba4f2f88),
	.w7(32'h3818cde1),
	.w8(32'hbade1d9c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b637367),
	.w1(32'h392ac8ce),
	.w2(32'h3af0b150),
	.w3(32'hbaf3f5c9),
	.w4(32'hba4e3197),
	.w5(32'h39a4f54b),
	.w6(32'hb9d6daec),
	.w7(32'h3a9e5dd3),
	.w8(32'h3aa8c5ee),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d62e7),
	.w1(32'h3b5e71a6),
	.w2(32'h3b141007),
	.w3(32'hbb96c9f0),
	.w4(32'h3b53fbb1),
	.w5(32'h3abe0fc7),
	.w6(32'hbb8ab8bb),
	.w7(32'h3b5d08e7),
	.w8(32'h3b57c9fa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a19bc),
	.w1(32'h3bd77e5f),
	.w2(32'h3afbefb7),
	.w3(32'h3ae01063),
	.w4(32'h3b1aade2),
	.w5(32'h3a8a9eb5),
	.w6(32'h3bedb669),
	.w7(32'h39b21cff),
	.w8(32'h38ec8dcc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01d55d),
	.w1(32'h3ad576e4),
	.w2(32'h3a4f33ef),
	.w3(32'hb95cd559),
	.w4(32'hb9d2eb05),
	.w5(32'h3bb874e2),
	.w6(32'h39b46771),
	.w7(32'hb8af1861),
	.w8(32'h3b826323),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed609f),
	.w1(32'h3a24b07e),
	.w2(32'hb99f9241),
	.w3(32'h3bf0ed2f),
	.w4(32'h3b287320),
	.w5(32'hbb24e4ab),
	.w6(32'h3b8ff8c6),
	.w7(32'h3bbf4a5a),
	.w8(32'h3b834f8e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbbaae),
	.w1(32'hbb2e0c1b),
	.w2(32'hbb33f852),
	.w3(32'h3ac3648b),
	.w4(32'hbc24d388),
	.w5(32'h3b001c9b),
	.w6(32'hba8783bf),
	.w7(32'hbbe61ef6),
	.w8(32'hbbba9360),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e3ffe),
	.w1(32'hb8a6a191),
	.w2(32'h3a7849ef),
	.w3(32'hbad63614),
	.w4(32'h3a4fb4bc),
	.w5(32'hbaf8e91e),
	.w6(32'h3abec001),
	.w7(32'h3a21ff01),
	.w8(32'h3b07f012),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebc57b),
	.w1(32'hb9649c14),
	.w2(32'h39ba36a8),
	.w3(32'h39bc34e9),
	.w4(32'hbaa79abb),
	.w5(32'hba97f3e8),
	.w6(32'hbadc8b7f),
	.w7(32'hb9f4d2bb),
	.w8(32'hbabf8bdc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa69985),
	.w1(32'h3a7afd04),
	.w2(32'h3b3f0b04),
	.w3(32'hbb279db7),
	.w4(32'h3ad29801),
	.w5(32'hba5c48f7),
	.w6(32'h39c8003f),
	.w7(32'h3a16c177),
	.w8(32'h3ac9e249),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20283c),
	.w1(32'h3b34ef83),
	.w2(32'h3b07a4c0),
	.w3(32'hba9583c5),
	.w4(32'h3a89635b),
	.w5(32'hbac34012),
	.w6(32'h39b4d88b),
	.w7(32'h3940b8cb),
	.w8(32'hb95ae8f6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06197),
	.w1(32'hbbe293b1),
	.w2(32'hba828b36),
	.w3(32'hbb230259),
	.w4(32'h3a3096c4),
	.w5(32'h390ea0f7),
	.w6(32'hbb914ea3),
	.w7(32'hba6206e6),
	.w8(32'h3b04e976),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f89f9),
	.w1(32'h3ae0a517),
	.w2(32'h3b2023ab),
	.w3(32'h3b0becee),
	.w4(32'hba19b05b),
	.w5(32'h3a97fe3b),
	.w6(32'h3b09aea6),
	.w7(32'h3ae2a0c0),
	.w8(32'hb8c4a30e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d3ec8),
	.w1(32'h3b7c600f),
	.w2(32'h3b7f108a),
	.w3(32'hb8f19500),
	.w4(32'h3ae33380),
	.w5(32'h39b1c59f),
	.w6(32'hbafd2e32),
	.w7(32'hbad9c122),
	.w8(32'hbb416ea7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96bf31),
	.w1(32'hb8684902),
	.w2(32'hbb43be39),
	.w3(32'hba189770),
	.w4(32'hba8e2994),
	.w5(32'hbb801f72),
	.w6(32'hbaa4c729),
	.w7(32'hb96431cd),
	.w8(32'hba0756a6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae86841),
	.w1(32'hbbe77219),
	.w2(32'hbbad098c),
	.w3(32'h3ae2dda8),
	.w4(32'hbc04ed71),
	.w5(32'h39f022a9),
	.w6(32'h3a903e9e),
	.w7(32'hbb6ac455),
	.w8(32'h3b17b9f1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0abbb1),
	.w1(32'h3b492437),
	.w2(32'h3a71ff87),
	.w3(32'hbb126b3d),
	.w4(32'h3a9af32d),
	.w5(32'hbb32e3da),
	.w6(32'hbb671b85),
	.w7(32'hbb01c270),
	.w8(32'hba962467),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe232b),
	.w1(32'h3a923769),
	.w2(32'hbb82e87f),
	.w3(32'h3b8362aa),
	.w4(32'hb9ab0f58),
	.w5(32'h3a4c6c95),
	.w6(32'h3b6981eb),
	.w7(32'hb96779a3),
	.w8(32'h39cb9714),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8e334),
	.w1(32'h3be4f489),
	.w2(32'hbb341198),
	.w3(32'h3b74494e),
	.w4(32'h3b7514f8),
	.w5(32'h3968747b),
	.w6(32'h3afa00c5),
	.w7(32'h3aed10f4),
	.w8(32'h3adf471b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f104),
	.w1(32'h38444547),
	.w2(32'h3ad3b7f2),
	.w3(32'h3a1571a5),
	.w4(32'h393fd257),
	.w5(32'h3a32d261),
	.w6(32'h3b0e1c07),
	.w7(32'h3b0b118c),
	.w8(32'h3aff6f8f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a165e6a),
	.w1(32'h387da354),
	.w2(32'hbb067c5d),
	.w3(32'h3b0c6a16),
	.w4(32'hb969b534),
	.w5(32'hbac8d757),
	.w6(32'h3b948042),
	.w7(32'hb980a886),
	.w8(32'h39bab574),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cd817),
	.w1(32'h3b1c31b6),
	.w2(32'h3bd30ad7),
	.w3(32'h3b80bae9),
	.w4(32'hba46615c),
	.w5(32'h3b329522),
	.w6(32'h3b5a7721),
	.w7(32'h3b5b3181),
	.w8(32'h3a72d7f6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995a112),
	.w1(32'hba82eaa0),
	.w2(32'h3a15a31b),
	.w3(32'h39a306df),
	.w4(32'hba94f33e),
	.w5(32'h3ae5bc7a),
	.w6(32'hba71d329),
	.w7(32'hba9f570b),
	.w8(32'h3b310792),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd3cdf),
	.w1(32'hba85ff29),
	.w2(32'hb9f00877),
	.w3(32'h3aee88dd),
	.w4(32'hbacb90c0),
	.w5(32'h3b378399),
	.w6(32'hbaa9e71b),
	.w7(32'hbb6156d3),
	.w8(32'h3bbc574e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831ac8),
	.w1(32'h3b9aab17),
	.w2(32'h3b8284d9),
	.w3(32'hb9b3abb6),
	.w4(32'hbb2bd219),
	.w5(32'h3864a3cc),
	.w6(32'hbaf02208),
	.w7(32'hbab008a5),
	.w8(32'hbb39fde3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb3fb),
	.w1(32'hb9dd1b11),
	.w2(32'hbb09bd9c),
	.w3(32'h39a7ad46),
	.w4(32'h3a98a42e),
	.w5(32'hbb8861e8),
	.w6(32'h3a36573f),
	.w7(32'h39cd2a56),
	.w8(32'hbb3baf7a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb6811),
	.w1(32'hb99a2053),
	.w2(32'hbb10f02f),
	.w3(32'h38947c9e),
	.w4(32'hbb0d29a5),
	.w5(32'hba864a7a),
	.w6(32'hbac5abbc),
	.w7(32'hb9646f0b),
	.w8(32'hb9a67019),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1e166),
	.w1(32'h3a416ea1),
	.w2(32'h3a725dc7),
	.w3(32'h3ba22189),
	.w4(32'h3a82410d),
	.w5(32'h3b2e648c),
	.w6(32'h3b3ca69b),
	.w7(32'h3ab51955),
	.w8(32'hbaf6124c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71147e),
	.w1(32'h3ada7981),
	.w2(32'h3b0c8994),
	.w3(32'hbb41a3d6),
	.w4(32'h3a8a6805),
	.w5(32'hba1464ce),
	.w6(32'hb8a289bb),
	.w7(32'h3b124b5c),
	.w8(32'h393d523d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5f16a),
	.w1(32'h3a002739),
	.w2(32'hbad913cf),
	.w3(32'h3a3103cd),
	.w4(32'hbabb73ee),
	.w5(32'hba0f3c69),
	.w6(32'h3b0b5068),
	.w7(32'h3a59edc5),
	.w8(32'hbb97699c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1fbfc),
	.w1(32'h3bace33d),
	.w2(32'h39dddbc6),
	.w3(32'h3ba1fd09),
	.w4(32'h3b20043c),
	.w5(32'hba921441),
	.w6(32'h3bf12813),
	.w7(32'h3bd987e0),
	.w8(32'h3bbabd4b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4743c4),
	.w1(32'hbac41573),
	.w2(32'hba6d493f),
	.w3(32'h39be18a2),
	.w4(32'h38c3d58c),
	.w5(32'hbb269ec2),
	.w6(32'hbb189f92),
	.w7(32'hb9212de4),
	.w8(32'hbb6b9571),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc004),
	.w1(32'h3afe7a83),
	.w2(32'hbbd52d26),
	.w3(32'hbb218a13),
	.w4(32'hbbcad832),
	.w5(32'hbb85e17f),
	.w6(32'h3c2aedee),
	.w7(32'hbc244110),
	.w8(32'hbbeba0a4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad98df9),
	.w1(32'hba8b8c73),
	.w2(32'hb9db5e8d),
	.w3(32'hba00ed6a),
	.w4(32'h39d40e95),
	.w5(32'h3b1e98f1),
	.w6(32'hbb0b8420),
	.w7(32'h398e0675),
	.w8(32'h3ada7d73),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1edc02),
	.w1(32'h3aa1c64d),
	.w2(32'h3ad07349),
	.w3(32'h39f326ad),
	.w4(32'h3adde7e6),
	.w5(32'hbbb3e910),
	.w6(32'h3836822c),
	.w7(32'h397170cb),
	.w8(32'hbb72fd6b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2c11),
	.w1(32'hba89dc0f),
	.w2(32'h3b2001a0),
	.w3(32'hbc6ed65c),
	.w4(32'h3b4c1505),
	.w5(32'hbad7b2ec),
	.w6(32'h3a7c56ed),
	.w7(32'h3abec64b),
	.w8(32'h3b5ff5ab),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999e77d),
	.w1(32'h3b6f4c9d),
	.w2(32'hbbabfb6d),
	.w3(32'h3b99b6db),
	.w4(32'h3a91563e),
	.w5(32'hbb6c9d69),
	.w6(32'h3c23111d),
	.w7(32'h3b90adc0),
	.w8(32'hba454030),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca67ed),
	.w1(32'hb9e073a0),
	.w2(32'hbb201bb4),
	.w3(32'hbbd1355c),
	.w4(32'h3b9e9412),
	.w5(32'hbb12e95f),
	.w6(32'h3ab11628),
	.w7(32'h3b70b84a),
	.w8(32'hbaf2733c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae89660),
	.w1(32'hbb588b8a),
	.w2(32'hb78bc018),
	.w3(32'hbb5283b2),
	.w4(32'hba595aa3),
	.w5(32'h394a9f58),
	.w6(32'hbb867311),
	.w7(32'hb9968355),
	.w8(32'h3a7bb788),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa58fb),
	.w1(32'hba367a2b),
	.w2(32'h3b8c8352),
	.w3(32'hbb34bb28),
	.w4(32'hbb717a65),
	.w5(32'h3b27bb92),
	.w6(32'hbb13cd3a),
	.w7(32'hbb3c32e1),
	.w8(32'hb9303b68),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e3674),
	.w1(32'hb95f440d),
	.w2(32'hbb2c263a),
	.w3(32'hba62dae9),
	.w4(32'hbb0cfbd6),
	.w5(32'hba9e678c),
	.w6(32'h3a16b2bc),
	.w7(32'hbb2b58f4),
	.w8(32'hb9f92fc9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932ff5),
	.w1(32'hbb9fe1d9),
	.w2(32'hba5598f5),
	.w3(32'hbb4b8cf8),
	.w4(32'hbb939a55),
	.w5(32'hb9189ae0),
	.w6(32'h3a954276),
	.w7(32'hbb9842b5),
	.w8(32'h3a3ba8b7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74a4bcc),
	.w1(32'hbb12806b),
	.w2(32'hbb752211),
	.w3(32'hba90b1d4),
	.w4(32'hb9c8d99a),
	.w5(32'h3bf0a0f8),
	.w6(32'hbbafcbfd),
	.w7(32'hba1b07bc),
	.w8(32'h3bb411a2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939657d),
	.w1(32'h38ff6f43),
	.w2(32'h3b80d21d),
	.w3(32'h3aef25b2),
	.w4(32'h3a7483c3),
	.w5(32'hba98bb88),
	.w6(32'hbac984a2),
	.w7(32'h3b344189),
	.w8(32'hba369a2c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc554),
	.w1(32'hbb19ae36),
	.w2(32'h393002ae),
	.w3(32'hbba08971),
	.w4(32'hbaf7a9c0),
	.w5(32'h3b2489d8),
	.w6(32'hbb261be2),
	.w7(32'hbb16e3d0),
	.w8(32'h3a893935),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbad00),
	.w1(32'h3b641170),
	.w2(32'h39f135cf),
	.w3(32'h3a86f273),
	.w4(32'h3b2671cd),
	.w5(32'h3aae5064),
	.w6(32'h3a89df83),
	.w7(32'h3a9fd053),
	.w8(32'h3baf419d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dafde),
	.w1(32'h3acf78c7),
	.w2(32'hb830a65f),
	.w3(32'h3b0b2702),
	.w4(32'h3b57775c),
	.w5(32'hbb7fa757),
	.w6(32'h3a8098b3),
	.w7(32'h3a8c60d0),
	.w8(32'hbb4e5195),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d6983),
	.w1(32'h3acb5bfa),
	.w2(32'h3a04f1ec),
	.w3(32'hbac66f70),
	.w4(32'hb993d6ff),
	.w5(32'hba0164a5),
	.w6(32'hbafa57e4),
	.w7(32'hba65352b),
	.w8(32'hb8e69dd0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab541db),
	.w1(32'h3b3f8749),
	.w2(32'hbb0b8288),
	.w3(32'h3b121eba),
	.w4(32'h3ba6bcbe),
	.w5(32'hbb37a7e8),
	.w6(32'h3bcee509),
	.w7(32'h3c0e6ec4),
	.w8(32'h3ba59887),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14f52e),
	.w1(32'h3b1ec1a0),
	.w2(32'hba5ca665),
	.w3(32'h3a74f3cd),
	.w4(32'h3abb6e77),
	.w5(32'hbb62e33e),
	.w6(32'h3b34e09d),
	.w7(32'h3b082612),
	.w8(32'h3a33ed94),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b94c1),
	.w1(32'hba4f6230),
	.w2(32'hba15868b),
	.w3(32'hba4d4f95),
	.w4(32'hbab03a1a),
	.w5(32'h3bebc8f8),
	.w6(32'hb9fc55e9),
	.w7(32'hbb25adbc),
	.w8(32'h3bbbf062),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34fec6),
	.w1(32'h3b382062),
	.w2(32'hb7d2f9a8),
	.w3(32'h3bcc8317),
	.w4(32'h3a9594e7),
	.w5(32'hbad7b09c),
	.w6(32'h3c037be2),
	.w7(32'h3b2ff684),
	.w8(32'hb9ca2cff),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c441),
	.w1(32'hbab27362),
	.w2(32'h3a86a9f3),
	.w3(32'hbab868a6),
	.w4(32'hbb2de194),
	.w5(32'h3a390919),
	.w6(32'hbb6afc33),
	.w7(32'h3a480157),
	.w8(32'h3a87b183),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398428d1),
	.w1(32'h3a6e91e7),
	.w2(32'h3a30c06a),
	.w3(32'h3a85254d),
	.w4(32'h3a7a9a85),
	.w5(32'hba4928b1),
	.w6(32'h3a9a7046),
	.w7(32'h3ab2ace7),
	.w8(32'hb98abdec),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19f0cf),
	.w1(32'h3983a02e),
	.w2(32'hba2a4e48),
	.w3(32'h39e734ec),
	.w4(32'h3a5d3728),
	.w5(32'h3a011b0a),
	.w6(32'h3998febe),
	.w7(32'hb942c7c8),
	.w8(32'hba05a857),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ab7cd),
	.w1(32'hb85fbe79),
	.w2(32'h3ad93e4a),
	.w3(32'hb8ae33b4),
	.w4(32'h39e967a5),
	.w5(32'hbb218746),
	.w6(32'hba07bd51),
	.w7(32'h39c67f87),
	.w8(32'hbad60028),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7dc46),
	.w1(32'hb9bf028a),
	.w2(32'h3ac06814),
	.w3(32'hbabe2d50),
	.w4(32'hbb014468),
	.w5(32'hb9dd234b),
	.w6(32'hb9463a99),
	.w7(32'hba5a1a49),
	.w8(32'hba819e04),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc4c9b),
	.w1(32'hba73959b),
	.w2(32'hbb3cd886),
	.w3(32'hb9b9f2fb),
	.w4(32'hbb49e8d4),
	.w5(32'h39ace113),
	.w6(32'h39a30ccc),
	.w7(32'hb9804bd3),
	.w8(32'hbbd2a064),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57d90e),
	.w1(32'h3ab83259),
	.w2(32'hbb159cd3),
	.w3(32'h3b452252),
	.w4(32'hb9676253),
	.w5(32'hbb384ebb),
	.w6(32'h3b8101d9),
	.w7(32'hba2e66a8),
	.w8(32'hba46d97f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a814a09),
	.w1(32'hbb52bcec),
	.w2(32'hbbe6f4b4),
	.w3(32'h3b19343b),
	.w4(32'hbb0b96b3),
	.w5(32'hbb37857a),
	.w6(32'h3afd49ab),
	.w7(32'hba3fd5d9),
	.w8(32'hbb6e909a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ee386),
	.w1(32'hba715cc0),
	.w2(32'hbb093527),
	.w3(32'h3710581f),
	.w4(32'h3a033cec),
	.w5(32'hbaf7df0e),
	.w6(32'h3ab3c06f),
	.w7(32'hbab078f7),
	.w8(32'hbac70dfd),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6efbbc),
	.w1(32'h3b1293c9),
	.w2(32'h3b0a9a6e),
	.w3(32'hba8f050b),
	.w4(32'h39fe5337),
	.w5(32'h3ab0022b),
	.w6(32'hbb032e39),
	.w7(32'h3a7327fc),
	.w8(32'h3b19c16d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70c7a2),
	.w1(32'h3a2f9818),
	.w2(32'h39f1e7d5),
	.w3(32'h3a7573de),
	.w4(32'hba008430),
	.w5(32'hbae2db5b),
	.w6(32'h3ae72b1e),
	.w7(32'h397aa3de),
	.w8(32'hb9997045),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29dae2),
	.w1(32'h397a6933),
	.w2(32'h3a9c0b73),
	.w3(32'hb71177a0),
	.w4(32'h3a0a5c3a),
	.w5(32'hbad8f6d4),
	.w6(32'h3acf0940),
	.w7(32'h3a9a51ca),
	.w8(32'hba3a66dd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42bea6),
	.w1(32'h39d643a7),
	.w2(32'hbb469b7b),
	.w3(32'h3b3fc14a),
	.w4(32'h3abd1879),
	.w5(32'hbb3d2c38),
	.w6(32'h3b2d9e74),
	.w7(32'h3a2edb11),
	.w8(32'h393a456a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e371fc),
	.w1(32'hba98eae1),
	.w2(32'hbb23d8a8),
	.w3(32'hbb63a21e),
	.w4(32'hbabfdcb8),
	.w5(32'hba03494a),
	.w6(32'hbba32f2c),
	.w7(32'hbb92280c),
	.w8(32'hb9b4214c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f78be),
	.w1(32'hbb0e5639),
	.w2(32'h3990f3de),
	.w3(32'hbaf176e1),
	.w4(32'hb88618f4),
	.w5(32'h3a18848f),
	.w6(32'hbb478664),
	.w7(32'hbac1611c),
	.w8(32'hbaf78ea2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c60af),
	.w1(32'h3b6047b0),
	.w2(32'h3b461042),
	.w3(32'h3b47da3b),
	.w4(32'h3a0aa9a4),
	.w5(32'h39fbc078),
	.w6(32'hb94334c2),
	.w7(32'h3a527c41),
	.w8(32'h3a9f6049),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8f235),
	.w1(32'h39b53621),
	.w2(32'hbb005c9d),
	.w3(32'h3a85e075),
	.w4(32'h38cf8cbf),
	.w5(32'h3b6cc85c),
	.w6(32'hba1c94fa),
	.w7(32'hba5084ac),
	.w8(32'hb9a3aa70),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3fb07),
	.w1(32'h3a806e08),
	.w2(32'h3afa7002),
	.w3(32'h3b3a3bda),
	.w4(32'hbaf1c101),
	.w5(32'hbb099df5),
	.w6(32'h3bb1211f),
	.w7(32'h3a276016),
	.w8(32'h3979fa25),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e94f2f),
	.w1(32'h3a8cef6f),
	.w2(32'hba96212a),
	.w3(32'h3a15ad36),
	.w4(32'h3aa85916),
	.w5(32'h3a83caf4),
	.w6(32'hb9f7bfa6),
	.w7(32'h3a02a1ff),
	.w8(32'hb9df2d3e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3aa1),
	.w1(32'hba3c72ae),
	.w2(32'hb93a419f),
	.w3(32'h3c2afc3d),
	.w4(32'h3b7c34ce),
	.w5(32'h3aeae0b4),
	.w6(32'h3c20dc17),
	.w7(32'h3b96591a),
	.w8(32'hbb3cf103),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5da2b),
	.w1(32'h3a8fba7c),
	.w2(32'h3ae9d152),
	.w3(32'h39e6dcf0),
	.w4(32'h3ae83b80),
	.w5(32'hbaa22a7e),
	.w6(32'h3a9fe14b),
	.w7(32'h3a7d7867),
	.w8(32'hba97757f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a9252),
	.w1(32'h3b39124f),
	.w2(32'h3b21fc0a),
	.w3(32'h3b490b6d),
	.w4(32'h3b0009cc),
	.w5(32'h3ad2712d),
	.w6(32'h3b6631a6),
	.w7(32'h3b0d00bf),
	.w8(32'h3bc7a0be),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule