module layer_8_featuremap_11(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccc8c3),
	.w1(32'hbc862675),
	.w2(32'hba4c144b),
	.w3(32'h3d0feae4),
	.w4(32'hbc2c8d8e),
	.w5(32'h3b8c0ac2),
	.w6(32'h3cce81b8),
	.w7(32'h3c193670),
	.w8(32'h3b2bb406),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6193fd),
	.w1(32'hbac9283e),
	.w2(32'h3b504f5d),
	.w3(32'h3afe8c58),
	.w4(32'h3a14b41f),
	.w5(32'h3bc290ac),
	.w6(32'h3b9af4e3),
	.w7(32'h3bacba41),
	.w8(32'h3ba8510f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66e382),
	.w1(32'h3ba12587),
	.w2(32'h3c1ce996),
	.w3(32'h3c15ee78),
	.w4(32'h3ba5289a),
	.w5(32'h3bc65503),
	.w6(32'h3c5e12bb),
	.w7(32'h3bd1cc0a),
	.w8(32'h3b032998),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913cda),
	.w1(32'h3bcaa609),
	.w2(32'h3c12bff6),
	.w3(32'hbb022f7c),
	.w4(32'h3c35680d),
	.w5(32'h3b31f36e),
	.w6(32'h3c6405bd),
	.w7(32'h3c88c849),
	.w8(32'h3a9c5bda),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd39e),
	.w1(32'h3b575740),
	.w2(32'h3b1ec9f4),
	.w3(32'hbb30a0b0),
	.w4(32'h3b4d6823),
	.w5(32'h3bc7f9c0),
	.w6(32'h3bb0bf2a),
	.w7(32'h3ba9d034),
	.w8(32'hba572fbd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130116),
	.w1(32'h3c84d8e9),
	.w2(32'h3c466a55),
	.w3(32'h3c08b7ca),
	.w4(32'h3c0f653e),
	.w5(32'h3c6c7eed),
	.w6(32'h3b2ce662),
	.w7(32'hbce476f5),
	.w8(32'hbc63116e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27bf02),
	.w1(32'hbbb69a05),
	.w2(32'hbc099407),
	.w3(32'h3c014b19),
	.w4(32'hbba2d5b1),
	.w5(32'hbb314a53),
	.w6(32'h3bd1786b),
	.w7(32'hbbcd10c9),
	.w8(32'hba0febfd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4580f8),
	.w1(32'h3b4ecb7c),
	.w2(32'h3baba0c6),
	.w3(32'hbc772ba0),
	.w4(32'h3a8dcca2),
	.w5(32'h3c936b01),
	.w6(32'h39ff9c65),
	.w7(32'hbb02553b),
	.w8(32'hbb6a801f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a2e61),
	.w1(32'h3c12e329),
	.w2(32'h3c18a4d4),
	.w3(32'h3b4360ba),
	.w4(32'h3c0e9397),
	.w5(32'h3bd5fb25),
	.w6(32'h3c8cfe1d),
	.w7(32'h3c099353),
	.w8(32'h3be2ed1b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef0368),
	.w1(32'h39d87945),
	.w2(32'hbc28c96e),
	.w3(32'h3c15b018),
	.w4(32'h3c3af03a),
	.w5(32'hbc01fee7),
	.w6(32'h3c4758a9),
	.w7(32'h3c4d1d89),
	.w8(32'hb9d8aa1a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfa9d6b),
	.w1(32'hba1f590b),
	.w2(32'h3bc98e8a),
	.w3(32'hbd1d981e),
	.w4(32'hbc4c15fb),
	.w5(32'hbb8cc5dd),
	.w6(32'hbcf84ec3),
	.w7(32'h3bbc0b90),
	.w8(32'h3b7b6f56),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa75e),
	.w1(32'hbc58550f),
	.w2(32'hbb85858d),
	.w3(32'h3ae1af19),
	.w4(32'hbb123d93),
	.w5(32'hbc11b4ab),
	.w6(32'h3c008600),
	.w7(32'hbc089ca0),
	.w8(32'hbbfaa5d4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8f93d),
	.w1(32'hbbca131b),
	.w2(32'hbc6a9947),
	.w3(32'hb957e6ed),
	.w4(32'h3cfdb592),
	.w5(32'h3c04dc3b),
	.w6(32'hba8f6747),
	.w7(32'h3c51d42f),
	.w8(32'h3ce4d359),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e13a9),
	.w1(32'h3a71ea5a),
	.w2(32'h3c5f9f22),
	.w3(32'hbd311ebb),
	.w4(32'hbc6331d7),
	.w5(32'hbcccaeee),
	.w6(32'hbbb13940),
	.w7(32'hb98ada61),
	.w8(32'hbcd4b742),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1970f3),
	.w1(32'h3b8b164d),
	.w2(32'h3b2a6b56),
	.w3(32'h3c68b251),
	.w4(32'h3c1a9721),
	.w5(32'h3c6f3694),
	.w6(32'hbbbadc96),
	.w7(32'h3bb4167c),
	.w8(32'h3c51a3b6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0427c1),
	.w1(32'h3b9651d1),
	.w2(32'h3c432965),
	.w3(32'h3b15b113),
	.w4(32'hba81006c),
	.w5(32'h3b933f82),
	.w6(32'h3c147267),
	.w7(32'h3bd8c456),
	.w8(32'h3be85076),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba76e9d),
	.w1(32'hbc40023d),
	.w2(32'h3ab39601),
	.w3(32'h3abc3319),
	.w4(32'hbc65e770),
	.w5(32'hbc950edc),
	.w6(32'h3b0f6325),
	.w7(32'h3a71449e),
	.w8(32'hbcaf0cfa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c147541),
	.w1(32'h3c10d57a),
	.w2(32'h3c88dfa8),
	.w3(32'h3d0dcbf2),
	.w4(32'h3c389446),
	.w5(32'h3c0036ec),
	.w6(32'h3d238522),
	.w7(32'h3c897c86),
	.w8(32'h3c0bf8f7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43705c),
	.w1(32'hbc810082),
	.w2(32'h3c27a917),
	.w3(32'hbd3d51a7),
	.w4(32'hbd1faead),
	.w5(32'h3d0dc5df),
	.w6(32'hbb752f63),
	.w7(32'h3d0c0424),
	.w8(32'h3d23ab89),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4b2d8),
	.w1(32'hbc133e6e),
	.w2(32'hbc5f388b),
	.w3(32'h3c9ae7ed),
	.w4(32'h3bba006a),
	.w5(32'h3beba87d),
	.w6(32'h3c2f47c6),
	.w7(32'hbbc20ab1),
	.w8(32'h3baab408),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf9bb8),
	.w1(32'h395be711),
	.w2(32'h3b863a82),
	.w3(32'hbb23bed5),
	.w4(32'hbc8d07ce),
	.w5(32'hbca45b1c),
	.w6(32'h39fad1db),
	.w7(32'hbc384fec),
	.w8(32'hbc6769b6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d004203),
	.w1(32'h3c7351fb),
	.w2(32'h3c063a14),
	.w3(32'h3cb59a83),
	.w4(32'hbb426b20),
	.w5(32'hbc3c9208),
	.w6(32'h3baec035),
	.w7(32'h39f0adfc),
	.w8(32'hbd1ece94),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf8d2e),
	.w1(32'h3c008371),
	.w2(32'h3d4cf475),
	.w3(32'hba9ead1b),
	.w4(32'h3ab14c1f),
	.w5(32'h3d8a94d9),
	.w6(32'hbc15b2ba),
	.w7(32'h3c195f1b),
	.w8(32'h3da2857d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933e31),
	.w1(32'h3a1b9f1d),
	.w2(32'h38bd4340),
	.w3(32'h3ca5cbd6),
	.w4(32'hb9beb7be),
	.w5(32'h3bcb6246),
	.w6(32'h3cff7ed1),
	.w7(32'hbc3a3a37),
	.w8(32'hbbb55f7a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364ca7),
	.w1(32'h3b5f4405),
	.w2(32'hbb8b7880),
	.w3(32'hb9af5898),
	.w4(32'h3b7fdd4a),
	.w5(32'hbb895f34),
	.w6(32'hb9d0b475),
	.w7(32'h39a74b2d),
	.w8(32'hbb5f1db9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3381a6),
	.w1(32'hba3ce7f4),
	.w2(32'h3bf27009),
	.w3(32'hbc998995),
	.w4(32'hbc5e6f1d),
	.w5(32'h3b9134ba),
	.w6(32'hbb055739),
	.w7(32'hbc9acf7b),
	.w8(32'hba4b81f1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb090e0),
	.w1(32'h3b8b18e6),
	.w2(32'h3b2b453b),
	.w3(32'h3bcb5461),
	.w4(32'h3b3fbe91),
	.w5(32'hbb297385),
	.w6(32'h3aed08ab),
	.w7(32'h3bfc4e32),
	.w8(32'h3a87b95e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c7136),
	.w1(32'hbcb4f0d2),
	.w2(32'hb9cf343c),
	.w3(32'hbd89def7),
	.w4(32'hbdbfce7a),
	.w5(32'hbd77950f),
	.w6(32'hbc104456),
	.w7(32'hbd8324f0),
	.w8(32'h3d49a633),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b2035),
	.w1(32'h3ad940e2),
	.w2(32'h3c8c11ed),
	.w3(32'hbc60ac81),
	.w4(32'h3b4fd780),
	.w5(32'h3c2ede1b),
	.w6(32'h3c8d4c97),
	.w7(32'h3c49a27b),
	.w8(32'h3ca1f1ec),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98d6cc),
	.w1(32'hbabd5cee),
	.w2(32'hb8578201),
	.w3(32'h3c70a79a),
	.w4(32'hb99e976d),
	.w5(32'hba6204cb),
	.w6(32'h3ca5197c),
	.w7(32'hba94a02f),
	.w8(32'h3affaa57),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8383bf),
	.w1(32'hbb5e496a),
	.w2(32'hbc6944c3),
	.w3(32'hbad34f6e),
	.w4(32'hbc1e4ab3),
	.w5(32'hbc6f0b8b),
	.w6(32'h3b17268d),
	.w7(32'hbc8bd900),
	.w8(32'hbc4ea43f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc091d94),
	.w1(32'hbaf2686f),
	.w2(32'h3b7768bc),
	.w3(32'hbc5c977b),
	.w4(32'hbbdd3442),
	.w5(32'h3b9defe2),
	.w6(32'hbc3ac8e5),
	.w7(32'hbc090168),
	.w8(32'h3b5e8d40),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2027c4),
	.w1(32'h3b1c9db1),
	.w2(32'h3b835e8b),
	.w3(32'h39b85dc7),
	.w4(32'hbaa7dfd0),
	.w5(32'hbb0f5fc1),
	.w6(32'h3aa50044),
	.w7(32'h3ae99815),
	.w8(32'hba8e780d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1747b7),
	.w1(32'h3bc3b596),
	.w2(32'h3ca60c54),
	.w3(32'h3b42f3ca),
	.w4(32'hbc57fa99),
	.w5(32'h3cf0bed6),
	.w6(32'h3ab7be37),
	.w7(32'hbcbd6e56),
	.w8(32'hba53e14b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb225c9),
	.w1(32'hbb8230a8),
	.w2(32'hba653504),
	.w3(32'h3cc29dbf),
	.w4(32'h3a83867b),
	.w5(32'h3a8367f8),
	.w6(32'h3b993363),
	.w7(32'hbc186647),
	.w8(32'hbbdd6432),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099837),
	.w1(32'hbc9dc4c1),
	.w2(32'hbb5723ab),
	.w3(32'hbc51b495),
	.w4(32'hbcc41b3c),
	.w5(32'h3b561760),
	.w6(32'hbbc1d178),
	.w7(32'hbc45334b),
	.w8(32'h3c39a078),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ba2d),
	.w1(32'hbc307ed5),
	.w2(32'hbc46605b),
	.w3(32'h3b923fe7),
	.w4(32'h3c7e3ad9),
	.w5(32'h3c30859e),
	.w6(32'h3bc8df50),
	.w7(32'h3cc48e80),
	.w8(32'h3cecea2d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91d160),
	.w1(32'hbc8a13bf),
	.w2(32'hbca769b2),
	.w3(32'hbd45423d),
	.w4(32'hbbf00ff8),
	.w5(32'hbce93793),
	.w6(32'hbc93a901),
	.w7(32'hb896f42f),
	.w8(32'hbccaf5e7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc558),
	.w1(32'hbb93a610),
	.w2(32'hbbb6cceb),
	.w3(32'hbc906518),
	.w4(32'h3c060964),
	.w5(32'h3c8d62e7),
	.w6(32'hbc32b66d),
	.w7(32'hbc31fd60),
	.w8(32'h3c9c97f5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d4fa2),
	.w1(32'hbbaf4207),
	.w2(32'hbc364dc8),
	.w3(32'hbbba759c),
	.w4(32'hbbb7f0b5),
	.w5(32'h3c135359),
	.w6(32'h3c934521),
	.w7(32'hbc9a3de8),
	.w8(32'h3c2514d1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83b044),
	.w1(32'h3cb88cda),
	.w2(32'h3cabf140),
	.w3(32'h3c2679db),
	.w4(32'h3cfc1e1e),
	.w5(32'h3c57514a),
	.w6(32'h3cfdfe05),
	.w7(32'h3d0e1d42),
	.w8(32'h3c707a79),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900dfb),
	.w1(32'hbb024f26),
	.w2(32'h3c28483c),
	.w3(32'hbc048252),
	.w4(32'hbc5d7f7f),
	.w5(32'hbc2b2769),
	.w6(32'hbbceedd4),
	.w7(32'h3a06bef6),
	.w8(32'hbbfe76bd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1fdd9),
	.w1(32'hbb7ac30a),
	.w2(32'hbb795b90),
	.w3(32'h3c2cecf9),
	.w4(32'hbba9b7b4),
	.w5(32'hbbd60b19),
	.w6(32'h3b28fcdd),
	.w7(32'hbbe772d7),
	.w8(32'hbbf073b8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b73b),
	.w1(32'hbb7a3000),
	.w2(32'h3b604181),
	.w3(32'hbbe6c9da),
	.w4(32'hbca68eb7),
	.w5(32'h3ca875d3),
	.w6(32'hba74b2b7),
	.w7(32'hbc36f86a),
	.w8(32'h3966c819),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89697b),
	.w1(32'h3bb07fb9),
	.w2(32'hbaf7ee29),
	.w3(32'hbc5ba758),
	.w4(32'hbb6e52da),
	.w5(32'hbbee9d44),
	.w6(32'h3ad0bf3c),
	.w7(32'h3cd755a1),
	.w8(32'h3d5a5243),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c56ab),
	.w1(32'hbc18660e),
	.w2(32'h399fb421),
	.w3(32'hbd0b96f0),
	.w4(32'hbc75bfed),
	.w5(32'h3c1264e2),
	.w6(32'hbba9de72),
	.w7(32'h3bc01a5d),
	.w8(32'h3ce10245),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5b32),
	.w1(32'hbb8164a7),
	.w2(32'h3bbab23a),
	.w3(32'hbc3904c4),
	.w4(32'hbb4397a0),
	.w5(32'h3b26bf0e),
	.w6(32'h3bcd4fae),
	.w7(32'hbc01a204),
	.w8(32'hbc93b440),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94d081),
	.w1(32'hbc82b7bc),
	.w2(32'h3ae237b2),
	.w3(32'hbc15205f),
	.w4(32'hbd5eb240),
	.w5(32'hbb8941fd),
	.w6(32'hba093ab2),
	.w7(32'hbd1fa2d3),
	.w8(32'h39d5c577),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc918660),
	.w1(32'h3bf26b04),
	.w2(32'h3b695752),
	.w3(32'hbc8a9021),
	.w4(32'h3c1024fa),
	.w5(32'h3c2b8a24),
	.w6(32'hbb0ddbb6),
	.w7(32'h3b9b4c24),
	.w8(32'h3c2ec14c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aa690),
	.w1(32'h3bbd41e3),
	.w2(32'h3c0eaa98),
	.w3(32'hbc443559),
	.w4(32'h3b9e3190),
	.w5(32'hbba12dd4),
	.w6(32'h3c2cdb53),
	.w7(32'h3cd6953e),
	.w8(32'h3bc7768f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f9037),
	.w1(32'h3bd23a7c),
	.w2(32'h3c6f0788),
	.w3(32'hbb8e6e0a),
	.w4(32'h3bfc1403),
	.w5(32'h3ca52a7f),
	.w6(32'hbc53595e),
	.w7(32'h3ba7146f),
	.w8(32'h3cb78e4c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba89c4a),
	.w1(32'hbb4a3963),
	.w2(32'h3c4bf32f),
	.w3(32'hbcbef7e3),
	.w4(32'hbd137620),
	.w5(32'hbc6ecfe9),
	.w6(32'h3c7bb885),
	.w7(32'h3ad9e70d),
	.w8(32'h3c4dfd31),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab05e55),
	.w1(32'hbb595742),
	.w2(32'h3a9a199d),
	.w3(32'h3a887ddd),
	.w4(32'hbc832f2a),
	.w5(32'hbc70f930),
	.w6(32'h3a29ad1b),
	.w7(32'hbc84380f),
	.w8(32'h3a403f0f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf2fd4a),
	.w1(32'hbc77c0e6),
	.w2(32'hbbffeec9),
	.w3(32'hbc99331c),
	.w4(32'h3c2a5087),
	.w5(32'h3ca4123d),
	.w6(32'h3ba35609),
	.w7(32'hbc479fa9),
	.w8(32'hbc429a39),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa64a5),
	.w1(32'h3a7645d9),
	.w2(32'hbbed4780),
	.w3(32'h3c9d2647),
	.w4(32'h3cf2ea69),
	.w5(32'h3cd35f6d),
	.w6(32'h3c4c3d61),
	.w7(32'h3c4e6ecc),
	.w8(32'h3cf401cd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd357219),
	.w1(32'hbc801f67),
	.w2(32'h3b92e632),
	.w3(32'hbd148ba3),
	.w4(32'hbc832337),
	.w5(32'h3c2a0bc8),
	.w6(32'h3b81b96b),
	.w7(32'h3c9d83d4),
	.w8(32'h3c96e968),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c116851),
	.w1(32'h3b89fc1a),
	.w2(32'h3c615eb6),
	.w3(32'h3c0f7a6b),
	.w4(32'h3c3fa8a1),
	.w5(32'h3d09498e),
	.w6(32'h3c0a3281),
	.w7(32'h3c2fb224),
	.w8(32'h3cf2d4d5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59edc),
	.w1(32'hbab5d712),
	.w2(32'h3c43b1f3),
	.w3(32'h3c7f4b12),
	.w4(32'hbc12cbb6),
	.w5(32'h3bbe0dd4),
	.w6(32'h3cfb5a99),
	.w7(32'hbb224517),
	.w8(32'h3c77f866),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4947),
	.w1(32'hba64c012),
	.w2(32'h3c3d44e3),
	.w3(32'hbb7987c6),
	.w4(32'hbc217485),
	.w5(32'h3c2aa106),
	.w6(32'hba4aa3df),
	.w7(32'hbb06002a),
	.w8(32'h3c8310e0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b749522),
	.w1(32'h3c690a19),
	.w2(32'hbbdc7670),
	.w3(32'h3b9b7f89),
	.w4(32'hbbaca0b5),
	.w5(32'h3c75463a),
	.w6(32'h3bd3d0cd),
	.w7(32'hbb058586),
	.w8(32'h3c980e23),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5f6b),
	.w1(32'hbb66a8f2),
	.w2(32'hbb819efc),
	.w3(32'hbc98944c),
	.w4(32'hbba3a9c8),
	.w5(32'hbc81680d),
	.w6(32'h3b3b7aff),
	.w7(32'h3c8d5cfe),
	.w8(32'hbb9832cb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba744aa),
	.w1(32'hbc86ad23),
	.w2(32'hbb7de3b9),
	.w3(32'hbc163fdd),
	.w4(32'hbc1f009b),
	.w5(32'h3bd29024),
	.w6(32'hbbd942b2),
	.w7(32'hbcdaa5af),
	.w8(32'hbc964093),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce31a5d),
	.w1(32'hbb969130),
	.w2(32'h3b0e90d4),
	.w3(32'hbcad420e),
	.w4(32'h3bb1081a),
	.w5(32'h3c6d1dad),
	.w6(32'h3ac78623),
	.w7(32'h3cb3cfcf),
	.w8(32'h3c675347),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba109a59),
	.w1(32'h3c0b8288),
	.w2(32'h38052b17),
	.w3(32'h3a555f74),
	.w4(32'hba68f2eb),
	.w5(32'h3c40739f),
	.w6(32'h3aef65be),
	.w7(32'hbbd86220),
	.w8(32'h3bbfc98e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdab323),
	.w1(32'hbbeb1a5f),
	.w2(32'hbb02e7d0),
	.w3(32'h3b8aaf67),
	.w4(32'hbc206422),
	.w5(32'hbc438c24),
	.w6(32'h3c01b489),
	.w7(32'hbbec4e87),
	.w8(32'hbc231a26),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be620a5),
	.w1(32'h3c2d2979),
	.w2(32'hbb2c6d0f),
	.w3(32'hbb121451),
	.w4(32'h3bac5d84),
	.w5(32'hbbfe1d7d),
	.w6(32'h3a1b77e6),
	.w7(32'h3c7d48ea),
	.w8(32'hba08908c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0801),
	.w1(32'h3bb772b1),
	.w2(32'h3c0e1698),
	.w3(32'h3bf25750),
	.w4(32'h3b7a25bd),
	.w5(32'hbc04d701),
	.w6(32'h3bbbcf65),
	.w7(32'h3bc72479),
	.w8(32'hbc0da923),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280415),
	.w1(32'hbbefe587),
	.w2(32'hbb1b9aa7),
	.w3(32'hbc2cfdcd),
	.w4(32'hbc2b9929),
	.w5(32'hbc50bbbb),
	.w6(32'hbbeec047),
	.w7(32'hba622955),
	.w8(32'hbc42e3df),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc65b55),
	.w1(32'h3adb0db0),
	.w2(32'h3bbcf321),
	.w3(32'h3b3b86e1),
	.w4(32'hbb851a56),
	.w5(32'hbb78e7e2),
	.w6(32'h3b211817),
	.w7(32'hba053bf6),
	.w8(32'hbbd69b95),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10182b),
	.w1(32'h3b90503c),
	.w2(32'h3c489271),
	.w3(32'hbcbe00bf),
	.w4(32'hbd5bf95f),
	.w5(32'hbc8066e4),
	.w6(32'hbcba75fe),
	.w7(32'hbc87d3c3),
	.w8(32'h3c853843),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe2d14),
	.w1(32'h3ab3a4bb),
	.w2(32'h3ca3c13b),
	.w3(32'h3a2fb74b),
	.w4(32'h3c9c624f),
	.w5(32'h3d29bb41),
	.w6(32'hbad75fdc),
	.w7(32'h3c0bc8f6),
	.w8(32'h3cd4c6e1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fc525),
	.w1(32'hbb4444e0),
	.w2(32'h3bebe8eb),
	.w3(32'h3ccc35f9),
	.w4(32'hbc24913a),
	.w5(32'hbb11faa7),
	.w6(32'h3c74436e),
	.w7(32'hbc065412),
	.w8(32'hb73a9285),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d9f0c),
	.w1(32'hbb022e7c),
	.w2(32'hbaa495ca),
	.w3(32'h3bb118f7),
	.w4(32'h39016343),
	.w5(32'hba52887e),
	.w6(32'h3ad0a70d),
	.w7(32'hbaa7368d),
	.w8(32'hbb1141c9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3727d),
	.w1(32'hbb91a037),
	.w2(32'h3c3f1216),
	.w3(32'h3ba7cd20),
	.w4(32'h3c262dae),
	.w5(32'h3bc2af7e),
	.w6(32'h3c232de8),
	.w7(32'h3c3aac21),
	.w8(32'h3c0f7572),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dee2b9),
	.w1(32'hbbe42902),
	.w2(32'hbb2852b2),
	.w3(32'h390e06b2),
	.w4(32'hbb8050a9),
	.w5(32'hbaad2ebc),
	.w6(32'hbb8819fa),
	.w7(32'hbbb32a1f),
	.w8(32'hbb0ff339),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba618f2b),
	.w1(32'hbbc890a6),
	.w2(32'hbace8a0c),
	.w3(32'h37585557),
	.w4(32'hbbbbc950),
	.w5(32'h397619e6),
	.w6(32'hbb7d0db2),
	.w7(32'hbb30e9a5),
	.w8(32'h3b8e9cd5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72bd7c),
	.w1(32'hbbb84022),
	.w2(32'hbace37c7),
	.w3(32'h3b7d1345),
	.w4(32'hbc122ecb),
	.w5(32'hbc37e419),
	.w6(32'h3abb987f),
	.w7(32'hbbb393c8),
	.w8(32'hbc2931ca),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d4adc),
	.w1(32'h3c009f66),
	.w2(32'h3cc3bd59),
	.w3(32'hbc9fd7d0),
	.w4(32'h3c275923),
	.w5(32'h3d3072a5),
	.w6(32'hbc5f46fc),
	.w7(32'h3c85118f),
	.w8(32'h3d242f73),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8566c),
	.w1(32'hbcb4ff71),
	.w2(32'hbc03ec2a),
	.w3(32'h3c7069b4),
	.w4(32'hbcb51564),
	.w5(32'hbc03dc73),
	.w6(32'h3c5169c6),
	.w7(32'hbc6abf3f),
	.w8(32'hbc0dfee4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95a9c6),
	.w1(32'h3baa7f04),
	.w2(32'h3b8d04dd),
	.w3(32'hbcaaa22d),
	.w4(32'h3bc9384e),
	.w5(32'h3b9a98c3),
	.w6(32'hbccae1fb),
	.w7(32'hba82f838),
	.w8(32'hbb150ae7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d1e96),
	.w1(32'h37d2115b),
	.w2(32'hbab10aef),
	.w3(32'h3b85bc98),
	.w4(32'hbbe0fd6a),
	.w5(32'hbc319dba),
	.w6(32'hbae2d2c8),
	.w7(32'hbb093328),
	.w8(32'hbc2eb4e8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432041),
	.w1(32'h3b84a13c),
	.w2(32'h3c32b1d6),
	.w3(32'hbbfc2157),
	.w4(32'h3a1dd436),
	.w5(32'h3bfa5904),
	.w6(32'hbcc4e6d0),
	.w7(32'hbc60005a),
	.w8(32'h3b2ae9a9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a1f09),
	.w1(32'hbbf4e648),
	.w2(32'h3b119664),
	.w3(32'hbc91097d),
	.w4(32'hbcacca74),
	.w5(32'hbbdad05e),
	.w6(32'hbc325940),
	.w7(32'hbc4c794c),
	.w8(32'hbbc9b5a8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdab7f3),
	.w1(32'h3ca1c333),
	.w2(32'h3d1223b7),
	.w3(32'hbbf09c58),
	.w4(32'h3d302d65),
	.w5(32'h3d57dc37),
	.w6(32'h3c82fb83),
	.w7(32'h3d56f4d3),
	.w8(32'h3caedfb2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0894b2),
	.w1(32'hbc7e11bf),
	.w2(32'h3b0facf3),
	.w3(32'hbaef175c),
	.w4(32'hbd06cfcf),
	.w5(32'hbc507ccd),
	.w6(32'h3ca2510d),
	.w7(32'h3bb1e28a),
	.w8(32'h3c3bc62e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fbeeb),
	.w1(32'h3b717e2e),
	.w2(32'hb986c162),
	.w3(32'hbb98ab51),
	.w4(32'hbab07a3e),
	.w5(32'h39bdc88a),
	.w6(32'hbb3b4b1a),
	.w7(32'hbbb9826e),
	.w8(32'h3b732650),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6f522),
	.w1(32'hbc479431),
	.w2(32'hbc095467),
	.w3(32'hbb7c3843),
	.w4(32'h3aa5a54c),
	.w5(32'h3c0043e0),
	.w6(32'hbb1ba76c),
	.w7(32'hbaaed336),
	.w8(32'h3aa00610),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd29643),
	.w1(32'h3bfda1d2),
	.w2(32'h3cb0ade1),
	.w3(32'h3bd9ae7b),
	.w4(32'h3cb67e4f),
	.w5(32'h3d1c736d),
	.w6(32'hbb6dc267),
	.w7(32'h3c543b76),
	.w8(32'h3cda831d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bddff),
	.w1(32'h39fc052d),
	.w2(32'h3ae44b05),
	.w3(32'h3ccc452e),
	.w4(32'hbad67685),
	.w5(32'h3bb2a8de),
	.w6(32'h3c79c6f8),
	.w7(32'h3af7d2ac),
	.w8(32'hbb8ad59f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4166aa),
	.w1(32'hb825ac7d),
	.w2(32'h3a945eb7),
	.w3(32'hbbec8585),
	.w4(32'h3ac8563d),
	.w5(32'h3b98c0b8),
	.w6(32'hbc117665),
	.w7(32'h3a53bca9),
	.w8(32'h3bd27922),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc23e0),
	.w1(32'h3c6114a4),
	.w2(32'h3c5254bd),
	.w3(32'h3c46b21a),
	.w4(32'h3c0c0230),
	.w5(32'h3a1aed0e),
	.w6(32'h3c24f054),
	.w7(32'h3ba91dd9),
	.w8(32'h3b728817),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d40a1),
	.w1(32'h3c3efa4c),
	.w2(32'h3a5b1f54),
	.w3(32'h3ac57ba1),
	.w4(32'h3c0a178a),
	.w5(32'h3c01d14f),
	.w6(32'h3bae239c),
	.w7(32'hbba8c103),
	.w8(32'h3be06435),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf839c9),
	.w1(32'h3af474b8),
	.w2(32'h3ba531e6),
	.w3(32'h3c0f55cc),
	.w4(32'hbb151b64),
	.w5(32'hbb63051c),
	.w6(32'h3b6e334b),
	.w7(32'h3aecdf28),
	.w8(32'hb9ece174),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b704d48),
	.w1(32'h3b8cadd7),
	.w2(32'h3c8a1244),
	.w3(32'h3b5ef97b),
	.w4(32'h3c72a5e1),
	.w5(32'h3cdda1e2),
	.w6(32'h3bf7599d),
	.w7(32'h3c5f77f7),
	.w8(32'h3cb45b77),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b824cad),
	.w1(32'hbc1f7e9a),
	.w2(32'h3b8144a8),
	.w3(32'h3c7d6187),
	.w4(32'hbb26d08b),
	.w5(32'hbbcfe1a5),
	.w6(32'h3c3c8ef7),
	.w7(32'h3aeffcca),
	.w8(32'h3a99da55),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a94f5),
	.w1(32'h3b73ef8c),
	.w2(32'h3cc23cc3),
	.w3(32'hbcc35c5c),
	.w4(32'h3be395a5),
	.w5(32'h3ceaeec3),
	.w6(32'hbc0e6139),
	.w7(32'h3c0fb181),
	.w8(32'h3cbc906d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007a15),
	.w1(32'hbc52ff5d),
	.w2(32'h3c03a2f9),
	.w3(32'h3beb8373),
	.w4(32'h3c09c8f4),
	.w5(32'h3d0a7cda),
	.w6(32'h3a31bb2d),
	.w7(32'hb9bc8c71),
	.w8(32'h3c912a6a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f0e5c),
	.w1(32'hb7d28d93),
	.w2(32'h3bdb558a),
	.w3(32'h3c9ae93a),
	.w4(32'h3b024e84),
	.w5(32'h3c13b3bc),
	.w6(32'h3bb390d2),
	.w7(32'hba88e85d),
	.w8(32'h3b3629bb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af9dce),
	.w1(32'h3ac0e0fd),
	.w2(32'hba16ce3a),
	.w3(32'hbaa27af4),
	.w4(32'hba3e12e1),
	.w5(32'hbaf69c40),
	.w6(32'h3be69670),
	.w7(32'h3a50c7fb),
	.w8(32'hbacad81e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b121973),
	.w1(32'h3b4335c5),
	.w2(32'h3bea3892),
	.w3(32'hb90c407e),
	.w4(32'h3ba9dbaa),
	.w5(32'h3bda5953),
	.w6(32'h3a5b6728),
	.w7(32'h3c0b9e07),
	.w8(32'h3c1cd381),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1c319),
	.w1(32'h3b1d7503),
	.w2(32'h3c0083e7),
	.w3(32'h3b30b6e0),
	.w4(32'h3c2005f0),
	.w5(32'h3c0a918e),
	.w6(32'h3bc6e4fe),
	.w7(32'h3b556549),
	.w8(32'h3b3814ef),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977b43),
	.w1(32'h3bc55ca2),
	.w2(32'h3b5fbcb4),
	.w3(32'h3b3d7572),
	.w4(32'hbadad83c),
	.w5(32'hbb7a5921),
	.w6(32'hbb8114bc),
	.w7(32'h398f54a2),
	.w8(32'hbbf4eb19),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefc11d),
	.w1(32'hbbbdbb5c),
	.w2(32'hba2723bd),
	.w3(32'hbbfb5e60),
	.w4(32'h3a4e37ee),
	.w5(32'h3c229065),
	.w6(32'hbc0eda8f),
	.w7(32'h3b58953d),
	.w8(32'h3b99d920),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70dfec),
	.w1(32'hbb0466ff),
	.w2(32'h3c13434d),
	.w3(32'h3cbc9819),
	.w4(32'hba98a427),
	.w5(32'h3bd53423),
	.w6(32'h3b9e501d),
	.w7(32'hbc0fd425),
	.w8(32'hb99617b0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c000fd1),
	.w1(32'h3c028b81),
	.w2(32'h3c8c77da),
	.w3(32'h3c24da76),
	.w4(32'h3d000680),
	.w5(32'h3d4bc30a),
	.w6(32'h3c036bb1),
	.w7(32'h3c3772f4),
	.w8(32'h3cc4bd3a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3aa07),
	.w1(32'h3bb1c14a),
	.w2(32'h3c84f1f7),
	.w3(32'h3c11f40d),
	.w4(32'hbc1d5432),
	.w5(32'h3c61f4f0),
	.w6(32'h3a5ed5d0),
	.w7(32'h3af0ea84),
	.w8(32'h3cc289a5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48cbaa),
	.w1(32'hbb91195e),
	.w2(32'hbbc25c2f),
	.w3(32'h3c02a425),
	.w4(32'hbbb04d02),
	.w5(32'hbbfbe129),
	.w6(32'h3b6a6fa4),
	.w7(32'hbb807080),
	.w8(32'hbbbe4157),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b467aa5),
	.w1(32'hbb79ab15),
	.w2(32'h3ae639ea),
	.w3(32'h396bcf1d),
	.w4(32'h3b529845),
	.w5(32'hb9292307),
	.w6(32'hbb69a27e),
	.w7(32'hbb8cd361),
	.w8(32'h3bd03600),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc98fea),
	.w1(32'hbc0ddff9),
	.w2(32'hbbcb8a67),
	.w3(32'h3c123b40),
	.w4(32'hbc1751fa),
	.w5(32'h3b842e47),
	.w6(32'h3c26e1d6),
	.w7(32'h3b339638),
	.w8(32'h3c3c18f3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0048cf),
	.w1(32'hbb6d03b6),
	.w2(32'h3bde7f6f),
	.w3(32'h3bd6e556),
	.w4(32'h3add2d27),
	.w5(32'h3c1def2b),
	.w6(32'h3c2a72de),
	.w7(32'h3aa97950),
	.w8(32'h3c0184dc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf11aa8),
	.w1(32'hbc384665),
	.w2(32'hbc0f3a04),
	.w3(32'h3af29e02),
	.w4(32'hbc64549d),
	.w5(32'hbc2d304c),
	.w6(32'hbbbc87db),
	.w7(32'hbb73319c),
	.w8(32'hbb988ab3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7bfdc),
	.w1(32'hba6c3eba),
	.w2(32'h3818085f),
	.w3(32'h3bf69711),
	.w4(32'h3b2163b6),
	.w5(32'h3be64146),
	.w6(32'h3c335dcc),
	.w7(32'h3ac0f64f),
	.w8(32'h3bb40887),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70b5e9),
	.w1(32'h3c7c2e75),
	.w2(32'h3cd8d413),
	.w3(32'hba9b88e4),
	.w4(32'h3cd921e9),
	.w5(32'h3d19595b),
	.w6(32'hbac02455),
	.w7(32'h3cd30d55),
	.w8(32'h3d1392d8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6811d9),
	.w1(32'hbbba540a),
	.w2(32'hbb5fb04a),
	.w3(32'h3cd71df2),
	.w4(32'h399d4d20),
	.w5(32'h3b4136fa),
	.w6(32'h3cbfb61c),
	.w7(32'h3ab93448),
	.w8(32'h3bfcd29c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84478e),
	.w1(32'h3be17abc),
	.w2(32'h3c397963),
	.w3(32'h3a8ffd28),
	.w4(32'h3c45cd30),
	.w5(32'h3c9b93ee),
	.w6(32'h3c01096a),
	.w7(32'h3c5050c9),
	.w8(32'h3c908816),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66a596),
	.w1(32'hbbd26f6a),
	.w2(32'hbba368e5),
	.w3(32'h3c846710),
	.w4(32'hbb534148),
	.w5(32'hb9ed15cd),
	.w6(32'h3c63d329),
	.w7(32'hbb55c88b),
	.w8(32'hba348e98),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f022ba),
	.w1(32'hbbb96612),
	.w2(32'h3b50300e),
	.w3(32'h3b5e77b1),
	.w4(32'h3ae54963),
	.w5(32'h3bc6cffa),
	.w6(32'h3b26efce),
	.w7(32'h3b8ebe5d),
	.w8(32'h3c2862ab),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9100e),
	.w1(32'hbb1fd018),
	.w2(32'hba019f5f),
	.w3(32'hbbadcb09),
	.w4(32'hbb9d568e),
	.w5(32'h3ab010a4),
	.w6(32'h383b38b8),
	.w7(32'hbb2eb311),
	.w8(32'h3bd68bb8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb075c1b),
	.w1(32'hbb39019e),
	.w2(32'hbb6c9125),
	.w3(32'hbc18d65c),
	.w4(32'h3aa9e382),
	.w5(32'hbb72d9f0),
	.w6(32'hbc33f549),
	.w7(32'h3aa3d670),
	.w8(32'hbbe10390),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1a72b),
	.w1(32'hba9fe485),
	.w2(32'h3bd5b484),
	.w3(32'hbb8b7488),
	.w4(32'h3c03f79a),
	.w5(32'h3c6eb23a),
	.w6(32'hbc3b46f4),
	.w7(32'h3bd9a37e),
	.w8(32'h3c31c9e1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36d48c),
	.w1(32'h3c08c11c),
	.w2(32'h3c991554),
	.w3(32'h3c16eb29),
	.w4(32'h3cb2c604),
	.w5(32'h3d1296f7),
	.w6(32'hba69dae4),
	.w7(32'h3c93ef17),
	.w8(32'h3cddd2bd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f9875),
	.w1(32'h3920dfad),
	.w2(32'hba362311),
	.w3(32'h3cc19850),
	.w4(32'h3c1f165a),
	.w5(32'h3bfc1eb6),
	.w6(32'h3cc062a2),
	.w7(32'h3bdd9a1a),
	.w8(32'h3b1cc146),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e0cbc),
	.w1(32'hba8e422c),
	.w2(32'hbb1d0c01),
	.w3(32'h3be3da56),
	.w4(32'h39fa85d4),
	.w5(32'h3a9008f7),
	.w6(32'h3b962b20),
	.w7(32'h3b59b59d),
	.w8(32'h3b108206),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03959c),
	.w1(32'hbbc687b9),
	.w2(32'h3c14d3e3),
	.w3(32'h3b8a6b55),
	.w4(32'h3a9c6734),
	.w5(32'h3c1a6532),
	.w6(32'h3bbc9f12),
	.w7(32'hbbb00d3c),
	.w8(32'h3ae81953),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a330),
	.w1(32'h3ae349ee),
	.w2(32'h3b8ed8af),
	.w3(32'h3c0bf911),
	.w4(32'h3b65b64e),
	.w5(32'h3beb4c80),
	.w6(32'hb9831860),
	.w7(32'hbbbefb27),
	.w8(32'hbb4863bb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7adb00),
	.w1(32'hbb864c05),
	.w2(32'hb9c566d7),
	.w3(32'h3a38a21c),
	.w4(32'hbc264dea),
	.w5(32'hb9cd6f1e),
	.w6(32'hbc0ca02b),
	.w7(32'hbb74f701),
	.w8(32'h3b4cd0d4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca9eb5),
	.w1(32'h3c561454),
	.w2(32'h3cabf66e),
	.w3(32'hba55f373),
	.w4(32'h3ccbe4e8),
	.w5(32'h3cead9e0),
	.w6(32'hbacf8ee1),
	.w7(32'h3cdd7c16),
	.w8(32'h3cf24bf9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b741026),
	.w1(32'hbcc7e0c1),
	.w2(32'hbbd5d1da),
	.w3(32'h3bafa861),
	.w4(32'hbc95ec49),
	.w5(32'hba8bd151),
	.w6(32'h3c09e245),
	.w7(32'hbc71e6f8),
	.w8(32'h3bad66f3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule