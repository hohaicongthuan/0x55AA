module layer_8_featuremap_120(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c69ef),
	.w1(32'hb959e28d),
	.w2(32'h3c2ad67e),
	.w3(32'hb93fa206),
	.w4(32'h3b947db5),
	.w5(32'h3b4c8fcd),
	.w6(32'h3a53a8a9),
	.w7(32'h39b9889c),
	.w8(32'h3a7b637c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e22f8),
	.w1(32'h3b15b2a8),
	.w2(32'hbbb7ddf7),
	.w3(32'h3b851b0b),
	.w4(32'hba2f12ca),
	.w5(32'hbbfd22c3),
	.w6(32'h3adef657),
	.w7(32'hbaf328b8),
	.w8(32'hbc07aa8c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f11f),
	.w1(32'hbbd9b11c),
	.w2(32'h3b207203),
	.w3(32'hbc0b2e6e),
	.w4(32'hbb7328f8),
	.w5(32'h3a27f4bc),
	.w6(32'hbbf3aa3e),
	.w7(32'h3a00e219),
	.w8(32'h3afa6c60),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e747a),
	.w1(32'hb91f747c),
	.w2(32'h3ac3f696),
	.w3(32'hb8dee525),
	.w4(32'h3c17d085),
	.w5(32'h3c068c25),
	.w6(32'h39ac5b8d),
	.w7(32'h3c662cc9),
	.w8(32'h3bb87a30),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75b6e6),
	.w1(32'hbb37b03f),
	.w2(32'h3abdfe92),
	.w3(32'h3ba53279),
	.w4(32'hb948989a),
	.w5(32'hbb8ffe80),
	.w6(32'h3b74f46b),
	.w7(32'h3b63e539),
	.w8(32'hb9422e4f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf8aa4),
	.w1(32'hbb339b47),
	.w2(32'hbbd07421),
	.w3(32'hbb85d038),
	.w4(32'hbab500bb),
	.w5(32'hbbf6dfaa),
	.w6(32'hbb0b1ff1),
	.w7(32'h3bba261b),
	.w8(32'hbb730be5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099965),
	.w1(32'hbbbd6d21),
	.w2(32'hbb33b3d7),
	.w3(32'hbbfcd5fc),
	.w4(32'h3bfc0148),
	.w5(32'h3b78dff3),
	.w6(32'hbb145962),
	.w7(32'hba11ae5f),
	.w8(32'hbaa2034c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc02859),
	.w1(32'hbb29444c),
	.w2(32'hbb72852a),
	.w3(32'hbb1864c6),
	.w4(32'h3a9c7ea5),
	.w5(32'hbbe63e28),
	.w6(32'hbb9b01d3),
	.w7(32'h3afa739e),
	.w8(32'hba1d722f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c6e4),
	.w1(32'hbb383a49),
	.w2(32'hbc0822a5),
	.w3(32'hbb696eb6),
	.w4(32'h3c8b997d),
	.w5(32'h3bcf10d2),
	.w6(32'hbb285b7e),
	.w7(32'h39db6c2f),
	.w8(32'hbb7e7e39),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d475b9),
	.w1(32'h3b341c8d),
	.w2(32'h3c00f9e1),
	.w3(32'hbb261e54),
	.w4(32'hbc27499e),
	.w5(32'hbc279ee4),
	.w6(32'hbb2dd461),
	.w7(32'h3b8b0b2f),
	.w8(32'hbb88be84),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba528c4),
	.w1(32'h3b5d4183),
	.w2(32'hba2d898c),
	.w3(32'hbc4342cf),
	.w4(32'hbb7ad482),
	.w5(32'hbb376d8b),
	.w6(32'hbb07c81f),
	.w7(32'hbbf65cc0),
	.w8(32'hbc098dc5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9165e6),
	.w1(32'h39a9bbc7),
	.w2(32'hbbe75123),
	.w3(32'hbaf4efd9),
	.w4(32'hbb378da9),
	.w5(32'hbb7eb823),
	.w6(32'hbb21750d),
	.w7(32'hbb7c5f8f),
	.w8(32'hbbd68038),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe65781),
	.w1(32'hbc0eeaa3),
	.w2(32'hba7222ce),
	.w3(32'hbbdfd836),
	.w4(32'h3a78ff97),
	.w5(32'h39a4897c),
	.w6(32'hbc274c67),
	.w7(32'h3865e310),
	.w8(32'h3989f587),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3848e3cb),
	.w1(32'h39ac73d7),
	.w2(32'h39ea0703),
	.w3(32'h398eee82),
	.w4(32'h39ea0261),
	.w5(32'h3a36ec95),
	.w6(32'h390863de),
	.w7(32'h39cf4c44),
	.w8(32'h3a0d079a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d5d8ea),
	.w1(32'h36562c02),
	.w2(32'hb7a8f0c5),
	.w3(32'h3822acb0),
	.w4(32'h373247af),
	.w5(32'hb7b6cfd2),
	.w6(32'h3821dcdc),
	.w7(32'h37077e52),
	.w8(32'hb7d2d84a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8465e66),
	.w1(32'hb88f3703),
	.w2(32'hb81a426e),
	.w3(32'hb84caf23),
	.w4(32'hb79501b8),
	.w5(32'hb7aa2c0a),
	.w6(32'hb824b5bf),
	.w7(32'hb811af52),
	.w8(32'hb81d9fa0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2876c6),
	.w1(32'hb96de157),
	.w2(32'hba0eb29f),
	.w3(32'hb98fc6b1),
	.w4(32'h386351d5),
	.w5(32'hba12d9ba),
	.w6(32'hba59f3cb),
	.w7(32'hb961b8f4),
	.w8(32'hba2a28a1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bae266),
	.w1(32'h3708d98b),
	.w2(32'h38dfc371),
	.w3(32'hba1b0eff),
	.w4(32'h3a44b692),
	.w5(32'h3a252598),
	.w6(32'h39e9fca8),
	.w7(32'h3a434273),
	.w8(32'h399606f8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba974cae),
	.w1(32'hba8c2df3),
	.w2(32'hb9b031c4),
	.w3(32'hba282375),
	.w4(32'hbae10ca1),
	.w5(32'hbadb72c5),
	.w6(32'hb7d9c362),
	.w7(32'h38a926c0),
	.w8(32'hba3059b9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39823a7f),
	.w1(32'h3b17fa9c),
	.w2(32'h3b65f6f6),
	.w3(32'h3aedbecf),
	.w4(32'h3b9e1121),
	.w5(32'h3b8f8e4c),
	.w6(32'h3ad4582e),
	.w7(32'h3bbcb640),
	.w8(32'h3bbaffe8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e8bef),
	.w1(32'hb8837ec3),
	.w2(32'hb9313d08),
	.w3(32'hba87976c),
	.w4(32'hb7bc709c),
	.w5(32'h39822305),
	.w6(32'hba01cf3e),
	.w7(32'hb9693ca3),
	.w8(32'h39214597),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0fb0c),
	.w1(32'h3986459b),
	.w2(32'h3a855282),
	.w3(32'hb9cb18e9),
	.w4(32'h3a2df6a3),
	.w5(32'h3aa8d0af),
	.w6(32'hb9ff2d2e),
	.w7(32'h3a3138bc),
	.w8(32'h3a70562b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a669f4),
	.w1(32'h3b8dbcbf),
	.w2(32'h3b909bdc),
	.w3(32'h3acb7b64),
	.w4(32'h3bbb592f),
	.w5(32'h3bb0ecc9),
	.w6(32'h3ad17311),
	.w7(32'h3b9ff59e),
	.w8(32'h3b96f50f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8ae53),
	.w1(32'h3aa168c3),
	.w2(32'h3a93e674),
	.w3(32'h39a933cd),
	.w4(32'h3aa335f1),
	.w5(32'h3b05d2eb),
	.w6(32'h3a248146),
	.w7(32'h3ab2845a),
	.w8(32'h3b0ab0f9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9013cbd),
	.w1(32'h38bd4357),
	.w2(32'hb96a819e),
	.w3(32'hb854a3e9),
	.w4(32'h399992ec),
	.w5(32'h381ad760),
	.w6(32'hb8f7b105),
	.w7(32'h3976bd88),
	.w8(32'hb8f0ae68),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397cb0da),
	.w1(32'h3a804334),
	.w2(32'h3a649cf7),
	.w3(32'h37369805),
	.w4(32'h3ae99593),
	.w5(32'h3b235d7a),
	.w6(32'h3a746263),
	.w7(32'h3af0d353),
	.w8(32'h3b0fe4f4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d8fb1),
	.w1(32'hb9aaf649),
	.w2(32'hba0b793d),
	.w3(32'hb9857d43),
	.w4(32'hb75263f8),
	.w5(32'hb95e8e89),
	.w6(32'hb968a0a9),
	.w7(32'h38b7abb3),
	.w8(32'hb8c61125),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9d74),
	.w1(32'h3b08a313),
	.w2(32'h3c5e2f26),
	.w3(32'hbb69ebff),
	.w4(32'hbbb52e57),
	.w5(32'h3b0e561b),
	.w6(32'hbbe36cce),
	.w7(32'hbb375326),
	.w8(32'hbb29a0e2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828d13b),
	.w1(32'h39d32773),
	.w2(32'h399835db),
	.w3(32'h39b1614e),
	.w4(32'h3a03ba8d),
	.w5(32'h39974575),
	.w6(32'h3980fcb7),
	.w7(32'h3a25eed4),
	.w8(32'h39d545d3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65c7b4),
	.w1(32'hb9beab73),
	.w2(32'hb91d0bef),
	.w3(32'hba563e0a),
	.w4(32'hb9641909),
	.w5(32'hb96f7ebb),
	.w6(32'hba717ed9),
	.w7(32'hb9dcadbb),
	.w8(32'hb9a56b97),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00cc64),
	.w1(32'hbad2765f),
	.w2(32'hbb2cf285),
	.w3(32'hbab0844d),
	.w4(32'hba5ebe1b),
	.w5(32'hbb09552e),
	.w6(32'hbaa4232f),
	.w7(32'hba71c0ae),
	.w8(32'hbb0d3062),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe27fe),
	.w1(32'hba9b2304),
	.w2(32'hba981a56),
	.w3(32'hba61267a),
	.w4(32'hb93f1e4b),
	.w5(32'h3759f2dc),
	.w6(32'hba6e7804),
	.w7(32'hb9d0ae0a),
	.w8(32'hb8a8da16),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83e063a),
	.w1(32'hb906f40f),
	.w2(32'hb9296042),
	.w3(32'hb85c037e),
	.w4(32'hb717d56b),
	.w5(32'hb5aff3cf),
	.w6(32'h392e1ea6),
	.w7(32'hb816e9fd),
	.w8(32'h3855f7d4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3fb60),
	.w1(32'h3814eb7d),
	.w2(32'h38288a5b),
	.w3(32'h39039514),
	.w4(32'h3889e594),
	.w5(32'h38146853),
	.w6(32'h39047822),
	.w7(32'h38260268),
	.w8(32'h38d6bac0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dfefd),
	.w1(32'h3a486428),
	.w2(32'h3a2569ea),
	.w3(32'h39213732),
	.w4(32'h3a38b741),
	.w5(32'h3ac1d112),
	.w6(32'h38333e18),
	.w7(32'h3a8800db),
	.w8(32'h3ad282ec),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b7f16),
	.w1(32'hba3add4e),
	.w2(32'hb9ffa78d),
	.w3(32'hba8c88fb),
	.w4(32'hbaa14a67),
	.w5(32'hba5e34c9),
	.w6(32'hb9ab3f6e),
	.w7(32'hb95965b9),
	.w8(32'hb807f119),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892327f),
	.w1(32'h377f3382),
	.w2(32'hb7d33efa),
	.w3(32'h37dac34a),
	.w4(32'h38abe51c),
	.w5(32'h381982e1),
	.w6(32'h3719b8ee),
	.w7(32'h38a7cf90),
	.w8(32'h3865e956),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7451f),
	.w1(32'hba1990a4),
	.w2(32'hb8de5824),
	.w3(32'hba56371e),
	.w4(32'h39b08c2f),
	.w5(32'h3a348a95),
	.w6(32'hba8789fc),
	.w7(32'hb8cb43c2),
	.w8(32'hb8f33c45),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86678df),
	.w1(32'hb903aebb),
	.w2(32'hb8c7d174),
	.w3(32'hb8e1cf95),
	.w4(32'hb7e81447),
	.w5(32'h39c2c07d),
	.w6(32'hb88e4960),
	.w7(32'h3909a5bb),
	.w8(32'h3a05b140),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882a964),
	.w1(32'h395e5395),
	.w2(32'h39b61546),
	.w3(32'h38648423),
	.w4(32'h38596b00),
	.w5(32'h3966ff19),
	.w6(32'h386026d8),
	.w7(32'hb8babb05),
	.w8(32'hb835555d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36133c),
	.w1(32'hbae35b6d),
	.w2(32'hba191211),
	.w3(32'hbb246714),
	.w4(32'hbaf59aa0),
	.w5(32'hb885920b),
	.w6(32'hbb15915c),
	.w7(32'hbb032e10),
	.w8(32'hba6ef5c5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9be718),
	.w1(32'hba17955a),
	.w2(32'hb9d3c99c),
	.w3(32'hba8939cc),
	.w4(32'hb9b50a8e),
	.w5(32'h397f11fd),
	.w6(32'hba18b681),
	.w7(32'hb89da147),
	.w8(32'hb9e1727f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2c44a),
	.w1(32'h39c8fb46),
	.w2(32'h39b45b65),
	.w3(32'h398bfb54),
	.w4(32'h39291f4f),
	.w5(32'h393b5d1a),
	.w6(32'h38942cdb),
	.w7(32'h391c9b4d),
	.w8(32'h39a70313),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba998cb6),
	.w1(32'hba0bc505),
	.w2(32'h38c968d6),
	.w3(32'hba1c6863),
	.w4(32'hb8189405),
	.w5(32'h3983c9d7),
	.w6(32'hba0029c7),
	.w7(32'hba0cb123),
	.w8(32'hb9fb0afc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17fe92),
	.w1(32'h3a381c82),
	.w2(32'h3a55dd68),
	.w3(32'hba5d888f),
	.w4(32'h39076014),
	.w5(32'hba8526f3),
	.w6(32'hba63bb39),
	.w7(32'h39163ac5),
	.w8(32'hba8018ac),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928fb8f),
	.w1(32'hb8a73697),
	.w2(32'hb9b59720),
	.w3(32'hb88641ca),
	.w4(32'hb9883e8f),
	.w5(32'hba09b306),
	.w6(32'hb982231a),
	.w7(32'hb93a9b21),
	.w8(32'hba053993),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38830d93),
	.w1(32'hb8b5b540),
	.w2(32'h38d87803),
	.w3(32'h391bc6de),
	.w4(32'h372cf3d0),
	.w5(32'h37ae15e4),
	.w6(32'h38bb0704),
	.w7(32'h3804567c),
	.w8(32'hb7ba5468),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90307),
	.w1(32'h3b139f7f),
	.w2(32'h3b44b894),
	.w3(32'h3b211c8a),
	.w4(32'h3b64cd31),
	.w5(32'h3b29c8e6),
	.w6(32'h3b175bd9),
	.w7(32'h3b82ead6),
	.w8(32'h3b0ca06a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8bdcb),
	.w1(32'h3a02034a),
	.w2(32'h3a0a8698),
	.w3(32'h37f87e1a),
	.w4(32'h3a206c1f),
	.w5(32'h3a0a9704),
	.w6(32'hb9049cfb),
	.w7(32'h3a1c2903),
	.w8(32'h39dc227e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0655b),
	.w1(32'h3a205182),
	.w2(32'hb901fb58),
	.w3(32'h3a138ae2),
	.w4(32'h3a9899a8),
	.w5(32'hb8093899),
	.w6(32'h39f596f2),
	.w7(32'h3a7bba68),
	.w8(32'hba00aa03),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdebee),
	.w1(32'hbade0bb9),
	.w2(32'hbac82da5),
	.w3(32'hbb210ffb),
	.w4(32'hbb14a7da),
	.w5(32'hbb2060a5),
	.w6(32'hbb2716a5),
	.w7(32'hbb23bea3),
	.w8(32'hbb43fa8b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79e22a),
	.w1(32'hbb1a74d7),
	.w2(32'h3a9a2375),
	.w3(32'hba589ee6),
	.w4(32'h3ac50578),
	.w5(32'h3a90cb0e),
	.w6(32'hbb1eec80),
	.w7(32'hb7d848d6),
	.w8(32'h39dd2061),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93db181),
	.w1(32'h3a496e3c),
	.w2(32'h3a783fa9),
	.w3(32'h3ab98985),
	.w4(32'h3b2f63ab),
	.w5(32'h3a48d0c5),
	.w6(32'h3a6df01b),
	.w7(32'h3b568a9b),
	.w8(32'h3b08cb4c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d06acd),
	.w1(32'h38362468),
	.w2(32'hb991d57a),
	.w3(32'hba10df8a),
	.w4(32'hb9513d59),
	.w5(32'hba1e0432),
	.w6(32'hba365789),
	.w7(32'h39a816df),
	.w8(32'h37704b02),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d4583),
	.w1(32'hb758d8d4),
	.w2(32'h38659d3d),
	.w3(32'h3893c310),
	.w4(32'hb72a08d3),
	.w5(32'hb6bef213),
	.w6(32'h38905b3c),
	.w7(32'h3809d375),
	.w8(32'hb86017ad),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145df8),
	.w1(32'hbafd90cc),
	.w2(32'hbb6548e3),
	.w3(32'hbaf4db4f),
	.w4(32'hbab2f016),
	.w5(32'hbb867848),
	.w6(32'h398280d1),
	.w7(32'h3895b43c),
	.w8(32'hbb5ded5a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d83cf),
	.w1(32'h3a58a6f1),
	.w2(32'h3a504d55),
	.w3(32'h39ad8c6b),
	.w4(32'h3a0ae209),
	.w5(32'h3a36c204),
	.w6(32'hb9214b15),
	.w7(32'h3a4d6240),
	.w8(32'h3a4d90c5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4c81),
	.w1(32'hba8726de),
	.w2(32'hba21be28),
	.w3(32'hbadb16be),
	.w4(32'hba7681ca),
	.w5(32'hbac8f366),
	.w6(32'hbab87800),
	.w7(32'hba348373),
	.w8(32'hba842d3a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dec1a2),
	.w1(32'h38ee8e67),
	.w2(32'h3a2fb9fc),
	.w3(32'hb9ae3d0a),
	.w4(32'h39128168),
	.w5(32'h39aba200),
	.w6(32'hb92fe870),
	.w7(32'hb9157ada),
	.w8(32'hb9ba1b0e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3849d3d6),
	.w1(32'h385bb1b9),
	.w2(32'hb91ada79),
	.w3(32'h397995a9),
	.w4(32'h3846e1de),
	.w5(32'h395d3ab7),
	.w6(32'h379b1b26),
	.w7(32'hb970b70e),
	.w8(32'hb9cd6028),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9030b45),
	.w1(32'hb9202310),
	.w2(32'hb6b6533e),
	.w3(32'hb81257cc),
	.w4(32'hb927e56e),
	.w5(32'hb8b8e28c),
	.w6(32'hb956e69e),
	.w7(32'h36c654d2),
	.w8(32'hb85d8f58),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849e584),
	.w1(32'hb8e6bd5a),
	.w2(32'h388cd9c2),
	.w3(32'hb95555e0),
	.w4(32'hb8f70eca),
	.w5(32'hb714fe2c),
	.w6(32'hb92e74da),
	.w7(32'hb925cd74),
	.w8(32'hb92af225),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74087b),
	.w1(32'hbb70f786),
	.w2(32'hbb309a32),
	.w3(32'hbb07a198),
	.w4(32'hbb034295),
	.w5(32'hbad71666),
	.w6(32'hbaccdeca),
	.w7(32'hba534b3d),
	.w8(32'hba3ed62b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21c7b8),
	.w1(32'hb9ca666d),
	.w2(32'h3958ff79),
	.w3(32'hb9e337c7),
	.w4(32'h39ac5e23),
	.w5(32'hb8a96656),
	.w6(32'h369da1ed),
	.w7(32'h3a5f8479),
	.w8(32'h3a959298),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c19af0),
	.w1(32'h395e4a5c),
	.w2(32'h399a1dad),
	.w3(32'hb91e4b4a),
	.w4(32'h38e152ae),
	.w5(32'h3a445348),
	.w6(32'h3904174d),
	.w7(32'h37e44b14),
	.w8(32'h3a425924),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba530d3a),
	.w1(32'hb9400d0a),
	.w2(32'hb74e7528),
	.w3(32'hb9c6b205),
	.w4(32'h389c1bc7),
	.w5(32'h3930cfc2),
	.w6(32'h39f941c9),
	.w7(32'h3a8bca04),
	.w8(32'h3a989b63),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5d63c),
	.w1(32'hba609997),
	.w2(32'hba80f208),
	.w3(32'hb9e94718),
	.w4(32'h3a47fa5c),
	.w5(32'h3a7ed8e3),
	.w6(32'h389d991b),
	.w7(32'h3a9648bb),
	.w8(32'h3ab1fbc3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984ead7),
	.w1(32'h39d3ce73),
	.w2(32'h3a18b692),
	.w3(32'hb9b8a098),
	.w4(32'hb8e6cebd),
	.w5(32'hb89a12a9),
	.w6(32'hb9eb52da),
	.w7(32'h3732f1a2),
	.w8(32'h387fd64e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912bb84),
	.w1(32'h3712e41b),
	.w2(32'h3942b060),
	.w3(32'hb922cc19),
	.w4(32'hb512aa93),
	.w5(32'h395ac3d1),
	.w6(32'hb8818966),
	.w7(32'h367b4c8d),
	.w8(32'h3917a408),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8de2c),
	.w1(32'hbb106859),
	.w2(32'h397349a8),
	.w3(32'hbba02b07),
	.w4(32'hba7817d7),
	.w5(32'h3ad7f974),
	.w6(32'hbba11c98),
	.w7(32'hbaa24910),
	.w8(32'h3a0d4526),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b5526c),
	.w1(32'h390f4a96),
	.w2(32'h39446e31),
	.w3(32'hb883e904),
	.w4(32'h38d00855),
	.w5(32'h38a1d009),
	.w6(32'hb8eddb80),
	.w7(32'h385cf333),
	.w8(32'h384c3123),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae819e6),
	.w1(32'hba0ce280),
	.w2(32'h3a3a2d5e),
	.w3(32'hba277d68),
	.w4(32'h3a3e2f7b),
	.w5(32'h3ae8551a),
	.w6(32'hb9d40559),
	.w7(32'h3a8afa18),
	.w8(32'h3adea922),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c0b71),
	.w1(32'hb92a49c1),
	.w2(32'hb9202e58),
	.w3(32'hb986d827),
	.w4(32'hb9982ccd),
	.w5(32'hb96269e0),
	.w6(32'hb96c1f5d),
	.w7(32'hb96e86d3),
	.w8(32'hb966c463),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997aee),
	.w1(32'hbb7baaee),
	.w2(32'hbb7179f1),
	.w3(32'hbb57e532),
	.w4(32'hbaec8f4a),
	.w5(32'hbb08250f),
	.w6(32'hbb2a3867),
	.w7(32'hbb1c6b2a),
	.w8(32'hbb00071d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3825ba1e),
	.w1(32'h373e6213),
	.w2(32'h3892531a),
	.w3(32'h38b92c42),
	.w4(32'h3899b4b1),
	.w5(32'h38b8e460),
	.w6(32'hb88371d6),
	.w7(32'h389e6157),
	.w8(32'hb8297f09),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10cb57),
	.w1(32'h3990e4ff),
	.w2(32'hba761d8c),
	.w3(32'hb9e800bd),
	.w4(32'h3a1bb2df),
	.w5(32'hb910b2c0),
	.w6(32'hba14c3a5),
	.w7(32'h390bd814),
	.w8(32'hba00f5e5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37782cda),
	.w1(32'hb7a9de02),
	.w2(32'hb9c5e704),
	.w3(32'hb7614c06),
	.w4(32'h3b8377a4),
	.w5(32'h3a98dcd6),
	.w6(32'hb8340501),
	.w7(32'h3b5821d7),
	.w8(32'h3b04f0b7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dcfd6),
	.w1(32'h3a3a8e40),
	.w2(32'hba608238),
	.w3(32'h3b8b2a78),
	.w4(32'hbb8cba78),
	.w5(32'hbb943956),
	.w6(32'h3bb4f2f6),
	.w7(32'hbb48e60d),
	.w8(32'hbc125ae7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4dc25),
	.w1(32'h3ba21971),
	.w2(32'hbbf6247e),
	.w3(32'h3ac1c745),
	.w4(32'hbc1b4a69),
	.w5(32'hbb7b4455),
	.w6(32'h3a91dae8),
	.w7(32'hbc3b3b52),
	.w8(32'hbbcacfc1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97f84),
	.w1(32'hba31c9a1),
	.w2(32'hbc9d930f),
	.w3(32'hbb3232fb),
	.w4(32'h3c52cb99),
	.w5(32'h3c1cc02e),
	.w6(32'hbb2dd431),
	.w7(32'hbb8f5693),
	.w8(32'h3cf61a6f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c234244),
	.w1(32'hbbe54b9a),
	.w2(32'h3cb0676c),
	.w3(32'hbcb91242),
	.w4(32'h3c52bc5d),
	.w5(32'hbc7d19a5),
	.w6(32'hbbf8bb08),
	.w7(32'h3d03f27e),
	.w8(32'hbcc5bf25),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd9f1e),
	.w1(32'hbbd0d03c),
	.w2(32'h3d115409),
	.w3(32'hbb93b2c0),
	.w4(32'h3ca348d9),
	.w5(32'hbc8df5b4),
	.w6(32'h3a87ec87),
	.w7(32'h3c753e26),
	.w8(32'hbd2eed6d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04e24e),
	.w1(32'h3cd73667),
	.w2(32'h3b80af6d),
	.w3(32'h3c28d2db),
	.w4(32'hbacdb499),
	.w5(32'h3b59b1bf),
	.w6(32'h3d388e0c),
	.w7(32'hbb82db29),
	.w8(32'hbb34b3a1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07e375),
	.w1(32'hbbc38e73),
	.w2(32'h3bb44282),
	.w3(32'h3a123eb4),
	.w4(32'hbc942daa),
	.w5(32'h3b252dd2),
	.w6(32'hbb8a9902),
	.w7(32'hbd06f7ae),
	.w8(32'h390426b1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b5a61),
	.w1(32'hba571e98),
	.w2(32'hbc691235),
	.w3(32'hbc170a90),
	.w4(32'h3b25a920),
	.w5(32'hbbaadd0b),
	.w6(32'h3c58ab51),
	.w7(32'hbc8cdb55),
	.w8(32'hbbc09b76),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c440011),
	.w1(32'h3b7ea05e),
	.w2(32'hbbc6b1db),
	.w3(32'hb892f657),
	.w4(32'hbb456cec),
	.w5(32'hbc4d8554),
	.w6(32'h3c615555),
	.w7(32'hbbe21387),
	.w8(32'h3b8f5562),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb011b6),
	.w1(32'hbc68ed42),
	.w2(32'hbd0013a1),
	.w3(32'hbc921716),
	.w4(32'hbc5c9327),
	.w5(32'hbb294cf5),
	.w6(32'hbc2007f4),
	.w7(32'hbcaa4919),
	.w8(32'hbb445527),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47f354),
	.w1(32'h3a94c097),
	.w2(32'h3b04199f),
	.w3(32'hbc258744),
	.w4(32'h3aa0257c),
	.w5(32'hbc2757ed),
	.w6(32'h3c1ea6d2),
	.w7(32'h3c1d8151),
	.w8(32'hb9411892),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0640ba),
	.w1(32'hbb6052af),
	.w2(32'hbb20d825),
	.w3(32'hba397339),
	.w4(32'h39c263cc),
	.w5(32'h3b9fffca),
	.w6(32'h3a02b6f1),
	.w7(32'hbb95d67f),
	.w8(32'hbb91a4e7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55353),
	.w1(32'hbb8a73b8),
	.w2(32'h3cbff6b1),
	.w3(32'hbbcbe98a),
	.w4(32'h3c6569a3),
	.w5(32'hbc998d2c),
	.w6(32'hbb2a4b00),
	.w7(32'h3d3a2593),
	.w8(32'hbbc936a7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9038e6),
	.w1(32'hbc962815),
	.w2(32'hbc2b2a98),
	.w3(32'h3b1d2816),
	.w4(32'h3a93cdd2),
	.w5(32'h3c3b80b0),
	.w6(32'hbb4bc06c),
	.w7(32'hbcc66276),
	.w8(32'h3c841cff),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0081da),
	.w1(32'hbbf1046c),
	.w2(32'hbcc03f01),
	.w3(32'hbc442d86),
	.w4(32'hbc653b48),
	.w5(32'hbcc4c0c6),
	.w6(32'hbbbbfa0f),
	.w7(32'hbcf62e86),
	.w8(32'hbc0f4a80),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c151495),
	.w1(32'h3cb41f3a),
	.w2(32'hba63485e),
	.w3(32'h3c045244),
	.w4(32'hbc511f00),
	.w5(32'hbbf8c95d),
	.w6(32'h3d0085a0),
	.w7(32'hbc892b3c),
	.w8(32'h3cd03649),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfc020a),
	.w1(32'hbb5bbba0),
	.w2(32'h3bc34609),
	.w3(32'hbbb32102),
	.w4(32'hbc045495),
	.w5(32'h3b1cd65b),
	.w6(32'hbb87d1dd),
	.w7(32'h3c70f683),
	.w8(32'hbbbd67f4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7cde3),
	.w1(32'hbba4d3e9),
	.w2(32'hb99ccfc4),
	.w3(32'hbc389992),
	.w4(32'hba53b756),
	.w5(32'h3b9b31dd),
	.w6(32'hbc55debc),
	.w7(32'h3b7ac626),
	.w8(32'h3c058694),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60f718),
	.w1(32'h3abedc65),
	.w2(32'hbd137d21),
	.w3(32'h3abaf2a0),
	.w4(32'hbc5a22cf),
	.w5(32'hbb3311d9),
	.w6(32'h3bb54738),
	.w7(32'hbd132792),
	.w8(32'h3c9eec26),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19730d),
	.w1(32'h3c912f2f),
	.w2(32'h3d07fe81),
	.w3(32'h3bc8e502),
	.w4(32'h3c722f25),
	.w5(32'hbc6b05bb),
	.w6(32'h3c770842),
	.w7(32'h3d4e6726),
	.w8(32'hbc7a0cb7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92d4ed),
	.w1(32'hbcc81e38),
	.w2(32'h3b2bf652),
	.w3(32'hbb042b23),
	.w4(32'hbb5486ba),
	.w5(32'h3c29f4ba),
	.w6(32'hbbfe5909),
	.w7(32'h3cfc6823),
	.w8(32'hbaa22dc0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2129ce),
	.w1(32'hbcbfc6a5),
	.w2(32'h3c6d5fd7),
	.w3(32'hbc3b3ae1),
	.w4(32'h3c6dc08c),
	.w5(32'h3b667c20),
	.w6(32'hbce3c94d),
	.w7(32'h3c7e524f),
	.w8(32'h3b0ab6e7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0ebfe),
	.w1(32'hbabea740),
	.w2(32'hba715e7a),
	.w3(32'h3a47bce4),
	.w4(32'h3bf1e33b),
	.w5(32'hbbe48805),
	.w6(32'hbb943aff),
	.w7(32'h3cafb75e),
	.w8(32'hbc3203f3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28647c),
	.w1(32'h3c54e5ab),
	.w2(32'hbd14dc3a),
	.w3(32'h3c8b9c55),
	.w4(32'hbc77acdf),
	.w5(32'hba1f8329),
	.w6(32'h3c16824c),
	.w7(32'hbd28dbd1),
	.w8(32'hbbb63ef0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051fbf),
	.w1(32'h3c7ec829),
	.w2(32'h3ba4a642),
	.w3(32'hbc4cc128),
	.w4(32'h3acd86dd),
	.w5(32'hbbaa2ac6),
	.w6(32'h3c81434b),
	.w7(32'h3d02dbac),
	.w8(32'hbc4ec2e8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc815e26),
	.w1(32'hbc968ba6),
	.w2(32'hbc0a1f5c),
	.w3(32'hbc5b3e73),
	.w4(32'hbb5c2984),
	.w5(32'hbbbbdb26),
	.w6(32'hbc801a34),
	.w7(32'hbc494fbc),
	.w8(32'h3bde4b26),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf517f),
	.w1(32'hbc35dcdc),
	.w2(32'hbb06d37d),
	.w3(32'hbb70b270),
	.w4(32'h3c0d7c45),
	.w5(32'h3c7a43a1),
	.w6(32'hba8bb7b1),
	.w7(32'hbc348cb6),
	.w8(32'h3c30208d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e5749),
	.w1(32'h3bda2bf4),
	.w2(32'hbc3b2f47),
	.w3(32'hbbbf18cb),
	.w4(32'hbc0a8175),
	.w5(32'h3bdad247),
	.w6(32'h3b622d84),
	.w7(32'hbccf1bd7),
	.w8(32'h3d0369b9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babdf1a),
	.w1(32'hbcc58906),
	.w2(32'hbd17a8ac),
	.w3(32'hbcb02d68),
	.w4(32'hbc4ffadc),
	.w5(32'h3c2beade),
	.w6(32'hbcc353c4),
	.w7(32'hbcf32dc3),
	.w8(32'h3c16bf96),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c7191),
	.w1(32'h3cb0bb6a),
	.w2(32'h3c588e7b),
	.w3(32'h3c2b10a1),
	.w4(32'h3c18a64d),
	.w5(32'hbb26b93f),
	.w6(32'h3cd370be),
	.w7(32'h3d12a50d),
	.w8(32'hbc392c7f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc442b0e),
	.w1(32'hbc337eee),
	.w2(32'h3a13aab5),
	.w3(32'hbb4af94c),
	.w4(32'h3b001afb),
	.w5(32'h3ab41e31),
	.w6(32'hbcb6b638),
	.w7(32'h3be2cae8),
	.w8(32'h3bcf75fc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3434e4),
	.w1(32'hbaa7c5f1),
	.w2(32'h3c22f9ea),
	.w3(32'hba3426a4),
	.w4(32'hbb56781b),
	.w5(32'hbc54b0c4),
	.w6(32'h3b40973e),
	.w7(32'h3baf90ca),
	.w8(32'hbc06c523),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b377712),
	.w1(32'hbc393215),
	.w2(32'hbcc20836),
	.w3(32'h3c0fdd4c),
	.w4(32'h3c0428df),
	.w5(32'hbb51bfa6),
	.w6(32'hbaa07739),
	.w7(32'hbc4871de),
	.w8(32'h3c06d52e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd7714),
	.w1(32'hbbf6d1f2),
	.w2(32'hba0fabb6),
	.w3(32'hbc38fd0e),
	.w4(32'hbc6f610a),
	.w5(32'hbbb0118c),
	.w6(32'hbc00e5e3),
	.w7(32'hbcf9bbeb),
	.w8(32'h3b1f2907),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f85bc),
	.w1(32'h3cd68267),
	.w2(32'h3a192f65),
	.w3(32'hbbce5df3),
	.w4(32'h3be40e4b),
	.w5(32'hbcaef58e),
	.w6(32'h3c678035),
	.w7(32'h3ccb574e),
	.w8(32'hbc592b39),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db2ae),
	.w1(32'hbae86ef0),
	.w2(32'hbccba386),
	.w3(32'h3ba2fb28),
	.w4(32'hbc5ab401),
	.w5(32'h3baef088),
	.w6(32'h3b824de1),
	.w7(32'hbd140b82),
	.w8(32'h3ce9c22a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90a2fe),
	.w1(32'hbbb1574d),
	.w2(32'hbcc7bf7d),
	.w3(32'hbc1e513b),
	.w4(32'hbca8e506),
	.w5(32'hbc38bade),
	.w6(32'h3b414ded),
	.w7(32'hbcea3c2f),
	.w8(32'h3ca52fff),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe35644),
	.w1(32'hbc742683),
	.w2(32'h3c98c848),
	.w3(32'hbcb1a8a6),
	.w4(32'h37667bd5),
	.w5(32'h3c7193c3),
	.w6(32'h3ab5c6cf),
	.w7(32'h3d519ddb),
	.w8(32'hbc77563f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd051fa5),
	.w1(32'hbc07e619),
	.w2(32'hbaabb718),
	.w3(32'hbbf6e54f),
	.w4(32'h3c52193d),
	.w5(32'hbc3b9398),
	.w6(32'hbcc2a766),
	.w7(32'hbb6b948c),
	.w8(32'hbce0d325),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f38a),
	.w1(32'h3ce2c042),
	.w2(32'hbb9c4b1e),
	.w3(32'h3c8a1d1b),
	.w4(32'hba5425e3),
	.w5(32'hbc7a9618),
	.w6(32'h3cbe5308),
	.w7(32'hbc132ca2),
	.w8(32'hbd02cfe0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc392f0c),
	.w1(32'h3ce0a2d5),
	.w2(32'h3a1fac68),
	.w3(32'h3c9b162f),
	.w4(32'hb9f23d9a),
	.w5(32'h38b77eac),
	.w6(32'h3c8f17a1),
	.w7(32'h3acd2853),
	.w8(32'hb96a82ed),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba850e9f),
	.w1(32'hba884bd1),
	.w2(32'hbb5e192d),
	.w3(32'h3a8f9764),
	.w4(32'hbca27b10),
	.w5(32'hbc4757b8),
	.w6(32'h3a9ed53e),
	.w7(32'hbcf9c941),
	.w8(32'hba5d8657),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06c813),
	.w1(32'hbb8882da),
	.w2(32'h3b3a8f97),
	.w3(32'h3bed7696),
	.w4(32'hbb894e8a),
	.w5(32'hbba10d66),
	.w6(32'h3c75b702),
	.w7(32'h3b424481),
	.w8(32'h3c8c9253),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ee14e),
	.w1(32'hbc9f5824),
	.w2(32'hbb29d69d),
	.w3(32'hbc9fb454),
	.w4(32'h3a830197),
	.w5(32'hbbe2a93a),
	.w6(32'hbc980be3),
	.w7(32'hbb41bfc8),
	.w8(32'hbb868e0f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f5f07),
	.w1(32'h3c0bdd09),
	.w2(32'h3cffa94c),
	.w3(32'hb9e70aa9),
	.w4(32'h3c8addb9),
	.w5(32'h3b6a90dc),
	.w6(32'h3c488205),
	.w7(32'h3d2695b5),
	.w8(32'hbc93b37c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83985e),
	.w1(32'hbc1c8461),
	.w2(32'hba93af57),
	.w3(32'hbbe2e26e),
	.w4(32'hbadf73ae),
	.w5(32'hba69bb79),
	.w6(32'hbce0657b),
	.w7(32'h3b9463b9),
	.w8(32'h3b6e6593),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd480d),
	.w1(32'hbad403ba),
	.w2(32'hbc2e9b60),
	.w3(32'hb9a7d885),
	.w4(32'h388180a0),
	.w5(32'hbb8ae32e),
	.w6(32'h3b0b70cb),
	.w7(32'hbb8a5b27),
	.w8(32'hbbf372b3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939e491),
	.w1(32'hbb9f8a33),
	.w2(32'h3ce4afa3),
	.w3(32'hbb3f37c6),
	.w4(32'hba94b27f),
	.w5(32'h3a0b359a),
	.w6(32'hbbb5dcd6),
	.w7(32'h3d1af455),
	.w8(32'hbc1315b2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19b3a9),
	.w1(32'h3adba53c),
	.w2(32'h3916f716),
	.w3(32'h3b73fa27),
	.w4(32'h3b21b9b9),
	.w5(32'hbb88d46e),
	.w6(32'h3b55aae6),
	.w7(32'h3b9f1d98),
	.w8(32'hbb97c108),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab16f),
	.w1(32'hbaf94c7b),
	.w2(32'hbc22682b),
	.w3(32'hbb09ec8e),
	.w4(32'hbc89389d),
	.w5(32'hbc5aeea4),
	.w6(32'h3b7e770f),
	.w7(32'hbac2a8c9),
	.w8(32'h3c852410),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9423d5),
	.w1(32'hbb903b34),
	.w2(32'h3b4bb693),
	.w3(32'h3c74a2c7),
	.w4(32'hbc0c126e),
	.w5(32'h3c63b9c4),
	.w6(32'h3bad5db4),
	.w7(32'hbc6713e6),
	.w8(32'h3cc8d5d5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule