module layer_10_featuremap_412(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb444813),
	.w1(32'h3ac28f54),
	.w2(32'hbb0d1c49),
	.w3(32'h3aa5f467),
	.w4(32'h3b83dcc3),
	.w5(32'h3b5be2d6),
	.w6(32'h3bfeeab2),
	.w7(32'h39fe69ac),
	.w8(32'hba5cff47),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942964),
	.w1(32'hb9c1c9e6),
	.w2(32'hbada4289),
	.w3(32'h3b132017),
	.w4(32'hbb32f6f2),
	.w5(32'hbb52b54d),
	.w6(32'hbb8c3e21),
	.w7(32'hbbe1727b),
	.w8(32'hbbb4c152),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec7b6),
	.w1(32'h3b496d5a),
	.w2(32'hba725042),
	.w3(32'hbaae766d),
	.w4(32'hb9aabb37),
	.w5(32'h3b4d5802),
	.w6(32'h3840a872),
	.w7(32'hbb1309ef),
	.w8(32'hbb8b2881),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4db99d),
	.w1(32'hbb46779e),
	.w2(32'hba46cc8d),
	.w3(32'h38840a62),
	.w4(32'hbaf1da36),
	.w5(32'h3b3aac8a),
	.w6(32'hba73008d),
	.w7(32'h3b63d842),
	.w8(32'hbb8b69f0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1b9f2),
	.w1(32'h3a276ed8),
	.w2(32'hbb595765),
	.w3(32'hbba60c88),
	.w4(32'h3bd2e255),
	.w5(32'h3c0be3a9),
	.w6(32'hbb6a33a5),
	.w7(32'h3b0ffd53),
	.w8(32'h3c211047),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80cbfc),
	.w1(32'h3c38dbdf),
	.w2(32'h3ca6d28e),
	.w3(32'h3b7eace7),
	.w4(32'h3caf5190),
	.w5(32'h3c971c73),
	.w6(32'h3af84ed3),
	.w7(32'h3bdc7539),
	.w8(32'hbb19e403),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab59b9d),
	.w1(32'hbc04663a),
	.w2(32'hbc593af5),
	.w3(32'h3c8c8544),
	.w4(32'hbc30bab2),
	.w5(32'h3aa08cc0),
	.w6(32'h3b943a51),
	.w7(32'hbb218366),
	.w8(32'hbb504ee1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a512b),
	.w1(32'hbac6850d),
	.w2(32'hbba536b7),
	.w3(32'hbc238d2b),
	.w4(32'hbc1c9f16),
	.w5(32'hbc54da25),
	.w6(32'hbc54c07b),
	.w7(32'hbb829c97),
	.w8(32'hba4271c0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945046c),
	.w1(32'h3ab04abc),
	.w2(32'hbb11b40c),
	.w3(32'hbb40655d),
	.w4(32'hbb9c6783),
	.w5(32'hba59578c),
	.w6(32'h3b8158eb),
	.w7(32'hbbb689e0),
	.w8(32'hbb9b674c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aeabe),
	.w1(32'h3bc199f6),
	.w2(32'h3b4ec036),
	.w3(32'h3aeb0f46),
	.w4(32'h3c630c4b),
	.w5(32'h3c0377e8),
	.w6(32'hbb9771a5),
	.w7(32'hbb98d16a),
	.w8(32'hbc53697f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7223e),
	.w1(32'hbb14683a),
	.w2(32'h3b749c49),
	.w3(32'hbae0fc66),
	.w4(32'h3a78f005),
	.w5(32'h3ba2f8dd),
	.w6(32'hbc33bd73),
	.w7(32'hbc1cc469),
	.w8(32'hbb432615),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba41e2d),
	.w1(32'hbc2a0b9a),
	.w2(32'hbbafb2fd),
	.w3(32'h39857e24),
	.w4(32'hbbff4b6c),
	.w5(32'hbbdca36b),
	.w6(32'hbbc9c2be),
	.w7(32'hbbae79af),
	.w8(32'h3a9ff4b7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f05c),
	.w1(32'h3b0b6c0c),
	.w2(32'hbacd21b2),
	.w3(32'hbbab2631),
	.w4(32'h3bd899a8),
	.w5(32'hbc14c9f9),
	.w6(32'hbbc97899),
	.w7(32'h3b60430b),
	.w8(32'h3bba1ea7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe90b4),
	.w1(32'hbb1e78d1),
	.w2(32'hbbc9e131),
	.w3(32'h3b7dfa27),
	.w4(32'hba80c0bf),
	.w5(32'hbaa6d731),
	.w6(32'h3b0b0072),
	.w7(32'hbacba4de),
	.w8(32'h3b4130f6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac2bb1),
	.w1(32'h3a0df5db),
	.w2(32'hbb0325c6),
	.w3(32'hbb4b782e),
	.w4(32'hbbd7f5d6),
	.w5(32'hba8e67eb),
	.w6(32'h3b530a4a),
	.w7(32'h3b73c53b),
	.w8(32'h3a216013),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6e7c),
	.w1(32'hbc1ea01f),
	.w2(32'hbc37be66),
	.w3(32'h3b5dabbd),
	.w4(32'hbbb0a333),
	.w5(32'hbbe22926),
	.w6(32'hb9c741b3),
	.w7(32'hbb836466),
	.w8(32'hbb6d8365),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf66447),
	.w1(32'h3c87974f),
	.w2(32'h3c0ee68e),
	.w3(32'hbbef08d5),
	.w4(32'hbb8234e1),
	.w5(32'hbc51b383),
	.w6(32'hb9df6987),
	.w7(32'hbb00ed68),
	.w8(32'hbbc23540),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a242),
	.w1(32'h3b2fbf26),
	.w2(32'h38844498),
	.w3(32'hbc3e202c),
	.w4(32'h3ad9fcfa),
	.w5(32'hbb8f9472),
	.w6(32'hbc685db0),
	.w7(32'hbbf812a0),
	.w8(32'hbb859310),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d1c30),
	.w1(32'h3ace63c0),
	.w2(32'hbb2ae90b),
	.w3(32'h3bb7a5c8),
	.w4(32'hbb7383ce),
	.w5(32'hbc19c801),
	.w6(32'hbb848578),
	.w7(32'hbbe90223),
	.w8(32'hbbd38cd8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabe5db),
	.w1(32'hbaec3b16),
	.w2(32'hbbc887d1),
	.w3(32'hbab34afd),
	.w4(32'hbb3fce41),
	.w5(32'hbc156791),
	.w6(32'hbbb86686),
	.w7(32'h3c05e8f1),
	.w8(32'hbb1512ba),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1af25d),
	.w1(32'h3c0c43a0),
	.w2(32'h3c2bd0d5),
	.w3(32'hbb6e123e),
	.w4(32'h3b2fb23e),
	.w5(32'hbb88ac14),
	.w6(32'hbc3e321d),
	.w7(32'hb95c19b8),
	.w8(32'hba3a7294),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ba533),
	.w1(32'h3c250c11),
	.w2(32'h3c0fb090),
	.w3(32'h3a0d164b),
	.w4(32'h3c038e19),
	.w5(32'hba264c12),
	.w6(32'hbb16cc05),
	.w7(32'h3c1e7257),
	.w8(32'h3a7a1c6d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1e79d),
	.w1(32'hbba50880),
	.w2(32'h3c320e82),
	.w3(32'hbbd14a1a),
	.w4(32'h3c83d742),
	.w5(32'h3d285cc4),
	.w6(32'hbb79b032),
	.w7(32'h3b82529f),
	.w8(32'hbc35da9e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ab5ad),
	.w1(32'h3b74d005),
	.w2(32'h3b1a8e82),
	.w3(32'h3b7168ce),
	.w4(32'hbb8b1e41),
	.w5(32'hbb3c55e8),
	.w6(32'h3bd98e35),
	.w7(32'hbbad79e1),
	.w8(32'hbb2bca55),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4e133),
	.w1(32'h3a2ced5c),
	.w2(32'hbb2c1bc4),
	.w3(32'hbc84d985),
	.w4(32'hbbd18673),
	.w5(32'h3bd2c4d9),
	.w6(32'hbc8af35d),
	.w7(32'h3bb60db5),
	.w8(32'hbb26770e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb223826),
	.w1(32'h3bda0d80),
	.w2(32'hba1864a8),
	.w3(32'hb811f30c),
	.w4(32'h3af77dd1),
	.w5(32'h3bcf3e1d),
	.w6(32'h3b98d662),
	.w7(32'h3bcbe9fd),
	.w8(32'h3b217116),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee3ed0),
	.w1(32'h3bd1173b),
	.w2(32'h3b9cce34),
	.w3(32'hbb964424),
	.w4(32'hba016161),
	.w5(32'hbc4e75d2),
	.w6(32'hbb7fb0b2),
	.w7(32'hbbf193ee),
	.w8(32'hbc2feb68),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60533e),
	.w1(32'h3ba9ee18),
	.w2(32'h3bc4ac27),
	.w3(32'hbc3dfd24),
	.w4(32'h3b99edfc),
	.w5(32'h3c77e1bf),
	.w6(32'hbc08d521),
	.w7(32'h3c318565),
	.w8(32'h3b99db4f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fdb8c),
	.w1(32'h3b1bf368),
	.w2(32'h3bb80c24),
	.w3(32'hbbf835a2),
	.w4(32'h3c105704),
	.w5(32'hbb2bb6e7),
	.w6(32'hbbc560fc),
	.w7(32'hbb25e8a6),
	.w8(32'hbb1e1071),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55d6c8),
	.w1(32'h3c270199),
	.w2(32'hba920e84),
	.w3(32'hbbc57f10),
	.w4(32'h3a2aae61),
	.w5(32'hbb62b7d3),
	.w6(32'h3ba56956),
	.w7(32'hbbe726a8),
	.w8(32'hbc109141),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970c74),
	.w1(32'h39cbdd44),
	.w2(32'h3b2a750f),
	.w3(32'h3bc2fddf),
	.w4(32'hba8d60ff),
	.w5(32'h3ba9108a),
	.w6(32'hbae4a4b0),
	.w7(32'hba8979a0),
	.w8(32'hbb902430),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6948df),
	.w1(32'h3b74029a),
	.w2(32'hbb1fbf3d),
	.w3(32'h3ae934d3),
	.w4(32'hbb1d3548),
	.w5(32'h3ae05ca5),
	.w6(32'hbb7bf7dc),
	.w7(32'hbb90762b),
	.w8(32'hbb15c6d6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ddb23d),
	.w1(32'h3aad6e05),
	.w2(32'hbb44b88b),
	.w3(32'h3b5b67a8),
	.w4(32'h3bbc0485),
	.w5(32'h3be74cd7),
	.w6(32'hba942eba),
	.w7(32'h3bc40d96),
	.w8(32'h3bf44d52),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074593),
	.w1(32'h3bb77951),
	.w2(32'hbb368a0f),
	.w3(32'h3c02082d),
	.w4(32'h3bb0683e),
	.w5(32'h3cc4cf96),
	.w6(32'h39bb8092),
	.w7(32'h3ac2883b),
	.w8(32'hbb7f93b2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad263c6),
	.w1(32'hbb8446f7),
	.w2(32'h3aa3baa1),
	.w3(32'h3c08ec84),
	.w4(32'h3b15d934),
	.w5(32'hbb9e5156),
	.w6(32'hbba07c89),
	.w7(32'hbc2850be),
	.w8(32'h3b0f1980),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28866b),
	.w1(32'hbbb23c93),
	.w2(32'hbbc4ade2),
	.w3(32'h3bade6ef),
	.w4(32'hba85a38b),
	.w5(32'h3b9251ff),
	.w6(32'h392956d9),
	.w7(32'h3a9ceeb9),
	.w8(32'h3aa32fc6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64de7e),
	.w1(32'hbc68fed0),
	.w2(32'hbb802b6f),
	.w3(32'h3bac261b),
	.w4(32'h39b7faca),
	.w5(32'h3a2375b7),
	.w6(32'hbb12471c),
	.w7(32'hbbc12414),
	.w8(32'hbc2644dc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40e3e6),
	.w1(32'h3af7335a),
	.w2(32'h3b9b4bdc),
	.w3(32'hbc73b111),
	.w4(32'hbb0c9ace),
	.w5(32'h3b056a5c),
	.w6(32'hbc55525c),
	.w7(32'hbb124221),
	.w8(32'hbc2836b1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e19fe),
	.w1(32'hba9f8683),
	.w2(32'hbb017347),
	.w3(32'hbb05d2c0),
	.w4(32'hbb13afd1),
	.w5(32'hbb2dc0e9),
	.w6(32'hbbc07b7d),
	.w7(32'hbbec58dd),
	.w8(32'hbc1832af),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7cfca),
	.w1(32'h3af4a011),
	.w2(32'h3b42c05b),
	.w3(32'hbbc54c27),
	.w4(32'hbaf46588),
	.w5(32'h3bac3ff5),
	.w6(32'hbc16d584),
	.w7(32'h3bfd9da7),
	.w8(32'h3aba5434),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01bf87),
	.w1(32'hb9c9d62c),
	.w2(32'hbb3ac3cb),
	.w3(32'hbb7ce388),
	.w4(32'hbb5e5cde),
	.w5(32'hb945759b),
	.w6(32'hbb979442),
	.w7(32'h39fa19d2),
	.w8(32'h3bf5a913),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c01c),
	.w1(32'hbafb9e56),
	.w2(32'hbba23ff8),
	.w3(32'h3b95587f),
	.w4(32'hbb9863f2),
	.w5(32'hbb94d2ea),
	.w6(32'h3bb80637),
	.w7(32'hbb505fee),
	.w8(32'hbab35782),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb780cdc),
	.w1(32'h39a49daf),
	.w2(32'hba797790),
	.w3(32'h3ab68bf3),
	.w4(32'h3b97ed3b),
	.w5(32'h3b3e2a5d),
	.w6(32'hbb199f0d),
	.w7(32'h3a93d734),
	.w8(32'h3a829f39),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb996e4d),
	.w1(32'hba792d6d),
	.w2(32'hbb44d5d4),
	.w3(32'h3b5dc857),
	.w4(32'hbaaf3ab3),
	.w5(32'hbbdd0d53),
	.w6(32'hbaf32460),
	.w7(32'hbb485f72),
	.w8(32'hbc125811),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3f770),
	.w1(32'h3b6f3fcb),
	.w2(32'h3ba96b42),
	.w3(32'hbbdd7dcc),
	.w4(32'h3b61b82e),
	.w5(32'h3b9be05e),
	.w6(32'hbbaef68f),
	.w7(32'h390c6694),
	.w8(32'hbac6d66a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f23ae),
	.w1(32'hbb9f4177),
	.w2(32'hbc48668b),
	.w3(32'hba5230f6),
	.w4(32'hbc3469d1),
	.w5(32'hbbed85b5),
	.w6(32'hbb614e7b),
	.w7(32'hbbdd5d43),
	.w8(32'hbb3d9c2c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc661523),
	.w1(32'h3bb53799),
	.w2(32'h3c08fc3b),
	.w3(32'hbc4b1fa9),
	.w4(32'h3b623614),
	.w5(32'hbbb39e57),
	.w6(32'hbb9c1ef1),
	.w7(32'h3bcf7234),
	.w8(32'h3c21814b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2471),
	.w1(32'h3ae81649),
	.w2(32'hbc1afac0),
	.w3(32'hbb12434c),
	.w4(32'h3ab872ae),
	.w5(32'hbbf412cc),
	.w6(32'hbb7531cf),
	.w7(32'h3a0b7f63),
	.w8(32'hbc70b039),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba022d3),
	.w1(32'hba70327d),
	.w2(32'h396fcd9c),
	.w3(32'hbc0491f7),
	.w4(32'hbaac8c0b),
	.w5(32'hbbced87f),
	.w6(32'hbbc63335),
	.w7(32'h3b20084f),
	.w8(32'h3c0337ad),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85cb46),
	.w1(32'h3ab2e2fe),
	.w2(32'hbbe1c4d0),
	.w3(32'h3baa2806),
	.w4(32'hbab678d6),
	.w5(32'hbad82d61),
	.w6(32'h3a1aa4e7),
	.w7(32'h3b1ab3ab),
	.w8(32'h3a140d59),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa109),
	.w1(32'h3a974ebd),
	.w2(32'hbb7767bf),
	.w3(32'h3b0b8947),
	.w4(32'hbb920dd1),
	.w5(32'hbbec9de2),
	.w6(32'h3aae0a99),
	.w7(32'hba575a2b),
	.w8(32'h3bce2a1d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99ad0b),
	.w1(32'h3ae1d35c),
	.w2(32'h3b369b97),
	.w3(32'hbb16689a),
	.w4(32'hbb9e72c3),
	.w5(32'hbbcb995c),
	.w6(32'h3b0bc9ec),
	.w7(32'hbc042bc2),
	.w8(32'hbb336be8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc67212),
	.w1(32'hbac89cf0),
	.w2(32'hbb36d7bd),
	.w3(32'hbbb69f6a),
	.w4(32'h3a81fc07),
	.w5(32'h3bb20af4),
	.w6(32'hbc088297),
	.w7(32'hbb68eb30),
	.w8(32'hbb5f97c1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7ae5f),
	.w1(32'h3ba90be7),
	.w2(32'h3b85ffbd),
	.w3(32'h3b2751e9),
	.w4(32'h3ba6cce0),
	.w5(32'hbadf6bb5),
	.w6(32'hbb15f24f),
	.w7(32'hbb1f327f),
	.w8(32'hbb4973d9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6c7d9),
	.w1(32'hbbb290b5),
	.w2(32'hbbcdc9f9),
	.w3(32'h3ab0c436),
	.w4(32'hbb2dd9ca),
	.w5(32'hbb8ae8c8),
	.w6(32'h3afe85cf),
	.w7(32'h3a3d0b31),
	.w8(32'hbaf01e89),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3c4d7),
	.w1(32'hb95ab972),
	.w2(32'h3ab8d2a4),
	.w3(32'hbb826dfb),
	.w4(32'hbb243345),
	.w5(32'hbbdd5d62),
	.w6(32'hbb2be2d8),
	.w7(32'hbb11438a),
	.w8(32'hbbb29e56),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7560),
	.w1(32'h3aa9725c),
	.w2(32'hba08e7a3),
	.w3(32'h3acc5e79),
	.w4(32'h3bc3f318),
	.w5(32'h3a3eddef),
	.w6(32'hbb17108f),
	.w7(32'h3bc33ec8),
	.w8(32'h3b26f8bf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b944),
	.w1(32'h3b837d8d),
	.w2(32'h39300886),
	.w3(32'h3b7b909d),
	.w4(32'h3b852f33),
	.w5(32'h3c87c544),
	.w6(32'h3bc5a06b),
	.w7(32'h3b43e5e8),
	.w8(32'h3bc6b4d6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad250cf),
	.w1(32'h3b118543),
	.w2(32'h3c3da3aa),
	.w3(32'hbb0a1293),
	.w4(32'h3b351e08),
	.w5(32'hbb049441),
	.w6(32'h3c2ddf25),
	.w7(32'h3ae45a30),
	.w8(32'h3bac9cc9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4c989),
	.w1(32'hbb0d51f4),
	.w2(32'hbbe63f11),
	.w3(32'hbaebf54f),
	.w4(32'h3aea3842),
	.w5(32'hbab9425f),
	.w6(32'h3bcfd7da),
	.w7(32'h3ae8442e),
	.w8(32'h3c303f38),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab46ab4),
	.w1(32'h3b798c5e),
	.w2(32'h3bc8f90c),
	.w3(32'hbba5441d),
	.w4(32'h3b1772ce),
	.w5(32'hbb01c3dd),
	.w6(32'hbae6f7a7),
	.w7(32'hbbe05cd4),
	.w8(32'h3bb3fb97),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2ecae),
	.w1(32'h3aab3386),
	.w2(32'h3a8bd104),
	.w3(32'hbbdecd2f),
	.w4(32'h3b3d41c4),
	.w5(32'hbba55437),
	.w6(32'h3836ea52),
	.w7(32'h3be0d24b),
	.w8(32'h3bde9bce),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ec94b),
	.w1(32'hbb87d828),
	.w2(32'h3ae0130e),
	.w3(32'h3b345fcb),
	.w4(32'hba86f1ef),
	.w5(32'hba9ac211),
	.w6(32'h3adb05cc),
	.w7(32'h3a6483b4),
	.w8(32'hbb6fb8bd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe8f40),
	.w1(32'h3a75d841),
	.w2(32'hbafd1dc2),
	.w3(32'hbb9ce89e),
	.w4(32'h3b5776a1),
	.w5(32'h39880a03),
	.w6(32'hbabfd565),
	.w7(32'h3b7a9210),
	.w8(32'h3c06424a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da2a8),
	.w1(32'h3b9fb8e2),
	.w2(32'h3c2d7794),
	.w3(32'hb9e62a9b),
	.w4(32'h3bb5d4de),
	.w5(32'h3abf1898),
	.w6(32'h3b19db06),
	.w7(32'h3bb41944),
	.w8(32'h3c2061b7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd95169),
	.w1(32'hbbad7fae),
	.w2(32'hba0e94d1),
	.w3(32'h3bf96e40),
	.w4(32'h3b4a09ec),
	.w5(32'h392f5348),
	.w6(32'h3c0fca4c),
	.w7(32'hba2b8ff9),
	.w8(32'hba273bcb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2db0c3),
	.w1(32'hbb13fc64),
	.w2(32'hbbd0e217),
	.w3(32'h3c229947),
	.w4(32'h3c13b4f1),
	.w5(32'h3badeb5d),
	.w6(32'hbba6c725),
	.w7(32'hba986300),
	.w8(32'hb95d6e3e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fdbb4),
	.w1(32'h3c772950),
	.w2(32'h3bb55f10),
	.w3(32'h3b1ec391),
	.w4(32'h3a896e82),
	.w5(32'h3b8395b7),
	.w6(32'hbbb237e8),
	.w7(32'hbbc57c87),
	.w8(32'h3b53595f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1ee1b),
	.w1(32'hbb9abf41),
	.w2(32'hbc2f863c),
	.w3(32'hba0b3bab),
	.w4(32'hba5be6bb),
	.w5(32'hbc826605),
	.w6(32'hbc170df9),
	.w7(32'hba6aab9e),
	.w8(32'hbc459ac4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21622d),
	.w1(32'h3b7808ad),
	.w2(32'hba2a85c9),
	.w3(32'hbc55ba4d),
	.w4(32'hbad01756),
	.w5(32'hbb1bb4d9),
	.w6(32'hbc73582f),
	.w7(32'hbb8486ea),
	.w8(32'hbb9e8049),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38098057),
	.w1(32'hbae74e5f),
	.w2(32'hbb03a3e4),
	.w3(32'h39a4fc1c),
	.w4(32'h3a2d442f),
	.w5(32'h39a588de),
	.w6(32'hba9b819d),
	.w7(32'h3a2b7c26),
	.w8(32'h3a5c8612),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4bfe0),
	.w1(32'h3b21b7bf),
	.w2(32'h3a7091f2),
	.w3(32'h3b2d322f),
	.w4(32'h39a7cc02),
	.w5(32'h3a403564),
	.w6(32'h3acb3259),
	.w7(32'hbb0a3a9c),
	.w8(32'hba83dc88),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba379791),
	.w1(32'hbb7891a9),
	.w2(32'hbb8ede31),
	.w3(32'hbae66484),
	.w4(32'hbb8402ba),
	.w5(32'hbb901ec0),
	.w6(32'hbb288533),
	.w7(32'hbb20d6b3),
	.w8(32'hbb152d3e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d8b8e),
	.w1(32'h3991abba),
	.w2(32'h3a8fa80a),
	.w3(32'hbb6101fe),
	.w4(32'h3920c8a5),
	.w5(32'h3a918c27),
	.w6(32'hbb440c38),
	.w7(32'h3a3fa737),
	.w8(32'hb9234ca7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0267dd),
	.w1(32'h3aa320ca),
	.w2(32'h3aa6dfca),
	.w3(32'h3a06573a),
	.w4(32'hbabc12f6),
	.w5(32'hb9bb8b28),
	.w6(32'hba2e28f8),
	.w7(32'hba5f0d52),
	.w8(32'h3a4c0351),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa33b0a),
	.w1(32'hbb80800a),
	.w2(32'hbb9ab6c1),
	.w3(32'hbb2ba525),
	.w4(32'hb8a43f35),
	.w5(32'h3a9ac9f4),
	.w6(32'hbb46aa04),
	.w7(32'hba51ec0d),
	.w8(32'hb9bb3d3a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d080c),
	.w1(32'hbbc3dc77),
	.w2(32'hbbe3da11),
	.w3(32'hbb08efbc),
	.w4(32'hbc04f037),
	.w5(32'hbbbf6eb1),
	.w6(32'hbbb4b267),
	.w7(32'hbbed430c),
	.w8(32'hbbe78166),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d074b),
	.w1(32'h3b8086df),
	.w2(32'h3a33251b),
	.w3(32'hbb00cde4),
	.w4(32'h3b4ecfe2),
	.w5(32'h3a3aff78),
	.w6(32'hbab0efd8),
	.w7(32'h3b57f90f),
	.w8(32'hbb09abd0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c8fe0),
	.w1(32'h3b406441),
	.w2(32'h3a8f81c6),
	.w3(32'hbaa65ef2),
	.w4(32'h3b96804f),
	.w5(32'h39b692ea),
	.w6(32'hbb3df567),
	.w7(32'h3a994755),
	.w8(32'hba56acc2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a133752),
	.w1(32'hbbe981c6),
	.w2(32'hbb8850e3),
	.w3(32'h3b9f9672),
	.w4(32'hbb345ade),
	.w5(32'hbb399798),
	.w6(32'hbab43c2f),
	.w7(32'hbbb2fd93),
	.w8(32'hbbad036a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f736),
	.w1(32'h3c14238c),
	.w2(32'h3bc787ad),
	.w3(32'hbb9f1113),
	.w4(32'h3bfe89e3),
	.w5(32'h3b9628a5),
	.w6(32'hbb6618eb),
	.w7(32'h3c045a66),
	.w8(32'h3b9396f6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf1dda),
	.w1(32'h3a850712),
	.w2(32'hba4df8ae),
	.w3(32'h3bf9a3e1),
	.w4(32'h3b299a97),
	.w5(32'hba8b57dd),
	.w6(32'h3b9a8b54),
	.w7(32'h3a7df542),
	.w8(32'hbb181111),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e58677),
	.w1(32'hba22e8f3),
	.w2(32'hb9ee96bf),
	.w3(32'h3a628d53),
	.w4(32'hba98b0f1),
	.w5(32'hba69b07d),
	.w6(32'h399f1801),
	.w7(32'hb9fba22c),
	.w8(32'hb9dc306d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebf28b),
	.w1(32'hbb1e033f),
	.w2(32'hbb8db0c1),
	.w3(32'hbaed987f),
	.w4(32'hbae86235),
	.w5(32'hba4cfe51),
	.w6(32'hba4a5fbb),
	.w7(32'h39b0122e),
	.w8(32'hbaa8233e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8464c5),
	.w1(32'hbab26168),
	.w2(32'hbad345fb),
	.w3(32'h3a26a8f6),
	.w4(32'hbb078d93),
	.w5(32'hbb83aa4a),
	.w6(32'hbb047cfa),
	.w7(32'hbadf8cfd),
	.w8(32'hbb0b7b35),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ff829),
	.w1(32'hbb1ea41c),
	.w2(32'hb8fbf2cd),
	.w3(32'hba8f0cc1),
	.w4(32'hbba98bdc),
	.w5(32'hba2892c8),
	.w6(32'hbb39d2c4),
	.w7(32'hbb21c996),
	.w8(32'hb9f38854),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98bed1),
	.w1(32'hb9e9911d),
	.w2(32'h38b0e7fc),
	.w3(32'hbb9320c6),
	.w4(32'h3a69ddbd),
	.w5(32'h38dd2af4),
	.w6(32'hbb68a109),
	.w7(32'h39b8fa24),
	.w8(32'hba5ed782),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afda1ef),
	.w1(32'h3b1be6e0),
	.w2(32'h3b33902b),
	.w3(32'hba8f89d3),
	.w4(32'h3b155d39),
	.w5(32'h3b243f70),
	.w6(32'hbb2fb4fb),
	.w7(32'h3b0210c3),
	.w8(32'hba819240),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56968f),
	.w1(32'h3a6fe16d),
	.w2(32'hb89032dc),
	.w3(32'h37ba265e),
	.w4(32'hbb29f93b),
	.w5(32'hbacee28f),
	.w6(32'hb8772d54),
	.w7(32'hbae67e55),
	.w8(32'hbb5858ae),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6e37d),
	.w1(32'hbbaea401),
	.w2(32'hbb81f351),
	.w3(32'hbb5b9dbe),
	.w4(32'hbb787383),
	.w5(32'hbb8a213e),
	.w6(32'hbbdb5644),
	.w7(32'hbb9d8a2a),
	.w8(32'hbb6ae2fe),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa648dc),
	.w1(32'hba233a8d),
	.w2(32'hbb41f792),
	.w3(32'hba271cc4),
	.w4(32'hbb783212),
	.w5(32'hbb759bea),
	.w6(32'hbae5232e),
	.w7(32'hba16824f),
	.w8(32'hbb5da355),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b1ac8),
	.w1(32'hbc3de17e),
	.w2(32'hbbc2c848),
	.w3(32'h3b0c83ef),
	.w4(32'h3b298eb1),
	.w5(32'h3ad7c87d),
	.w6(32'hbb92348e),
	.w7(32'hbbb6a854),
	.w8(32'hbb04f316),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a793c72),
	.w1(32'h3b05d3a4),
	.w2(32'h3ab6672f),
	.w3(32'h39977ffe),
	.w4(32'hbaed9574),
	.w5(32'hbae707e3),
	.w6(32'hbb187bed),
	.w7(32'hbbaf2b55),
	.w8(32'hbb693a58),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb383d8),
	.w1(32'h3aaa9469),
	.w2(32'h3ad9fde8),
	.w3(32'hbb3ff311),
	.w4(32'h3ba32cee),
	.w5(32'h3b58cc54),
	.w6(32'hbbd97c23),
	.w7(32'hbaa6f3f5),
	.w8(32'h3a1b5e2e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4cba8),
	.w1(32'hbbe8f824),
	.w2(32'hbbbfa717),
	.w3(32'h38cb9f92),
	.w4(32'hbb47c54d),
	.w5(32'hbb294cba),
	.w6(32'hb97398f3),
	.w7(32'hbbc3255d),
	.w8(32'hbc012a7c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4c1b5),
	.w1(32'h3b21b1ae),
	.w2(32'hba465a48),
	.w3(32'hbbb9cda3),
	.w4(32'hbb3a37bb),
	.w5(32'hbb5cbd7e),
	.w6(32'hbbc38f94),
	.w7(32'hbb9d92b3),
	.w8(32'hbaec382f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1acc),
	.w1(32'h3a9b51a5),
	.w2(32'h39fa6f30),
	.w3(32'hba98177a),
	.w4(32'h3ae9d704),
	.w5(32'hbab34ed0),
	.w6(32'hbb1e19ac),
	.w7(32'h3aa38d14),
	.w8(32'hbb2f33ea),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aced4),
	.w1(32'hbb06e40a),
	.w2(32'hbaf29680),
	.w3(32'hba3f66c5),
	.w4(32'h3a123513),
	.w5(32'hbabd857a),
	.w6(32'hbbbff819),
	.w7(32'hbb86d0b4),
	.w8(32'hbafc61fd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe3a9),
	.w1(32'hbbca3df7),
	.w2(32'hbbacfbf6),
	.w3(32'hba8808f1),
	.w4(32'h39f7cf1c),
	.w5(32'hbafc90b0),
	.w6(32'hbbd37eba),
	.w7(32'hba938c85),
	.w8(32'hbb90bbae),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc417bec),
	.w1(32'hbc542c5f),
	.w2(32'hbac9ed84),
	.w3(32'hbc4a5b06),
	.w4(32'hbace5820),
	.w5(32'hbb495a53),
	.w6(32'hbc0acece),
	.w7(32'hbc0f3454),
	.w8(32'hbb071c0e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc423c53),
	.w1(32'hbb4c5015),
	.w2(32'h39910c77),
	.w3(32'hbc0b4de3),
	.w4(32'h3b065392),
	.w5(32'h3bedab9c),
	.w6(32'hbc3fed89),
	.w7(32'h38325fae),
	.w8(32'h3a6f8a2b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aef551),
	.w1(32'h3bb08008),
	.w2(32'h3addddb2),
	.w3(32'hb9ec50ae),
	.w4(32'h3b63eb6b),
	.w5(32'h36d5b801),
	.w6(32'hbb1fc128),
	.w7(32'h3ab25647),
	.w8(32'hbb108c5c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7d880),
	.w1(32'hbc0b806c),
	.w2(32'hbbd00f9d),
	.w3(32'hbb0829cf),
	.w4(32'h3adba41e),
	.w5(32'h3b9fb914),
	.w6(32'hbbc56d7b),
	.w7(32'hbb2fb80a),
	.w8(32'hbb839bae),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9a8b0),
	.w1(32'hba2456a9),
	.w2(32'hb8ff2752),
	.w3(32'h3a39ce0f),
	.w4(32'hbac047a0),
	.w5(32'hbb4906be),
	.w6(32'h39d7186d),
	.w7(32'hb955de8f),
	.w8(32'hbb01c5dd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26f489),
	.w1(32'hbbef9e3a),
	.w2(32'hbb5b7ca3),
	.w3(32'hbb8d53dd),
	.w4(32'hbac820dc),
	.w5(32'hbb39435e),
	.w6(32'hbc2b6f27),
	.w7(32'hbb791f9b),
	.w8(32'hbb688575),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e45ce),
	.w1(32'h3aaf59a6),
	.w2(32'h3add8a11),
	.w3(32'hba994b78),
	.w4(32'hb990fdc2),
	.w5(32'h3ab8b491),
	.w6(32'h3aa739fd),
	.w7(32'hba02c9e5),
	.w8(32'hb9d649e5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a319c9b),
	.w1(32'hbac4eb6b),
	.w2(32'hb9b8d23e),
	.w3(32'h3a0b1f4f),
	.w4(32'h3a5a3243),
	.w5(32'h386db425),
	.w6(32'hb9378759),
	.w7(32'h3ac68122),
	.w8(32'h3a126c7a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcee43),
	.w1(32'hb8fe4fcf),
	.w2(32'hbb5933e2),
	.w3(32'hba98e75c),
	.w4(32'hbb68f77d),
	.w5(32'hbbc283ef),
	.w6(32'hb8b1ee9c),
	.w7(32'hbb809436),
	.w8(32'hbb7a2b31),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9288b),
	.w1(32'h3b8541a2),
	.w2(32'hb8970938),
	.w3(32'h3a866f2d),
	.w4(32'h3bcf11dd),
	.w5(32'h3aa73930),
	.w6(32'hbb652fd2),
	.w7(32'h3baf474c),
	.w8(32'hba7b4beb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9794),
	.w1(32'hbad56a7f),
	.w2(32'hbb9c6e47),
	.w3(32'hb9f7dc49),
	.w4(32'hba9654f3),
	.w5(32'hbb1def5f),
	.w6(32'hb9aed83e),
	.w7(32'hbb17d377),
	.w8(32'hbb3bd8b2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb845d4),
	.w1(32'h3a924e7b),
	.w2(32'h3afd1b38),
	.w3(32'hbbb13aee),
	.w4(32'h3b033ef8),
	.w5(32'h3b6a6016),
	.w6(32'hbb9e0109),
	.w7(32'hbaa1bd7f),
	.w8(32'hbac16d0f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a5e6a),
	.w1(32'hbb60d9a8),
	.w2(32'hbb5d8dee),
	.w3(32'h3a98d94c),
	.w4(32'hbad78353),
	.w5(32'hbb1caa48),
	.w6(32'hba84aa7e),
	.w7(32'hbb0d720c),
	.w8(32'hbb70a440),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa84f03),
	.w1(32'h3b9b36f8),
	.w2(32'h3bd911aa),
	.w3(32'hbb833506),
	.w4(32'hb857764c),
	.w5(32'h3ab92d0a),
	.w6(32'hbc09cc03),
	.w7(32'hba692da6),
	.w8(32'h3ad5b5cb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88854ef),
	.w1(32'hbbb70a1b),
	.w2(32'hbb85acde),
	.w3(32'h3b2f9ed3),
	.w4(32'h3b8f3b71),
	.w5(32'hbaf17747),
	.w6(32'h3b36a16f),
	.w7(32'h3aaefff3),
	.w8(32'h39f5456c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947586),
	.w1(32'h3b022532),
	.w2(32'hb9b1983c),
	.w3(32'hbb8c0379),
	.w4(32'h3a8e400b),
	.w5(32'hba9aca7f),
	.w6(32'hbbb90d04),
	.w7(32'hb9d0a953),
	.w8(32'hbb4a3954),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b8680),
	.w1(32'h3abb82b3),
	.w2(32'hbb178390),
	.w3(32'hba80527f),
	.w4(32'h397e6f2a),
	.w5(32'hbb58a64d),
	.w6(32'hba79e960),
	.w7(32'hba1a34cd),
	.w8(32'hbaf2688e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3be887),
	.w1(32'hb834ee81),
	.w2(32'hb9d8effc),
	.w3(32'h39d866c6),
	.w4(32'h3ab2eea5),
	.w5(32'h3aaa3b7d),
	.w6(32'h3a13c132),
	.w7(32'hba0d3d6b),
	.w8(32'h39c40252),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6fc76),
	.w1(32'hbae0cd35),
	.w2(32'hb9e5737d),
	.w3(32'h3a865436),
	.w4(32'hbb6a423a),
	.w5(32'hbb3062d4),
	.w6(32'h3b07b884),
	.w7(32'hbb50af87),
	.w8(32'hbac6fe6d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34019e),
	.w1(32'h3b461e89),
	.w2(32'h3b13a387),
	.w3(32'hbba844de),
	.w4(32'hb886c035),
	.w5(32'h3a1515fa),
	.w6(32'hbb7795c3),
	.w7(32'h3930e896),
	.w8(32'hba2ff1eb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a848946),
	.w1(32'h3b93f92e),
	.w2(32'hb8d1b875),
	.w3(32'hbb00365b),
	.w4(32'h3b1728ed),
	.w5(32'hba51e5bb),
	.w6(32'hbaba0fdf),
	.w7(32'h39c71138),
	.w8(32'hba5d2fbf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cca52),
	.w1(32'hbac64f4f),
	.w2(32'hbaf9705a),
	.w3(32'hbb0195ee),
	.w4(32'hba49aec1),
	.w5(32'hbb03972b),
	.w6(32'h3ac67c51),
	.w7(32'hbac8559c),
	.w8(32'hbb08e674),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8309d0),
	.w1(32'hba9faa7b),
	.w2(32'hbb30157f),
	.w3(32'h3a4eea42),
	.w4(32'hba736398),
	.w5(32'hbaf3cf82),
	.w6(32'hbaf190fc),
	.w7(32'h3ab6903e),
	.w8(32'h3a142260),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782b94),
	.w1(32'h3aea7f56),
	.w2(32'h3ac1f728),
	.w3(32'hb99b7449),
	.w4(32'h3b316f56),
	.w5(32'h3a859fa0),
	.w6(32'hb9b63591),
	.w7(32'h3ae5954e),
	.w8(32'hbb63fee4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a387343),
	.w1(32'h3a49847e),
	.w2(32'h3b51ef2e),
	.w3(32'h3a0e183f),
	.w4(32'h3adea788),
	.w5(32'h3b524dae),
	.w6(32'h3ab7721a),
	.w7(32'hb97c67cc),
	.w8(32'h3b0b4dc2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fd6e9),
	.w1(32'hba6ce8e7),
	.w2(32'hba78c2fe),
	.w3(32'h3b28040f),
	.w4(32'hbac2ff10),
	.w5(32'hb883318a),
	.w6(32'h3abcd118),
	.w7(32'hb9a1fa49),
	.w8(32'h39cb69e1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a48340),
	.w1(32'hbb2f03ff),
	.w2(32'hb9dc12e0),
	.w3(32'hba1edd0b),
	.w4(32'hbaad48b8),
	.w5(32'hba63083a),
	.w6(32'hba5c7509),
	.w7(32'hbb123a9f),
	.w8(32'hbaadbdf7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849937),
	.w1(32'hbbd9afe1),
	.w2(32'hbaeeb329),
	.w3(32'hbb475f7f),
	.w4(32'hbbb0ea6d),
	.w5(32'h3976d92f),
	.w6(32'hbba5252e),
	.w7(32'hbbd3718b),
	.w8(32'hbbb425f5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80e04e),
	.w1(32'hb9f7c59d),
	.w2(32'h3bc3c1a4),
	.w3(32'h3a783a15),
	.w4(32'hbac046b3),
	.w5(32'hbb21a2d9),
	.w6(32'hbbf2ba5a),
	.w7(32'hbbad6caa),
	.w8(32'hbb4c06da),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb076398),
	.w1(32'h3b01feef),
	.w2(32'h39abc810),
	.w3(32'h3a7277d1),
	.w4(32'h3b23dd77),
	.w5(32'h3a645c1e),
	.w6(32'hbae498d5),
	.w7(32'h3ac92e4b),
	.w8(32'hba4d17b9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba251dd4),
	.w1(32'hbb294017),
	.w2(32'hb9fdceb6),
	.w3(32'hb946bd3f),
	.w4(32'hbad06ce7),
	.w5(32'hba146912),
	.w6(32'hba076aed),
	.w7(32'hbb64c272),
	.w8(32'hbac91873),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a233),
	.w1(32'hbb6f4c60),
	.w2(32'hbbebe846),
	.w3(32'hbbb82943),
	.w4(32'hbba4b80b),
	.w5(32'hbbc6a0b2),
	.w6(32'hbbd89439),
	.w7(32'h39476e99),
	.w8(32'hbb8bc103),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb243896),
	.w1(32'h3a260ae2),
	.w2(32'hba361ff4),
	.w3(32'hbb99790d),
	.w4(32'h3a109514),
	.w5(32'hbb986aa6),
	.w6(32'hbb35fff0),
	.w7(32'hbad95313),
	.w8(32'hbab60f41),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd10c29),
	.w1(32'hbab6006c),
	.w2(32'hbadfc495),
	.w3(32'hbb5afeaa),
	.w4(32'h397b66ac),
	.w5(32'hb96dca23),
	.w6(32'hbb8ad756),
	.w7(32'h380e63c7),
	.w8(32'hba8ae2a0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4872),
	.w1(32'hbb1efd86),
	.w2(32'hbb9d317b),
	.w3(32'hba820d3e),
	.w4(32'h3a8475c0),
	.w5(32'h39acedb6),
	.w6(32'hbb42abc0),
	.w7(32'h3a6d3c0d),
	.w8(32'hbb12e553),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf6aa5),
	.w1(32'h3ac6e307),
	.w2(32'h3aaf4494),
	.w3(32'hbacdc305),
	.w4(32'h3bc57456),
	.w5(32'h3b7d9d17),
	.w6(32'hbba65a7b),
	.w7(32'hb8ee02bc),
	.w8(32'hba567264),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f972b),
	.w1(32'h3b878001),
	.w2(32'h39dc4572),
	.w3(32'h3a835c3b),
	.w4(32'h3b24c66b),
	.w5(32'hbb2088dd),
	.w6(32'hba3359e7),
	.w7(32'h3b2e7b25),
	.w8(32'h3974bdba),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c83b6),
	.w1(32'hba817274),
	.w2(32'h38d679e4),
	.w3(32'hba8521fd),
	.w4(32'h3b156e0a),
	.w5(32'h3a2ce8c1),
	.w6(32'hba892c91),
	.w7(32'hba00031a),
	.w8(32'hbab9b3cc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af77b),
	.w1(32'hbb4bdcf6),
	.w2(32'hbb6427f1),
	.w3(32'hb9560c2e),
	.w4(32'h3af21d1f),
	.w5(32'h3a20f79b),
	.w6(32'hbbc5dd61),
	.w7(32'h39e2eb69),
	.w8(32'hbb2c3463),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b91f8),
	.w1(32'h3b3427ae),
	.w2(32'h3b86160b),
	.w3(32'hbadbc100),
	.w4(32'hb7e469f5),
	.w5(32'h3903ef86),
	.w6(32'hbb60136c),
	.w7(32'hbb4dc9de),
	.w8(32'hbb09836c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d41ec),
	.w1(32'hba8d4bcf),
	.w2(32'hbac7f93f),
	.w3(32'h3a16123a),
	.w4(32'h3b22a7dc),
	.w5(32'h39fb3af7),
	.w6(32'hbb820d77),
	.w7(32'hbac0589b),
	.w8(32'hbb6eed4f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5ed9c),
	.w1(32'h3a74c30f),
	.w2(32'h3a3ae9a0),
	.w3(32'h3a29643c),
	.w4(32'h3b1bedaa),
	.w5(32'h3a9fbe31),
	.w6(32'h39b723e2),
	.w7(32'h3a930c06),
	.w8(32'h3b12217f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dfe0d),
	.w1(32'h3b90f4c2),
	.w2(32'h3b9bed7f),
	.w3(32'hbb3aa256),
	.w4(32'hbb1b6708),
	.w5(32'h3a7524c5),
	.w6(32'hbb4f389a),
	.w7(32'hbac54e45),
	.w8(32'hbb6b1c68),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24b67c),
	.w1(32'hbaab34f6),
	.w2(32'hbb1155ef),
	.w3(32'hbb2c1f92),
	.w4(32'hb98994b1),
	.w5(32'hbb120a54),
	.w6(32'hbb91c989),
	.w7(32'hbb33ef41),
	.w8(32'hbb305561),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39867192),
	.w1(32'h3925d11b),
	.w2(32'hba32c665),
	.w3(32'hbab50817),
	.w4(32'h3a22eb65),
	.w5(32'hb8c97344),
	.w6(32'hbad4c281),
	.w7(32'h3a9eb571),
	.w8(32'h3a850eac),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b5ca),
	.w1(32'hbb2c97ec),
	.w2(32'hba836f69),
	.w3(32'h3b155762),
	.w4(32'hbad03bec),
	.w5(32'hba58750b),
	.w6(32'h3b120b89),
	.w7(32'hbb3cce7e),
	.w8(32'hbb0d8b99),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacacd7c),
	.w1(32'h3a2eed37),
	.w2(32'h3a270900),
	.w3(32'hba8416ee),
	.w4(32'h3a8b7f21),
	.w5(32'h3a776b8f),
	.w6(32'hbb5248b0),
	.w7(32'h3a06523c),
	.w8(32'h39035400),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba4e7),
	.w1(32'h3ac1db49),
	.w2(32'h3ab769a3),
	.w3(32'hb9e79b2d),
	.w4(32'h3b2c222c),
	.w5(32'hbaba547c),
	.w6(32'hbb0b3d20),
	.w7(32'h392a3cdf),
	.w8(32'hbb71f6ee),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad3c87),
	.w1(32'hbb43fb3f),
	.w2(32'hbb7447bd),
	.w3(32'h39917f1e),
	.w4(32'h3a1908e6),
	.w5(32'hbb7510a8),
	.w6(32'hbb2d30cd),
	.w7(32'hbb486024),
	.w8(32'hbc0fecda),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca6907),
	.w1(32'h3a1f9a6a),
	.w2(32'h3ab49833),
	.w3(32'h3a9e6a21),
	.w4(32'h3b063a25),
	.w5(32'h3b484ace),
	.w6(32'hbb625ac2),
	.w7(32'h3b0e7caa),
	.w8(32'h3a57ea45),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5d0f),
	.w1(32'hbb33e5c0),
	.w2(32'hbab8058f),
	.w3(32'h3b4282e0),
	.w4(32'h3a2eb513),
	.w5(32'hb83384dc),
	.w6(32'hbaa5d2b8),
	.w7(32'hbb5fa6e8),
	.w8(32'hbaa5bb95),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2b278),
	.w1(32'hb9b33923),
	.w2(32'hbabfebd4),
	.w3(32'h3aaaa248),
	.w4(32'hba3e3d8c),
	.w5(32'h3b035517),
	.w6(32'hba1d15eb),
	.w7(32'h3ac0b4c3),
	.w8(32'hb8a51ea6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9c93),
	.w1(32'hbc06d7e3),
	.w2(32'hbc1ac10e),
	.w3(32'h3aff0649),
	.w4(32'h3961892e),
	.w5(32'hba7e5342),
	.w6(32'hbb5e0ca1),
	.w7(32'hbb5db8bf),
	.w8(32'hbbe3323d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71dd22),
	.w1(32'h3aac4da0),
	.w2(32'hbbaa251b),
	.w3(32'hbb52389b),
	.w4(32'h3a961606),
	.w5(32'hba60f43a),
	.w6(32'hbbf4c96d),
	.w7(32'hbac7f2e1),
	.w8(32'hbc05bad0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab83586),
	.w1(32'hbb2246a9),
	.w2(32'hbb2e5984),
	.w3(32'h39c87f18),
	.w4(32'hbb8b763f),
	.w5(32'hbb368a41),
	.w6(32'hbae36d6f),
	.w7(32'hbaaa40aa),
	.w8(32'hbb4e6612),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cf376),
	.w1(32'h3a8d3f72),
	.w2(32'h3aab9a94),
	.w3(32'h3a5e3d61),
	.w4(32'h3a8b776f),
	.w5(32'h3b451502),
	.w6(32'h39c76960),
	.w7(32'h3a87ec81),
	.w8(32'h3b7b7aa0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d6985),
	.w1(32'h3b7e4551),
	.w2(32'h3b04ed8c),
	.w3(32'h3b53e938),
	.w4(32'h3b10764b),
	.w5(32'h3aa59181),
	.w6(32'h3a83c379),
	.w7(32'h3ab041d0),
	.w8(32'hb93a210d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb583d9f),
	.w1(32'hbaff2a1b),
	.w2(32'hbb273e12),
	.w3(32'hba363a54),
	.w4(32'hb9fa715f),
	.w5(32'h3b537118),
	.w6(32'hbb113bcf),
	.w7(32'hba1e2296),
	.w8(32'hbaed46d0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad90471),
	.w1(32'hb6cc2a73),
	.w2(32'h3a8e2c2b),
	.w3(32'hbb5da4e7),
	.w4(32'h38df963d),
	.w5(32'h3a896dd8),
	.w6(32'hbbab7d15),
	.w7(32'h389d9109),
	.w8(32'hbac45c5e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7bc1b),
	.w1(32'hbb137b98),
	.w2(32'hba288e29),
	.w3(32'h3a4ad30e),
	.w4(32'hbb540494),
	.w5(32'h3a3d0140),
	.w6(32'hba75e2a6),
	.w7(32'hbb219c61),
	.w8(32'hbad02840),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac97f9e),
	.w1(32'h3aeec276),
	.w2(32'hba7a6a92),
	.w3(32'hb931ea78),
	.w4(32'h3b2e8f43),
	.w5(32'hba85f00a),
	.w6(32'hba0c6fb4),
	.w7(32'h3ad95ce4),
	.w8(32'h3a31b73a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64e656),
	.w1(32'h3a5f94ce),
	.w2(32'hb9d11806),
	.w3(32'hba0f9403),
	.w4(32'h3bb47a7f),
	.w5(32'h3c00a0e7),
	.w6(32'hbb2af419),
	.w7(32'h3b859496),
	.w8(32'h3b5417ac),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dc3e2),
	.w1(32'h3a17f0e0),
	.w2(32'h39c52ac4),
	.w3(32'h3b2caa6c),
	.w4(32'h3a09bf00),
	.w5(32'h3a963330),
	.w6(32'h3a936b6d),
	.w7(32'h3ab2c8fb),
	.w8(32'hbab28eb1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd5f26),
	.w1(32'h3b2d339d),
	.w2(32'h3b21226c),
	.w3(32'hba669535),
	.w4(32'h386d6196),
	.w5(32'hbb2c8f08),
	.w6(32'hbb38f806),
	.w7(32'hb82013fb),
	.w8(32'hbb384981),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79e2e5),
	.w1(32'h3a9e0ad2),
	.w2(32'h39bff16b),
	.w3(32'hbaa4e35e),
	.w4(32'h3ad1d1ba),
	.w5(32'hba866081),
	.w6(32'hbaa828e3),
	.w7(32'h3a5d5656),
	.w8(32'h38a7fe4b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb909c),
	.w1(32'h3b3c7c8a),
	.w2(32'h3b3e7e4e),
	.w3(32'hb7570188),
	.w4(32'h3a3a23aa),
	.w5(32'h3a75d388),
	.w6(32'hbb4a348f),
	.w7(32'hbb92196c),
	.w8(32'hbaa945fb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab37a6a),
	.w1(32'h3b1aca50),
	.w2(32'h39d2234f),
	.w3(32'h3b119073),
	.w4(32'h3af33e1e),
	.w5(32'hb9a61b84),
	.w6(32'h3acd67c9),
	.w7(32'h3b0f76eb),
	.w8(32'h3b2617b1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc4e1),
	.w1(32'h3a3e13cc),
	.w2(32'hbb22578f),
	.w3(32'hba6892e6),
	.w4(32'hbb006baf),
	.w5(32'hbb4f4c5a),
	.w6(32'h3a6788de),
	.w7(32'hbaebf407),
	.w8(32'hba9dcba7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbbcef),
	.w1(32'h3baa14b3),
	.w2(32'h3a233d1d),
	.w3(32'hbab30ea7),
	.w4(32'h3b58dba0),
	.w5(32'hba22c686),
	.w6(32'hbb600e86),
	.w7(32'h3ad8008a),
	.w8(32'h392c7e8d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d0f41),
	.w1(32'h3b209f52),
	.w2(32'hb9b9c2e8),
	.w3(32'hbac06fc1),
	.w4(32'hbaddf660),
	.w5(32'hbb370ade),
	.w6(32'hbbc2f623),
	.w7(32'hbbc7556d),
	.w8(32'hbbd433b4),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba195d1),
	.w1(32'hb965565a),
	.w2(32'h3a4609b6),
	.w3(32'hbb1c5e1e),
	.w4(32'h399b4922),
	.w5(32'hba19e9c8),
	.w6(32'h3a888f1f),
	.w7(32'hba8d2ceb),
	.w8(32'hb91943b2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba312857),
	.w1(32'h3b157c62),
	.w2(32'hba3aa84d),
	.w3(32'hba98d3aa),
	.w4(32'h3b33e7dc),
	.w5(32'hbb871459),
	.w6(32'hbab3c0ef),
	.w7(32'h39a1771a),
	.w8(32'hb9b0f5c1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395980d0),
	.w1(32'h3b790eed),
	.w2(32'h3a4c48a8),
	.w3(32'h3aab49f2),
	.w4(32'h3b3f22d9),
	.w5(32'hb933336a),
	.w6(32'hba9c7857),
	.w7(32'h388530ec),
	.w8(32'hbaa8703c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09aa49),
	.w1(32'hbb96784c),
	.w2(32'hbbc7f52f),
	.w3(32'hbb91ab3e),
	.w4(32'hbaa65148),
	.w5(32'hbb35a8a6),
	.w6(32'hbbcefa74),
	.w7(32'hbb890b81),
	.w8(32'hbb873e15),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbaf7e),
	.w1(32'hbb936bc9),
	.w2(32'hbbb0f9fd),
	.w3(32'hbab7b232),
	.w4(32'hbacacc8a),
	.w5(32'hbad1cc35),
	.w6(32'hbb943859),
	.w7(32'hbb10ba90),
	.w8(32'hbb8113a6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cf7da),
	.w1(32'hba74d96e),
	.w2(32'h3a43a20c),
	.w3(32'hb9a3b48d),
	.w4(32'hba0ec796),
	.w5(32'hb9360857),
	.w6(32'hbb7f3fc4),
	.w7(32'hbb06da54),
	.w8(32'hbb4aac5c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba873bc5),
	.w1(32'hb9a24833),
	.w2(32'hbb38d4b2),
	.w3(32'hb80ff457),
	.w4(32'hba9726ea),
	.w5(32'hbb26cf39),
	.w6(32'h3a3726df),
	.w7(32'h3913d67d),
	.w8(32'hba8a5c81),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47ece7),
	.w1(32'h3adea64e),
	.w2(32'h3ad58fa5),
	.w3(32'hbad800c7),
	.w4(32'h3b8ebe7e),
	.w5(32'h3b755e1e),
	.w6(32'hbb34d22c),
	.w7(32'h3a3b7f8a),
	.w8(32'h38ccc337),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd9cf9),
	.w1(32'h3b312826),
	.w2(32'h3ab69485),
	.w3(32'h3b84282e),
	.w4(32'h3b66f508),
	.w5(32'h3af4348b),
	.w6(32'h3aceefb8),
	.w7(32'h3aba29e1),
	.w8(32'h3ae8bf84),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937ceaf),
	.w1(32'hba94945a),
	.w2(32'hba7c74e3),
	.w3(32'h3a51c2a9),
	.w4(32'hba8b18c8),
	.w5(32'h3a3c51dd),
	.w6(32'h3b7cfc26),
	.w7(32'hba1bac4f),
	.w8(32'hbb382e85),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3ab7c),
	.w1(32'hbbbf5ea8),
	.w2(32'hbb725896),
	.w3(32'hbb59f136),
	.w4(32'hbb9da63c),
	.w5(32'hbbb39e22),
	.w6(32'hbb090297),
	.w7(32'hbbbc1015),
	.w8(32'hbb06c9ed),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7f22),
	.w1(32'hba542036),
	.w2(32'hbb0a991c),
	.w3(32'hbb76c225),
	.w4(32'h3ae8e264),
	.w5(32'h3b045451),
	.w6(32'hbb99c107),
	.w7(32'hba397d5a),
	.w8(32'hbaf6b3b5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab97ee),
	.w1(32'hba98f274),
	.w2(32'hba7e6445),
	.w3(32'h3aac62c3),
	.w4(32'h3aba9e88),
	.w5(32'hba8773c3),
	.w6(32'h39b4a0aa),
	.w7(32'h3b508721),
	.w8(32'h3a89b4c5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62b92e),
	.w1(32'h3a8ae743),
	.w2(32'hba4a0f1e),
	.w3(32'hba632f5c),
	.w4(32'hba1d5f2d),
	.w5(32'hbb62f48e),
	.w6(32'h393a6ea1),
	.w7(32'hb66d2547),
	.w8(32'hba83e3ec),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e12d9),
	.w1(32'h3b1543cb),
	.w2(32'h3767bd40),
	.w3(32'h3a826bf8),
	.w4(32'h396ae4c0),
	.w5(32'hbb1eaf67),
	.w6(32'h39cc5021),
	.w7(32'h3ab14801),
	.w8(32'h39c42f2a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834649),
	.w1(32'h396c9ac9),
	.w2(32'h3b8003bc),
	.w3(32'hbb04b3f0),
	.w4(32'h3b079986),
	.w5(32'h3ae7bfde),
	.w6(32'hbb6b7836),
	.w7(32'h3a63eb09),
	.w8(32'hb9da9989),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029b6b),
	.w1(32'hbbcd2f56),
	.w2(32'hbb006e53),
	.w3(32'hba057672),
	.w4(32'hba94e778),
	.w5(32'h3b38eafb),
	.w6(32'hbb1f6ab7),
	.w7(32'hbb7b1401),
	.w8(32'h3b193214),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e50e7),
	.w1(32'hbb5ea451),
	.w2(32'hbb47f42b),
	.w3(32'hba4e0851),
	.w4(32'hbb016368),
	.w5(32'hbbac79fb),
	.w6(32'hba311308),
	.w7(32'hbb58cb47),
	.w8(32'hbae9fd2c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb562d2f),
	.w1(32'h3b13c788),
	.w2(32'hbb8bed01),
	.w3(32'h3a365b3d),
	.w4(32'h3a0a090c),
	.w5(32'hbc031072),
	.w6(32'hbba8ea28),
	.w7(32'hbae04771),
	.w8(32'hbc161ea3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc381c5),
	.w1(32'hbba465f1),
	.w2(32'hbbad5c23),
	.w3(32'hbac15cf0),
	.w4(32'h3aaa603a),
	.w5(32'h3b6fccf5),
	.w6(32'hbbfca382),
	.w7(32'hba30b733),
	.w8(32'hbb83bbda),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10b34f),
	.w1(32'hba91416c),
	.w2(32'hbb1266e6),
	.w3(32'hba560d38),
	.w4(32'hbac455d9),
	.w5(32'hbb04ca58),
	.w6(32'hbb4892ed),
	.w7(32'hbae72eec),
	.w8(32'hbb13bf9b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a394cd0),
	.w1(32'hba42d529),
	.w2(32'hbb416fe6),
	.w3(32'h3818fce1),
	.w4(32'hb9f7f789),
	.w5(32'hbb80847f),
	.w6(32'h39396dc4),
	.w7(32'hba121015),
	.w8(32'hb8857dad),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ea6d3),
	.w1(32'hb89f4f12),
	.w2(32'h3a248580),
	.w3(32'hba7cf984),
	.w4(32'hbad0d8d7),
	.w5(32'hbb0fbd04),
	.w6(32'hba8c177f),
	.w7(32'hba44fd8d),
	.w8(32'hbb1268e2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e05e1),
	.w1(32'h3b9e5fe8),
	.w2(32'h3b8101a3),
	.w3(32'hb95c80dd),
	.w4(32'h3b84211b),
	.w5(32'h3b122a69),
	.w6(32'h3a4eb0e1),
	.w7(32'h3b8d63a3),
	.w8(32'h3b5a60aa),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bdfcb),
	.w1(32'h3afb34cd),
	.w2(32'h3b2f941e),
	.w3(32'h3b82ba60),
	.w4(32'h3b5c4ad6),
	.w5(32'h3afcf221),
	.w6(32'h3b16088d),
	.w7(32'hbadbcfba),
	.w8(32'h3ad0090b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ed77),
	.w1(32'h3adce504),
	.w2(32'h3b87679f),
	.w3(32'h3a48fa4e),
	.w4(32'h3b48f194),
	.w5(32'h3b903097),
	.w6(32'hba9a699b),
	.w7(32'hb997505b),
	.w8(32'hbb61d95d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b497884),
	.w1(32'h3b086028),
	.w2(32'h3a822934),
	.w3(32'h3ba47483),
	.w4(32'h3b0d69f2),
	.w5(32'h39888e7e),
	.w6(32'h3a09fe2d),
	.w7(32'h3bcacc3f),
	.w8(32'h3a884429),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ec048),
	.w1(32'hba27d894),
	.w2(32'hbb0dcd00),
	.w3(32'hbadb03da),
	.w4(32'hba5f3fec),
	.w5(32'hba6b859a),
	.w6(32'hba02a581),
	.w7(32'hba7dd35e),
	.w8(32'hbb271c84),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c38dd),
	.w1(32'h3bab257c),
	.w2(32'h3aece818),
	.w3(32'hba4bbc79),
	.w4(32'h3c13a7a8),
	.w5(32'h3bdcabc0),
	.w6(32'hbbad4e12),
	.w7(32'h3b585dc2),
	.w8(32'h3986a77f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d1684),
	.w1(32'h3c086133),
	.w2(32'h3c1b130a),
	.w3(32'h3c1832db),
	.w4(32'h3b8fbf3b),
	.w5(32'hba96c701),
	.w6(32'h3bf9194d),
	.w7(32'hb8d94564),
	.w8(32'hbbfefdd9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c9029),
	.w1(32'hba009e6b),
	.w2(32'hbb8ed2ab),
	.w3(32'hbbec5f52),
	.w4(32'hb7aae9ce),
	.w5(32'hbb60b26b),
	.w6(32'hbc0c96d9),
	.w7(32'hbaa9c2b4),
	.w8(32'h39ebc50d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8fac4),
	.w1(32'h3b03b0d3),
	.w2(32'h3aa19624),
	.w3(32'h3c34195b),
	.w4(32'h3bdb5c6f),
	.w5(32'h38ba61a7),
	.w6(32'h3bedd87c),
	.w7(32'h3891fcd9),
	.w8(32'h3ace6ac4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e2b5ee),
	.w1(32'hbaa47d21),
	.w2(32'hb98a484e),
	.w3(32'hbab82ee0),
	.w4(32'hba3f5c3b),
	.w5(32'hba807261),
	.w6(32'h3b26c7d8),
	.w7(32'hbb363d12),
	.w8(32'hbb22ff98),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fe4e5),
	.w1(32'h3ae0cc1b),
	.w2(32'hbb77aecc),
	.w3(32'hbb77068e),
	.w4(32'h3b8bde00),
	.w5(32'h3b0d1e09),
	.w6(32'hbbeaedbe),
	.w7(32'h3ad70c6d),
	.w8(32'hbb68f962),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaea4fd),
	.w1(32'h39ae827a),
	.w2(32'h3acd1032),
	.w3(32'hbc17052b),
	.w4(32'hba12e957),
	.w5(32'hba73a3e3),
	.w6(32'hbc7a5902),
	.w7(32'hbb8335d5),
	.w8(32'h3714a298),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0d87e),
	.w1(32'h3b984be8),
	.w2(32'h3af2c9f1),
	.w3(32'hbb106310),
	.w4(32'h3b07e196),
	.w5(32'h37625ab3),
	.w6(32'hbb56fc6b),
	.w7(32'h3b55b7d9),
	.w8(32'hbab334ff),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87cb71),
	.w1(32'h3b584cb8),
	.w2(32'h3b388a04),
	.w3(32'h3bbf0e21),
	.w4(32'h3aa8dde8),
	.w5(32'h3b801d82),
	.w6(32'h39fe1509),
	.w7(32'hbbb69bf7),
	.w8(32'h3ab3db00),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85aaa5),
	.w1(32'hb99f9403),
	.w2(32'hba027a7b),
	.w3(32'hba88c319),
	.w4(32'hbb009f38),
	.w5(32'hbb2deada),
	.w6(32'h38586c01),
	.w7(32'hbb232d51),
	.w8(32'hbbc43c91),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965e067),
	.w1(32'h3a76b1aa),
	.w2(32'h3bb6d2bd),
	.w3(32'h378b4ea5),
	.w4(32'h3bc71e0d),
	.w5(32'h3b73ec5e),
	.w6(32'h3aa04032),
	.w7(32'h39c9d876),
	.w8(32'h3b861355),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf007a),
	.w1(32'h3b52cc62),
	.w2(32'hba265a5e),
	.w3(32'h3b7fe552),
	.w4(32'h3acbb959),
	.w5(32'h3b6e5718),
	.w6(32'h3a822a18),
	.w7(32'hbb287d46),
	.w8(32'hbbc0ba91),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74aba9),
	.w1(32'hb9430caa),
	.w2(32'hbb8c8cff),
	.w3(32'hbb84387a),
	.w4(32'hba8cbc44),
	.w5(32'hbb8cd59f),
	.w6(32'hbad18343),
	.w7(32'hbb084184),
	.w8(32'hbb232e99),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0409bb),
	.w1(32'h3b09236e),
	.w2(32'h3a5730fd),
	.w3(32'hbad6814f),
	.w4(32'hbab29b84),
	.w5(32'hb9ebf703),
	.w6(32'hba1f8e22),
	.w7(32'hbbba6c02),
	.w8(32'hbb88d74b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f60112),
	.w1(32'h3b18da0e),
	.w2(32'h3c3754fc),
	.w3(32'hbaf357a8),
	.w4(32'h39d124f4),
	.w5(32'h3c52e78e),
	.w6(32'hbc2b0efc),
	.w7(32'h3afa89ba),
	.w8(32'h3b99bf9b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d659),
	.w1(32'hba8d4c35),
	.w2(32'hbbcabce4),
	.w3(32'hba58c8d9),
	.w4(32'hbac5dd3f),
	.w5(32'hbc37cac2),
	.w6(32'hbb5e4ce6),
	.w7(32'hbacd65eb),
	.w8(32'hbbee8d3e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb854990),
	.w1(32'h3ba81ab5),
	.w2(32'h3bb0d52e),
	.w3(32'hbba6dac9),
	.w4(32'h3c0a64a4),
	.w5(32'h3c39414b),
	.w6(32'hbbaf1134),
	.w7(32'hb9dfc854),
	.w8(32'hbba8c525),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dfae6),
	.w1(32'hbc4fd273),
	.w2(32'hbb9ab918),
	.w3(32'h3bc02fed),
	.w4(32'hbbcd2d9a),
	.w5(32'h39b16905),
	.w6(32'h3af8aad9),
	.w7(32'hbc2db6e4),
	.w8(32'hbb6b0138),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec28a),
	.w1(32'hba754faf),
	.w2(32'hba531ed4),
	.w3(32'h3971b32e),
	.w4(32'hbb1e4495),
	.w5(32'hbbcc5056),
	.w6(32'h3b9a2680),
	.w7(32'hbc3b4dd7),
	.w8(32'hbbd1fadf),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4549),
	.w1(32'h3983d779),
	.w2(32'hb9ec7f13),
	.w3(32'hbb697ebb),
	.w4(32'hbba88d16),
	.w5(32'hbbd090cb),
	.w6(32'hbbbe781f),
	.w7(32'h3b5d0561),
	.w8(32'h3b7f6da7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ba8f1),
	.w1(32'h3b42a3a1),
	.w2(32'hbaffea80),
	.w3(32'hbb0abe22),
	.w4(32'h3b64a612),
	.w5(32'hbb91edde),
	.w6(32'hbb06f854),
	.w7(32'hbadb0932),
	.w8(32'h3b7a1a5a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dfb68),
	.w1(32'h3b42d5d2),
	.w2(32'hbb8182b2),
	.w3(32'hbbf1a83d),
	.w4(32'h3a9a0de8),
	.w5(32'hbc5f64a8),
	.w6(32'hbc084537),
	.w7(32'hbb55bd19),
	.w8(32'hbc1e586f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9ad79),
	.w1(32'hbab982fd),
	.w2(32'h3b7b4eb4),
	.w3(32'hbbac1585),
	.w4(32'h3bb13f7e),
	.w5(32'h3c0d5ee4),
	.w6(32'hbc3d04ce),
	.w7(32'hbb2881d7),
	.w8(32'hbbcb3720),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea47bc),
	.w1(32'hbb926e0f),
	.w2(32'hbb346441),
	.w3(32'hba9d2c81),
	.w4(32'hbbc42ccd),
	.w5(32'h3aa5b06a),
	.w6(32'hbafb4276),
	.w7(32'hbbc7924b),
	.w8(32'hbbed1526),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4f8d5),
	.w1(32'hbb50ff98),
	.w2(32'hbba42882),
	.w3(32'hbb6f01af),
	.w4(32'h3b4339fa),
	.w5(32'h3be0398e),
	.w6(32'hbb303d93),
	.w7(32'hbbb7a221),
	.w8(32'hbb8b8ab1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeee347),
	.w1(32'h3b9f6974),
	.w2(32'h3be888e2),
	.w3(32'h39466d4b),
	.w4(32'h3c30ff85),
	.w5(32'h3c06bbc5),
	.w6(32'h3b1ee1ec),
	.w7(32'h3c2f9847),
	.w8(32'h3bfe3abe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b545726),
	.w1(32'hbab0db31),
	.w2(32'h3b0ad0ff),
	.w3(32'h3b85dbb9),
	.w4(32'h3ae7f0aa),
	.w5(32'h3bd93b29),
	.w6(32'h3c0a3b7d),
	.w7(32'hb8d519a0),
	.w8(32'h3b481f1b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11d699),
	.w1(32'h3b7198e5),
	.w2(32'hba52d075),
	.w3(32'h3705faf6),
	.w4(32'h3b299a3a),
	.w5(32'hbaf67f59),
	.w6(32'hbbadd754),
	.w7(32'hbb7a097d),
	.w8(32'hbc076ae5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb310d79),
	.w1(32'h3ad801ca),
	.w2(32'h3abec23e),
	.w3(32'hbb3521c1),
	.w4(32'h3b8a87a2),
	.w5(32'h3a24aaef),
	.w6(32'hbb223a70),
	.w7(32'h3b82af87),
	.w8(32'h3ae3a860),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa2ed1),
	.w1(32'hba6665e3),
	.w2(32'hbb8d95da),
	.w3(32'h3bfa64a9),
	.w4(32'h3a8aaf13),
	.w5(32'hbc15b469),
	.w6(32'hbb39c090),
	.w7(32'h3a130f85),
	.w8(32'h3b72933d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c08290),
	.w1(32'h3b9607b1),
	.w2(32'h3b89206b),
	.w3(32'hbbac4254),
	.w4(32'h3babe5c8),
	.w5(32'h3c6df4e8),
	.w6(32'hb98f7c87),
	.w7(32'h3bd254e1),
	.w8(32'h3c31c190),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2249aa),
	.w1(32'h3b02a46f),
	.w2(32'h3a1af730),
	.w3(32'h3bff6ff0),
	.w4(32'hba8a6e45),
	.w5(32'hbb104c5a),
	.w6(32'h3c0dd9ea),
	.w7(32'hbad09302),
	.w8(32'hbb155a6f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae72c2e),
	.w1(32'hbb76142e),
	.w2(32'hbbe4c0d5),
	.w3(32'hbb446920),
	.w4(32'hb7c3be08),
	.w5(32'hbb5786b4),
	.w6(32'h39eb840e),
	.w7(32'hbae0408b),
	.w8(32'hbc10ab88),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34c494),
	.w1(32'h3ba941eb),
	.w2(32'h3bc7b836),
	.w3(32'hbbc01dbb),
	.w4(32'h3b13097f),
	.w5(32'h394d3309),
	.w6(32'hbc7cf74b),
	.w7(32'hbba6782c),
	.w8(32'hbc33ae7b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fabae),
	.w1(32'hbb5d15c5),
	.w2(32'hbbc1e390),
	.w3(32'hb9c840dc),
	.w4(32'hbb3ad4ca),
	.w5(32'hbad55bd7),
	.w6(32'hbb684f26),
	.w7(32'hbbd62cbf),
	.w8(32'hbbd277d6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176a61),
	.w1(32'hbb7479f6),
	.w2(32'hbb6b6e62),
	.w3(32'hbb870474),
	.w4(32'hbb88712f),
	.w5(32'hba0a6d43),
	.w6(32'h3a0bcb61),
	.w7(32'hbacc4f57),
	.w8(32'h3b0358d9),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f6e2),
	.w1(32'hb91eb686),
	.w2(32'hbba0f8fa),
	.w3(32'h3aeaabed),
	.w4(32'h3adcc1c1),
	.w5(32'hbb634833),
	.w6(32'hba68e9d8),
	.w7(32'h3ac15e33),
	.w8(32'hb88f1d03),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba597c9f),
	.w1(32'h3b0660c4),
	.w2(32'h3be4677f),
	.w3(32'hb961c619),
	.w4(32'h3b4b7a92),
	.w5(32'h3c05284e),
	.w6(32'h3a6168ef),
	.w7(32'hbba950ca),
	.w8(32'hbb6fa79c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27c1d4),
	.w1(32'hbb687abc),
	.w2(32'hba6b7943),
	.w3(32'hbbaecc46),
	.w4(32'hbb2f0b1c),
	.w5(32'hbb18a495),
	.w6(32'hbbe14cdf),
	.w7(32'hbb86242b),
	.w8(32'hbb29e085),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995a535),
	.w1(32'hbb39f500),
	.w2(32'hbb8fb4f5),
	.w3(32'hbab00d5f),
	.w4(32'hb88ec704),
	.w5(32'hbb0f8b4a),
	.w6(32'hbb999bd5),
	.w7(32'hb902d6bc),
	.w8(32'h3b69bf91),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b82ba),
	.w1(32'h3b1968ac),
	.w2(32'h3b25eea5),
	.w3(32'h3b8274b5),
	.w4(32'h3b5dd8d9),
	.w5(32'h3c243578),
	.w6(32'h3b0b5263),
	.w7(32'h3b7269f3),
	.w8(32'h3b56252d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54a66d),
	.w1(32'h3a1926a2),
	.w2(32'h3b69c9ef),
	.w3(32'h3bcba8fe),
	.w4(32'hba12befb),
	.w5(32'hbc6aa201),
	.w6(32'h3b8712a2),
	.w7(32'h3b2f3990),
	.w8(32'h3b1d081c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85495d),
	.w1(32'h3c119113),
	.w2(32'hbaba44ea),
	.w3(32'hbb14e84b),
	.w4(32'h3c61fdc4),
	.w5(32'hbb372243),
	.w6(32'h3b4b85ac),
	.w7(32'h3be4f0c8),
	.w8(32'hbbb60a67),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75123e),
	.w1(32'h3bfad92b),
	.w2(32'h3b801c34),
	.w3(32'hbb4b170e),
	.w4(32'h3c27d447),
	.w5(32'h3ad654fa),
	.w6(32'hbc0007bd),
	.w7(32'h3ad9ddad),
	.w8(32'hbb0d002d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e4fb8),
	.w1(32'h3a74b278),
	.w2(32'h3b12f456),
	.w3(32'h3a5e130d),
	.w4(32'h39fea69c),
	.w5(32'h3c0e278b),
	.w6(32'hbacdec30),
	.w7(32'hbb4ee8a5),
	.w8(32'hbbe8f984),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11647e),
	.w1(32'hba66d2a5),
	.w2(32'hbb9b2bc5),
	.w3(32'hb944a16c),
	.w4(32'hbaca0de4),
	.w5(32'hbb954671),
	.w6(32'h3bd42a2f),
	.w7(32'hbb5182ee),
	.w8(32'hbb9d6a3e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4242b3),
	.w1(32'h3b9c2752),
	.w2(32'h3b8548ce),
	.w3(32'h3b67d475),
	.w4(32'h3beead55),
	.w5(32'h3bf93206),
	.w6(32'h3b843532),
	.w7(32'h3bd6da0e),
	.w8(32'h3b5c88f1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ae92),
	.w1(32'h3aecf7f6),
	.w2(32'h3a38edd6),
	.w3(32'h3ba87ae6),
	.w4(32'hba80141e),
	.w5(32'hbb40ad24),
	.w6(32'hbae1171b),
	.w7(32'hbabc5fd3),
	.w8(32'hb9efb76c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50137),
	.w1(32'hbac4ffed),
	.w2(32'hbabc2ce9),
	.w3(32'hbae6fbac),
	.w4(32'h3b7268fa),
	.w5(32'hbba680eb),
	.w6(32'hbb6662b0),
	.w7(32'hbbbb2e2f),
	.w8(32'hbb31dd0e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0165ba),
	.w1(32'hbb49aa2b),
	.w2(32'hbb8a07a1),
	.w3(32'hbb18f807),
	.w4(32'h3a08a144),
	.w5(32'hbb46a07f),
	.w6(32'hbb7fa008),
	.w7(32'hbbd1e245),
	.w8(32'hbbadfc01),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae79dec),
	.w1(32'hbac0466c),
	.w2(32'h3b827018),
	.w3(32'hbb3de595),
	.w4(32'hbb4395c9),
	.w5(32'hbb4b8a73),
	.w6(32'hbb101850),
	.w7(32'hbabe0f52),
	.w8(32'hba27b853),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5433ed),
	.w1(32'hba073e1d),
	.w2(32'hbad97320),
	.w3(32'h3b10062a),
	.w4(32'h3ab2d746),
	.w5(32'h3a22d6f4),
	.w6(32'h39a04f5b),
	.w7(32'hba78c39e),
	.w8(32'hba9f4bfe),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d69b8),
	.w1(32'h390981b7),
	.w2(32'h3bc97d40),
	.w3(32'hba0d997f),
	.w4(32'hba2d1472),
	.w5(32'hbb0b081d),
	.w6(32'h39fd8645),
	.w7(32'hb875e898),
	.w8(32'h3aef67b3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59a0a2),
	.w1(32'h3b8ac0ee),
	.w2(32'h3bb5985c),
	.w3(32'hbb46e6a2),
	.w4(32'h3b82fdfa),
	.w5(32'h3bae42d2),
	.w6(32'hbaa86b49),
	.w7(32'hba6a3ffa),
	.w8(32'hba5976e0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05575f),
	.w1(32'h3b385770),
	.w2(32'h3a0ee675),
	.w3(32'h3b3182b2),
	.w4(32'h3b5cf81b),
	.w5(32'hbae53706),
	.w6(32'hbb652488),
	.w7(32'h3b3e1537),
	.w8(32'hbb311716),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e23d9),
	.w1(32'hbb19cdb5),
	.w2(32'hbb956a71),
	.w3(32'hbc2b3d61),
	.w4(32'h3b8d0b8b),
	.w5(32'h3b135fa4),
	.w6(32'hbad24817),
	.w7(32'hbb5039e5),
	.w8(32'hbb437c28),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58f7ef),
	.w1(32'hbbd284b2),
	.w2(32'hbb7e3ebf),
	.w3(32'h3ad69751),
	.w4(32'h3c55c11c),
	.w5(32'h3c49dcd6),
	.w6(32'hbb9915d0),
	.w7(32'h3b56e258),
	.w8(32'hbaf56004),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed9957),
	.w1(32'hbb29b0e9),
	.w2(32'hbb4bcfe8),
	.w3(32'h3aac0682),
	.w4(32'hbbb5c3aa),
	.w5(32'hbb81be03),
	.w6(32'h3bb6c172),
	.w7(32'hbc6afaf7),
	.w8(32'hbc725a56),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbece6f3),
	.w1(32'hb8bbbafb),
	.w2(32'hbb208464),
	.w3(32'hbc789c9e),
	.w4(32'hbba6a3eb),
	.w5(32'h39cef3f2),
	.w6(32'hbc9dc3f5),
	.w7(32'hbaf7233c),
	.w8(32'hbab3315e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule