module layer_10_featuremap_483(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eefcfb),
	.w1(32'h3afe2d40),
	.w2(32'hba84d857),
	.w3(32'hbbb83c81),
	.w4(32'h3be9cd1a),
	.w5(32'hbc14d09b),
	.w6(32'hbb6fe7e0),
	.w7(32'h3be5a24a),
	.w8(32'h3bb2e984),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e25b),
	.w1(32'hbb9bb7db),
	.w2(32'h3b2e4ee7),
	.w3(32'h3c0f316e),
	.w4(32'h3be3337a),
	.w5(32'h3c819fc9),
	.w6(32'h3a756ed0),
	.w7(32'hbb1920dc),
	.w8(32'h3a7d0abb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaed545),
	.w1(32'h3c15f483),
	.w2(32'hbbcc0aac),
	.w3(32'hbbf9f10e),
	.w4(32'h3c22983e),
	.w5(32'h3c508af3),
	.w6(32'hbc2f2e01),
	.w7(32'hb9918b97),
	.w8(32'h3aba1783),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b691e),
	.w1(32'hba37cceb),
	.w2(32'h3bb02bec),
	.w3(32'h3a518ec8),
	.w4(32'hbc03114a),
	.w5(32'hbac21965),
	.w6(32'h3b0c006a),
	.w7(32'hbba2e016),
	.w8(32'h3b4a8a49),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74a1a1),
	.w1(32'h39bf7474),
	.w2(32'h3b0a9228),
	.w3(32'h3a1fc8cc),
	.w4(32'h3b8005c4),
	.w5(32'h3a8a1642),
	.w6(32'h3c1510d8),
	.w7(32'h3c064a7c),
	.w8(32'h3b7ed76d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b387c),
	.w1(32'hbad65f1d),
	.w2(32'hbade2012),
	.w3(32'h3a9e9047),
	.w4(32'h3b6510c2),
	.w5(32'h3b17ef89),
	.w6(32'hb939af0f),
	.w7(32'h3bb0ab8e),
	.w8(32'h3bb30a51),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b864282),
	.w1(32'hb84ce854),
	.w2(32'h3aa7315f),
	.w3(32'hbac10b63),
	.w4(32'hbc1bb42b),
	.w5(32'hbbcea4f9),
	.w6(32'hbbabaa52),
	.w7(32'h3a87799d),
	.w8(32'h3adf3b0d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c5649),
	.w1(32'h3b442b6a),
	.w2(32'hbbc97d0a),
	.w3(32'hbc481033),
	.w4(32'hbb8a7048),
	.w5(32'hbc2a283a),
	.w6(32'hbc16b646),
	.w7(32'h39c9c491),
	.w8(32'hbbdb362b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdefabd),
	.w1(32'hbacb91fc),
	.w2(32'h3c213e21),
	.w3(32'h3a38849d),
	.w4(32'hbb5e681a),
	.w5(32'hbb464af1),
	.w6(32'hbb808d0d),
	.w7(32'h3ac5c9cf),
	.w8(32'h3bae512d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b96e2),
	.w1(32'hba0722a5),
	.w2(32'h3b0ea96c),
	.w3(32'hbb4917a3),
	.w4(32'hbb2d93c7),
	.w5(32'hbb1d7084),
	.w6(32'h3ac27854),
	.w7(32'hba77135e),
	.w8(32'h3bb51086),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6bab8),
	.w1(32'h3c77ce18),
	.w2(32'h3bde7b1b),
	.w3(32'hbb08762c),
	.w4(32'h3c21b09a),
	.w5(32'h3ce04892),
	.w6(32'h37d7f2f2),
	.w7(32'hbbb1ae03),
	.w8(32'h3a0397a7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9f49),
	.w1(32'hbb47d23a),
	.w2(32'h3b4f055a),
	.w3(32'h3b9e918a),
	.w4(32'hbbfd198f),
	.w5(32'hbb9a4160),
	.w6(32'h3b8184f9),
	.w7(32'hbb44c20a),
	.w8(32'hbc23e307),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd77653),
	.w1(32'hbbba8de8),
	.w2(32'h39ae20fd),
	.w3(32'h3b0a169d),
	.w4(32'hbbca4beb),
	.w5(32'hbbca03a2),
	.w6(32'hbc104e89),
	.w7(32'hbbc69177),
	.w8(32'hbc6edf45),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1581b5),
	.w1(32'h3b2e59e4),
	.w2(32'h3b1e57b4),
	.w3(32'hbc14f945),
	.w4(32'h3b3f9e8a),
	.w5(32'h3c81a4b4),
	.w6(32'hbbb12d75),
	.w7(32'hba93baa8),
	.w8(32'h3b9bc64c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed8fa3),
	.w1(32'h3b65d095),
	.w2(32'hbbc20398),
	.w3(32'h3ae420b7),
	.w4(32'h3b4abf49),
	.w5(32'hbbc457d8),
	.w6(32'h3b6b6468),
	.w7(32'h3bb2109d),
	.w8(32'h3ba9c958),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda60be),
	.w1(32'hbb3076a8),
	.w2(32'hbb2f9215),
	.w3(32'hbbf861ae),
	.w4(32'hba9d7c59),
	.w5(32'hbc6727cb),
	.w6(32'hbb7f23f2),
	.w7(32'h3ad1c41e),
	.w8(32'hbbfe5f72),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f7776),
	.w1(32'h3b38569a),
	.w2(32'h3aff384b),
	.w3(32'hbaf3ac55),
	.w4(32'h3b9f4f58),
	.w5(32'h3a9e8b4c),
	.w6(32'hbc2d3a43),
	.w7(32'h3b3f4325),
	.w8(32'h3c08632e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3192bf),
	.w1(32'h3b804ce8),
	.w2(32'hbb4d8677),
	.w3(32'hbb464305),
	.w4(32'h3c030162),
	.w5(32'hbbf764b9),
	.w6(32'hb8abc39e),
	.w7(32'h3b6ccbc2),
	.w8(32'h3b283410),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45891a),
	.w1(32'hba1176c0),
	.w2(32'h3ae7f7d0),
	.w3(32'hbbb5978c),
	.w4(32'h3be82fdc),
	.w5(32'hba99f4af),
	.w6(32'hbab5d064),
	.w7(32'h3c1041e0),
	.w8(32'h3ace8e18),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea426),
	.w1(32'h3c1479a6),
	.w2(32'hbc44f8e8),
	.w3(32'h3a867e8b),
	.w4(32'h3c325602),
	.w5(32'hbb6adb08),
	.w6(32'hbb568e6d),
	.w7(32'h3a8a8198),
	.w8(32'hbb642c10),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0321a5),
	.w1(32'hbbf7aa18),
	.w2(32'hbb8014ed),
	.w3(32'hbbc40e0d),
	.w4(32'hbbcba1e2),
	.w5(32'hbb79752a),
	.w6(32'hbb26d774),
	.w7(32'hbace75ab),
	.w8(32'hbbd0f382),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e5e40),
	.w1(32'hba47505c),
	.w2(32'hbbd66354),
	.w3(32'hbbf165b9),
	.w4(32'hbba45a64),
	.w5(32'hbad2d2f3),
	.w6(32'hbb8dc101),
	.w7(32'hbc1136c0),
	.w8(32'hbc0b9978),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10ab44),
	.w1(32'h3bdcf8ae),
	.w2(32'h3b44350e),
	.w3(32'hbc0e401a),
	.w4(32'hbab80eff),
	.w5(32'hbc02c22e),
	.w6(32'hbb82e493),
	.w7(32'hbb6125f5),
	.w8(32'hbb2417af),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99393d),
	.w1(32'h3b0f6c78),
	.w2(32'hbb7fc0ef),
	.w3(32'hba8975ac),
	.w4(32'hbb0447ca),
	.w5(32'hbc65633f),
	.w6(32'h3c12699b),
	.w7(32'h396428a1),
	.w8(32'hbbe362ec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104d28),
	.w1(32'hbba36e94),
	.w2(32'hbbd05d6c),
	.w3(32'hbbb99dd1),
	.w4(32'hbc583492),
	.w5(32'h3b7a3d54),
	.w6(32'hb7e84252),
	.w7(32'hbc6ca2b1),
	.w8(32'h3b444e8f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55d9ea),
	.w1(32'hba9d6191),
	.w2(32'hbba0272f),
	.w3(32'hbc1225ff),
	.w4(32'hbb468eb5),
	.w5(32'h3bb27ca4),
	.w6(32'hbb83e739),
	.w7(32'hbbadd4dc),
	.w8(32'hbbfca66e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029ce6),
	.w1(32'hbb8fd3db),
	.w2(32'hbb6abed4),
	.w3(32'h391fbe94),
	.w4(32'hbbe26bcb),
	.w5(32'hbc56317c),
	.w6(32'h3bb54d71),
	.w7(32'h3a52059f),
	.w8(32'hbc2d1b0e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af914),
	.w1(32'hbb737ce6),
	.w2(32'hbc0ed72f),
	.w3(32'hbc081272),
	.w4(32'hbbc6ffaa),
	.w5(32'hbb21d711),
	.w6(32'hbc1a57ab),
	.w7(32'hbb3f65de),
	.w8(32'hba5c1edf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1ee42),
	.w1(32'hbba3314a),
	.w2(32'hbc1d2977),
	.w3(32'hbbbef549),
	.w4(32'hbc035502),
	.w5(32'hbbadd830),
	.w6(32'hbbc5f84e),
	.w7(32'h3b75e485),
	.w8(32'h3b9eda7b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8fc01),
	.w1(32'hbb3d238e),
	.w2(32'h3b781142),
	.w3(32'h3b52c2de),
	.w4(32'hbc11a850),
	.w5(32'h3b8efcdf),
	.w6(32'h3bed73af),
	.w7(32'hbc28e6c7),
	.w8(32'hbb072555),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf318a),
	.w1(32'h3b2fdf30),
	.w2(32'hbb7493e3),
	.w3(32'hba960e7e),
	.w4(32'h3aa074e8),
	.w5(32'hbbc779af),
	.w6(32'hba680d57),
	.w7(32'hbb4074a4),
	.w8(32'h3aecdd4b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00579),
	.w1(32'h3bb312fd),
	.w2(32'h3b2ef73a),
	.w3(32'hbb33d0f6),
	.w4(32'hbb7bdf0d),
	.w5(32'h3b7e25f4),
	.w6(32'h3b9f9e0b),
	.w7(32'h3b40d408),
	.w8(32'h3bcb04b7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996f4f),
	.w1(32'h3c1b1d41),
	.w2(32'h3c0eaf42),
	.w3(32'hbad22521),
	.w4(32'h3b132fd1),
	.w5(32'h3b6f8360),
	.w6(32'h3b58f0f5),
	.w7(32'h3ab33cbf),
	.w8(32'h3c0f16f5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47892a),
	.w1(32'h3aad42d9),
	.w2(32'hbb28c660),
	.w3(32'h3b92cb11),
	.w4(32'h3aadbbdf),
	.w5(32'h3bd93457),
	.w6(32'hbb3e8e7f),
	.w7(32'hba2dc6a8),
	.w8(32'hbb80e352),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81873e),
	.w1(32'h3bc46794),
	.w2(32'h3b70ab64),
	.w3(32'h3b917b9e),
	.w4(32'h3babec87),
	.w5(32'hbb4ccd11),
	.w6(32'h3af57dac),
	.w7(32'h3bac764c),
	.w8(32'hbc06f386),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db1a0),
	.w1(32'h3bdad3f2),
	.w2(32'h3bb402e9),
	.w3(32'h3ba6469e),
	.w4(32'h3ba1eb5a),
	.w5(32'h3b343412),
	.w6(32'hbbc143b1),
	.w7(32'h3bb311de),
	.w8(32'h3b6fb20d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fef3e),
	.w1(32'h3b3e7ef1),
	.w2(32'hbbca93ff),
	.w3(32'h39e5adc2),
	.w4(32'hbb993980),
	.w5(32'h3c87c792),
	.w6(32'h3ba59d46),
	.w7(32'hbc1289ad),
	.w8(32'h3ab27b29),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc336698),
	.w1(32'h3a71d667),
	.w2(32'hb9cdce8d),
	.w3(32'hbbcbfb21),
	.w4(32'hbb3d2e11),
	.w5(32'h3bcbdb75),
	.w6(32'h3c0abd3f),
	.w7(32'hbb4b6a3c),
	.w8(32'hbac1e250),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89d0bd),
	.w1(32'h3b70de71),
	.w2(32'h3c265699),
	.w3(32'hbb7826fa),
	.w4(32'h39a449d8),
	.w5(32'hba56ca3f),
	.w6(32'hbba985cf),
	.w7(32'hbaa1fd40),
	.w8(32'h3aeb7769),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22fbb6),
	.w1(32'hbad7bad0),
	.w2(32'hbba0f3bd),
	.w3(32'h3c1be6f0),
	.w4(32'hbac7e337),
	.w5(32'hba2f891e),
	.w6(32'h3c0e08f6),
	.w7(32'hbb8a2333),
	.w8(32'hbbccbffe),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffb701),
	.w1(32'h3a2e0259),
	.w2(32'h3c71c035),
	.w3(32'hbb71e04d),
	.w4(32'h3a1e0bc3),
	.w5(32'h3b709351),
	.w6(32'hba03023d),
	.w7(32'h3a8e2ed1),
	.w8(32'h3c08e608),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f9bbb),
	.w1(32'h3b73b7fc),
	.w2(32'h39e2ab38),
	.w3(32'h3b13d083),
	.w4(32'hbbb12580),
	.w5(32'h38e3880e),
	.w6(32'h3bcf923f),
	.w7(32'h3abf401f),
	.w8(32'hbb6cdc7f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009ab9),
	.w1(32'h3af7d49b),
	.w2(32'h3bb100a8),
	.w3(32'h3ad2b043),
	.w4(32'hbb41f052),
	.w5(32'h3be31c8c),
	.w6(32'hbbc4abf4),
	.w7(32'hbb9c1a0e),
	.w8(32'h3c0070d6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb347417),
	.w1(32'h39dc81e7),
	.w2(32'hbb2aa4ca),
	.w3(32'h3971724f),
	.w4(32'hbb308c3d),
	.w5(32'h39d93a23),
	.w6(32'h3bbd7ffd),
	.w7(32'hbb58faed),
	.w8(32'hbb5b0774),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d876f),
	.w1(32'hbb9dba86),
	.w2(32'hbb7bf05c),
	.w3(32'hbbbb54d5),
	.w4(32'h3b051c4c),
	.w5(32'hbb876891),
	.w6(32'hbb3f9272),
	.w7(32'h3bae345f),
	.w8(32'h3be7cf8f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78652d),
	.w1(32'hbaca30a4),
	.w2(32'h3c0c292b),
	.w3(32'h39b99876),
	.w4(32'hba54498b),
	.w5(32'hbbf1c797),
	.w6(32'hba62675d),
	.w7(32'h3bb69e10),
	.w8(32'hbc08f909),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92e93f),
	.w1(32'hb7fbd3c3),
	.w2(32'h38980dfb),
	.w3(32'h3bcb7f05),
	.w4(32'hbc0f8b54),
	.w5(32'hbbc49ec1),
	.w6(32'hbc07aefd),
	.w7(32'hbc32fea6),
	.w8(32'hbc5e7224),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4978ae),
	.w1(32'h3b1a02f7),
	.w2(32'h3c270d41),
	.w3(32'hbbe9c8db),
	.w4(32'hbb352f06),
	.w5(32'h3bfd1617),
	.w6(32'hbc33e6b1),
	.w7(32'hbb373954),
	.w8(32'h3bb9a3a7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ab192),
	.w1(32'h3b50585d),
	.w2(32'h3c027e33),
	.w3(32'h3c0d891c),
	.w4(32'h3a45a24c),
	.w5(32'hba8be698),
	.w6(32'h3ba0c363),
	.w7(32'h3aeeb5cc),
	.w8(32'h3b0b1757),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef2cfc),
	.w1(32'h3bd24559),
	.w2(32'h3b61e56e),
	.w3(32'h3aaabdbc),
	.w4(32'hb9a35f94),
	.w5(32'hbb54a83a),
	.w6(32'hbbbf3595),
	.w7(32'h3bd7e686),
	.w8(32'h3c0320fe),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a82d5),
	.w1(32'h3af339ea),
	.w2(32'h3b945d66),
	.w3(32'hb928cbe5),
	.w4(32'h3ba1bff8),
	.w5(32'hbbf23327),
	.w6(32'hbb6f4626),
	.w7(32'h3a9608d8),
	.w8(32'h3b2ef5b4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b754333),
	.w1(32'h3be46547),
	.w2(32'h3bc9d3a5),
	.w3(32'hbaad5b3d),
	.w4(32'hba44cdd0),
	.w5(32'h3b2078ef),
	.w6(32'hbc030b7f),
	.w7(32'h3b13535e),
	.w8(32'hbbd029ff),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee5541),
	.w1(32'h3aad489f),
	.w2(32'h3999c679),
	.w3(32'h3ad130bd),
	.w4(32'h38f1f14a),
	.w5(32'hbb364782),
	.w6(32'h3a9b9107),
	.w7(32'hbad68fc7),
	.w8(32'h3a9edb62),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a242e1f),
	.w1(32'hba48260e),
	.w2(32'hba8e362a),
	.w3(32'h3ac0aac7),
	.w4(32'hbc0ea2f2),
	.w5(32'h3b6aa8fc),
	.w6(32'h3abb7add),
	.w7(32'h3af26229),
	.w8(32'hbc1b9951),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e957),
	.w1(32'hbc11058d),
	.w2(32'hbc1998d4),
	.w3(32'hba489222),
	.w4(32'hbc15efc5),
	.w5(32'hb9bdbe2a),
	.w6(32'h3ba7d3e3),
	.w7(32'hbc4fd57c),
	.w8(32'hbba812d8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b04f),
	.w1(32'hba285a34),
	.w2(32'h3c2ba305),
	.w3(32'hbc000da0),
	.w4(32'hbba58775),
	.w5(32'h3c2efa64),
	.w6(32'hbb1952f0),
	.w7(32'hbbce34db),
	.w8(32'h39c56d96),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18123c),
	.w1(32'hbb23769b),
	.w2(32'h3ad1afa2),
	.w3(32'hbb73f14b),
	.w4(32'hbb212299),
	.w5(32'h3bba175f),
	.w6(32'h3b07bf9c),
	.w7(32'h3b16c96c),
	.w8(32'hbbdf22b1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43d7f2),
	.w1(32'h3a4a2fd6),
	.w2(32'hbb911ad1),
	.w3(32'hbb0c2d2f),
	.w4(32'h3ab8c551),
	.w5(32'h3b0fde4f),
	.w6(32'hbbca2e7c),
	.w7(32'h3aa8b75d),
	.w8(32'hbbb67f4b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38a241),
	.w1(32'hbb6d69bf),
	.w2(32'hba0c1eff),
	.w3(32'hbb8829d8),
	.w4(32'hb782fdb5),
	.w5(32'h3b68d488),
	.w6(32'hbb4ff7dd),
	.w7(32'h3bb85f86),
	.w8(32'h3b14d64a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8511d),
	.w1(32'h3c5b9748),
	.w2(32'h3c8c8df1),
	.w3(32'hb7801b0b),
	.w4(32'h3c0da9ca),
	.w5(32'h3d01c735),
	.w6(32'h3af43559),
	.w7(32'h3b94e483),
	.w8(32'hbb53c87a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacc084),
	.w1(32'h3ba6cfbd),
	.w2(32'h3c384fe7),
	.w3(32'h3c931de7),
	.w4(32'hbb972711),
	.w5(32'hbc50d654),
	.w6(32'h3c4f6e1c),
	.w7(32'hbba85d3d),
	.w8(32'hba9c2d8d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c362055),
	.w1(32'hbbe0b338),
	.w2(32'hbb546022),
	.w3(32'hbc150764),
	.w4(32'hbbd76071),
	.w5(32'hba3f079e),
	.w6(32'hba8a4772),
	.w7(32'h3b66972c),
	.w8(32'h3bf23a59),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcecc9e),
	.w1(32'hbb94965e),
	.w2(32'hbb7365f9),
	.w3(32'hb9da0276),
	.w4(32'hbc55dbf0),
	.w5(32'h3b17ca56),
	.w6(32'h3b235e44),
	.w7(32'hbc6b3d0c),
	.w8(32'h3adcad4a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2734cd),
	.w1(32'hbadba14a),
	.w2(32'h39995d1e),
	.w3(32'hbbf3bcc9),
	.w4(32'h3ba935a5),
	.w5(32'hbbaa8277),
	.w6(32'h3b80a827),
	.w7(32'h3bd9b2f4),
	.w8(32'h3900db26),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27499d),
	.w1(32'h3bd5e7ac),
	.w2(32'h3b4781d8),
	.w3(32'h3bb8a859),
	.w4(32'h3bb6c20b),
	.w5(32'hbbcd6ae0),
	.w6(32'hbb48efca),
	.w7(32'h3c152729),
	.w8(32'hba0e4e0e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf5576),
	.w1(32'hba975e2d),
	.w2(32'hbb84b4bc),
	.w3(32'h3ba74be4),
	.w4(32'hbb925787),
	.w5(32'h38afb98f),
	.w6(32'h3ba2780e),
	.w7(32'hbbd5698a),
	.w8(32'hbbe44d07),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc915c63),
	.w1(32'hbbd40f6d),
	.w2(32'hbbbefb05),
	.w3(32'hbc34d703),
	.w4(32'h3b8e80db),
	.w5(32'h3a520306),
	.w6(32'hba098d69),
	.w7(32'hbae00e9a),
	.w8(32'hbb918291),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b514c),
	.w1(32'hbb3b73cf),
	.w2(32'hbc152fe5),
	.w3(32'hbbc2ffd5),
	.w4(32'h38be2741),
	.w5(32'h3a4ac145),
	.w6(32'hbc36980f),
	.w7(32'h3b743179),
	.w8(32'h3c98eed0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba461aa),
	.w1(32'hba97d6b2),
	.w2(32'h3cd7d9e9),
	.w3(32'hbb648f5a),
	.w4(32'h3c05e186),
	.w5(32'h3c5d9185),
	.w6(32'h3bf03e1e),
	.w7(32'h3bfc28af),
	.w8(32'h3cb3c695),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1415cc),
	.w1(32'hbc09a6d6),
	.w2(32'hbb827fd1),
	.w3(32'hbb397edb),
	.w4(32'h3a208ed7),
	.w5(32'hbac5f01c),
	.w6(32'h3a7becec),
	.w7(32'h3be9f5e0),
	.w8(32'h3b8f8422),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11644),
	.w1(32'hbb0590e3),
	.w2(32'hba65c2e9),
	.w3(32'hbbe5de5b),
	.w4(32'hba9c8c1b),
	.w5(32'hbb980f77),
	.w6(32'hbb9ca360),
	.w7(32'hbaa6958e),
	.w8(32'hbbb96434),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8ce31),
	.w1(32'h3c27a84a),
	.w2(32'hba361111),
	.w3(32'hbbef59de),
	.w4(32'hb8a564dd),
	.w5(32'h3b9e07a2),
	.w6(32'hbbd65d1d),
	.w7(32'hb9ea7cd0),
	.w8(32'hbbe6e42a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca1813),
	.w1(32'h3b1ec7c1),
	.w2(32'hba275943),
	.w3(32'h3b904afa),
	.w4(32'h3a1f4555),
	.w5(32'h3c1d0e2e),
	.w6(32'h3a873ede),
	.w7(32'h3baedd71),
	.w8(32'h3be98df0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c5e07),
	.w1(32'h3a958812),
	.w2(32'h3b731a7e),
	.w3(32'hba45dc15),
	.w4(32'h3abfd790),
	.w5(32'hbb246c09),
	.w6(32'h3b64c77b),
	.w7(32'hba1170fa),
	.w8(32'hb92ea5f8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d5d32),
	.w1(32'h381b1e9e),
	.w2(32'hba590cde),
	.w3(32'hbadbe06f),
	.w4(32'hbb19ffb0),
	.w5(32'h3b356a88),
	.w6(32'h3b257010),
	.w7(32'hbb336e94),
	.w8(32'hbb54ec6b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01af73),
	.w1(32'h3bb63066),
	.w2(32'h3bec05b0),
	.w3(32'hbb5ac80e),
	.w4(32'h3b0beceb),
	.w5(32'h3af7e61a),
	.w6(32'h3b074093),
	.w7(32'hbb3b0680),
	.w8(32'h3bbb08d1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b1772),
	.w1(32'h3a09d032),
	.w2(32'hbb5dd9fc),
	.w3(32'hba323ba3),
	.w4(32'h3c010c4d),
	.w5(32'hbbc2b254),
	.w6(32'h3b957a9c),
	.w7(32'h3b9eb63d),
	.w8(32'h3baeaf1f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd21182),
	.w1(32'h3b1c740b),
	.w2(32'h3bee06fe),
	.w3(32'hbbf95a4f),
	.w4(32'hbbd02322),
	.w5(32'h3c209a32),
	.w6(32'hb8ba622d),
	.w7(32'hbbb3ff0e),
	.w8(32'hbc1ce8c4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5452f),
	.w1(32'hbafd303d),
	.w2(32'h39f6d459),
	.w3(32'h3c513eaa),
	.w4(32'hb9fdb98f),
	.w5(32'h3b31d0e4),
	.w6(32'h3b737323),
	.w7(32'hbacb45e9),
	.w8(32'hbb8f978e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae125f5),
	.w1(32'h3a5abeea),
	.w2(32'h3a8e3483),
	.w3(32'h3bcc1cc4),
	.w4(32'hbb80446b),
	.w5(32'hbbba15ff),
	.w6(32'h39f131d5),
	.w7(32'hbb706b67),
	.w8(32'h3ac8395d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a595b),
	.w1(32'h3b7467b8),
	.w2(32'h3a2f8eea),
	.w3(32'hbbcd2f03),
	.w4(32'h3b2e7ba9),
	.w5(32'hbb451066),
	.w6(32'hbb66faa3),
	.w7(32'h3aea77e2),
	.w8(32'hbb77f056),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0c496),
	.w1(32'hbb9f0d72),
	.w2(32'hbb8b41cd),
	.w3(32'h3b60a3fc),
	.w4(32'hbbaa199d),
	.w5(32'hbb85b0b6),
	.w6(32'h3b999b31),
	.w7(32'hbb2878e7),
	.w8(32'hbb0ccc08),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab19fbf),
	.w1(32'h3ba46806),
	.w2(32'h3a607921),
	.w3(32'hbb5caca7),
	.w4(32'h3a955648),
	.w5(32'h3be7562d),
	.w6(32'hba0538a0),
	.w7(32'h39187b70),
	.w8(32'h39cd852e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba951f42),
	.w1(32'h397edbf7),
	.w2(32'h3b3ca8e8),
	.w3(32'hbb0a80b6),
	.w4(32'h39b7c044),
	.w5(32'hba285b8b),
	.w6(32'h3bd00391),
	.w7(32'hba9aa42b),
	.w8(32'hbb01bdad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fb76d),
	.w1(32'h3be20ee1),
	.w2(32'h3bfabdbe),
	.w3(32'hbb167469),
	.w4(32'hbba383ba),
	.w5(32'h3c68f692),
	.w6(32'hbb1084ed),
	.w7(32'hbb206840),
	.w8(32'hbb5fdd6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3214f5),
	.w1(32'h39fd3791),
	.w2(32'h3b2a6d17),
	.w3(32'h3c3af826),
	.w4(32'hbaf9d4ce),
	.w5(32'hbb7c0e0f),
	.w6(32'h39db064e),
	.w7(32'hbb62f8f5),
	.w8(32'h3b837fbb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34532032),
	.w1(32'h3b84da6a),
	.w2(32'h3baeedd9),
	.w3(32'h3ae1f6de),
	.w4(32'hb9826099),
	.w5(32'h3c8ebed1),
	.w6(32'hbbb00908),
	.w7(32'hbb4e6944),
	.w8(32'hbaaf24c5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aa9d6),
	.w1(32'h3aed3e6c),
	.w2(32'hb88359bf),
	.w3(32'h3bd91922),
	.w4(32'h3bd69310),
	.w5(32'h3c3f13f7),
	.w6(32'hbb504baa),
	.w7(32'hbb8068d4),
	.w8(32'hbb45ee66),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9344d8),
	.w1(32'hbaa58ddc),
	.w2(32'hb97807b7),
	.w3(32'hb9df4bc5),
	.w4(32'h3b9bf1dc),
	.w5(32'h3acd66df),
	.w6(32'h3a2bf370),
	.w7(32'h3b0bc299),
	.w8(32'h3be3cdf3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf38de8),
	.w1(32'h3ad73a1c),
	.w2(32'h3a8b21d6),
	.w3(32'hbbb84fc2),
	.w4(32'h3a9a9055),
	.w5(32'h3c264d40),
	.w6(32'h3a357242),
	.w7(32'hb9a406a2),
	.w8(32'h3bc0f93c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb038af9),
	.w1(32'hbb4e685c),
	.w2(32'hbb4e416b),
	.w3(32'h3b3641dc),
	.w4(32'hbb8548e0),
	.w5(32'hbb8cf869),
	.w6(32'h3b172f5f),
	.w7(32'h3a9bf88a),
	.w8(32'hba1627f1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61fc1c),
	.w1(32'hba1e2ecd),
	.w2(32'hbb16c6ba),
	.w3(32'hbb83485a),
	.w4(32'hbab3372e),
	.w5(32'hbaa0f841),
	.w6(32'hb882eddf),
	.w7(32'hbb03d72c),
	.w8(32'h3a1aa4ee),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d55b1),
	.w1(32'hbb1dfcd3),
	.w2(32'hbbd89a57),
	.w3(32'h3a30c61a),
	.w4(32'hbb88fe73),
	.w5(32'hbb381000),
	.w6(32'hbbcfa5f9),
	.w7(32'h3b6b9253),
	.w8(32'h389d4c44),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030ae4),
	.w1(32'hbb46b474),
	.w2(32'hba9235a5),
	.w3(32'hbbdfea00),
	.w4(32'hbb5125ef),
	.w5(32'hbc4e519c),
	.w6(32'hbb2fcf5c),
	.w7(32'h3b093cf7),
	.w8(32'hba8543f0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1461c3),
	.w1(32'hb9db9102),
	.w2(32'hb9677091),
	.w3(32'hbbc0a989),
	.w4(32'h3a5d88f9),
	.w5(32'hba968e5c),
	.w6(32'hbbaac558),
	.w7(32'hbbf1027f),
	.w8(32'hbbc7560d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf670b8),
	.w1(32'hbb05162d),
	.w2(32'h3bb42579),
	.w3(32'h3b35a70c),
	.w4(32'hbb832d65),
	.w5(32'hbbc05a71),
	.w6(32'hbba534b4),
	.w7(32'hbc0bcf27),
	.w8(32'hbb59fd16),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8375f1b),
	.w1(32'hbb8e8c18),
	.w2(32'hbbf275d6),
	.w3(32'hbb1fcf5d),
	.w4(32'hbb88d4a1),
	.w5(32'hbc129f7a),
	.w6(32'hbb84df02),
	.w7(32'hba2ecf18),
	.w8(32'hbbbccc56),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56cea),
	.w1(32'h3836ae60),
	.w2(32'h3ac050b8),
	.w3(32'hbbc1d011),
	.w4(32'hbb0f1613),
	.w5(32'h3c112e23),
	.w6(32'hbaa4c2d8),
	.w7(32'h3b067af9),
	.w8(32'h3b8ea2ce),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b38f1),
	.w1(32'hbac3cc7a),
	.w2(32'hbba9c62f),
	.w3(32'hbaba0eb3),
	.w4(32'hbab2e4b3),
	.w5(32'h3ab02525),
	.w6(32'h3ba16227),
	.w7(32'h3a529aca),
	.w8(32'h3a1e813d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42762a),
	.w1(32'h3b66494d),
	.w2(32'hbc01f914),
	.w3(32'hbbd0347a),
	.w4(32'hbb283adf),
	.w5(32'h3b426c2a),
	.w6(32'hbb7e5165),
	.w7(32'hba1f84b9),
	.w8(32'hbbb8a476),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a2ac),
	.w1(32'hbb8f9254),
	.w2(32'h3a9503d9),
	.w3(32'hbb9a500d),
	.w4(32'hbb8c27a8),
	.w5(32'hbbd91da8),
	.w6(32'h3ba08e9b),
	.w7(32'hbbafd672),
	.w8(32'hbb8e3e15),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829ebc),
	.w1(32'hbb6e16d3),
	.w2(32'hbb87e960),
	.w3(32'hbbab6202),
	.w4(32'hbc007d6a),
	.w5(32'hba99a892),
	.w6(32'hbc1aa779),
	.w7(32'hba5daf76),
	.w8(32'hbb62cb87),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998c06),
	.w1(32'h3a9a557c),
	.w2(32'hbc032c6c),
	.w3(32'hba6ef06c),
	.w4(32'h3c0f7ca3),
	.w5(32'h3c25b09b),
	.w6(32'hbae656c0),
	.w7(32'hbbac9cd6),
	.w8(32'hbc19e0bd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473fc5),
	.w1(32'h3b8aec1c),
	.w2(32'h38c4087b),
	.w3(32'hbbe7a478),
	.w4(32'hbbe98474),
	.w5(32'h3ca999c8),
	.w6(32'hbbe18d31),
	.w7(32'hbc45755f),
	.w8(32'hbc25fb3c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb064),
	.w1(32'h3b71a5b3),
	.w2(32'h39d5dac5),
	.w3(32'h3c1fbfdd),
	.w4(32'h3a08818e),
	.w5(32'h3b310daa),
	.w6(32'hbab8e3c9),
	.w7(32'h3b690608),
	.w8(32'hbb4a9882),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e9475),
	.w1(32'hba41fc1f),
	.w2(32'hbb290446),
	.w3(32'hba406172),
	.w4(32'hbacf019f),
	.w5(32'hba8e042d),
	.w6(32'hbc01d9d2),
	.w7(32'h3a044968),
	.w8(32'hbb01a73b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb234910),
	.w1(32'h3ada25eb),
	.w2(32'h39c27b33),
	.w3(32'h3ac011ba),
	.w4(32'h3b1cb538),
	.w5(32'hbb6598f9),
	.w6(32'hbb280112),
	.w7(32'h3b171d21),
	.w8(32'h3b392953),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0567fd),
	.w1(32'h3aafc38f),
	.w2(32'hbae81f43),
	.w3(32'h3b399049),
	.w4(32'h3b97cfbf),
	.w5(32'h3b4e1de2),
	.w6(32'h39c0854b),
	.w7(32'h3bacdfee),
	.w8(32'h3b012e6a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb295982),
	.w1(32'h3b1dbdd3),
	.w2(32'hbb48cff5),
	.w3(32'hbb856665),
	.w4(32'h39bddd47),
	.w5(32'h3c522fee),
	.w6(32'hba0145d9),
	.w7(32'h3940f70d),
	.w8(32'h3a02c5ba),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31b73a),
	.w1(32'hbb0a6b38),
	.w2(32'h3b450fdb),
	.w3(32'h39dc3fd5),
	.w4(32'hbbfcd087),
	.w5(32'h3a017471),
	.w6(32'hbb4fa11a),
	.w7(32'hbbee69a4),
	.w8(32'hbbdb7a81),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57691d),
	.w1(32'hbb6b0f64),
	.w2(32'h3ad09ff4),
	.w3(32'h3a82b19a),
	.w4(32'hbb0f1f11),
	.w5(32'hba9558bb),
	.w6(32'hbb8ef2e9),
	.w7(32'hbac3aa3b),
	.w8(32'h3aabb949),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2554c5),
	.w1(32'hbb8c2d93),
	.w2(32'hb9a608f5),
	.w3(32'hbb6e0554),
	.w4(32'hbb9efc9f),
	.w5(32'hbbea58df),
	.w6(32'hbbfa1e15),
	.w7(32'hbaf29364),
	.w8(32'hbb45464d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e127d),
	.w1(32'h3b13590b),
	.w2(32'h3abaf451),
	.w3(32'hbb3c77d9),
	.w4(32'h3a61d405),
	.w5(32'hbae0b1af),
	.w6(32'hbb1f8c99),
	.w7(32'h3aee929d),
	.w8(32'h3bac999f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799ff4),
	.w1(32'h3a96b881),
	.w2(32'h3ab28e2a),
	.w3(32'hbb0a132a),
	.w4(32'hbbd0a11d),
	.w5(32'hbc8d1907),
	.w6(32'hb8821908),
	.w7(32'hbb328b27),
	.w8(32'h3b907731),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842679),
	.w1(32'hba8dc2ab),
	.w2(32'hbbca59b4),
	.w3(32'h3b758ef3),
	.w4(32'h3baaeeca),
	.w5(32'hbb7df401),
	.w6(32'h3b9ac36c),
	.w7(32'h3a9d0223),
	.w8(32'h3b70a0b2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab224b),
	.w1(32'h3b5b2305),
	.w2(32'h3b8ff2ad),
	.w3(32'h3af0e41c),
	.w4(32'h38de20c1),
	.w5(32'h3b3f25c9),
	.w6(32'hbb5ac25d),
	.w7(32'hba1c362a),
	.w8(32'hb9767481),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900907),
	.w1(32'hb9b8dacb),
	.w2(32'h3b461226),
	.w3(32'h3a35c530),
	.w4(32'hba079087),
	.w5(32'hb94571f1),
	.w6(32'h3ae86a3a),
	.w7(32'h3901ea0c),
	.w8(32'h3bdce59a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f9bd4),
	.w1(32'hbace9059),
	.w2(32'hbbbe32d5),
	.w3(32'h3c2da1ae),
	.w4(32'hba3577fc),
	.w5(32'hbbd80d49),
	.w6(32'h3bc19b30),
	.w7(32'h3af57201),
	.w8(32'hbb871e97),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99a168),
	.w1(32'hba2f1c78),
	.w2(32'h3b096a7b),
	.w3(32'hbb837aa0),
	.w4(32'hba815a1a),
	.w5(32'h3b06ea5b),
	.w6(32'hbc035798),
	.w7(32'hbb914b92),
	.w8(32'h3a56e1aa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4d86),
	.w1(32'hbac3926e),
	.w2(32'hbb3d31cc),
	.w3(32'h3a6b6207),
	.w4(32'h3b63919e),
	.w5(32'hbb829a54),
	.w6(32'h3a1dafc9),
	.w7(32'hbabc0afe),
	.w8(32'h3aec6558),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad429c2),
	.w1(32'hbb8c6bd2),
	.w2(32'h3b0db248),
	.w3(32'h3a178e66),
	.w4(32'hb9c4d27e),
	.w5(32'hbac645f0),
	.w6(32'h3b689b78),
	.w7(32'hbbb0c154),
	.w8(32'h3b53cee7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121e31),
	.w1(32'hbb9a32f1),
	.w2(32'hba1eb710),
	.w3(32'hba02decf),
	.w4(32'h3b9be854),
	.w5(32'h3b60dff6),
	.w6(32'h3ae9b25c),
	.w7(32'h370a2db4),
	.w8(32'h3a291382),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a257c),
	.w1(32'h3b64ebaa),
	.w2(32'hbaf45be2),
	.w3(32'h3ad747e5),
	.w4(32'h3b84143c),
	.w5(32'h3b051743),
	.w6(32'hbb1f8e0d),
	.w7(32'h3a0394e5),
	.w8(32'hbb2a4374),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39559ea1),
	.w1(32'h3a74050d),
	.w2(32'h3b1e1357),
	.w3(32'h3b200be0),
	.w4(32'h3970504a),
	.w5(32'hbb4e4419),
	.w6(32'h3b6780fe),
	.w7(32'hb9c09b0d),
	.w8(32'hbb1e1291),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00659f),
	.w1(32'h3bdec79f),
	.w2(32'h3bdf5da0),
	.w3(32'h39e1a00e),
	.w4(32'hba411c5b),
	.w5(32'h3c04b409),
	.w6(32'h3b62f9fe),
	.w7(32'hbb179db0),
	.w8(32'hba5731df),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c8677),
	.w1(32'h3a823cd4),
	.w2(32'hbaea1f7b),
	.w3(32'h3bf50725),
	.w4(32'hbb52535b),
	.w5(32'hbc005f9a),
	.w6(32'h3a769197),
	.w7(32'hbbb21f3c),
	.w8(32'hbbcd2880),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba105b0d),
	.w1(32'hbad0e484),
	.w2(32'hbc1f4001),
	.w3(32'hbbe00856),
	.w4(32'hbbb17184),
	.w5(32'hbbd90d29),
	.w6(32'hbbfe996f),
	.w7(32'hbb94f165),
	.w8(32'hbbb2483c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc305d41),
	.w1(32'hbaf9be2f),
	.w2(32'hbaa11fdb),
	.w3(32'hbc2b81d0),
	.w4(32'h3bbdbefb),
	.w5(32'hb95fbd72),
	.w6(32'hbc03ff54),
	.w7(32'h3b7d731b),
	.w8(32'hba175093),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36eccc),
	.w1(32'hbadb067a),
	.w2(32'hba4214b4),
	.w3(32'hbaa0d6b8),
	.w4(32'hbb6f7176),
	.w5(32'hbbabe4b0),
	.w6(32'h39bc1a94),
	.w7(32'hbb7f859e),
	.w8(32'hbbe3256f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4037e5),
	.w1(32'h3ad8a211),
	.w2(32'h3a975972),
	.w3(32'hbb44231b),
	.w4(32'hbb26e545),
	.w5(32'h3b0f0f99),
	.w6(32'hbbeac78d),
	.w7(32'hbae39e18),
	.w8(32'h3b8bd11c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f2dc),
	.w1(32'hbb7bd5a1),
	.w2(32'hbaa313aa),
	.w3(32'h3c24b8bd),
	.w4(32'hbaa34175),
	.w5(32'h3b736830),
	.w6(32'hb8130d80),
	.w7(32'hbbcaf29c),
	.w8(32'h39008c22),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be66830),
	.w1(32'hba2f8a2e),
	.w2(32'hba583f35),
	.w3(32'hbb498aca),
	.w4(32'hbaab245b),
	.w5(32'hbae63fcd),
	.w6(32'hb9b5c266),
	.w7(32'hba3515d6),
	.w8(32'h3b260c9c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1e7f),
	.w1(32'hba8aa300),
	.w2(32'hbb8ca930),
	.w3(32'h3b410891),
	.w4(32'hbb288ee8),
	.w5(32'h3b5e1dd7),
	.w6(32'h3bb5c0de),
	.w7(32'hbb265ba7),
	.w8(32'hbb8a67b2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb484443),
	.w1(32'h3b480b57),
	.w2(32'h38509734),
	.w3(32'hbad283db),
	.w4(32'h3a8373a1),
	.w5(32'hbc02ef56),
	.w6(32'hbb245d3f),
	.w7(32'h3b3b0002),
	.w8(32'hb8632a70),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86861e),
	.w1(32'h3bb50ff9),
	.w2(32'h3c34caaf),
	.w3(32'hbb5b0f41),
	.w4(32'hbab580ad),
	.w5(32'h3afdfcf1),
	.w6(32'hbbe138af),
	.w7(32'hba1c8e71),
	.w8(32'hbb25ccc8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9aeee),
	.w1(32'hbb836657),
	.w2(32'hbafc3e92),
	.w3(32'h39b9d553),
	.w4(32'hb9fddfa5),
	.w5(32'hbc2e4e9b),
	.w6(32'h3b635482),
	.w7(32'h36fec967),
	.w8(32'hbb44e284),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1a6f8),
	.w1(32'h3abef00c),
	.w2(32'hbbfe6cfc),
	.w3(32'hbb335ff6),
	.w4(32'hba9caa69),
	.w5(32'h3b41cb20),
	.w6(32'hbb3f21f3),
	.w7(32'h3b89f009),
	.w8(32'h3b889fec),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46e846),
	.w1(32'h3bcbaca1),
	.w2(32'h3a83a4cf),
	.w3(32'h3bad334f),
	.w4(32'h39f431cf),
	.w5(32'hba076cf4),
	.w6(32'h3bbfabf4),
	.w7(32'hbac5d4a9),
	.w8(32'hbbcd6210),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a9898),
	.w1(32'h3bc44355),
	.w2(32'h3bcf58fd),
	.w3(32'hbb5a13a9),
	.w4(32'hbbb7ecdb),
	.w5(32'h3ae47e2e),
	.w6(32'hbc19bc6a),
	.w7(32'hbb125676),
	.w8(32'hbbc17fbd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5d2c6),
	.w1(32'hbaad0601),
	.w2(32'h3a896e33),
	.w3(32'h3b8f0453),
	.w4(32'h3aa43e2f),
	.w5(32'hbb3e5083),
	.w6(32'hbb53e2ca),
	.w7(32'hba7d5f29),
	.w8(32'hbb8a7129),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad528e4),
	.w1(32'hbb84261b),
	.w2(32'h3b0a0d18),
	.w3(32'hb98525b9),
	.w4(32'hbba31f96),
	.w5(32'hbb8d065e),
	.w6(32'hbb016c97),
	.w7(32'hbb53f2d4),
	.w8(32'hbad1a64d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37c9d2),
	.w1(32'h39caff36),
	.w2(32'hbb43abdb),
	.w3(32'hba251cfd),
	.w4(32'h3b1d9c0f),
	.w5(32'h3d1a2f82),
	.w6(32'hbb51ad09),
	.w7(32'hbb85a591),
	.w8(32'hbbca2b07),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974e145),
	.w1(32'h3bc3a5ca),
	.w2(32'h3bc4eb9a),
	.w3(32'h3c560c9f),
	.w4(32'h3b9fa86c),
	.w5(32'h3c1ee4ce),
	.w6(32'hb9799e50),
	.w7(32'h3b66b61d),
	.w8(32'h3be20507),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b316c49),
	.w1(32'hb976a471),
	.w2(32'h3b800fc4),
	.w3(32'h3bec8142),
	.w4(32'h3b6d7f98),
	.w5(32'h3b81421d),
	.w6(32'h3b9cb491),
	.w7(32'hb9ff2a5a),
	.w8(32'h3b80051f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6cd23),
	.w1(32'h3bf8756a),
	.w2(32'h3c63a4a9),
	.w3(32'h3b8f2594),
	.w4(32'h3979958f),
	.w5(32'h3b8f6eb9),
	.w6(32'h3bee53fa),
	.w7(32'hba4e992a),
	.w8(32'hbb2ea6fc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2edb11),
	.w1(32'h3b9e44b7),
	.w2(32'hba143c32),
	.w3(32'h3c51380c),
	.w4(32'h3b5b0958),
	.w5(32'hbbb23ca9),
	.w6(32'hb99d4d7f),
	.w7(32'hbb82033a),
	.w8(32'h3b576b1e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917bc77),
	.w1(32'hba2d5ee1),
	.w2(32'h3b9397f9),
	.w3(32'hbba13c2b),
	.w4(32'hbbddfe1e),
	.w5(32'hbbbb91ac),
	.w6(32'hb9d27274),
	.w7(32'hbb0982a9),
	.w8(32'hbb901a73),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f04b0),
	.w1(32'hbb452102),
	.w2(32'hbaf31d36),
	.w3(32'h3bd4d818),
	.w4(32'hbb63917d),
	.w5(32'hb9484a7e),
	.w6(32'h3af9826e),
	.w7(32'h3a4e21e3),
	.w8(32'hbc190c2d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc199922),
	.w1(32'h3b025a56),
	.w2(32'hbaa934a0),
	.w3(32'hbbb4fdd4),
	.w4(32'h3a86ede1),
	.w5(32'hbb51c287),
	.w6(32'hbb202d7a),
	.w7(32'h3ae891f3),
	.w8(32'hbbc4b8e2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e9b29),
	.w1(32'h3ae05dbf),
	.w2(32'h38517a72),
	.w3(32'h3b97e956),
	.w4(32'hbb5abe3c),
	.w5(32'h3a7e7ef4),
	.w6(32'hbb8d430f),
	.w7(32'h3b7b1f9d),
	.w8(32'h3b1fd5ff),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb505b),
	.w1(32'h399ccd4d),
	.w2(32'hb9907d52),
	.w3(32'hbb92a26b),
	.w4(32'h3a69c4be),
	.w5(32'hbb417d09),
	.w6(32'hb974cad4),
	.w7(32'hba89eeb9),
	.w8(32'hbb343ad7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f1253),
	.w1(32'hba5661e9),
	.w2(32'hbabb8a81),
	.w3(32'h3aa62307),
	.w4(32'h3a871130),
	.w5(32'hbaa83615),
	.w6(32'hb99d29a9),
	.w7(32'h39b3789c),
	.w8(32'hbaa2a773),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7984ff),
	.w1(32'h3be62b6b),
	.w2(32'h3ba1dc01),
	.w3(32'h39398cbc),
	.w4(32'h3b0e64f6),
	.w5(32'h3c4b3be5),
	.w6(32'hbade8970),
	.w7(32'h3b505135),
	.w8(32'h3af54d60),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb78a08),
	.w1(32'h3a6656d4),
	.w2(32'hbbb87d40),
	.w3(32'h387239b0),
	.w4(32'h3be9203a),
	.w5(32'h3b159339),
	.w6(32'h3b465f0b),
	.w7(32'h3bc7822c),
	.w8(32'h3c22f926),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862131),
	.w1(32'hbbbbd191),
	.w2(32'hbb304624),
	.w3(32'hbaccd881),
	.w4(32'h3b7c6272),
	.w5(32'hbb98b982),
	.w6(32'h3ba9e5d9),
	.w7(32'h3b5a764a),
	.w8(32'hbb5d79d8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9d2f5),
	.w1(32'h3afa9e47),
	.w2(32'hb6bdb783),
	.w3(32'hbbb1e11c),
	.w4(32'h3b0551ef),
	.w5(32'hbb1c6079),
	.w6(32'h392c9997),
	.w7(32'h3b8c7d15),
	.w8(32'h3b55ce47),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a517e9c),
	.w1(32'hba9c02df),
	.w2(32'hbbf3e3f5),
	.w3(32'hb92ca483),
	.w4(32'h3b8d0a7c),
	.w5(32'hbb246fa7),
	.w6(32'hbb25ee79),
	.w7(32'h3b23360d),
	.w8(32'h39032a07),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb263a),
	.w1(32'hbbd581ec),
	.w2(32'hbbb616fc),
	.w3(32'hbbab8851),
	.w4(32'h3a94e651),
	.w5(32'hbba454c7),
	.w6(32'hbb53a598),
	.w7(32'h3b63c6e6),
	.w8(32'hba668724),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdfbe1),
	.w1(32'h3ba379fb),
	.w2(32'h3a0bb587),
	.w3(32'hbb3951e6),
	.w4(32'hbacc8bb3),
	.w5(32'h3a73fb39),
	.w6(32'hbad78fc7),
	.w7(32'h3a084114),
	.w8(32'h3b041b0d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345b6a),
	.w1(32'hbbe099d0),
	.w2(32'hbb9109ba),
	.w3(32'h3b4c6bf4),
	.w4(32'hbada2d5d),
	.w5(32'hba2b096b),
	.w6(32'hbac378e6),
	.w7(32'h3a5f73b0),
	.w8(32'h3b841f66),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976007),
	.w1(32'h39839bf7),
	.w2(32'hb9ce8250),
	.w3(32'hbac99762),
	.w4(32'h3a8eedcb),
	.w5(32'h3cac55b4),
	.w6(32'h3a763436),
	.w7(32'hbb7384ec),
	.w8(32'hbc5f29cc),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c405f7),
	.w1(32'h38022c59),
	.w2(32'hbad60dfa),
	.w3(32'h3a6f0905),
	.w4(32'hbab8786d),
	.w5(32'hbb5f27d6),
	.w6(32'hbb71564d),
	.w7(32'h3b8ec796),
	.w8(32'hbb5d6fa4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b6720),
	.w1(32'h3bbe9e12),
	.w2(32'h3bf5bba7),
	.w3(32'hbbb39f61),
	.w4(32'hbbd89fb6),
	.w5(32'h3be59b76),
	.w6(32'hbbc37d87),
	.w7(32'h3bc22613),
	.w8(32'h3b09ecf8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f16f9),
	.w1(32'h3be2b050),
	.w2(32'h3aec7e2a),
	.w3(32'hbb12eed5),
	.w4(32'h3b06b3ad),
	.w5(32'hbb8bba6a),
	.w6(32'h3af9bc31),
	.w7(32'h3b3ac0e1),
	.w8(32'hbaae70d1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928348),
	.w1(32'h399f2b3f),
	.w2(32'h3b38a7e1),
	.w3(32'h3c054549),
	.w4(32'h3ba1a817),
	.w5(32'h3c1f4fa6),
	.w6(32'h3ad5958b),
	.w7(32'h3bc2de3c),
	.w8(32'h3a871bb9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62914f),
	.w1(32'hbabaa520),
	.w2(32'h3b62a548),
	.w3(32'h3c732543),
	.w4(32'hbb18a251),
	.w5(32'h3b906ffa),
	.w6(32'h3c520293),
	.w7(32'hbb5bf563),
	.w8(32'h3af5f3eb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6cb8ab),
	.w1(32'hbafdd8f0),
	.w2(32'h39b327d2),
	.w3(32'h3c19fdc7),
	.w4(32'hbc0f3ebf),
	.w5(32'hbba000e5),
	.w6(32'hba2634fb),
	.w7(32'hbbe46b44),
	.w8(32'hbbeacb3a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab511ad),
	.w1(32'hb99c1e3d),
	.w2(32'hbb6768a4),
	.w3(32'h3a44d5fc),
	.w4(32'h3abe4322),
	.w5(32'h3b62b17f),
	.w6(32'hbbe83aef),
	.w7(32'hb93c66ec),
	.w8(32'hba21bd41),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb518250),
	.w1(32'hbc160137),
	.w2(32'hbc6e9c9c),
	.w3(32'h3b11c459),
	.w4(32'h3c3afe21),
	.w5(32'h3c70b266),
	.w6(32'hbb6c3a5d),
	.w7(32'hbc47a77d),
	.w8(32'hbaaf27ec),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a676c),
	.w1(32'hbbc61e0b),
	.w2(32'hbc14031a),
	.w3(32'hbbecdc54),
	.w4(32'hbaa545a3),
	.w5(32'hbb0031b7),
	.w6(32'h3beb3f04),
	.w7(32'hbb10c164),
	.w8(32'hbb175460),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178d31),
	.w1(32'hbb3b48d4),
	.w2(32'hb9b43839),
	.w3(32'hbb8ae538),
	.w4(32'hbb93d9a7),
	.w5(32'hbbd5acd0),
	.w6(32'h3aa05316),
	.w7(32'hbae64f20),
	.w8(32'hba961775),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe140f6),
	.w1(32'hbb4a1c1a),
	.w2(32'h3aeedad4),
	.w3(32'hbb857ea8),
	.w4(32'hbb284bf6),
	.w5(32'hbb514a11),
	.w6(32'hb883f855),
	.w7(32'hbb615805),
	.w8(32'h3ad29032),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45155e),
	.w1(32'h3b7684cd),
	.w2(32'h3ac8d778),
	.w3(32'h3b058933),
	.w4(32'h3b909229),
	.w5(32'h3b5cea31),
	.w6(32'h394647e3),
	.w7(32'h3a940282),
	.w8(32'h3b8cb29c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57e3da),
	.w1(32'hbaaf323a),
	.w2(32'hbb90dd6b),
	.w3(32'hbb68630b),
	.w4(32'h3aee44cd),
	.w5(32'hbb8298b8),
	.w6(32'h3ab74bd7),
	.w7(32'hb9810fcd),
	.w8(32'hbad193a0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cc9e4),
	.w1(32'h39f18227),
	.w2(32'hbbb30f5f),
	.w3(32'hbb762741),
	.w4(32'hbaa1f50d),
	.w5(32'hbbbdce6d),
	.w6(32'h384553ba),
	.w7(32'hbb4f59a8),
	.w8(32'hbbce7cd8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac38fa3),
	.w1(32'h3ab2b643),
	.w2(32'h3a945cfa),
	.w3(32'hbb843897),
	.w4(32'hbb865afb),
	.w5(32'hbb03dd5d),
	.w6(32'hbbbeac62),
	.w7(32'h3abfceaa),
	.w8(32'h3a467eaf),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2fad8),
	.w1(32'h3999f177),
	.w2(32'hbacde8ee),
	.w3(32'h3afa6304),
	.w4(32'h3bcb17d6),
	.w5(32'h3ba50a62),
	.w6(32'hba971c04),
	.w7(32'h3b215c7e),
	.w8(32'hbc030ca5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2307ac),
	.w1(32'hbb84bebb),
	.w2(32'hbb95bf12),
	.w3(32'h3ba2371f),
	.w4(32'h3b0774e6),
	.w5(32'hbc0c3bbb),
	.w6(32'hbb2a2b5e),
	.w7(32'hbbd516a4),
	.w8(32'hbb983b13),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a0b6f),
	.w1(32'h3b5b791b),
	.w2(32'hbaca9cbe),
	.w3(32'hbb600269),
	.w4(32'h3a151032),
	.w5(32'h3aadb346),
	.w6(32'h3a54ec16),
	.w7(32'hbb2ac451),
	.w8(32'h3b856eeb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874a18),
	.w1(32'h3b1450cc),
	.w2(32'h3b7fdd31),
	.w3(32'hbb079c80),
	.w4(32'hbb9645d0),
	.w5(32'h3b8c7bcc),
	.w6(32'hbb938fbd),
	.w7(32'hbabdfc25),
	.w8(32'hbb21d6dc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4e31),
	.w1(32'hbb035426),
	.w2(32'h39088462),
	.w3(32'h3b8b8bde),
	.w4(32'h3ab6747c),
	.w5(32'hbaab0425),
	.w6(32'h3babe081),
	.w7(32'h3abc2f80),
	.w8(32'h3a938292),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67a3cd),
	.w1(32'h3bc1dfae),
	.w2(32'h3b8f07ea),
	.w3(32'h389d6861),
	.w4(32'h3b651899),
	.w5(32'h3c0a8a44),
	.w6(32'h3b7bcde3),
	.w7(32'h3c0b1a4e),
	.w8(32'h3b95d063),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94529d6),
	.w1(32'h3a4572cd),
	.w2(32'hba0b7824),
	.w3(32'h3b221a99),
	.w4(32'h3ab4f00b),
	.w5(32'h3b9a863d),
	.w6(32'hbac5048f),
	.w7(32'hba9c7bf1),
	.w8(32'hb7e1dce7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d6f6c),
	.w1(32'h3ac863a9),
	.w2(32'hbb802f8d),
	.w3(32'hbb9b09b3),
	.w4(32'hbbc13418),
	.w5(32'h3c6afb76),
	.w6(32'hbb93ac40),
	.w7(32'h3a7b53b5),
	.w8(32'h38d26386),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9076ae),
	.w1(32'hbb918ca6),
	.w2(32'hbb4ab331),
	.w3(32'hba4751db),
	.w4(32'hbb069658),
	.w5(32'hbb89138e),
	.w6(32'hbb84b157),
	.w7(32'hb98b29cb),
	.w8(32'hbb4477e7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34f4f8),
	.w1(32'hb9ee9cc2),
	.w2(32'hbb797fe5),
	.w3(32'hbae4d6d3),
	.w4(32'hbbb2eb66),
	.w5(32'hbbcc18d5),
	.w6(32'hbba19532),
	.w7(32'hbbca220e),
	.w8(32'hbb0e356c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36b855),
	.w1(32'hbb85672f),
	.w2(32'hbb9daa17),
	.w3(32'hbbe0f55e),
	.w4(32'hbb7c9ed1),
	.w5(32'hbba35dfb),
	.w6(32'hba842596),
	.w7(32'hbaa9945c),
	.w8(32'hbb7ed05a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8830d7),
	.w1(32'h3c299acb),
	.w2(32'hba9de9e6),
	.w3(32'hbbd09aeb),
	.w4(32'h3b293d4f),
	.w5(32'h3bd7d6c3),
	.w6(32'hbb7f2356),
	.w7(32'hbac69771),
	.w8(32'hbc193426),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c2ecc),
	.w1(32'hbb92595a),
	.w2(32'hbbdec778),
	.w3(32'h3b34fbd9),
	.w4(32'h3a4102b0),
	.w5(32'hbb4ffe4a),
	.w6(32'h3b0966ad),
	.w7(32'h3a99735b),
	.w8(32'h3bc0772e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc368dc2),
	.w1(32'h3a826ef8),
	.w2(32'hba41e862),
	.w3(32'hbc08e253),
	.w4(32'h3b1008f1),
	.w5(32'h3a8ae683),
	.w6(32'hbbae5257),
	.w7(32'h3b0a3064),
	.w8(32'h3b274c04),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2875db),
	.w1(32'hb8b25a42),
	.w2(32'hba63f5f7),
	.w3(32'h3b0317b7),
	.w4(32'hb95053d1),
	.w5(32'hbae95b6c),
	.w6(32'h3a2f79fd),
	.w7(32'hbbcc888f),
	.w8(32'h3aa9408b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46a54),
	.w1(32'h3b176c56),
	.w2(32'hbad23145),
	.w3(32'hba7ae045),
	.w4(32'hbad7ab5a),
	.w5(32'h39a1a1fa),
	.w6(32'h3ac96aa5),
	.w7(32'h3a5e2786),
	.w8(32'hbb3f5f68),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dafd6),
	.w1(32'h3b6abc88),
	.w2(32'h3af84108),
	.w3(32'hbb5dbd07),
	.w4(32'hba9ed53d),
	.w5(32'h3b35bcaf),
	.w6(32'hbb9346f3),
	.w7(32'hbb82dd9e),
	.w8(32'hbb5d59fe),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fb251),
	.w1(32'h3b874679),
	.w2(32'h3bea225c),
	.w3(32'h3b8ecb03),
	.w4(32'hba9531d8),
	.w5(32'hbb2be613),
	.w6(32'hba6db100),
	.w7(32'h3a5d61f3),
	.w8(32'hbb5ea021),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba880bfd),
	.w1(32'hba5b3c54),
	.w2(32'h3aedfc84),
	.w3(32'hb9d25628),
	.w4(32'hb85172e2),
	.w5(32'h3b9c6285),
	.w6(32'hbb8f2205),
	.w7(32'hbbe251bb),
	.w8(32'hbada83ff),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b941a26),
	.w1(32'hbb4c4a08),
	.w2(32'hbc07e0c8),
	.w3(32'h3b53579f),
	.w4(32'hbb976f9f),
	.w5(32'hbbc62c5a),
	.w6(32'hb9e248e0),
	.w7(32'hbae973f5),
	.w8(32'hb878af13),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe97f7c),
	.w1(32'hbb9daf6c),
	.w2(32'hbb9370d0),
	.w3(32'hbbf9a082),
	.w4(32'hbc101401),
	.w5(32'hbaef671f),
	.w6(32'hbb2cdac3),
	.w7(32'hbb58b198),
	.w8(32'h3ae28f9d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab23c9c),
	.w1(32'hbb0b03ce),
	.w2(32'hb9e573c7),
	.w3(32'hbbb5e591),
	.w4(32'hbb2f05cd),
	.w5(32'hbae47b10),
	.w6(32'hbbaf0af2),
	.w7(32'hbb0ec7fc),
	.w8(32'hbb0e85ab),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06c478),
	.w1(32'hba031d98),
	.w2(32'hba5b2e0b),
	.w3(32'hba6aa372),
	.w4(32'hba0b66c7),
	.w5(32'hba272a6f),
	.w6(32'hba92d750),
	.w7(32'hba6d949d),
	.w8(32'hbab4aa43),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c6e82),
	.w1(32'hb9f26e50),
	.w2(32'hba747502),
	.w3(32'hba87dba1),
	.w4(32'hba9124fe),
	.w5(32'hba6a39a0),
	.w6(32'hba9b7470),
	.w7(32'hba023984),
	.w8(32'hbaa0d066),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba570cb6),
	.w1(32'h38c39896),
	.w2(32'h398220ae),
	.w3(32'hb9b4741e),
	.w4(32'hb9a7ef96),
	.w5(32'hb88e64f8),
	.w6(32'hba388121),
	.w7(32'hba1fc901),
	.w8(32'hba200e8c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f35a0c),
	.w1(32'h39f35a5e),
	.w2(32'h39bc5b8b),
	.w3(32'h39a1255e),
	.w4(32'hb9a3ea75),
	.w5(32'h382e89e8),
	.w6(32'h3a203a7e),
	.w7(32'hb99a878a),
	.w8(32'h3918656b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1e2bb),
	.w1(32'hb9d6c798),
	.w2(32'h39f7c6fc),
	.w3(32'hba0534d4),
	.w4(32'h39c58be4),
	.w5(32'h3a8bbf05),
	.w6(32'hb731c4a6),
	.w7(32'hb970dfc7),
	.w8(32'h3973a693),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399af5d5),
	.w1(32'h3a30b633),
	.w2(32'h39c3d848),
	.w3(32'h3a5ebf27),
	.w4(32'h3a2d4df0),
	.w5(32'h3a012f26),
	.w6(32'h3aaef0f5),
	.w7(32'h3a2d3064),
	.w8(32'h3a5fa738),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f414),
	.w1(32'h3a9b5d1d),
	.w2(32'h3aa5b353),
	.w3(32'hb92407dd),
	.w4(32'h3a396176),
	.w5(32'h3a185cfe),
	.w6(32'h398dd44c),
	.w7(32'h3a54cdd2),
	.w8(32'h3a73d304),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d32292),
	.w1(32'h395f61a2),
	.w2(32'hba032312),
	.w3(32'h39274c00),
	.w4(32'hb7e8b13b),
	.w5(32'hb99d4900),
	.w6(32'h37c66734),
	.w7(32'hb9c95671),
	.w8(32'hba580660),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3e8cd),
	.w1(32'h3a6aa133),
	.w2(32'h3a294b1d),
	.w3(32'hba8c13ec),
	.w4(32'h3a573024),
	.w5(32'h3a016029),
	.w6(32'hba26f065),
	.w7(32'h39fc53a3),
	.w8(32'h3a07f1eb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b128b),
	.w1(32'hb9eeea66),
	.w2(32'hba4a7729),
	.w3(32'h3a75088a),
	.w4(32'hba96f3e8),
	.w5(32'hba319fa5),
	.w6(32'h3a516171),
	.w7(32'hba954eeb),
	.w8(32'hba4a4fb9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbc82a),
	.w1(32'h3b25ce1a),
	.w2(32'h3b45f6fd),
	.w3(32'hbab1f469),
	.w4(32'h3b0ff0af),
	.w5(32'h3b482451),
	.w6(32'hba926bcc),
	.w7(32'h3b1c3ec1),
	.w8(32'h3b2d6619),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b224a24),
	.w1(32'h3a02c2f5),
	.w2(32'h3a153ec2),
	.w3(32'h3b1ea73a),
	.w4(32'h3a181326),
	.w5(32'h3a10b6e7),
	.w6(32'h3b000f74),
	.w7(32'h399eef46),
	.w8(32'h39212b5a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fbf16),
	.w1(32'hb9cbe541),
	.w2(32'h38dc27e7),
	.w3(32'h392d3238),
	.w4(32'hb9d6f323),
	.w5(32'hba3ca97f),
	.w6(32'h37e0968b),
	.w7(32'hba02aee0),
	.w8(32'hb969c6e5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919effa),
	.w1(32'hb9c6a0a3),
	.w2(32'h3a3e6844),
	.w3(32'hbad012af),
	.w4(32'h3ac85376),
	.w5(32'h3b2734c0),
	.w6(32'hba1c27a3),
	.w7(32'h3a1fe8af),
	.w8(32'h3a972eb2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fcd5f),
	.w1(32'h3a9826e5),
	.w2(32'h3aad7a33),
	.w3(32'h3a571416),
	.w4(32'h3a647afb),
	.w5(32'h3abc47ca),
	.w6(32'h3a922365),
	.w7(32'h3a99b4b5),
	.w8(32'h3a87f6df),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c4a74),
	.w1(32'hba64f4ff),
	.w2(32'hbac7f4df),
	.w3(32'h39e59cb1),
	.w4(32'hba3edb36),
	.w5(32'hbacd7bfd),
	.w6(32'h3a4c1314),
	.w7(32'hb9d8ef82),
	.w8(32'hba627684),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac94642),
	.w1(32'h39148913),
	.w2(32'hb8adcba0),
	.w3(32'hba0130b5),
	.w4(32'h3904b733),
	.w5(32'h393adfa4),
	.w6(32'hb93f5082),
	.w7(32'h3a170204),
	.w8(32'hba10dd88),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df12bd),
	.w1(32'h39b62222),
	.w2(32'h3937ffa9),
	.w3(32'hba022a1a),
	.w4(32'hb995d154),
	.w5(32'h39b195f9),
	.w6(32'hba0ce842),
	.w7(32'hb9adfc38),
	.w8(32'hb8c9a15e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee9166),
	.w1(32'hb98793c7),
	.w2(32'h3a246b8d),
	.w3(32'hb9f4a353),
	.w4(32'h3a799882),
	.w5(32'h3aea88f0),
	.w6(32'hb9a6a05f),
	.w7(32'h3a39f24d),
	.w8(32'h3a7f2eaa),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57efbd),
	.w1(32'hbabcad27),
	.w2(32'h3953aa75),
	.w3(32'h3a106f78),
	.w4(32'hbacfc1c1),
	.w5(32'h39cc4681),
	.w6(32'h39de30a9),
	.w7(32'hbacc1a0c),
	.w8(32'hb9628fbf),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac49071),
	.w1(32'hbb369c64),
	.w2(32'hbad97333),
	.w3(32'hba1356a8),
	.w4(32'hbb3cc69d),
	.w5(32'hbb22070c),
	.w6(32'hba0c45aa),
	.w7(32'hbb30f50c),
	.w8(32'hbb4587b9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb282fff),
	.w1(32'h38dc32d3),
	.w2(32'h37fde472),
	.w3(32'hbb5b3683),
	.w4(32'h398f45e5),
	.w5(32'h390cfe4a),
	.w6(32'hbb4e4cd0),
	.w7(32'hba02278e),
	.w8(32'hb9ad6061),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dcc79),
	.w1(32'h3a6a6ab9),
	.w2(32'h3ac9a2d5),
	.w3(32'h39d43fc5),
	.w4(32'h39af3cc1),
	.w5(32'h39f133c3),
	.w6(32'h388d0d5c),
	.w7(32'h3a8611dc),
	.w8(32'h3aaa42ed),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac93ea),
	.w1(32'h378b439e),
	.w2(32'h3a433189),
	.w3(32'hb8c6503e),
	.w4(32'hba137ed4),
	.w5(32'h39b426db),
	.w6(32'h3a0b5b68),
	.w7(32'hb8ea962d),
	.w8(32'h3a8b92ca),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c640ce),
	.w1(32'h38c2d6e3),
	.w2(32'hb910419e),
	.w3(32'h39402a5a),
	.w4(32'h3a4e575a),
	.w5(32'h3a0b0633),
	.w6(32'h39384437),
	.w7(32'hba2e77aa),
	.w8(32'h391672a4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a008073),
	.w1(32'h38ac0fd0),
	.w2(32'hb96ad90a),
	.w3(32'h3a805f2a),
	.w4(32'hba1a21ed),
	.w5(32'hba45297e),
	.w6(32'h3ac35f1e),
	.w7(32'h3899c63d),
	.w8(32'hba62fa4b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b79ab),
	.w1(32'h397f0c74),
	.w2(32'hb9ec4ae7),
	.w3(32'hb8b6c7a7),
	.w4(32'h3835f250),
	.w5(32'hb9985f38),
	.w6(32'hba64664b),
	.w7(32'hba2c0fcc),
	.w8(32'hba327264),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9854766),
	.w1(32'hba7cb1bd),
	.w2(32'hb7a7994e),
	.w3(32'hb979dde3),
	.w4(32'hba678a11),
	.w5(32'h38fa1663),
	.w6(32'h38b7c083),
	.w7(32'hba84796a),
	.w8(32'hba442530),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47c5ec),
	.w1(32'hba8b3fe9),
	.w2(32'hba289afe),
	.w3(32'h38a5ad19),
	.w4(32'hb9d4e35e),
	.w5(32'hba011503),
	.w6(32'hb754c51b),
	.w7(32'hba927129),
	.w8(32'hba984ffd),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0600fe),
	.w1(32'hb9d0bd9d),
	.w2(32'h39f0165a),
	.w3(32'hbaf2f7ae),
	.w4(32'h390a54c4),
	.w5(32'h3a016f14),
	.w6(32'hbb0f1791),
	.w7(32'h3793ce21),
	.w8(32'h35d374cc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a565894),
	.w1(32'hb96b7cab),
	.w2(32'hba1b416a),
	.w3(32'h39d0fe20),
	.w4(32'hba117199),
	.w5(32'hb94edc4c),
	.w6(32'h3a68f714),
	.w7(32'hba3cb09b),
	.w8(32'hb9ce6454),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d76be8),
	.w1(32'h3a8b858f),
	.w2(32'hb848bc21),
	.w3(32'hb9a82df9),
	.w4(32'h3a168672),
	.w5(32'hba483466),
	.w6(32'hb9722466),
	.w7(32'h3aa42f0e),
	.w8(32'hb9b369ea),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff8346),
	.w1(32'hba9b0b50),
	.w2(32'hba7ec127),
	.w3(32'hba39e737),
	.w4(32'hb983ff38),
	.w5(32'hb9e80335),
	.w6(32'hba1223d0),
	.w7(32'hba6aa346),
	.w8(32'hba93b703),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae448c5),
	.w1(32'h3ac9c490),
	.w2(32'h3aaa8c37),
	.w3(32'hbb05e288),
	.w4(32'h3aa52b65),
	.w5(32'h3abfec6d),
	.w6(32'hbac1b24f),
	.w7(32'h3abcc723),
	.w8(32'h3ac7be8a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a970ad3),
	.w1(32'hba14d9cc),
	.w2(32'h38f8fadd),
	.w3(32'h3a9dcf73),
	.w4(32'hb9cb8249),
	.w5(32'h38e3d859),
	.w6(32'h3aef6e6e),
	.w7(32'hba1099f9),
	.w8(32'h3907ced7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d09d9),
	.w1(32'h39988b2e),
	.w2(32'h3a6000a4),
	.w3(32'hba9d10db),
	.w4(32'h3a15fd96),
	.w5(32'h3a2c9d11),
	.w6(32'hba80d224),
	.w7(32'h3814279b),
	.w8(32'h39206734),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4af1b9),
	.w1(32'h38471327),
	.w2(32'h3942cce2),
	.w3(32'h3a329b90),
	.w4(32'h38e82763),
	.w5(32'hb93c22e2),
	.w6(32'h39cddf37),
	.w7(32'h389061ad),
	.w8(32'h39c13dec),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9807588),
	.w1(32'hba4abf67),
	.w2(32'hb9e89539),
	.w3(32'hb9e4f475),
	.w4(32'hba5c1ca8),
	.w5(32'hb9f74388),
	.w6(32'hb90161d2),
	.w7(32'hb9698b25),
	.w8(32'h384cb758),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93cd9b),
	.w1(32'h39ad39ed),
	.w2(32'h39ae9db0),
	.w3(32'hbac141ea),
	.w4(32'hb9482b04),
	.w5(32'hb8daf37d),
	.w6(32'hba9573dc),
	.w7(32'hb9b72a8d),
	.w8(32'hb986989b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f0054),
	.w1(32'hba1a24be),
	.w2(32'h38731c0a),
	.w3(32'hba56aa05),
	.w4(32'hba8f2190),
	.w5(32'hba9a379b),
	.w6(32'hba00b3ad),
	.w7(32'h3986aaaf),
	.w8(32'hb99c4b40),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9565088),
	.w1(32'h392e8989),
	.w2(32'h3943d49f),
	.w3(32'hba8de5d7),
	.w4(32'hb9e13003),
	.w5(32'h39a67497),
	.w6(32'hba1883f9),
	.w7(32'hba98dfb8),
	.w8(32'hb956d36e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d2e26),
	.w1(32'hba285b1c),
	.w2(32'hba4c5225),
	.w3(32'h39c26acc),
	.w4(32'hbabe4fd1),
	.w5(32'hb9b10fe2),
	.w6(32'h387f79fc),
	.w7(32'hba5d8fb4),
	.w8(32'hba69f7f8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a14ad6),
	.w1(32'h3978e008),
	.w2(32'h39c6b739),
	.w3(32'hb7f072b5),
	.w4(32'hb9618925),
	.w5(32'h396820de),
	.w6(32'hb835c600),
	.w7(32'hb9cf00c1),
	.w8(32'hba159e48),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33063e),
	.w1(32'h39d91407),
	.w2(32'hb9f576ab),
	.w3(32'hba6e5602),
	.w4(32'hb955cf06),
	.w5(32'hba32dc98),
	.w6(32'hbaa0fdd0),
	.w7(32'hb9ac7315),
	.w8(32'hb9bf4902),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d3277),
	.w1(32'hb8de3d32),
	.w2(32'h383e1cb1),
	.w3(32'hba556f06),
	.w4(32'hba053c7a),
	.w5(32'hba0ab552),
	.w6(32'hb96c1ed3),
	.w7(32'hb9fe02bc),
	.w8(32'hba1398c7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b27c6),
	.w1(32'h3a9c0c14),
	.w2(32'h3a3f3860),
	.w3(32'h38bca1a2),
	.w4(32'h3a879a27),
	.w5(32'h3a5d5b98),
	.w6(32'hb9b94d39),
	.w7(32'h3a376a54),
	.w8(32'h3a68f03d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a737392),
	.w1(32'hb9af440d),
	.w2(32'h38a37abe),
	.w3(32'h39f2f993),
	.w4(32'hb9d44068),
	.w5(32'hb98282ef),
	.w6(32'h3a174013),
	.w7(32'h3937dac0),
	.w8(32'hb8ec37a2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af1bfb),
	.w1(32'h3a96d590),
	.w2(32'h3aabc18e),
	.w3(32'hb931f922),
	.w4(32'h38265f65),
	.w5(32'h3a1b3ae6),
	.w6(32'h38a46a4e),
	.w7(32'h3a08a3bf),
	.w8(32'h3ab2cfb3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f6856),
	.w1(32'hba2ed269),
	.w2(32'hba11f6e5),
	.w3(32'h393f9dec),
	.w4(32'hba5f2489),
	.w5(32'hb8a7cb8c),
	.w6(32'h3a20b846),
	.w7(32'hba78badf),
	.w8(32'hba0dd933),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cca874),
	.w1(32'h3a14aab9),
	.w2(32'h3a5f9af7),
	.w3(32'hbaa0e0e4),
	.w4(32'h3992a720),
	.w5(32'h3aaaf54a),
	.w6(32'hba5f9bd8),
	.w7(32'h39ac53c0),
	.w8(32'h3a8de8bd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d72f09),
	.w1(32'h3922b8ba),
	.w2(32'h39af2dbf),
	.w3(32'h3a109a9f),
	.w4(32'h392d0cfd),
	.w5(32'hb901d9ee),
	.w6(32'h39c88f37),
	.w7(32'h3a2c72a9),
	.w8(32'h3a1c1b53),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57b73d),
	.w1(32'hba47579d),
	.w2(32'hb7cd96f6),
	.w3(32'hba4fd648),
	.w4(32'h3a22e79d),
	.w5(32'h3aae70a8),
	.w6(32'hb8951418),
	.w7(32'h39656a66),
	.w8(32'h3a62dcb4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be5929),
	.w1(32'hb904a5d6),
	.w2(32'hb9ba89b2),
	.w3(32'hba00faf6),
	.w4(32'h392cb2a6),
	.w5(32'h39a919aa),
	.w6(32'hb9039a51),
	.w7(32'hba16ba5a),
	.w8(32'hb814b625),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849327),
	.w1(32'h3aa19cfa),
	.w2(32'h3aaba314),
	.w3(32'hba16193c),
	.w4(32'h3a92ec29),
	.w5(32'h3ab1ec1d),
	.w6(32'h392adcba),
	.w7(32'h3a7f8fd5),
	.w8(32'h3aa0910f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a750d8e),
	.w1(32'h3a5cd4bf),
	.w2(32'h3a82df80),
	.w3(32'h39c61264),
	.w4(32'h39a48b91),
	.w5(32'h3a81f487),
	.w6(32'h3a0b3814),
	.w7(32'h3aa0319f),
	.w8(32'h3a8b76c4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adfb87),
	.w1(32'hb8c70938),
	.w2(32'hba0bd4a6),
	.w3(32'h3946e1fc),
	.w4(32'hba3b8576),
	.w5(32'hba218c48),
	.w6(32'h3a1730ca),
	.w7(32'hb815d16d),
	.w8(32'hb9f0ab3d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba415c81),
	.w1(32'hbb329f98),
	.w2(32'hbb03f3b6),
	.w3(32'hbaa14611),
	.w4(32'hbb470435),
	.w5(32'hbb1e2142),
	.w6(32'hba0af1a4),
	.w7(32'hbb1dee55),
	.w8(32'hbb3c5260),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb016535),
	.w1(32'h3a1cec7d),
	.w2(32'h3a24bbdc),
	.w3(32'hbb44464a),
	.w4(32'h3a36167d),
	.w5(32'h39844b1f),
	.w6(32'hbb387cf1),
	.w7(32'h3a050841),
	.w8(32'hb9d0e42e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule