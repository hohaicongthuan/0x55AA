module layer_10_featuremap_216(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb55a6d49),
	.w1(32'h37360bac),
	.w2(32'h376ce3a3),
	.w3(32'hb69c44a3),
	.w4(32'hb622bd03),
	.w5(32'h37a5a704),
	.w6(32'hb7bd8104),
	.w7(32'hb7ad40ee),
	.w8(32'h37393515),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99ceda),
	.w1(32'h39795165),
	.w2(32'h3a0bb408),
	.w3(32'hbb1feafd),
	.w4(32'h3acb383d),
	.w5(32'h3aa62ac0),
	.w6(32'hbb6813c5),
	.w7(32'h3a6c0ae1),
	.w8(32'h3b172372),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34169cc2),
	.w1(32'h364d550c),
	.w2(32'h36e8279d),
	.w3(32'hb59a9760),
	.w4(32'h3592640b),
	.w5(32'h3687986a),
	.w6(32'h35b5086f),
	.w7(32'h3619178e),
	.w8(32'h356a9171),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387dcb23),
	.w1(32'hba799105),
	.w2(32'hba53d5c9),
	.w3(32'h3a8d3dae),
	.w4(32'hb897e72f),
	.w5(32'hba444f0d),
	.w6(32'h3aadd90d),
	.w7(32'h39f71f9e),
	.w8(32'hba1e8460),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398525a6),
	.w1(32'h390a0420),
	.w2(32'h36d51698),
	.w3(32'h399771c5),
	.w4(32'h396dcc5a),
	.w5(32'h38d65358),
	.w6(32'h398b98e2),
	.w7(32'h3980f747),
	.w8(32'h39048804),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3603c971),
	.w1(32'h36cde969),
	.w2(32'h37463c89),
	.w3(32'h35bcccb9),
	.w4(32'h35bcf237),
	.w5(32'h373b8729),
	.w6(32'hb611cfab),
	.w7(32'h35ce6244),
	.w8(32'h37501ae6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2d13a),
	.w1(32'hbb3989f4),
	.w2(32'h3aca8cd4),
	.w3(32'hbaa07ae3),
	.w4(32'hbbc1f830),
	.w5(32'h3a3e49dc),
	.w6(32'h3b8ae861),
	.w7(32'h3b22bcd1),
	.w8(32'h3ac88adb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf005f1),
	.w1(32'h3a15e28e),
	.w2(32'h3c06af87),
	.w3(32'h3c07c6f4),
	.w4(32'h3c396b08),
	.w5(32'h3b79fa09),
	.w6(32'h3cafad5c),
	.w7(32'h3c1fcb71),
	.w8(32'h3c29a84f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca8270),
	.w1(32'h398420e9),
	.w2(32'hba24fdf6),
	.w3(32'h3a03b238),
	.w4(32'h39770223),
	.w5(32'hb9ac8026),
	.w6(32'h39dd7344),
	.w7(32'h3959b04b),
	.w8(32'hb9b44e89),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b17be),
	.w1(32'h3a86b124),
	.w2(32'h3ab4cb4b),
	.w3(32'h3942cdee),
	.w4(32'hbacb892f),
	.w5(32'h3acd2548),
	.w6(32'h3abeda0f),
	.w7(32'h3a8ceb82),
	.w8(32'h3a86c2db),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a42c17),
	.w1(32'hb9d4b57f),
	.w2(32'h38187c75),
	.w3(32'hb9b164b5),
	.w4(32'hb9a2ea69),
	.w5(32'h39833d4c),
	.w6(32'hb9a0162e),
	.w7(32'hb95af92c),
	.w8(32'h3a025c39),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6609),
	.w1(32'hbbd957b2),
	.w2(32'hbbb07f0a),
	.w3(32'h3b822e79),
	.w4(32'hbc2672ee),
	.w5(32'hbbdd96e9),
	.w6(32'h3bb3fbff),
	.w7(32'h3a09c47f),
	.w8(32'hbb62e702),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87de0b),
	.w1(32'h3ac13c24),
	.w2(32'h383b0767),
	.w3(32'h3b73ebe2),
	.w4(32'hb7b38cf7),
	.w5(32'h3abda0d1),
	.w6(32'h3bb5c115),
	.w7(32'h3b1f37c5),
	.w8(32'h3a9bba97),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf4a1),
	.w1(32'hbad088ff),
	.w2(32'h3b0c998b),
	.w3(32'hba9902d9),
	.w4(32'h38eb0f84),
	.w5(32'h3b022c0a),
	.w6(32'hba41451b),
	.w7(32'h3a26717f),
	.w8(32'h3b1c7425),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a32988),
	.w1(32'h3ad5e2a9),
	.w2(32'h38cc8138),
	.w3(32'hbae0e09b),
	.w4(32'h3a792298),
	.w5(32'h3a4a08db),
	.w6(32'hbb322481),
	.w7(32'h39f8fdd5),
	.w8(32'h3af8623f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0170d),
	.w1(32'h3a425a68),
	.w2(32'h3a1d7318),
	.w3(32'h3b1a82f7),
	.w4(32'h3b491ea4),
	.w5(32'h3b1f13e8),
	.w6(32'hb9d8fe85),
	.w7(32'h3bbd9b46),
	.w8(32'h3b90d9cb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10ed49),
	.w1(32'h394eb8f1),
	.w2(32'h385d7105),
	.w3(32'h394a603c),
	.w4(32'h39437abe),
	.w5(32'h3926dda4),
	.w6(32'hb901c79f),
	.w7(32'hb7e3f8f5),
	.w8(32'h391e1316),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c9958),
	.w1(32'h3a244d7f),
	.w2(32'h3be15ca3),
	.w3(32'h3b9ca210),
	.w4(32'h3a31908c),
	.w5(32'h3b7f9c07),
	.w6(32'h3c430926),
	.w7(32'h3b8ca8c4),
	.w8(32'hba80b20e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabfe6a),
	.w1(32'h3a41af20),
	.w2(32'h3aef6151),
	.w3(32'h3b518ea4),
	.w4(32'h38a08c24),
	.w5(32'h3a1af343),
	.w6(32'h3bdef1e7),
	.w7(32'h3b31f2cf),
	.w8(32'hba27e16b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39664020),
	.w1(32'hb6807a7b),
	.w2(32'hb84d3ad5),
	.w3(32'hb79de427),
	.w4(32'h3809fb33),
	.w5(32'hb8b6f72a),
	.w6(32'hb98b6730),
	.w7(32'h392f6ff9),
	.w8(32'h38d61069),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a78dad),
	.w1(32'h3867ab51),
	.w2(32'h391f9083),
	.w3(32'h388de959),
	.w4(32'h390b37f4),
	.w5(32'h390210bd),
	.w6(32'h386b879f),
	.w7(32'h379b142b),
	.w8(32'h38a4c52e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983061d),
	.w1(32'h3a207268),
	.w2(32'h3a1cbc6d),
	.w3(32'hba26bd47),
	.w4(32'h3a5e3677),
	.w5(32'h3a9051a5),
	.w6(32'hba99e556),
	.w7(32'h39f61a77),
	.w8(32'h3aaceb60),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb037754),
	.w1(32'h3b773013),
	.w2(32'h3b752680),
	.w3(32'h3c0f034b),
	.w4(32'h3a0c191e),
	.w5(32'hb9081f54),
	.w6(32'h3aa3be62),
	.w7(32'h3bd0dc96),
	.w8(32'hba175c43),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9171929),
	.w1(32'hba18eff2),
	.w2(32'hbab3ed52),
	.w3(32'hba336118),
	.w4(32'hbab4dcd1),
	.w5(32'hbab32dbc),
	.w6(32'hba25262f),
	.w7(32'h399b682a),
	.w8(32'h39130ba1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ffd8),
	.w1(32'h3a9520e8),
	.w2(32'hbb4eccc4),
	.w3(32'hbb79dc51),
	.w4(32'h3b2b13ae),
	.w5(32'hba3d4a23),
	.w6(32'hbc0c9216),
	.w7(32'h3aa1b103),
	.w8(32'h3b429b86),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39265bf7),
	.w1(32'h39b397e8),
	.w2(32'h39a916ac),
	.w3(32'h39226b6e),
	.w4(32'h39ad6b44),
	.w5(32'h39c8a4e8),
	.w6(32'h37a19f6e),
	.w7(32'h39422940),
	.w8(32'h39a0f78d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363c6fd4),
	.w1(32'hb8158952),
	.w2(32'hb88d4fd3),
	.w3(32'hb7079377),
	.w4(32'hb78f3093),
	.w5(32'hb83527f1),
	.w6(32'hb85fbb98),
	.w7(32'hb7c36cdf),
	.w8(32'hb74debaf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91e67e),
	.w1(32'hbb15611e),
	.w2(32'hb9e08660),
	.w3(32'hbbd9f640),
	.w4(32'hbbad2a19),
	.w5(32'h3a220bf3),
	.w6(32'hbba7e1ef),
	.w7(32'hbb928300),
	.w8(32'hba52998a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afacdf),
	.w1(32'hba2b2257),
	.w2(32'h39c142ea),
	.w3(32'hb9b65b28),
	.w4(32'hba537a54),
	.w5(32'h39507957),
	.w6(32'hb974befb),
	.w7(32'hb9f6d290),
	.w8(32'h396619cb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0c76),
	.w1(32'hb97f4f37),
	.w2(32'hbb01c058),
	.w3(32'hbc09bb3b),
	.w4(32'h3a9add55),
	.w5(32'h3a9b9140),
	.w6(32'hbc3cfe4a),
	.w7(32'hb96cf527),
	.w8(32'h3b58cfbb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b43590),
	.w1(32'h353d9ad4),
	.w2(32'h3784d5f8),
	.w3(32'h36ecef1a),
	.w4(32'hb7467290),
	.w5(32'h372260cb),
	.w6(32'hb66e18dc),
	.w7(32'hb707ed3b),
	.w8(32'h37476d53),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7862efb),
	.w1(32'hb80f90c2),
	.w2(32'h3804ec54),
	.w3(32'hb814b66d),
	.w4(32'hb8a1ba7a),
	.w5(32'h390d6ec9),
	.w6(32'hb86d7af6),
	.w7(32'hb88cebfd),
	.w8(32'h39437fd4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee6fdc),
	.w1(32'h39bc6f73),
	.w2(32'h3a2cae74),
	.w3(32'h3a74a183),
	.w4(32'hb9a13b41),
	.w5(32'hb9cea911),
	.w6(32'h3b412771),
	.w7(32'h3ae8a101),
	.w8(32'hb8970944),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5cc11),
	.w1(32'h390cdbdd),
	.w2(32'hba020725),
	.w3(32'hbb08e8cf),
	.w4(32'h396fedd2),
	.w5(32'h3922be0e),
	.w6(32'hbb2c82a9),
	.w7(32'hb98e9503),
	.w8(32'h39dbc4b2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a4bf3),
	.w1(32'hb905fe24),
	.w2(32'hb96f1482),
	.w3(32'hb8c8d90e),
	.w4(32'hba6f3aff),
	.w5(32'hba51652d),
	.w6(32'h39e3d19a),
	.w7(32'h39c682f5),
	.w8(32'hb94ba9eb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b78ecd),
	.w1(32'hbb067baa),
	.w2(32'hbac396ea),
	.w3(32'h3b4afaad),
	.w4(32'hbb37ba20),
	.w5(32'hbb03b8e9),
	.w6(32'h3bb15cb8),
	.w7(32'h3ae03484),
	.w8(32'h3a7b003b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c916440),
	.w1(32'h3aa85a2e),
	.w2(32'hbc0d9c59),
	.w3(32'h3ca18e43),
	.w4(32'h3b143d4c),
	.w5(32'hbae0c59c),
	.w6(32'h3b77d759),
	.w7(32'h3aff3630),
	.w8(32'hbbb722a5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fc32c),
	.w1(32'h3b23b4bf),
	.w2(32'hbaa447db),
	.w3(32'hbbf4592b),
	.w4(32'h3b008a6c),
	.w5(32'h3ade16e4),
	.w6(32'hbc334708),
	.w7(32'h3b249e9d),
	.w8(32'h3be3a248),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb613f48),
	.w1(32'h3b446f89),
	.w2(32'h3b6b606b),
	.w3(32'hbc0d0e9e),
	.w4(32'hbb1e9deb),
	.w5(32'h3b895b03),
	.w6(32'hbc1769ea),
	.w7(32'hba49c8b6),
	.w8(32'h3b96b42b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a2253),
	.w1(32'h39aad5ac),
	.w2(32'hba0adf46),
	.w3(32'hb981e946),
	.w4(32'h3a4916b6),
	.w5(32'h398e36ac),
	.w6(32'hba4bf3f7),
	.w7(32'h3a8d7489),
	.w8(32'h3aa06768),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a29bcd),
	.w1(32'hb888ee31),
	.w2(32'h379cc25c),
	.w3(32'hb7fa9794),
	.w4(32'hb81ac06d),
	.w5(32'h3891d209),
	.w6(32'hb564ade1),
	.w7(32'h3888a405),
	.w8(32'h391e98b7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0097c),
	.w1(32'hb8dd29ca),
	.w2(32'hb96ef4d2),
	.w3(32'hb7db01da),
	.w4(32'hb831422e),
	.w5(32'hb948b5f7),
	.w6(32'hb8b17024),
	.w7(32'hb8d74fb7),
	.w8(32'hb95c8c87),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9873532),
	.w1(32'hb9eb45bb),
	.w2(32'h39184d20),
	.w3(32'hba0cad9c),
	.w4(32'hba206781),
	.w5(32'h398b2bc9),
	.w6(32'hb9ddd5ee),
	.w7(32'hba3ff17d),
	.w8(32'h397b54ef),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b263576),
	.w1(32'hbb2764fa),
	.w2(32'h3bbe147d),
	.w3(32'h3b74e564),
	.w4(32'hbb1c43d9),
	.w5(32'h3b784ebe),
	.w6(32'h3bc09e62),
	.w7(32'h3ad103bb),
	.w8(32'h3aa744ad),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae4ed),
	.w1(32'h3a005733),
	.w2(32'hbb7a642b),
	.w3(32'hbafc78cf),
	.w4(32'h3ac9b0de),
	.w5(32'hbacf6278),
	.w6(32'hbb8afa7e),
	.w7(32'h3785a302),
	.w8(32'hb9ad91fe),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48037e),
	.w1(32'hba9950ac),
	.w2(32'hbb98625e),
	.w3(32'h3a933452),
	.w4(32'h3975b1ef),
	.w5(32'hbaeaea3d),
	.w6(32'h3ad888a2),
	.w7(32'h3acb821c),
	.w8(32'h3992aee9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc6577),
	.w1(32'h3af35728),
	.w2(32'hba101076),
	.w3(32'hb9721efc),
	.w4(32'h3ae1665b),
	.w5(32'hba53cb72),
	.w6(32'h3a8f0881),
	.w7(32'h3a3d9d54),
	.w8(32'hba800084),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44a2a),
	.w1(32'hba13c1a9),
	.w2(32'h3b434fff),
	.w3(32'h3c12ec03),
	.w4(32'hb90659b1),
	.w5(32'h3a601ef2),
	.w6(32'h3c910605),
	.w7(32'h3c01da1a),
	.w8(32'hbae6825f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a42e97),
	.w1(32'hb9f74db5),
	.w2(32'hb955064d),
	.w3(32'hb99a24b9),
	.w4(32'hb981c8eb),
	.w5(32'hb96cb501),
	.w6(32'hb909b91f),
	.w7(32'h375ce968),
	.w8(32'hb954eeb3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f4dc6),
	.w1(32'h398492c2),
	.w2(32'hb793b1fc),
	.w3(32'hb88b0136),
	.w4(32'h39c11c68),
	.w5(32'h376bad50),
	.w6(32'h362d8736),
	.w7(32'h3919609b),
	.w8(32'hba1c844a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d27c9d),
	.w1(32'hb9b32f85),
	.w2(32'hb94d7fef),
	.w3(32'hb9378ef8),
	.w4(32'h37a0107f),
	.w5(32'hb8e564fe),
	.w6(32'hb96e5354),
	.w7(32'hb86a0d0d),
	.w8(32'hb79494a6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f79327),
	.w1(32'h3a3d07fe),
	.w2(32'h3a920bf4),
	.w3(32'h3a885ad8),
	.w4(32'h3ac0a2b7),
	.w5(32'h3b0ce64a),
	.w6(32'hbac5122e),
	.w7(32'h3b1f7d94),
	.w8(32'h3b264d98),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aad1a5),
	.w1(32'hb92bcb1e),
	.w2(32'h38db56fa),
	.w3(32'h39f91737),
	.w4(32'h39261c01),
	.w5(32'hb94ebc8b),
	.w6(32'h3a7e069c),
	.w7(32'h3a0a5a43),
	.w8(32'hb80b5f2c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a790d20),
	.w1(32'hbaf572f7),
	.w2(32'h3b49090d),
	.w3(32'h3b07c2a7),
	.w4(32'hbb585237),
	.w5(32'hb9b88eae),
	.w6(32'h3c3a18de),
	.w7(32'h3b659a31),
	.w8(32'hbb5ac61e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914f530),
	.w1(32'hba37062b),
	.w2(32'hb99e5b7c),
	.w3(32'hba47ecda),
	.w4(32'hba5d64e6),
	.w5(32'h3724f7e2),
	.w6(32'h399eb2a4),
	.w7(32'h38fe12f1),
	.w8(32'h399f6201),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90acf05),
	.w1(32'h3929b911),
	.w2(32'h38a7447c),
	.w3(32'hb973766d),
	.w4(32'h386bfe23),
	.w5(32'h38b74a83),
	.w6(32'hb9b4a983),
	.w7(32'hb8743279),
	.w8(32'h38a69170),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a521e),
	.w1(32'h35e4b33e),
	.w2(32'hb7c45a38),
	.w3(32'h37276820),
	.w4(32'h37fda34d),
	.w5(32'h356fc78a),
	.w6(32'hb7d7ea99),
	.w7(32'h37a7c867),
	.w8(32'h36f8c682),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43531c),
	.w1(32'hb94db180),
	.w2(32'hb8d5e841),
	.w3(32'hba7774a4),
	.w4(32'hba084a77),
	.w5(32'h39975baf),
	.w6(32'hba951638),
	.w7(32'hb981b65f),
	.w8(32'h3a0ff204),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c78021),
	.w1(32'h3988cb06),
	.w2(32'h38f10215),
	.w3(32'h3982bf81),
	.w4(32'h397650cc),
	.w5(32'h3893190f),
	.w6(32'h391d92df),
	.w7(32'h387502fe),
	.w8(32'hb7adfe4f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a35e0),
	.w1(32'h390e10b4),
	.w2(32'hb8b28dca),
	.w3(32'h38a1a8d5),
	.w4(32'hb9ed262a),
	.w5(32'hb9619eb9),
	.w6(32'h38fddb9d),
	.w7(32'hb9b1fba0),
	.w8(32'hb9f6c089),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a604b3a),
	.w1(32'hb9b99acc),
	.w2(32'h3a67375e),
	.w3(32'h3b16972e),
	.w4(32'hb9dfd6a1),
	.w5(32'hb98ff4c1),
	.w6(32'h3b4d7342),
	.w7(32'h3abf54f7),
	.w8(32'hb96b78cf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b685b6e),
	.w1(32'h3b86ee35),
	.w2(32'h3b939087),
	.w3(32'h3adb18b3),
	.w4(32'h3bbf4ccd),
	.w5(32'h3b80cf43),
	.w6(32'hbb0834ed),
	.w7(32'h3a960a1e),
	.w8(32'h3a7f6626),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83fffe0),
	.w1(32'hb79aed90),
	.w2(32'h360ece05),
	.w3(32'h36b5359c),
	.w4(32'h382be001),
	.w5(32'h3815b3d9),
	.w6(32'hb65db893),
	.w7(32'h3811e48a),
	.w8(32'h37ec29af),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3696b375),
	.w1(32'h3719c7d0),
	.w2(32'hb79f80c0),
	.w3(32'hb7191dc1),
	.w4(32'h370649b6),
	.w5(32'hb61501ca),
	.w6(32'hb80a66f2),
	.w7(32'hb6f1936d),
	.w8(32'hb6be2c36),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82334c4),
	.w1(32'hb84e1960),
	.w2(32'h38943059),
	.w3(32'hb7ae6cf2),
	.w4(32'hb8ca0f6b),
	.w5(32'h37fe54c9),
	.w6(32'h37c331ec),
	.w7(32'hb84b2ac9),
	.w8(32'h37a32448),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fc8fa5),
	.w1(32'hb8048ba1),
	.w2(32'hb82c2a03),
	.w3(32'h3791c812),
	.w4(32'h35b3da89),
	.w5(32'hb7b5de96),
	.w6(32'hb4a6d772),
	.w7(32'h37591b94),
	.w8(32'hb71633d3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b8c5f),
	.w1(32'h3acdb482),
	.w2(32'h3be1c44b),
	.w3(32'hbaab19e6),
	.w4(32'hbb71140e),
	.w5(32'h3bc55da6),
	.w6(32'h3c03b0ce),
	.w7(32'h3a44ca21),
	.w8(32'h3a8f4bbc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35c48c),
	.w1(32'hbb3f110e),
	.w2(32'hbbc39b01),
	.w3(32'h3bbc229b),
	.w4(32'h3aeac959),
	.w5(32'h3b225ffd),
	.w6(32'h3c510530),
	.w7(32'h3c2ec4fc),
	.w8(32'h3bfa8d7c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0f2d4),
	.w1(32'h39dd1621),
	.w2(32'h3af26e49),
	.w3(32'h3a5e3325),
	.w4(32'h3a296296),
	.w5(32'h3b14f4f9),
	.w6(32'h3ad325a2),
	.w7(32'h3b19faf7),
	.w8(32'h3a87804d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88225a),
	.w1(32'hbae43783),
	.w2(32'hbbf39b59),
	.w3(32'hbba390ea),
	.w4(32'hba3a719d),
	.w5(32'hbb9eb428),
	.w6(32'hbc0dc239),
	.w7(32'h3ab21235),
	.w8(32'h3b4c110c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3819d8be),
	.w1(32'hb7b3105a),
	.w2(32'hb81ba712),
	.w3(32'h388ec15b),
	.w4(32'hb7295052),
	.w5(32'hb7f7992e),
	.w6(32'h381e673a),
	.w7(32'hb6e2aeee),
	.w8(32'h37a0c61f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fab7f6),
	.w1(32'hb77092be),
	.w2(32'hb7afbedf),
	.w3(32'hb72fab26),
	.w4(32'h381bd723),
	.w5(32'h37328432),
	.w6(32'hb8630d97),
	.w7(32'h36842671),
	.w8(32'h35680828),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38037742),
	.w1(32'h382be18b),
	.w2(32'h335e5790),
	.w3(32'h384cd427),
	.w4(32'h38635eba),
	.w5(32'h35ead28d),
	.w6(32'hb798a1cb),
	.w7(32'h383743ae),
	.w8(32'h381674ec),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d45ce),
	.w1(32'hb81d9e17),
	.w2(32'h3a06b4fa),
	.w3(32'h3a5fdede),
	.w4(32'hb9085603),
	.w5(32'h3a192b51),
	.w6(32'h3b3f861a),
	.w7(32'h3ac55a93),
	.w8(32'h3a697635),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83042c1),
	.w1(32'hb8749937),
	.w2(32'hb89e5e29),
	.w3(32'h38b8e35a),
	.w4(32'h37fabcc0),
	.w5(32'hb886c533),
	.w6(32'h389e0627),
	.w7(32'h375118cb),
	.w8(32'hb8bea4f3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9894bf),
	.w1(32'hb7ee8ca4),
	.w2(32'h3a536628),
	.w3(32'h3b4ac271),
	.w4(32'hba1e1769),
	.w5(32'hbaba915f),
	.w6(32'h3b9c59af),
	.w7(32'h3acb88f2),
	.w8(32'hbad48f9d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89004e),
	.w1(32'h3a43689b),
	.w2(32'h3b7302e5),
	.w3(32'h3c01c9c5),
	.w4(32'h3af9a93e),
	.w5(32'hbaaf9ced),
	.w6(32'h3c50be6e),
	.w7(32'h3be7cd43),
	.w8(32'h3b0ea41e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879f037),
	.w1(32'h3b1b0cad),
	.w2(32'hba85dcc3),
	.w3(32'hb9e0ea48),
	.w4(32'h3b8f6c86),
	.w5(32'h3b2a23b9),
	.w6(32'hbb8980b8),
	.w7(32'h3aa362c5),
	.w8(32'h3afc846f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91a8d3),
	.w1(32'hba518e64),
	.w2(32'h3b0fe4ac),
	.w3(32'hbabc7b1e),
	.w4(32'hbaa6e6dd),
	.w5(32'h3ab5f9d2),
	.w6(32'h3a537918),
	.w7(32'hb9f2525c),
	.w8(32'h3a206261),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4c1ab),
	.w1(32'hba74f733),
	.w2(32'hbb027d91),
	.w3(32'hb9bb3d2b),
	.w4(32'hbb5a2aa7),
	.w5(32'hbacf9db6),
	.w6(32'h39933f46),
	.w7(32'hbae95294),
	.w8(32'hba0e561f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba376b54),
	.w1(32'hb941bb26),
	.w2(32'hba629a65),
	.w3(32'hbb10b9b2),
	.w4(32'hb9f48977),
	.w5(32'hb966c93d),
	.w6(32'hbb108cb5),
	.w7(32'hbaa8e98c),
	.w8(32'hba3f534c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af82397),
	.w1(32'hb9e5d506),
	.w2(32'h3a017bfc),
	.w3(32'h3b26b729),
	.w4(32'hba3ea316),
	.w5(32'hb9f6df7b),
	.w6(32'h3b99e14b),
	.w7(32'h3ad1ec7d),
	.w8(32'hbaafa573),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb643dfcb),
	.w1(32'h368c9cc9),
	.w2(32'h379434a0),
	.w3(32'h36afa954),
	.w4(32'h37525d8c),
	.w5(32'h374aaa69),
	.w6(32'h36e2595c),
	.w7(32'h3658975e),
	.w8(32'hb4692624),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37df32a9),
	.w1(32'h3836d7ae),
	.w2(32'h38067f15),
	.w3(32'hb510e3cc),
	.w4(32'h383a87d5),
	.w5(32'h387669f9),
	.w6(32'hb803fd0b),
	.w7(32'hb5b90798),
	.w8(32'h3802b2b0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a432f0),
	.w1(32'h371be825),
	.w2(32'hb703c93e),
	.w3(32'h373fdd83),
	.w4(32'h37d084b3),
	.w5(32'h376af2d6),
	.w6(32'hb79514cd),
	.w7(32'hb7b064f2),
	.w8(32'h3731eac2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ca95b),
	.w1(32'hba126d59),
	.w2(32'h392afdd5),
	.w3(32'hba5c3d56),
	.w4(32'hba39010d),
	.w5(32'h39b132c6),
	.w6(32'hba6b0699),
	.w7(32'hb9cc6a1c),
	.w8(32'h39fa021f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a018f24),
	.w1(32'h38bcfd4b),
	.w2(32'hbb299516),
	.w3(32'hbac93677),
	.w4(32'h3a9d3427),
	.w5(32'hbaaf04fe),
	.w6(32'hbb5573a9),
	.w7(32'h3a3affac),
	.w8(32'h3a4f18fa),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990f2e8),
	.w1(32'h39b2fec0),
	.w2(32'h3946718e),
	.w3(32'h39a4769d),
	.w4(32'h39b227a0),
	.w5(32'h394bc2d0),
	.w6(32'h397568ce),
	.w7(32'h3992598d),
	.w8(32'h393360a0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e861ce),
	.w1(32'hba3df199),
	.w2(32'hbb8cfa00),
	.w3(32'h3ad8eadc),
	.w4(32'h3a98659a),
	.w5(32'hbb0d2408),
	.w6(32'h3a6d95f6),
	.w7(32'h3aeefbe2),
	.w8(32'h3946466e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395545e7),
	.w1(32'hbab49431),
	.w2(32'h3bb2506e),
	.w3(32'h3b1927f0),
	.w4(32'hbb09ac87),
	.w5(32'h39b46b20),
	.w6(32'h3bdf8235),
	.w7(32'h3b70b2c1),
	.w8(32'hbb027823),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb488fa8),
	.w1(32'h39a9812f),
	.w2(32'hba99c15a),
	.w3(32'hbb97ca94),
	.w4(32'hba453a64),
	.w5(32'h39845cc8),
	.w6(32'hbb89caa8),
	.w7(32'hb95c30a7),
	.w8(32'h3ae3dc23),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66c883),
	.w1(32'h3a569249),
	.w2(32'hbba9fa40),
	.w3(32'h3c5de377),
	.w4(32'h3ad124e8),
	.w5(32'hbb169d9c),
	.w6(32'h3be396b5),
	.w7(32'h3b9b104a),
	.w8(32'hbb4371de),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bc96e),
	.w1(32'hbb0c1d2c),
	.w2(32'hbb15b152),
	.w3(32'hbb7dba4c),
	.w4(32'hbb07f7e4),
	.w5(32'h3a9a8966),
	.w6(32'hbb7d19e9),
	.w7(32'hba05c8fe),
	.w8(32'h3ac9399b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ae4b0),
	.w1(32'hbb9b5f86),
	.w2(32'h3b860fb0),
	.w3(32'hbb90456d),
	.w4(32'hbb6ed819),
	.w5(32'h3a08482a),
	.w6(32'hba9f9d36),
	.w7(32'hb91c498f),
	.w8(32'hba073903),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cb88f),
	.w1(32'hbb2a882a),
	.w2(32'hbb1b9740),
	.w3(32'hbb6b4881),
	.w4(32'hbb37ace2),
	.w5(32'hb77ea936),
	.w6(32'hbba07a44),
	.w7(32'hbb180f8c),
	.w8(32'hb97878b5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165fdb),
	.w1(32'h3a11f950),
	.w2(32'hba48721f),
	.w3(32'hbb88ec23),
	.w4(32'h3b0d50c9),
	.w5(32'h3accc822),
	.w6(32'hbba0304a),
	.w7(32'h3affa9dc),
	.w8(32'h3b8c54a3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aab51d),
	.w1(32'h37e80578),
	.w2(32'hba2a7bd1),
	.w3(32'hb9f0a2f8),
	.w4(32'hba08e2f3),
	.w5(32'hba70795d),
	.w6(32'hb9dcbf82),
	.w7(32'hba4db371),
	.w8(32'hba984ec6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75ead8),
	.w1(32'h368b2944),
	.w2(32'h3aab458d),
	.w3(32'h3a8caa78),
	.w4(32'hbaa2afa2),
	.w5(32'hba8f3639),
	.w6(32'h3bac986d),
	.w7(32'h3ab728d9),
	.w8(32'hbafcd62b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dd3a3),
	.w1(32'hbb3f1f51),
	.w2(32'hbb1cb17e),
	.w3(32'h3acc7f41),
	.w4(32'hbbc8db0e),
	.w5(32'hbaa6432e),
	.w6(32'h3a31435a),
	.w7(32'hbb2b1215),
	.w8(32'hbba5da9c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69efc4),
	.w1(32'h3abeffe2),
	.w2(32'h39ddeb96),
	.w3(32'h3cc3f246),
	.w4(32'h3b8b7fc5),
	.w5(32'h392fc832),
	.w6(32'h3c3131f5),
	.w7(32'h3c7a9912),
	.w8(32'h3b2b0525),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb271659),
	.w1(32'hba477075),
	.w2(32'hba7fa9c1),
	.w3(32'hbb9f88b3),
	.w4(32'h3a8073a6),
	.w5(32'h3b35ffd3),
	.w6(32'hbbb441db),
	.w7(32'h3ab4c383),
	.w8(32'h3b810c64),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e96fd),
	.w1(32'hba6ad37d),
	.w2(32'hbba273d0),
	.w3(32'hbb4add3f),
	.w4(32'hb970c1d1),
	.w5(32'hbb170b4e),
	.w6(32'hbbb2fc94),
	.w7(32'h3a113cde),
	.w8(32'h3a81baa9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d1578),
	.w1(32'hbb9c6cd8),
	.w2(32'hbb8bb1a9),
	.w3(32'h3b9f1881),
	.w4(32'hbc04d7f5),
	.w5(32'hbbb43796),
	.w6(32'h3b317bf3),
	.w7(32'h3a985602),
	.w8(32'hbc054d44),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba574bc2),
	.w1(32'hba8d7e57),
	.w2(32'hbae83b8e),
	.w3(32'hba2d1d95),
	.w4(32'hba62a536),
	.w5(32'hbad2b5e0),
	.w6(32'hb9b96d82),
	.w7(32'hba2af218),
	.w8(32'hbadc2240),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ea077),
	.w1(32'hb9f37fe4),
	.w2(32'h3bedd246),
	.w3(32'h3c54e6f8),
	.w4(32'h3b85f68d),
	.w5(32'h3ae63189),
	.w6(32'h3b8ee606),
	.w7(32'h3c0babf3),
	.w8(32'h3b27b7df),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7649ed),
	.w1(32'hb980e25b),
	.w2(32'h398d4b52),
	.w3(32'h3b99ec86),
	.w4(32'hbb1a9e1a),
	.w5(32'hbb6c5e2a),
	.w6(32'h3b98a1bf),
	.w7(32'h3af9ffa5),
	.w8(32'hbaf8c681),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ce9bcd),
	.w1(32'h39455d4c),
	.w2(32'hb7bfa3d8),
	.w3(32'h370c00ec),
	.w4(32'h39b0b919),
	.w5(32'h3967e2b1),
	.w6(32'hb9838c6b),
	.w7(32'h37994c93),
	.w8(32'h39473b0e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39220713),
	.w1(32'h3a4b0573),
	.w2(32'h39806f6f),
	.w3(32'h3a636d49),
	.w4(32'h3aba567f),
	.w5(32'h3ac525db),
	.w6(32'hb9e2cebe),
	.w7(32'h3b10bce8),
	.w8(32'h3b28f4ee),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade0284),
	.w1(32'hb87a73cd),
	.w2(32'h3a68ae96),
	.w3(32'h3b1ebc32),
	.w4(32'hb9c9a34d),
	.w5(32'h3a415820),
	.w6(32'h3b71d9d9),
	.w7(32'h3ae9b90c),
	.w8(32'h3a5eea86),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6777),
	.w1(32'h39b6c1ae),
	.w2(32'hbab3d810),
	.w3(32'hbb03e116),
	.w4(32'h3a51e8f3),
	.w5(32'hba0b672f),
	.w6(32'hbb65f2a2),
	.w7(32'h3a72690e),
	.w8(32'h3aacc7d3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ba5c6),
	.w1(32'h3bcd3b8a),
	.w2(32'h3bc22e93),
	.w3(32'hbaabbb83),
	.w4(32'h3b06c524),
	.w5(32'h3bef5d72),
	.w6(32'hbafe4788),
	.w7(32'h3b34b315),
	.w8(32'h3b9b795c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafefb8f),
	.w1(32'h3984f997),
	.w2(32'hba3fc804),
	.w3(32'hbb54d136),
	.w4(32'h39ef20ae),
	.w5(32'hb8a24ccd),
	.w6(32'hbb952e6b),
	.w7(32'hbac73825),
	.w8(32'h39b53acd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace2da4),
	.w1(32'hbb8f021d),
	.w2(32'hbc647bdf),
	.w3(32'h3be07306),
	.w4(32'h3ac15fc3),
	.w5(32'hbc13f6d7),
	.w6(32'h3c2ec9d0),
	.w7(32'h3be05071),
	.w8(32'h3ac38f9a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab4cb2),
	.w1(32'hba24de42),
	.w2(32'h3a7d3dd6),
	.w3(32'h38867340),
	.w4(32'h3a5ec743),
	.w5(32'h3a9d630c),
	.w6(32'hbb302bbb),
	.w7(32'h3ae14b6a),
	.w8(32'h37bedbb0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3e2e9),
	.w1(32'hb9c716b9),
	.w2(32'hbae544ef),
	.w3(32'hb9f8f4b5),
	.w4(32'hb925befd),
	.w5(32'hba15ea41),
	.w6(32'hba929e65),
	.w7(32'hb94854c7),
	.w8(32'hb9a193a3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8f2d1),
	.w1(32'h389cfd77),
	.w2(32'h3683e091),
	.w3(32'h3831b5f2),
	.w4(32'h38c05bac),
	.w5(32'hb67760cc),
	.w6(32'h3634067c),
	.w7(32'h364e522c),
	.w8(32'hb7e4d78a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3542df),
	.w1(32'h396cf825),
	.w2(32'hba0727b7),
	.w3(32'hb931272b),
	.w4(32'h39d0b939),
	.w5(32'hb9f8b068),
	.w6(32'hba1e336d),
	.w7(32'hba13f893),
	.w8(32'hb9c2876e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ad201),
	.w1(32'hb73155c2),
	.w2(32'h37cd33a7),
	.w3(32'h377d27b7),
	.w4(32'h36e3ee43),
	.w5(32'h377624ad),
	.w6(32'h37c67850),
	.w7(32'h379dbc19),
	.w8(32'h361c48d6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982a456),
	.w1(32'h39f5b3b3),
	.w2(32'h3a0b9bf4),
	.w3(32'h3940ddf1),
	.w4(32'h39e11131),
	.w5(32'h39e6d783),
	.w6(32'h397a1d2e),
	.w7(32'h39a2803a),
	.w8(32'h3888fe3b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ce434e),
	.w1(32'hb99f650e),
	.w2(32'hbb176941),
	.w3(32'hba09dc34),
	.w4(32'hba09a42b),
	.w5(32'hba8c2940),
	.w6(32'hbaf06cf7),
	.w7(32'hba8a7c9b),
	.w8(32'hba926cb8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6da39),
	.w1(32'h3813604e),
	.w2(32'hb906e6de),
	.w3(32'h389c9236),
	.w4(32'h38243fd3),
	.w5(32'h391e806d),
	.w6(32'hb9a76e9d),
	.w7(32'h388d4d47),
	.w8(32'h39580821),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc1582),
	.w1(32'hba807b73),
	.w2(32'hbacdf8ce),
	.w3(32'h3b20c555),
	.w4(32'hbafd95c9),
	.w5(32'hbb3994fb),
	.w6(32'h3b9dbed4),
	.w7(32'h39c9f3b1),
	.w8(32'hbb09f65b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfa612),
	.w1(32'h3b0e6fc5),
	.w2(32'h3a710357),
	.w3(32'hbb794bb0),
	.w4(32'h3b6fa971),
	.w5(32'h3b1b2469),
	.w6(32'hbbc3c338),
	.w7(32'h3b0be7f5),
	.w8(32'h3ba68e6d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80dc9a9),
	.w1(32'hb76020bf),
	.w2(32'h38a297d5),
	.w3(32'hb872ad16),
	.w4(32'h38328ef3),
	.w5(32'h38ef02a3),
	.w6(32'hb8e95c03),
	.w7(32'h36dea95e),
	.w8(32'h38f4561c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38216523),
	.w1(32'hb79cead9),
	.w2(32'hb8890eb2),
	.w3(32'h38c3e575),
	.w4(32'h377dcd21),
	.w5(32'hb83cddae),
	.w6(32'h38890e9d),
	.w7(32'hb80ee0f1),
	.w8(32'hb853940f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787bbaa),
	.w1(32'h37993f5b),
	.w2(32'h389159ef),
	.w3(32'h37b620bf),
	.w4(32'h37a0152c),
	.w5(32'h387e9077),
	.w6(32'h368284c2),
	.w7(32'hb70a3472),
	.w8(32'h38788d1b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38425ba3),
	.w1(32'h3a1328a7),
	.w2(32'h39ae9a80),
	.w3(32'h39e6fea4),
	.w4(32'h3a75c331),
	.w5(32'h3a1369d9),
	.w6(32'h39aff959),
	.w7(32'h3a3a225a),
	.w8(32'h39fa1166),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a495393),
	.w1(32'hbbbf0bfd),
	.w2(32'hbbbff924),
	.w3(32'h3befc575),
	.w4(32'hbac35910),
	.w5(32'h3a72cc23),
	.w6(32'h3c413c66),
	.w7(32'h3c35ef4a),
	.w8(32'h3c008be7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39971905),
	.w1(32'h398c1ef0),
	.w2(32'h3a629bfb),
	.w3(32'h390e625c),
	.w4(32'hbacdeda8),
	.w5(32'h3b0d4cee),
	.w6(32'h3c07774a),
	.w7(32'h3b2a8b58),
	.w8(32'h39a27a86),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c31dea),
	.w1(32'hba78bc3d),
	.w2(32'h3a265953),
	.w3(32'hb98f9a9c),
	.w4(32'hbae8e02f),
	.w5(32'hba5ffa43),
	.w6(32'hb9b99a01),
	.w7(32'hba373fda),
	.w8(32'hbabba0b6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea4247),
	.w1(32'hb84868dc),
	.w2(32'h3a77fb0f),
	.w3(32'h39bee95e),
	.w4(32'h38c5d64d),
	.w5(32'hb8dfbe04),
	.w6(32'h3a69b00a),
	.w7(32'h3a9d159a),
	.w8(32'h3a3055c2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaff61d),
	.w1(32'hba4dcbda),
	.w2(32'hbb166ef1),
	.w3(32'hbb0194e3),
	.w4(32'hba67ef0a),
	.w5(32'hba8c591c),
	.w6(32'hbb006f9e),
	.w7(32'hb9f03bea),
	.w8(32'hb9a131c8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1754dd),
	.w1(32'h39d25205),
	.w2(32'h3a35cb32),
	.w3(32'hbb163006),
	.w4(32'h3a2ba18a),
	.w5(32'h3a8b5816),
	.w6(32'h3a935298),
	.w7(32'h39f90993),
	.w8(32'h39a5696e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61b9c6),
	.w1(32'hbb1c286d),
	.w2(32'hbb17fff8),
	.w3(32'hbbb60739),
	.w4(32'hbaad0c04),
	.w5(32'hbab5c477),
	.w6(32'hbc0192be),
	.w7(32'hbace209a),
	.w8(32'hbaa62852),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1049f3),
	.w1(32'hba253567),
	.w2(32'h3af838f5),
	.w3(32'h3b0234b6),
	.w4(32'hbb9ee541),
	.w5(32'hba41cb71),
	.w6(32'h3c10660f),
	.w7(32'h3b0e98a7),
	.w8(32'hbb24dc94),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82d693),
	.w1(32'h39d12276),
	.w2(32'hbae3822d),
	.w3(32'hbad785ca),
	.w4(32'h3a96e1d6),
	.w5(32'hb943bfc3),
	.w6(32'hbb4e289a),
	.w7(32'h3a82aa15),
	.w8(32'h3a8cd826),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b1288),
	.w1(32'h3a7bdeb7),
	.w2(32'hba8d2c7c),
	.w3(32'h3a603df0),
	.w4(32'hb9dae30d),
	.w5(32'hb9bd8fb9),
	.w6(32'hbaa762ae),
	.w7(32'h3ad1e88a),
	.w8(32'h399ab8bf),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebe0b4),
	.w1(32'hbb70b033),
	.w2(32'h39dcdb6c),
	.w3(32'h3ad9a423),
	.w4(32'hbbbf5f7f),
	.w5(32'hbb74f6ee),
	.w6(32'h3bef342a),
	.w7(32'hb808581c),
	.w8(32'hbb9b58b4),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f4e7),
	.w1(32'hba90940b),
	.w2(32'hbba5071c),
	.w3(32'h3b867012),
	.w4(32'h3ac07ad1),
	.w5(32'hbb3ebfeb),
	.w6(32'h3aab559e),
	.w7(32'h3b32b8b7),
	.w8(32'h3a8311bc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa446),
	.w1(32'h3aabc697),
	.w2(32'hba05c2f7),
	.w3(32'h3a5ebe91),
	.w4(32'h39e003d1),
	.w5(32'hb89269b7),
	.w6(32'h3a3779b5),
	.w7(32'hba50189f),
	.w8(32'hbab7ee7d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb5436),
	.w1(32'h39b31bae),
	.w2(32'hb9db5301),
	.w3(32'h3945e843),
	.w4(32'h3a22fac9),
	.w5(32'h39b13506),
	.w6(32'h39de4bad),
	.w7(32'h3a13e2a8),
	.w8(32'h39dd84ec),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e7b5),
	.w1(32'h3acf4eb3),
	.w2(32'hbb00ddc1),
	.w3(32'hbbc01765),
	.w4(32'h3b1c6f47),
	.w5(32'h3b3a9e65),
	.w6(32'hbc09d16a),
	.w7(32'h3858b649),
	.w8(32'h3b537477),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61d89d),
	.w1(32'h3a3c8b1f),
	.w2(32'hba099c85),
	.w3(32'hba9df4d3),
	.w4(32'h3a2f4857),
	.w5(32'h37f9f0b0),
	.w6(32'h3ab06a90),
	.w7(32'h3a859821),
	.w8(32'h39da44a2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39549079),
	.w1(32'hb9f28104),
	.w2(32'h38e28b7d),
	.w3(32'h3987c782),
	.w4(32'hba2d6625),
	.w5(32'hb98d1a9b),
	.w6(32'hba14f8d9),
	.w7(32'hb8d7460b),
	.w8(32'hb80efec3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db7c39),
	.w1(32'h3a85902c),
	.w2(32'h3a25e759),
	.w3(32'hb9db48db),
	.w4(32'h39d91d1c),
	.w5(32'h3a34f11d),
	.w6(32'h3a85ca77),
	.w7(32'h3a8ea783),
	.w8(32'h388cbcb3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b026e),
	.w1(32'h3a835157),
	.w2(32'h3a4e74e4),
	.w3(32'h3b422433),
	.w4(32'hba14b5e8),
	.w5(32'hba1736fe),
	.w6(32'h3ac2fe86),
	.w7(32'h3ace25b2),
	.w8(32'hb9050ef7),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4b1c2),
	.w1(32'h3a6b5828),
	.w2(32'hb7b918f6),
	.w3(32'hba3cd874),
	.w4(32'h3a5e2753),
	.w5(32'hba25df8d),
	.w6(32'hbb4103b9),
	.w7(32'h39ae0b28),
	.w8(32'hb9779c0b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06489b),
	.w1(32'h3ac5ff97),
	.w2(32'h3a8a303e),
	.w3(32'h3b24072f),
	.w4(32'h3acaf6c1),
	.w5(32'h3b253327),
	.w6(32'h3b3f7550),
	.w7(32'h3b1d729e),
	.w8(32'h3b1c4430),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901c03d),
	.w1(32'h38a5095e),
	.w2(32'h39f83126),
	.w3(32'hb851ef86),
	.w4(32'hb9e9060b),
	.w5(32'hb9e18594),
	.w6(32'h39401ef8),
	.w7(32'h3977d2bd),
	.w8(32'hb904ecad),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af58154),
	.w1(32'h3a9c8c6f),
	.w2(32'h3a0eb319),
	.w3(32'hb90124de),
	.w4(32'hbb16082a),
	.w5(32'h378b7992),
	.w6(32'h3b454efe),
	.w7(32'hba573b74),
	.w8(32'hbb0212ff),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1fb8e),
	.w1(32'h3a6df6cd),
	.w2(32'hb999071f),
	.w3(32'hbb168a70),
	.w4(32'h39e100f8),
	.w5(32'hb8d0e9f1),
	.w6(32'h3a289d1c),
	.w7(32'h3b067353),
	.w8(32'h3a81c6fa),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3520),
	.w1(32'hbabe754a),
	.w2(32'hba2aa33b),
	.w3(32'h3b6c42ac),
	.w4(32'hbb124769),
	.w5(32'hba94dbf2),
	.w6(32'h3bca22f9),
	.w7(32'h3a915f31),
	.w8(32'hbb1c297c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1473a),
	.w1(32'h3b9ea3b7),
	.w2(32'hbb2ac32e),
	.w3(32'hbbf2c377),
	.w4(32'h3ab4af16),
	.w5(32'h39a97531),
	.w6(32'hbbce7f3b),
	.w7(32'hbb151f3f),
	.w8(32'h39e5e08b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b38a8),
	.w1(32'hb99991e9),
	.w2(32'hba5e67c7),
	.w3(32'hbaef0e26),
	.w4(32'hba9c2cff),
	.w5(32'hba957746),
	.w6(32'hbb048d0b),
	.w7(32'hba29a200),
	.w8(32'h394bcbe3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9005ec),
	.w1(32'hba9e289b),
	.w2(32'hba8f2f64),
	.w3(32'hba78f443),
	.w4(32'hba654a9d),
	.w5(32'hba127277),
	.w6(32'hba322153),
	.w7(32'hba3cd9a3),
	.w8(32'hba6362df),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b716f),
	.w1(32'h3ae45994),
	.w2(32'hbb03c67e),
	.w3(32'h39b4bea2),
	.w4(32'h3ace3b74),
	.w5(32'hba8f8c52),
	.w6(32'h362d5f4e),
	.w7(32'h3a8b163e),
	.w8(32'hb926aa98),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1a08d),
	.w1(32'h395aa2ce),
	.w2(32'hba935145),
	.w3(32'hbafb5267),
	.w4(32'hba0fc2c2),
	.w5(32'hba7bedc7),
	.w6(32'hbb983f29),
	.w7(32'hbae1de0a),
	.w8(32'hbaa15451),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388bd1ee),
	.w1(32'h39dde126),
	.w2(32'h39902e42),
	.w3(32'hba4a45c3),
	.w4(32'hb9dd6a19),
	.w5(32'h399bf01b),
	.w6(32'hbb34e4dc),
	.w7(32'hb9dfce42),
	.w8(32'h3a7aeaa7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a028c78),
	.w1(32'hb84513a4),
	.w2(32'h3a17a0ef),
	.w3(32'h39e9198e),
	.w4(32'hbac131b0),
	.w5(32'hba5b88d5),
	.w6(32'h3aa090ab),
	.w7(32'hb9526b94),
	.w8(32'hbabaa9ca),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbc652),
	.w1(32'hb4d6898d),
	.w2(32'h39c5e70d),
	.w3(32'hba0c68bb),
	.w4(32'hba04b605),
	.w5(32'h39b50e47),
	.w6(32'hb96a882a),
	.w7(32'h390854d7),
	.w8(32'h399bd4a5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a972d63),
	.w1(32'h3abb28e5),
	.w2(32'h3b17cd4c),
	.w3(32'h3af48eaa),
	.w4(32'hb9278464),
	.w5(32'h3a0d387b),
	.w6(32'h3b6c8cbc),
	.w7(32'h3b3278f3),
	.w8(32'hb92ba44a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec5126),
	.w1(32'hba5edade),
	.w2(32'hb929ff70),
	.w3(32'h3a554c28),
	.w4(32'hb9c96b75),
	.w5(32'h3787f84a),
	.w6(32'hb9178039),
	.w7(32'h38ba1bcf),
	.w8(32'h3a75d824),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ae99a),
	.w1(32'h39a90048),
	.w2(32'hba860871),
	.w3(32'hba01d8d9),
	.w4(32'h39885060),
	.w5(32'hb988cc20),
	.w6(32'hbb2ea668),
	.w7(32'h3abb0a05),
	.w8(32'h3a316aef),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ed45e),
	.w1(32'h38f2d95f),
	.w2(32'h39420228),
	.w3(32'h3a218156),
	.w4(32'hb7982905),
	.w5(32'h38c8179a),
	.w6(32'h3a012ddd),
	.w7(32'h3a23030d),
	.w8(32'h39d428b1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b147d6),
	.w1(32'hba0609ba),
	.w2(32'h3b2dbbbe),
	.w3(32'h3abe677e),
	.w4(32'hbaff18fb),
	.w5(32'h3abca09e),
	.w6(32'h3b709a4e),
	.w7(32'h3b067a8e),
	.w8(32'h3b16a47c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2ddb5),
	.w1(32'hba68a78a),
	.w2(32'h38587078),
	.w3(32'hb8e42e2f),
	.w4(32'hbab834b4),
	.w5(32'hba6d22d2),
	.w6(32'hbaa3b28d),
	.w7(32'hba78abe5),
	.w8(32'hba90b281),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74df28),
	.w1(32'hba3b453c),
	.w2(32'hb991e39d),
	.w3(32'hba4e76a1),
	.w4(32'hba126b01),
	.w5(32'hb9cf2fca),
	.w6(32'hba737b35),
	.w7(32'hba5c09cc),
	.w8(32'hb9a3c3b6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1947e8),
	.w1(32'hb988f875),
	.w2(32'hb9b294aa),
	.w3(32'hbb6cd5dd),
	.w4(32'hb9a320fc),
	.w5(32'h394caea0),
	.w6(32'hbb86990f),
	.w7(32'hba80c66e),
	.w8(32'h3a27cffb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b956),
	.w1(32'hba9a9004),
	.w2(32'hbb390e07),
	.w3(32'h3bcddb28),
	.w4(32'hba87cff5),
	.w5(32'hbaa7dba1),
	.w6(32'h3c2b78f5),
	.w7(32'h3bde15be),
	.w8(32'h3b21bbf5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47eaa9),
	.w1(32'hba7569a1),
	.w2(32'hb91b5175),
	.w3(32'hba016b39),
	.w4(32'hba65e003),
	.w5(32'hba050059),
	.w6(32'hba0b4c84),
	.w7(32'hba319ab4),
	.w8(32'hba75f6f7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cffb2),
	.w1(32'hbacb8a52),
	.w2(32'hbb149a4f),
	.w3(32'hbb4d5c7c),
	.w4(32'h3830cf77),
	.w5(32'hb844cee8),
	.w6(32'hbb5fc824),
	.w7(32'hba9b4216),
	.w8(32'h3a63b50a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e830a),
	.w1(32'h3b186413),
	.w2(32'hba0bd1f7),
	.w3(32'hba659bbd),
	.w4(32'h3a464ca9),
	.w5(32'h3ab0f000),
	.w6(32'hb90198a4),
	.w7(32'hba0a168c),
	.w8(32'h3745c588),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b4e1),
	.w1(32'h39ecded0),
	.w2(32'h3b922584),
	.w3(32'h3b2327bd),
	.w4(32'hbaf0e9b1),
	.w5(32'h3bcc2552),
	.w6(32'h3b1aa413),
	.w7(32'hba10a346),
	.w8(32'h3b628280),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c44dd),
	.w1(32'hbaca6870),
	.w2(32'h38f11a56),
	.w3(32'hba9bede2),
	.w4(32'hba908c7f),
	.w5(32'hba8038b1),
	.w6(32'h391ae10d),
	.w7(32'hb9f016e5),
	.w8(32'h38e2f184),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887c72),
	.w1(32'hb80bafae),
	.w2(32'h3a9e9ff2),
	.w3(32'h3911866e),
	.w4(32'hba9e1847),
	.w5(32'h399be6dc),
	.w6(32'h3b8b2207),
	.w7(32'h3ac77ff9),
	.w8(32'hbb04f342),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9313887),
	.w1(32'h3a8d8306),
	.w2(32'h3af79e5d),
	.w3(32'h399303f2),
	.w4(32'h39984dd6),
	.w5(32'h3a962b92),
	.w6(32'hb9a396ce),
	.w7(32'h3a75a659),
	.w8(32'h391c41e0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8a39),
	.w1(32'hbaccca38),
	.w2(32'hba860808),
	.w3(32'hbb41d8e6),
	.w4(32'hbb12a2c0),
	.w5(32'hb9e55b1d),
	.w6(32'hba6497ea),
	.w7(32'hbb214f16),
	.w8(32'hbaf1105f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39394d2f),
	.w1(32'hb95eb043),
	.w2(32'hb981e376),
	.w3(32'h38e111ce),
	.w4(32'hb8a4e9cb),
	.w5(32'hb9ad7b32),
	.w6(32'hb9624a79),
	.w7(32'hb9b57d5a),
	.w8(32'hba108495),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb0432),
	.w1(32'h398b4301),
	.w2(32'hb8c7c7ca),
	.w3(32'hb9ad667e),
	.w4(32'hb9e02a65),
	.w5(32'hba2e4850),
	.w6(32'h3a266eb7),
	.w7(32'h3a0254b0),
	.w8(32'h3a39cc12),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392df3a4),
	.w1(32'h3af56b10),
	.w2(32'hb947c57a),
	.w3(32'hbaaacdcf),
	.w4(32'h3ae7e14f),
	.w5(32'h3a69fae4),
	.w6(32'hb9991c0c),
	.w7(32'h3af388e5),
	.w8(32'h3ac6d7ad),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf949d),
	.w1(32'hbb039231),
	.w2(32'h3ad49be0),
	.w3(32'hba75d324),
	.w4(32'hbadb14e2),
	.w5(32'h3abc71df),
	.w6(32'hbb50ee0e),
	.w7(32'hb959c910),
	.w8(32'h3ae03e5b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa80647),
	.w1(32'h390ffbf7),
	.w2(32'hb9e4bc88),
	.w3(32'hbaac11e8),
	.w4(32'hba085caf),
	.w5(32'hba699006),
	.w6(32'h39d62b3e),
	.w7(32'hb29a95b0),
	.w8(32'hb9d13a90),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c1f50),
	.w1(32'h39ae9393),
	.w2(32'h392346dc),
	.w3(32'hb9e7afea),
	.w4(32'h394f464e),
	.w5(32'h37c19c52),
	.w6(32'h38c5febb),
	.w7(32'h380bdf76),
	.w8(32'h37c5c6b6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9919f),
	.w1(32'hba5debd5),
	.w2(32'hbaee0ce9),
	.w3(32'hba201cdc),
	.w4(32'hba34b3e0),
	.w5(32'hba97b019),
	.w6(32'hba7a39c1),
	.w7(32'h39553872),
	.w8(32'h3887064a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab62e92),
	.w1(32'hba8dceb7),
	.w2(32'hbb13ebf9),
	.w3(32'hb962d2f3),
	.w4(32'hbb241f13),
	.w5(32'hbaa28324),
	.w6(32'hbaa12f54),
	.w7(32'hba75b4cb),
	.w8(32'hbacb9419),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eef71),
	.w1(32'h39ec03e9),
	.w2(32'hbb3a2ff6),
	.w3(32'h3ba4266b),
	.w4(32'hb98fe664),
	.w5(32'hb9ab7396),
	.w6(32'h3bcd4575),
	.w7(32'h3b433628),
	.w8(32'h39567d2e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d41a1),
	.w1(32'hba381a6a),
	.w2(32'hb9191ec8),
	.w3(32'hba6d71e8),
	.w4(32'hba912b88),
	.w5(32'hba3cd283),
	.w6(32'hb9ce9dbd),
	.w7(32'hba2a1ef1),
	.w8(32'hb9d51e39),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99df7b),
	.w1(32'h3a03ec47),
	.w2(32'h3a4f91bf),
	.w3(32'h3bde7bdf),
	.w4(32'hba1397a1),
	.w5(32'h393d2e1d),
	.w6(32'h3c29b110),
	.w7(32'h3b311b63),
	.w8(32'hb9e7a23d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba686e91),
	.w1(32'h3ab22a99),
	.w2(32'hbb8f0b0b),
	.w3(32'hbc009dd3),
	.w4(32'hbb1f4043),
	.w5(32'hbb632766),
	.w6(32'hbc030ae3),
	.w7(32'hbbc0d145),
	.w8(32'hb9e95be9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2531d),
	.w1(32'h384a14dd),
	.w2(32'hba609e32),
	.w3(32'h39e70a9e),
	.w4(32'hb94bcdd3),
	.w5(32'hba1fa0b1),
	.w6(32'h3b102233),
	.w7(32'h378b3249),
	.w8(32'hb994cee2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9961b9e),
	.w1(32'h3a51d195),
	.w2(32'hba8244d2),
	.w3(32'hb9a2d8ec),
	.w4(32'h3a63a45d),
	.w5(32'hb93854db),
	.w6(32'h3a984510),
	.w7(32'h3872ea44),
	.w8(32'hba5d41ae),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882d745),
	.w1(32'h39bdf70f),
	.w2(32'h3a3bd6a7),
	.w3(32'hb9f5810a),
	.w4(32'h3a118bfb),
	.w5(32'h3a1a225a),
	.w6(32'h3a3539fd),
	.w7(32'h3a27af52),
	.w8(32'h3a3278cf),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcc8bf),
	.w1(32'hb79e2475),
	.w2(32'h3858085a),
	.w3(32'h39f460b7),
	.w4(32'hb99fae89),
	.w5(32'h398910dc),
	.w6(32'hb7bf8428),
	.w7(32'h3992af32),
	.w8(32'h3958792f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fd035),
	.w1(32'hbb0716ef),
	.w2(32'hbb49897b),
	.w3(32'h3aebe8a4),
	.w4(32'hbadc6b04),
	.w5(32'hba74880f),
	.w6(32'h3b9c8d3f),
	.w7(32'h3b4eb174),
	.w8(32'h393cfab0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae15dc8),
	.w1(32'hbb205616),
	.w2(32'hba7d9748),
	.w3(32'hb93a986e),
	.w4(32'hbb2696a4),
	.w5(32'hbab9659d),
	.w6(32'hba2e9aef),
	.w7(32'hba8a0ab6),
	.w8(32'hbacc29a9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c8d53),
	.w1(32'h3af92993),
	.w2(32'hba5a5015),
	.w3(32'hbb080661),
	.w4(32'h3b329467),
	.w5(32'h3a75c90e),
	.w6(32'hbb179e84),
	.w7(32'h3b3e80e0),
	.w8(32'h3b61e12b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e6b37),
	.w1(32'hba3ecd39),
	.w2(32'hba052c63),
	.w3(32'hba394e02),
	.w4(32'hba3611e7),
	.w5(32'hba6fa313),
	.w6(32'hba923339),
	.w7(32'h37ed83e1),
	.w8(32'hb88d1ec1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ae25c),
	.w1(32'h3a83d098),
	.w2(32'h3ab9b3d5),
	.w3(32'h3b61ffe1),
	.w4(32'h3a437e4a),
	.w5(32'h3af2c645),
	.w6(32'h3be4ca93),
	.w7(32'h3b9e8691),
	.w8(32'h3b4b4217),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b576e47),
	.w1(32'h39f7d244),
	.w2(32'hba273907),
	.w3(32'h3b8d132a),
	.w4(32'hba00d297),
	.w5(32'hbb17d02a),
	.w6(32'h3b0afae5),
	.w7(32'h39e47779),
	.w8(32'hbab16a8b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c63ba),
	.w1(32'hb9a18aac),
	.w2(32'hb8ab5b39),
	.w3(32'hb96a00e1),
	.w4(32'hb9cbbaca),
	.w5(32'hb9e86a61),
	.w6(32'hb8f07949),
	.w7(32'hb9a3152d),
	.w8(32'hb96991f6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c0773),
	.w1(32'hbaa4bd7c),
	.w2(32'h39a6b63e),
	.w3(32'h3a466c91),
	.w4(32'hba1ab154),
	.w5(32'hba26ee1d),
	.w6(32'h391b1bbd),
	.w7(32'h39e6e3de),
	.w8(32'h3a2b7f1d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba429962),
	.w1(32'h38a2c3dd),
	.w2(32'h39ad11c9),
	.w3(32'hba269d71),
	.w4(32'h36576c7b),
	.w5(32'h38686a06),
	.w6(32'h3959842c),
	.w7(32'h39e60865),
	.w8(32'h38f30e4d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f5c36),
	.w1(32'h37fa46fd),
	.w2(32'h3aa8a714),
	.w3(32'h3a975c08),
	.w4(32'hba35820d),
	.w5(32'h3958b1ae),
	.w6(32'h3aca4c3a),
	.w7(32'h3adf8a36),
	.w8(32'h3a44a9a4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee1b42),
	.w1(32'h3b0481cf),
	.w2(32'hbb8d5b1a),
	.w3(32'hbb427871),
	.w4(32'hb8ecd4ac),
	.w5(32'hbb818858),
	.w6(32'hbb8170a3),
	.w7(32'hb8df5f9d),
	.w8(32'hba0cc6b9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e74db),
	.w1(32'hba80945f),
	.w2(32'hbb532c21),
	.w3(32'hbb1a2199),
	.w4(32'hb9c545ea),
	.w5(32'hbac14e81),
	.w6(32'hbb057566),
	.w7(32'hb9bfa9cf),
	.w8(32'hba2bfe1e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f10325),
	.w1(32'hbaa71c53),
	.w2(32'hba8b0ba8),
	.w3(32'hb9ec3b8d),
	.w4(32'hbabfc5f1),
	.w5(32'hbac3b90c),
	.w6(32'hba8d7d76),
	.w7(32'hba9cd371),
	.w8(32'hba8a56af),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be6fa),
	.w1(32'h3ab3f326),
	.w2(32'hbb39aa6d),
	.w3(32'hbb6c1c88),
	.w4(32'h3b632e86),
	.w5(32'h3a7f0670),
	.w6(32'hbb86454f),
	.w7(32'h3a223fc0),
	.w8(32'h3ab73d39),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9fe9),
	.w1(32'h3a0b9457),
	.w2(32'h3ae8bd52),
	.w3(32'h3b36bd91),
	.w4(32'hb9bc216e),
	.w5(32'h3a8b2924),
	.w6(32'h3ad6f1cf),
	.w7(32'h3a9c1c16),
	.w8(32'h396d4a37),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b598791),
	.w1(32'h3ada97b2),
	.w2(32'h39935227),
	.w3(32'h3b1a176d),
	.w4(32'h3ad1340b),
	.w5(32'h3a8217da),
	.w6(32'h3b0361db),
	.w7(32'h3af5c471),
	.w8(32'h3a4fca94),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56699e),
	.w1(32'hba83f07c),
	.w2(32'h39d20c50),
	.w3(32'hba2430db),
	.w4(32'hbabb391d),
	.w5(32'hba789ad4),
	.w6(32'hba7ccad7),
	.w7(32'hb9e82de7),
	.w8(32'hba796c01),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b2387),
	.w1(32'h3a2eeab5),
	.w2(32'h3a3f2b27),
	.w3(32'hbab10175),
	.w4(32'h393ba150),
	.w5(32'h3a249a02),
	.w6(32'hba6949a8),
	.w7(32'h392e822d),
	.w8(32'h39038d4e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238845),
	.w1(32'hbb57c2ff),
	.w2(32'hbbe0ce6a),
	.w3(32'h3bd7c6b8),
	.w4(32'hbb1abb38),
	.w5(32'hbb4db869),
	.w6(32'h3c0ecc45),
	.w7(32'h3b92baab),
	.w8(32'h3b02cafd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba772511),
	.w1(32'hba9e8cd5),
	.w2(32'hba0ce34c),
	.w3(32'h3aa939b3),
	.w4(32'hba2c5748),
	.w5(32'hb845153f),
	.w6(32'h3b874a09),
	.w7(32'h3b16c2c0),
	.w8(32'h39efec21),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39954e63),
	.w1(32'hba877487),
	.w2(32'hbb243452),
	.w3(32'h38a825ae),
	.w4(32'hba47020d),
	.w5(32'hbaf1b15c),
	.w6(32'hbb0a9069),
	.w7(32'hb969c8f2),
	.w8(32'hba7228be),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72ac6e),
	.w1(32'hbb8004c5),
	.w2(32'hbbeb85e2),
	.w3(32'h3a439274),
	.w4(32'hbbe57f2e),
	.w5(32'hbbadd728),
	.w6(32'hba50075a),
	.w7(32'hbb6ce111),
	.w8(32'hbb58277c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5353a),
	.w1(32'hb91c55f6),
	.w2(32'h3a74fc3e),
	.w3(32'hb9f207ad),
	.w4(32'hb9370994),
	.w5(32'h3a055cb8),
	.w6(32'hb865036f),
	.w7(32'h39f1f98f),
	.w8(32'h3a063235),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad109f0),
	.w1(32'hba47a205),
	.w2(32'h3a9ae428),
	.w3(32'hb9d79c23),
	.w4(32'h39cf4b85),
	.w5(32'h3a25e590),
	.w6(32'h3a2afa1a),
	.w7(32'h3a17e9df),
	.w8(32'h3ac1f784),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e69b2),
	.w1(32'hb9ea3e8b),
	.w2(32'hbc056733),
	.w3(32'h3c8b39d4),
	.w4(32'hbb709db4),
	.w5(32'hbbcb42e3),
	.w6(32'h3c85d74a),
	.w7(32'h3c6a07d5),
	.w8(32'h3a4e75c7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ad439),
	.w1(32'hb7126d54),
	.w2(32'h3abfa2c8),
	.w3(32'h3bd2bf49),
	.w4(32'hbafa944c),
	.w5(32'hb9c10f54),
	.w6(32'h3c22cddd),
	.w7(32'h3b3521db),
	.w8(32'hba0ec117),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1ee81),
	.w1(32'hbb20bece),
	.w2(32'hb9374473),
	.w3(32'h3c0a292c),
	.w4(32'hbb3f7a7d),
	.w5(32'hbb4ff8cc),
	.w6(32'h3c2258d7),
	.w7(32'h3bdad333),
	.w8(32'hbb0363a7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf3193),
	.w1(32'hba3efa20),
	.w2(32'hba92ce3a),
	.w3(32'hbb330166),
	.w4(32'hb970f949),
	.w5(32'hba0699a8),
	.w6(32'hbb82a564),
	.w7(32'hb9ff7f2d),
	.w8(32'h3a98e569),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49cb38),
	.w1(32'h3a16accc),
	.w2(32'hbb011fe6),
	.w3(32'hbbd453ad),
	.w4(32'hb6b7680e),
	.w5(32'hb9a8bf1a),
	.w6(32'hbc04bc91),
	.w7(32'hba9c372f),
	.w8(32'h3ac3a13a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f26dc2),
	.w1(32'hba0e4caa),
	.w2(32'hb770c84d),
	.w3(32'hb9aeddfd),
	.w4(32'hba4ecc8d),
	.w5(32'hba2bd50a),
	.w6(32'hba4273c7),
	.w7(32'hba38464e),
	.w8(32'hba8d4444),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ac669),
	.w1(32'hba984ada),
	.w2(32'hba336df9),
	.w3(32'hba7d63d9),
	.w4(32'hba83d192),
	.w5(32'hb9123a27),
	.w6(32'hba9511cd),
	.w7(32'hbac4ef62),
	.w8(32'hba969b94),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c36b21),
	.w1(32'h3963e667),
	.w2(32'h3a40d05d),
	.w3(32'h3828b489),
	.w4(32'hb811afa0),
	.w5(32'h39005b7c),
	.w6(32'h3b7d94f0),
	.w7(32'h3b3c7295),
	.w8(32'h3b56d106),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99c0ad),
	.w1(32'h39fe2f50),
	.w2(32'hba73f023),
	.w3(32'h3a87810b),
	.w4(32'h392c8f1e),
	.w5(32'hb97a583f),
	.w6(32'h39fd84e8),
	.w7(32'hb974b06c),
	.w8(32'h38c5df84),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95cb20a),
	.w1(32'hbb44a531),
	.w2(32'h3a417b7b),
	.w3(32'hb989748e),
	.w4(32'hbb3287b4),
	.w5(32'hb9e2455a),
	.w6(32'h3ac608fc),
	.w7(32'hba3282d3),
	.w8(32'hb952f588),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23369e),
	.w1(32'hbaf99980),
	.w2(32'h3a78616d),
	.w3(32'h3a4da960),
	.w4(32'hbaf33c33),
	.w5(32'h3a50819c),
	.w6(32'hba4d882a),
	.w7(32'h3b34a9f4),
	.w8(32'h3adcb17a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d5393),
	.w1(32'h3ac52725),
	.w2(32'hba92f4ff),
	.w3(32'hb839a40c),
	.w4(32'h3a6dcac3),
	.w5(32'h39963e69),
	.w6(32'h3b062b8c),
	.w7(32'h3b122657),
	.w8(32'h3a7453ee),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66d359),
	.w1(32'h3837a00c),
	.w2(32'hbafc467e),
	.w3(32'h395e2d28),
	.w4(32'hb915cc15),
	.w5(32'hba483eb3),
	.w6(32'h3aa1d043),
	.w7(32'h382a49b1),
	.w8(32'hba17f0be),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73f6e),
	.w1(32'hbb7afed1),
	.w2(32'hbb6a7c43),
	.w3(32'h3c2f1ae7),
	.w4(32'hbb8f70d6),
	.w5(32'hbbd3a87a),
	.w6(32'h3c885fa5),
	.w7(32'h3b9cc5a7),
	.w8(32'hbb74a3e9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0d8ec),
	.w1(32'hb6664a66),
	.w2(32'h3ab3f537),
	.w3(32'h3ab5a406),
	.w4(32'hba52c4ec),
	.w5(32'hb9b299ce),
	.w6(32'h3b3b8b57),
	.w7(32'h3a2ec821),
	.w8(32'hba27333b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c1b1e),
	.w1(32'hb920fead),
	.w2(32'hb9c4d1bd),
	.w3(32'hba36a5e3),
	.w4(32'h38d04509),
	.w5(32'hb89f9b98),
	.w6(32'hb82be7f8),
	.w7(32'hb921082e),
	.w8(32'hb90cf492),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ee12e),
	.w1(32'hb8e6abb9),
	.w2(32'h38a13e99),
	.w3(32'h3b764ecc),
	.w4(32'hb93ab36e),
	.w5(32'hba30b413),
	.w6(32'h3bd7cf5f),
	.w7(32'h3b5255ff),
	.w8(32'h397756e6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb605e),
	.w1(32'hba487681),
	.w2(32'hb97ab178),
	.w3(32'h38de6e50),
	.w4(32'hbab54cae),
	.w5(32'hba95180c),
	.w6(32'hbabded5d),
	.w7(32'hbaa4848b),
	.w8(32'hbac946e9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cafc2),
	.w1(32'hb99aa040),
	.w2(32'h3949a765),
	.w3(32'hba4432bb),
	.w4(32'hb9ca7057),
	.w5(32'hba284d2b),
	.w6(32'h38d71334),
	.w7(32'hb801081f),
	.w8(32'hba6c6ebe),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc71dc),
	.w1(32'hb97bc01f),
	.w2(32'hb9ee07c6),
	.w3(32'hba0eea82),
	.w4(32'hb6e73a9d),
	.w5(32'hb9abae84),
	.w6(32'hb88fb07d),
	.w7(32'hb9955f75),
	.w8(32'hb9bf9108),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9faa55f),
	.w1(32'hba80c9ac),
	.w2(32'hbada3bb2),
	.w3(32'hb9e1f88e),
	.w4(32'hbaace808),
	.w5(32'hbaf1cdc8),
	.w6(32'hba27e574),
	.w7(32'hba697a33),
	.w8(32'hba4d6d5f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06d38f),
	.w1(32'hbac42b16),
	.w2(32'hbb1a1707),
	.w3(32'hbb520900),
	.w4(32'hbae3c360),
	.w5(32'hbac68e88),
	.w6(32'hbb312c81),
	.w7(32'hba96ec54),
	.w8(32'hba2f483a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972a88a),
	.w1(32'hba9a9243),
	.w2(32'h39166572),
	.w3(32'hbb2ae6d2),
	.w4(32'hbb547c39),
	.w5(32'h3b2fd479),
	.w6(32'h3a5d6bc2),
	.w7(32'hba8850c2),
	.w8(32'h3ae92602),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e2e06),
	.w1(32'hbb00f5e2),
	.w2(32'h39930181),
	.w3(32'h3b1a8776),
	.w4(32'hbb597b62),
	.w5(32'hbb032417),
	.w6(32'h3b76868d),
	.w7(32'h39ee4655),
	.w8(32'hbb1958d4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34640b),
	.w1(32'hbaa6c543),
	.w2(32'h3ab5f922),
	.w3(32'hb9c2731a),
	.w4(32'hbb6ee57b),
	.w5(32'h389f5d31),
	.w6(32'h3b5788eb),
	.w7(32'h39b9bab6),
	.w8(32'hba36114f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ce0ec),
	.w1(32'h3a275c9c),
	.w2(32'h394c0e84),
	.w3(32'hbaabd0a4),
	.w4(32'h3a09e3b6),
	.w5(32'h390af67f),
	.w6(32'h395ab120),
	.w7(32'h3800c7a8),
	.w8(32'hb924c45a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a63da8),
	.w1(32'hba123919),
	.w2(32'hba117590),
	.w3(32'h38d2141a),
	.w4(32'h39222784),
	.w5(32'hb9acb2f5),
	.w6(32'h38fb2282),
	.w7(32'hb9340add),
	.w8(32'hb915395f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5857ff),
	.w1(32'hba705d75),
	.w2(32'hba3135a1),
	.w3(32'hba2a24b9),
	.w4(32'hba3bec0e),
	.w5(32'hba178a85),
	.w6(32'hba383c7a),
	.w7(32'hba369898),
	.w8(32'hba235433),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47a246),
	.w1(32'hba46c952),
	.w2(32'hba2d798b),
	.w3(32'hba2bf789),
	.w4(32'hba11ec6c),
	.w5(32'hb9f7c282),
	.w6(32'hba1df219),
	.w7(32'hba29e7c4),
	.w8(32'hba36b377),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c34a8),
	.w1(32'hb847d385),
	.w2(32'h3b7cfcc1),
	.w3(32'hbb20f222),
	.w4(32'h3a1edbed),
	.w5(32'h3af60a6d),
	.w6(32'h3ab737b8),
	.w7(32'h39dd0baf),
	.w8(32'hb9c83d0c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39495091),
	.w1(32'h3a62ae54),
	.w2(32'h3a053767),
	.w3(32'hb9944370),
	.w4(32'h39e2b547),
	.w5(32'h39e969d9),
	.w6(32'h39eed373),
	.w7(32'h3a636efb),
	.w8(32'h39675f07),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b47fa),
	.w1(32'hb83209df),
	.w2(32'h3a87a1b7),
	.w3(32'h3a0b0114),
	.w4(32'h3998ce79),
	.w5(32'h3a6cd944),
	.w6(32'h3a1b0565),
	.w7(32'h3a4ad950),
	.w8(32'h3a25895c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3a6cd),
	.w1(32'h3ae2af9d),
	.w2(32'h3ac9ff92),
	.w3(32'h3adda8b2),
	.w4(32'h3afcd4b4),
	.w5(32'h3a662c2b),
	.w6(32'h3ab933c7),
	.w7(32'h3add7a03),
	.w8(32'h3ad824ec),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39798992),
	.w1(32'hb9e1ba15),
	.w2(32'hba076f59),
	.w3(32'h399361c7),
	.w4(32'hb9621d09),
	.w5(32'hba092b68),
	.w6(32'hb9afcb2d),
	.w7(32'hb9e58463),
	.w8(32'hba1d1edb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985a39a),
	.w1(32'hb986324b),
	.w2(32'h38c1b2e2),
	.w3(32'h397c45a4),
	.w4(32'h377a4cb0),
	.w5(32'hb813789e),
	.w6(32'h3b2c4bb8),
	.w7(32'h3aaf831d),
	.w8(32'h35d10264),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9727af),
	.w1(32'hbaf0a6d5),
	.w2(32'h39a2a92a),
	.w3(32'hba690aa4),
	.w4(32'hbb06af3f),
	.w5(32'hba9a07f1),
	.w6(32'hbb40f5a5),
	.w7(32'hbb24493e),
	.w8(32'hbac5e7a1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a492d03),
	.w1(32'h3acb7edc),
	.w2(32'h3be7cb8c),
	.w3(32'hbb2bf3d4),
	.w4(32'h3ae0c584),
	.w5(32'h3bf37a37),
	.w6(32'h3b0d8558),
	.w7(32'h3b55df96),
	.w8(32'h3b8e199f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8ee88),
	.w1(32'h38c96856),
	.w2(32'h397adff4),
	.w3(32'hb98a0a97),
	.w4(32'h394a7e84),
	.w5(32'h385457c1),
	.w6(32'h3928246f),
	.w7(32'h392aac7d),
	.w8(32'h389ce597),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a312da6),
	.w1(32'hbad310ed),
	.w2(32'hbba1fc90),
	.w3(32'h3b34283c),
	.w4(32'hbab39c5a),
	.w5(32'hbb4af9eb),
	.w6(32'h3b3df5d2),
	.w7(32'h3addd688),
	.w8(32'h39bf3f81),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule