module layer_10_featuremap_416(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b343100),
	.w1(32'h3b7166a6),
	.w2(32'h3a399c1c),
	.w3(32'h3c1adeea),
	.w4(32'h3bd904eb),
	.w5(32'h3b66a7cc),
	.w6(32'h38ba7618),
	.w7(32'hb8d05950),
	.w8(32'h3b65351c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45429b),
	.w1(32'hbc854a12),
	.w2(32'hbbecaeea),
	.w3(32'hbb00e085),
	.w4(32'hbc853aa2),
	.w5(32'h3cfd7225),
	.w6(32'h3b263747),
	.w7(32'hbc44c22d),
	.w8(32'hbb7120fe),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c5fd),
	.w1(32'hbc2d1747),
	.w2(32'hbc5cf113),
	.w3(32'h3c130bae),
	.w4(32'hbc006bc0),
	.w5(32'hbc17a53e),
	.w6(32'h3af935a1),
	.w7(32'hbc674b61),
	.w8(32'h3bf2c837),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c5575),
	.w1(32'h381db65a),
	.w2(32'hbc77b95d),
	.w3(32'hba20e3ec),
	.w4(32'hb910b949),
	.w5(32'h3bebe286),
	.w6(32'hbb6eac9b),
	.w7(32'hbc47eda8),
	.w8(32'hbc263aca),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2caabc),
	.w1(32'h3c212e9f),
	.w2(32'hbbae11d2),
	.w3(32'h3bcc2ddc),
	.w4(32'h3c750255),
	.w5(32'hbca05185),
	.w6(32'h3bdf2b3a),
	.w7(32'h3bec4c13),
	.w8(32'h3b9048cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebec6f),
	.w1(32'h3b3a969d),
	.w2(32'hbae0a5a2),
	.w3(32'hbc02a749),
	.w4(32'hbb846205),
	.w5(32'hbba383b1),
	.w6(32'hbb0aa94d),
	.w7(32'hbbb35ac8),
	.w8(32'hbc473396),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe012d3),
	.w1(32'hbb2b8a7e),
	.w2(32'h3be3e8d0),
	.w3(32'hbb99cf20),
	.w4(32'hbacf2647),
	.w5(32'hbc0bbf0e),
	.w6(32'hbb3ca58c),
	.w7(32'h3b3eba26),
	.w8(32'h39314a4e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95ba1b),
	.w1(32'h3c9181ca),
	.w2(32'hbbc8cf7c),
	.w3(32'h3abfa6f0),
	.w4(32'h3c389407),
	.w5(32'hbc2823c6),
	.w6(32'h3b9f60b5),
	.w7(32'h3b10c382),
	.w8(32'hbb1302a5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c6748),
	.w1(32'hbbe76167),
	.w2(32'hbbc281a4),
	.w3(32'hba20a41b),
	.w4(32'hba59ad3b),
	.w5(32'h3bcfc6fc),
	.w6(32'hb9af4450),
	.w7(32'hbb6ea481),
	.w8(32'hbb86e4c9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3d58),
	.w1(32'h38c1dcf9),
	.w2(32'hbb302e8c),
	.w3(32'hbba2f607),
	.w4(32'h3b9306ae),
	.w5(32'h3adfc123),
	.w6(32'hbc110ba5),
	.w7(32'hbbb43a1a),
	.w8(32'h3bd870fd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf73bdc),
	.w1(32'hbb7ce355),
	.w2(32'hbbc6ffa9),
	.w3(32'hbc7bc07e),
	.w4(32'h3ba504a5),
	.w5(32'hbaafbfda),
	.w6(32'h3be947dd),
	.w7(32'hb9cff8f8),
	.w8(32'h3c052d06),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5459a5),
	.w1(32'h3bedf256),
	.w2(32'h3b19fb9c),
	.w3(32'hbad7e146),
	.w4(32'h3ab90efd),
	.w5(32'hbbdee355),
	.w6(32'hbae7422f),
	.w7(32'h3a32f1ed),
	.w8(32'hba86ff8f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb5e23),
	.w1(32'hbc3fe815),
	.w2(32'hbc1b6a96),
	.w3(32'h3851f29f),
	.w4(32'hbc3e87c7),
	.w5(32'h3ce0a158),
	.w6(32'h3b47d225),
	.w7(32'hbc7a4b58),
	.w8(32'h3b6e326e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf85c82),
	.w1(32'h3a8db4df),
	.w2(32'hbc43bd4e),
	.w3(32'hbb983903),
	.w4(32'h3bb5013e),
	.w5(32'hbc96b339),
	.w6(32'h3a2877b2),
	.w7(32'hbaa76ea0),
	.w8(32'h3b040186),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bab95),
	.w1(32'h3c024d28),
	.w2(32'h3c5b7d3b),
	.w3(32'hb9b260e4),
	.w4(32'h3babc0da),
	.w5(32'hbb973410),
	.w6(32'hbc2c12bb),
	.w7(32'h3b118f7d),
	.w8(32'h3c0ff0a1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1001fe),
	.w1(32'h3c35701c),
	.w2(32'h3b69579a),
	.w3(32'h3c7e6aee),
	.w4(32'h3c3fcb11),
	.w5(32'hbc40f3e3),
	.w6(32'h3c174510),
	.w7(32'h3c1d9275),
	.w8(32'h3b22bd23),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be49d0a),
	.w1(32'hbb324b0a),
	.w2(32'h3bef1c7b),
	.w3(32'h396e379c),
	.w4(32'hbb91566a),
	.w5(32'h3b29818c),
	.w6(32'h3bce2bc3),
	.w7(32'hbc06b365),
	.w8(32'hbbde8c74),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f3d1c),
	.w1(32'h3bf9baac),
	.w2(32'h3b29880e),
	.w3(32'h3c56c7cf),
	.w4(32'h3c068970),
	.w5(32'h3c5009f7),
	.w6(32'h3be27ebf),
	.w7(32'h3b35d375),
	.w8(32'h3b2197a5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003807),
	.w1(32'h3b7c9f91),
	.w2(32'hba68dd45),
	.w3(32'h399ff1cb),
	.w4(32'h3b1f8223),
	.w5(32'hbc90a0cb),
	.w6(32'h3a8a0f85),
	.w7(32'h3b210603),
	.w8(32'h3b60ee8b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80dd88),
	.w1(32'h3c015603),
	.w2(32'hbb299d94),
	.w3(32'h3bfa6aa2),
	.w4(32'hbb242d2d),
	.w5(32'hbb0b1db5),
	.w6(32'h3a695efa),
	.w7(32'h394b628c),
	.w8(32'h3bdf67da),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb113d86),
	.w1(32'h3b3c7dc5),
	.w2(32'h3b97984b),
	.w3(32'h3aa4c655),
	.w4(32'h3b8246a6),
	.w5(32'hbc1abda2),
	.w6(32'h398a5220),
	.w7(32'hb99a9e9b),
	.w8(32'h3bdcddb1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17c890),
	.w1(32'hbc3972ae),
	.w2(32'h3a391559),
	.w3(32'hbb9a8141),
	.w4(32'hbc850e58),
	.w5(32'hbb8141de),
	.w6(32'h3b93c29a),
	.w7(32'hbc5d469a),
	.w8(32'hbb2fb0b4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2358af),
	.w1(32'h3c748fb2),
	.w2(32'hba9f7f59),
	.w3(32'h3bd023bf),
	.w4(32'h3b6fd3a6),
	.w5(32'hbbc647e0),
	.w6(32'h3badab97),
	.w7(32'hba8a16ea),
	.w8(32'h3afeca0a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb982121),
	.w1(32'h3ae0615a),
	.w2(32'h3c4942a2),
	.w3(32'hbb729b61),
	.w4(32'hbbbf2fb6),
	.w5(32'h3b05dfc4),
	.w6(32'hbbe3be36),
	.w7(32'h3b3eca38),
	.w8(32'h3c638c7e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b119d92),
	.w1(32'h3a3b0c4d),
	.w2(32'hbbd0c2f8),
	.w3(32'hbc1ba1ef),
	.w4(32'hbb4824ae),
	.w5(32'hbc63f173),
	.w6(32'h3b979367),
	.w7(32'h3a177355),
	.w8(32'h398db9aa),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05955c),
	.w1(32'h3b768482),
	.w2(32'hb8ae2a17),
	.w3(32'h3c2d7d92),
	.w4(32'h3bb8e27e),
	.w5(32'hbc2015a7),
	.w6(32'hba227cb1),
	.w7(32'h3bd30d93),
	.w8(32'h3a8deafb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf4a3),
	.w1(32'h3b4b9cb1),
	.w2(32'h3c1681aa),
	.w3(32'hbb439095),
	.w4(32'hbb403f99),
	.w5(32'hbbd64c98),
	.w6(32'h3ac648a6),
	.w7(32'h3af14b6b),
	.w8(32'h3c13fa37),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fa874),
	.w1(32'hbbc6f8c9),
	.w2(32'hbb9d0e2b),
	.w3(32'hbb99234b),
	.w4(32'hbb523ebf),
	.w5(32'hbb8b6881),
	.w6(32'hbbe509c8),
	.w7(32'hbb89b929),
	.w8(32'h3aed9868),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7376),
	.w1(32'hbb885f37),
	.w2(32'hbc8584dc),
	.w3(32'h3c2c658b),
	.w4(32'hbc84e12c),
	.w5(32'hbb112fcc),
	.w6(32'h3b8e6fd6),
	.w7(32'hbc45590f),
	.w8(32'hbb968431),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67fcab),
	.w1(32'hbb690c3e),
	.w2(32'hbb42a685),
	.w3(32'hbc84ad6e),
	.w4(32'hbb63c976),
	.w5(32'hbb900010),
	.w6(32'hbb9cba09),
	.w7(32'hbb3c8a3f),
	.w8(32'hbb842dba),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe544),
	.w1(32'hbbb81713),
	.w2(32'hbb8ce193),
	.w3(32'hbc133685),
	.w4(32'h3aafac7f),
	.w5(32'hbaa4ee41),
	.w6(32'hbb121d20),
	.w7(32'h39ea7c0d),
	.w8(32'hbb90ef7d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49b5ee),
	.w1(32'hbc2a13e6),
	.w2(32'hbbd95a69),
	.w3(32'hbb3a399b),
	.w4(32'hbc273646),
	.w5(32'h3c441e9b),
	.w6(32'hbbebddaa),
	.w7(32'hbc5f2037),
	.w8(32'hb91461e2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20b999),
	.w1(32'hbbc44964),
	.w2(32'h3b6c4e79),
	.w3(32'hbaf87b4c),
	.w4(32'hbc32c779),
	.w5(32'h3b015000),
	.w6(32'hbb03fb71),
	.w7(32'hbab138f6),
	.w8(32'h3baeb566),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aa7a8),
	.w1(32'hbc12a99b),
	.w2(32'hbb641a1f),
	.w3(32'h3b25cce5),
	.w4(32'hbc514f3b),
	.w5(32'hbc3e6218),
	.w6(32'h3c58f591),
	.w7(32'hbb3fed27),
	.w8(32'h3b0ea4cb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37241c),
	.w1(32'hbb62b553),
	.w2(32'hbc6a3e51),
	.w3(32'h3c711063),
	.w4(32'hba6d9c17),
	.w5(32'hbc39e0e9),
	.w6(32'h3c1a2b15),
	.w7(32'hba3d75fa),
	.w8(32'hba76d900),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83f0f2),
	.w1(32'hbbdfaa38),
	.w2(32'h3bd6ba05),
	.w3(32'h3ba4d0b2),
	.w4(32'h3b6dafdc),
	.w5(32'h3d3177ec),
	.w6(32'h3b268eaa),
	.w7(32'hba23c797),
	.w8(32'h3be1e9f0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30455e),
	.w1(32'h3bbdcadc),
	.w2(32'h3bdbfec9),
	.w3(32'hbb5bb7e7),
	.w4(32'h3c13d0e9),
	.w5(32'h3c3eaeb9),
	.w6(32'hbb96c2a7),
	.w7(32'h3c1c67e2),
	.w8(32'h3c497914),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7eba1),
	.w1(32'hbbce73ce),
	.w2(32'h3b66beff),
	.w3(32'hbbd32b85),
	.w4(32'hbc3a3ddc),
	.w5(32'h3d4d7a43),
	.w6(32'h3ba53493),
	.w7(32'hbc6b452d),
	.w8(32'h3b55fd24),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3637c5),
	.w1(32'hbbc2c0df),
	.w2(32'hbbb21b26),
	.w3(32'hbc72d3e7),
	.w4(32'hbb9e859b),
	.w5(32'hbcc1877a),
	.w6(32'hbc1ff413),
	.w7(32'h39ae6123),
	.w8(32'hbb0a4cab),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73adce),
	.w1(32'h3b2c8703),
	.w2(32'h3b5fd01a),
	.w3(32'h3c1c5ed3),
	.w4(32'h3c49dba8),
	.w5(32'h3c543524),
	.w6(32'hbbe67f94),
	.w7(32'h3b057d2e),
	.w8(32'hbb1aef14),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02e4f8),
	.w1(32'h3b91249b),
	.w2(32'hbae83572),
	.w3(32'hbb6dc067),
	.w4(32'hbc25cb87),
	.w5(32'h3c103fb2),
	.w6(32'h3c0a9016),
	.w7(32'hbbec0359),
	.w8(32'hbb3718b1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3587af),
	.w1(32'hbbaae85e),
	.w2(32'h3bc12625),
	.w3(32'hbba5a9cc),
	.w4(32'hbc3f36ca),
	.w5(32'h3b3f844c),
	.w6(32'h3b624321),
	.w7(32'hbac16427),
	.w8(32'h38aac1f5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a782030),
	.w1(32'hbc8d24e9),
	.w2(32'hbc9a73b9),
	.w3(32'hbc1f09cc),
	.w4(32'hbca5c606),
	.w5(32'h3cf63647),
	.w6(32'hbc0f2262),
	.w7(32'hbca59e66),
	.w8(32'hbb920c28),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12e347),
	.w1(32'h3b051747),
	.w2(32'hbbe1aec2),
	.w3(32'h3c3781a8),
	.w4(32'h3c8460c7),
	.w5(32'hbc97589c),
	.w6(32'h3be185f7),
	.w7(32'h3c509fc5),
	.w8(32'hbacfe28a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0470f1),
	.w1(32'h399b7fcc),
	.w2(32'h3bd89f4a),
	.w3(32'h3bd716a9),
	.w4(32'h3b46fe15),
	.w5(32'hbafab4ed),
	.w6(32'h3beff7d2),
	.w7(32'h3bf93099),
	.w8(32'h3c37ec99),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fcf3a),
	.w1(32'h3b50b8d5),
	.w2(32'hbb66a069),
	.w3(32'h3c08d76e),
	.w4(32'h3b660dbe),
	.w5(32'hbbd563d7),
	.w6(32'h3b523d6f),
	.w7(32'h39138e2d),
	.w8(32'hbb4c6dda),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fd78d),
	.w1(32'h3afcde6a),
	.w2(32'h3af8ece2),
	.w3(32'hbb429dcd),
	.w4(32'hbbd3cf3c),
	.w5(32'h3b3aaaf3),
	.w6(32'h3b8fce36),
	.w7(32'hbbc40d1b),
	.w8(32'h3b60666a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37df68),
	.w1(32'h3c381398),
	.w2(32'h3c260e0a),
	.w3(32'h3b6073b9),
	.w4(32'h3bde8f7f),
	.w5(32'h3c306508),
	.w6(32'h3b9a5b1c),
	.w7(32'h3be19d80),
	.w8(32'h3c20989c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e45315),
	.w1(32'h3ba77ab9),
	.w2(32'h388c3ced),
	.w3(32'hbaf060c7),
	.w4(32'h3c061ade),
	.w5(32'hbc256602),
	.w6(32'hbb00c54b),
	.w7(32'h3b78ec4e),
	.w8(32'h38a2287b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889bead),
	.w1(32'h3ad67bc5),
	.w2(32'hb82803e8),
	.w3(32'h3bae2a24),
	.w4(32'hbbfb2c31),
	.w5(32'h3c6876de),
	.w6(32'hbc0ddfb4),
	.w7(32'hba72e4e5),
	.w8(32'h381823ff),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3788dd),
	.w1(32'hba08f32f),
	.w2(32'h3ae501fc),
	.w3(32'hbb9b6685),
	.w4(32'hbc188c7e),
	.w5(32'h3b0a07b1),
	.w6(32'hbb5848a0),
	.w7(32'hbb2723c8),
	.w8(32'h3bc44eed),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b950a7c),
	.w1(32'h3b02e417),
	.w2(32'hbac92d70),
	.w3(32'hba5c84af),
	.w4(32'h3b81f19c),
	.w5(32'hbb897958),
	.w6(32'h3bc0fb0b),
	.w7(32'hba0cf9f6),
	.w8(32'hbba4039e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9865c6),
	.w1(32'h3bcf1705),
	.w2(32'h3b7e524d),
	.w3(32'hbb207fa9),
	.w4(32'hbb990da7),
	.w5(32'hbc436094),
	.w6(32'h3afb858f),
	.w7(32'hbac47538),
	.w8(32'hbb03fb22),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea0fc8),
	.w1(32'h3c1764b6),
	.w2(32'h3a859351),
	.w3(32'h3b8edb20),
	.w4(32'h3bae7b86),
	.w5(32'h3c2ae817),
	.w6(32'h3bc87c82),
	.w7(32'hbb0663b8),
	.w8(32'h3c2c4615),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1d747),
	.w1(32'hbc1a59b0),
	.w2(32'hbc40ff16),
	.w3(32'hbaa4917b),
	.w4(32'hbbb34e12),
	.w5(32'hbb17f1dc),
	.w6(32'h3c64a147),
	.w7(32'hbb977e37),
	.w8(32'hbc911bc3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be72bee),
	.w1(32'hbc976829),
	.w2(32'hbb86a3a4),
	.w3(32'hbc15374a),
	.w4(32'hbc25a1bd),
	.w5(32'h3d23c1a0),
	.w6(32'hbb91907d),
	.w7(32'hbc501b31),
	.w8(32'hbc16afbf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfd0f6),
	.w1(32'h3bc7d15b),
	.w2(32'h3a9f7a16),
	.w3(32'h3bf2a699),
	.w4(32'h3c4d2940),
	.w5(32'hbca4e085),
	.w6(32'hbba2bd5e),
	.w7(32'h3b7ce3a2),
	.w8(32'h3ba5a11a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181055),
	.w1(32'h3baa0b96),
	.w2(32'h3c1e0eb1),
	.w3(32'h3b4b67d8),
	.w4(32'h3c0eff83),
	.w5(32'h3c1bd2ff),
	.w6(32'h3c115188),
	.w7(32'h3b1aea36),
	.w8(32'h3c033e7e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33d1d3),
	.w1(32'hbc96a02b),
	.w2(32'hbc8c0d50),
	.w3(32'hbbc66566),
	.w4(32'hbc5dbbc8),
	.w5(32'hbc94d577),
	.w6(32'h3b97eb8d),
	.w7(32'hbc80cbd6),
	.w8(32'hbc85714c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404578),
	.w1(32'hbb081e60),
	.w2(32'h3bb58418),
	.w3(32'hb9bd2451),
	.w4(32'h3c3b408f),
	.w5(32'hbbece50d),
	.w6(32'hbbd1303d),
	.w7(32'h3b36e840),
	.w8(32'hbad0a630),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e75f8),
	.w1(32'hba51143d),
	.w2(32'h3bd2fc64),
	.w3(32'h396edf8e),
	.w4(32'h3bc6a1e2),
	.w5(32'hbb9ee5c5),
	.w6(32'h3b5fd053),
	.w7(32'h3a3f710b),
	.w8(32'h3b8941b6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d0574),
	.w1(32'h3bc5e0c2),
	.w2(32'h3be90204),
	.w3(32'hbc462a45),
	.w4(32'h3bcf2fdf),
	.w5(32'hbc5c4bf2),
	.w6(32'h3b732cee),
	.w7(32'h3c129311),
	.w8(32'h3c29f12d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d898),
	.w1(32'hbc924a82),
	.w2(32'hbcbdfc95),
	.w3(32'h3c91c00f),
	.w4(32'hbc43b71e),
	.w5(32'hba8dfeb7),
	.w6(32'h3a6827d0),
	.w7(32'hbcb836bc),
	.w8(32'hbc689d72),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc667819),
	.w1(32'h3c127ac8),
	.w2(32'hbb850ad7),
	.w3(32'hbb1b33a5),
	.w4(32'h3ba58843),
	.w5(32'hbc6c00ac),
	.w6(32'h3ad27be6),
	.w7(32'h3b3aadba),
	.w8(32'h3bdb4101),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b631d02),
	.w1(32'h3c573e5c),
	.w2(32'h3a8eea5c),
	.w3(32'h3af900c7),
	.w4(32'h3c80fb2e),
	.w5(32'hb94e70c6),
	.w6(32'h3b88db4c),
	.w7(32'h3c3b539c),
	.w8(32'h3b1b45dc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4adac2),
	.w1(32'hba5d3a69),
	.w2(32'hbc161b66),
	.w3(32'hbc7093d8),
	.w4(32'hba80144f),
	.w5(32'hbcc21fd0),
	.w6(32'hbaa24f06),
	.w7(32'hb8a906a7),
	.w8(32'hbc36976f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51f02a),
	.w1(32'hbc5f46fd),
	.w2(32'h3bbebd16),
	.w3(32'h3c18bf9a),
	.w4(32'hbc63d4b4),
	.w5(32'h3c19837b),
	.w6(32'hbc075f9a),
	.w7(32'h3b4d2959),
	.w8(32'h3b83b17f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31fd62),
	.w1(32'hbc84cc2c),
	.w2(32'hbba0e9bf),
	.w3(32'h3c760c58),
	.w4(32'hbce05045),
	.w5(32'h3bc9607e),
	.w6(32'h3b94bf5e),
	.w7(32'hbbb5a7b3),
	.w8(32'hb961e61e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27126a),
	.w1(32'h3a620833),
	.w2(32'hbb9583ea),
	.w3(32'h3bb1cd23),
	.w4(32'hbc09e7ea),
	.w5(32'h3c8294bc),
	.w6(32'h3bd6d6ac),
	.w7(32'h3b8ef973),
	.w8(32'h3b661a54),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b850b35),
	.w1(32'hbb40faa2),
	.w2(32'hba8a3b9c),
	.w3(32'hbbf44067),
	.w4(32'hbb200049),
	.w5(32'h3acd0a5d),
	.w6(32'hbb7d79cb),
	.w7(32'hbb2f6844),
	.w8(32'h3a8ec8a0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c7f594),
	.w1(32'hb72d95d3),
	.w2(32'hb7a3f139),
	.w3(32'hb7a90339),
	.w4(32'h37cfd080),
	.w5(32'h3735f24d),
	.w6(32'hb544e96b),
	.w7(32'h37783ec7),
	.w8(32'hb7670b26),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e9dd7c),
	.w1(32'h37eced99),
	.w2(32'hb836ad7e),
	.w3(32'hb7bde445),
	.w4(32'h378a1910),
	.w5(32'hb8219a35),
	.w6(32'hb83fc84c),
	.w7(32'hb7830ec4),
	.w8(32'hb85fdf3a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85fe0e4),
	.w1(32'h379af968),
	.w2(32'h37133956),
	.w3(32'hb7f04e62),
	.w4(32'h37fda7ab),
	.w5(32'h37f0cfa7),
	.w6(32'hb823db7a),
	.w7(32'h35dc1a45),
	.w8(32'hb80c7d6c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288244),
	.w1(32'h3a90f5ce),
	.w2(32'h3a89f030),
	.w3(32'h3a354e3d),
	.w4(32'h3a8b0d66),
	.w5(32'h3a3e088d),
	.w6(32'h3a619b3d),
	.w7(32'h3a6a9266),
	.w8(32'h3a4c1127),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62a3f70),
	.w1(32'h3824d73f),
	.w2(32'hb785956e),
	.w3(32'hb84666a8),
	.w4(32'hb7ac1190),
	.w5(32'hb8355cb7),
	.w6(32'hb82031bd),
	.w7(32'hb857e04e),
	.w8(32'hb8867666),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae232c1),
	.w1(32'h3bc75af7),
	.w2(32'h3b40db45),
	.w3(32'h3b629800),
	.w4(32'h3bbf8b4b),
	.w5(32'h3a91020c),
	.w6(32'h3b992aae),
	.w7(32'h3b0623e0),
	.w8(32'h39e7e48e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b413eac),
	.w1(32'h3bfa90c2),
	.w2(32'h3bc22aca),
	.w3(32'h3b4fe3b0),
	.w4(32'h3c127553),
	.w5(32'h3b62c553),
	.w6(32'h3bf02853),
	.w7(32'h3bbadc0f),
	.w8(32'h3b4de4c8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95450fa),
	.w1(32'hbb3b1088),
	.w2(32'h3961a48a),
	.w3(32'hbaeab30c),
	.w4(32'hbb161456),
	.w5(32'h3ad66a64),
	.w6(32'hbb14b14a),
	.w7(32'hbaebf13a),
	.w8(32'h3ad36e40),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb11b3),
	.w1(32'h3a824a31),
	.w2(32'h3980d6a7),
	.w3(32'h3b03ece6),
	.w4(32'h3a8ad76b),
	.w5(32'hb831d279),
	.w6(32'h3b0d692d),
	.w7(32'h3a63419c),
	.w8(32'h39712399),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f58a8c),
	.w1(32'h389c41f5),
	.w2(32'h39000cfd),
	.w3(32'h393e4758),
	.w4(32'hb95af4ae),
	.w5(32'hb9e08b8f),
	.w6(32'h3ab5277f),
	.w7(32'h3a483395),
	.w8(32'h3a6654f1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a228fb2),
	.w1(32'hba0c5b05),
	.w2(32'h388f1e3d),
	.w3(32'h39697a81),
	.w4(32'hba12ddc2),
	.w5(32'h39d2cbfb),
	.w6(32'h38ac32c8),
	.w7(32'hb9d91fe7),
	.w8(32'h39aea39b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2534b1),
	.w1(32'h3b89e7e4),
	.w2(32'h3b36ae87),
	.w3(32'h3b6af31a),
	.w4(32'h3b72ce35),
	.w5(32'h3aca1681),
	.w6(32'h3b58cc68),
	.w7(32'h3b2d5523),
	.w8(32'h3a8452d6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc10f1),
	.w1(32'h37e45d9b),
	.w2(32'h36ccbe6a),
	.w3(32'h3801633f),
	.w4(32'h38043cb5),
	.w5(32'h37b94520),
	.w6(32'h36a3579e),
	.w7(32'h374f4014),
	.w8(32'h368792e5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0588d),
	.w1(32'hb7233b51),
	.w2(32'h3492e14a),
	.w3(32'hb73551ad),
	.w4(32'h36db71a6),
	.w5(32'h3819fea5),
	.w6(32'hb65e3832),
	.w7(32'hb419fae0),
	.w8(32'hb6af54be),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb762244f),
	.w1(32'hb9967432),
	.w2(32'hb95f31e5),
	.w3(32'hb951ac0c),
	.w4(32'hb9b8a0bf),
	.w5(32'hb7b20018),
	.w6(32'hb9906b99),
	.w7(32'hb97eb57d),
	.w8(32'hb87f0c76),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fe0647),
	.w1(32'hb8646c91),
	.w2(32'hb7606765),
	.w3(32'hb716b9e8),
	.w4(32'hb825b6e5),
	.w5(32'hb7f8f3de),
	.w6(32'h36794897),
	.w7(32'hb868be4a),
	.w8(32'hb8830671),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06a06b),
	.w1(32'hbb16d708),
	.w2(32'hba99c6ab),
	.w3(32'hbb06323d),
	.w4(32'hbb2fe928),
	.w5(32'hb9840389),
	.w6(32'hbadd7db4),
	.w7(32'hbaf48cdc),
	.w8(32'hb8e17af6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8b24f),
	.w1(32'h3812a194),
	.w2(32'h38bbe06f),
	.w3(32'hb97b80a4),
	.w4(32'hb8215208),
	.w5(32'h38a32329),
	.w6(32'hb907c81d),
	.w7(32'hb94ec7ef),
	.w8(32'hb930ceb3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbe20f),
	.w1(32'hb9d414aa),
	.w2(32'hb9449f8f),
	.w3(32'h393c47c7),
	.w4(32'hb8ea6706),
	.w5(32'h3932d95e),
	.w6(32'h3a978457),
	.w7(32'h3966e048),
	.w8(32'h37c941ff),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe03e4),
	.w1(32'h3c145e07),
	.w2(32'h3a7ebe0d),
	.w3(32'h3c2ae81f),
	.w4(32'h3c182917),
	.w5(32'hb9df2a5f),
	.w6(32'h3c36871f),
	.w7(32'h3bc604dd),
	.w8(32'h3a88f761),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c3a9d),
	.w1(32'hba8493bc),
	.w2(32'h3a0690bb),
	.w3(32'hbae39d44),
	.w4(32'hba3e912b),
	.w5(32'hb9043ee8),
	.w6(32'hbabd9a41),
	.w7(32'hba69edc0),
	.w8(32'hb936434d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9324974),
	.w1(32'h3b486c4a),
	.w2(32'h3b0315c8),
	.w3(32'h3b14ae51),
	.w4(32'h3b39cf78),
	.w5(32'h3b347943),
	.w6(32'h3ac43866),
	.w7(32'h3b0d9d01),
	.w8(32'h3b078270),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d42779),
	.w1(32'hbb33241b),
	.w2(32'hbb009ff0),
	.w3(32'hba552f85),
	.w4(32'hbb233fb0),
	.w5(32'hba8a0f8a),
	.w6(32'hba6b6b0b),
	.w7(32'hbb195981),
	.w8(32'hba87b611),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbe8e5),
	.w1(32'h39f65fd6),
	.w2(32'h3a60fab3),
	.w3(32'h3b309b86),
	.w4(32'h3a71563b),
	.w5(32'h3986a470),
	.w6(32'h3b3dc403),
	.w7(32'h3a896201),
	.w8(32'h3a06de05),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c7bcf),
	.w1(32'hba8a3bf9),
	.w2(32'hba02c59e),
	.w3(32'h3909abab),
	.w4(32'hbadf8d9d),
	.w5(32'hba1c222b),
	.w6(32'hb9ad017c),
	.w7(32'hba99892b),
	.w8(32'hba0066ef),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a832),
	.w1(32'hbb219709),
	.w2(32'hb8e4d3b2),
	.w3(32'hbae79f52),
	.w4(32'hbb0d0460),
	.w5(32'h3930ba16),
	.w6(32'hbaff0604),
	.w7(32'hbb0c6a7e),
	.w8(32'hba07424a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35169805),
	.w1(32'h39262fc5),
	.w2(32'h37b10e76),
	.w3(32'hb9a97484),
	.w4(32'h390706a0),
	.w5(32'h390a6cb4),
	.w6(32'hba0f3df1),
	.w7(32'h36bfd120),
	.w8(32'hb8bb4068),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeedb65),
	.w1(32'h3a8e8a79),
	.w2(32'h3adbd885),
	.w3(32'h3b0635cc),
	.w4(32'h3aa9527a),
	.w5(32'h3ad7c36c),
	.w6(32'h3af7b361),
	.w7(32'h3ad2be94),
	.w8(32'h3b0ab887),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd6d5),
	.w1(32'hb9863bd4),
	.w2(32'hb9e20458),
	.w3(32'hb9984093),
	.w4(32'hbb1eba19),
	.w5(32'hba2f8fb4),
	.w6(32'hb94784cc),
	.w7(32'hbac451ac),
	.w8(32'h39055b8c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5da6fc),
	.w1(32'h3c2810e2),
	.w2(32'h3b8e0694),
	.w3(32'h3bdebe36),
	.w4(32'h3c1f8252),
	.w5(32'h3b1f6b06),
	.w6(32'h3c09e386),
	.w7(32'h3bb51614),
	.w8(32'h3b1de404),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be8828),
	.w1(32'hbb3ca7ce),
	.w2(32'hba60c152),
	.w3(32'hbad449f3),
	.w4(32'hbb4c7275),
	.w5(32'h3a20d3bc),
	.w6(32'hbb6a1554),
	.w7(32'hbb161d4f),
	.w8(32'hb9b02baa),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940c5a6),
	.w1(32'hbb3956fe),
	.w2(32'hba8a2c57),
	.w3(32'hbadd7d48),
	.w4(32'hbaabdb62),
	.w5(32'h3a28009c),
	.w6(32'hba9874ba),
	.w7(32'hba8f75a4),
	.w8(32'h3aad3a37),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1bcde),
	.w1(32'h3b5fa161),
	.w2(32'h3adca585),
	.w3(32'h3b374347),
	.w4(32'h3b1765fc),
	.w5(32'h39f6ce0d),
	.w6(32'h3b5c0258),
	.w7(32'h3b263cc6),
	.w8(32'h3ad3ec9a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e76c1),
	.w1(32'hb93938d2),
	.w2(32'hba591d34),
	.w3(32'h39cca386),
	.w4(32'hb8019346),
	.w5(32'hba6002ec),
	.w6(32'h38b70c07),
	.w7(32'h3934bf33),
	.w8(32'hba56a7a2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9447d7),
	.w1(32'h3c681d4c),
	.w2(32'h3c174d77),
	.w3(32'h3bb4d444),
	.w4(32'h3c3d93fd),
	.w5(32'h3ba1f721),
	.w6(32'h3c12ebe8),
	.w7(32'h3bec385e),
	.w8(32'h3b6e9a31),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1e477),
	.w1(32'hba88041e),
	.w2(32'h3a895d56),
	.w3(32'hbada1f50),
	.w4(32'hba4680d5),
	.w5(32'h3b08aabf),
	.w6(32'hba85d21e),
	.w7(32'hba94fff1),
	.w8(32'h3a659fb5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846c924),
	.w1(32'hb864fe26),
	.w2(32'hb91a60fd),
	.w3(32'h35cbecf3),
	.w4(32'hb92474e6),
	.w5(32'hb8b94890),
	.w6(32'hb8a7e61c),
	.w7(32'hb8c33aa7),
	.w8(32'hb8494e53),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14429c),
	.w1(32'hb7978ea4),
	.w2(32'hb99c2c5d),
	.w3(32'h3a80c52f),
	.w4(32'h38f1a90c),
	.w5(32'hb8a0627c),
	.w6(32'h39ad5ea1),
	.w7(32'h3964c5dc),
	.w8(32'h3900e2c8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2e205),
	.w1(32'hbafaef34),
	.w2(32'hb88398cf),
	.w3(32'hb9bfdbe5),
	.w4(32'hba6ed985),
	.w5(32'h3a383f7e),
	.w6(32'h398c01e2),
	.w7(32'hb9cb5e0c),
	.w8(32'h3aaa0197),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c784f),
	.w1(32'hbb30baf3),
	.w2(32'h37a8ed8c),
	.w3(32'hbae3c37d),
	.w4(32'hbb058efb),
	.w5(32'h3a4d367a),
	.w6(32'hbafe6622),
	.w7(32'hbac88b1e),
	.w8(32'h3a86626e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce9005),
	.w1(32'hba0b99d2),
	.w2(32'h39ab6666),
	.w3(32'hb97f89de),
	.w4(32'hbb14510f),
	.w5(32'h3a005bc3),
	.w6(32'hb9de4ded),
	.w7(32'hbacf753b),
	.w8(32'hb9819c7b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16469c),
	.w1(32'hba3bb04c),
	.w2(32'h3673197a),
	.w3(32'h3a2fb779),
	.w4(32'hba0cefc4),
	.w5(32'h39a5463c),
	.w6(32'h39990580),
	.w7(32'hb9793fb7),
	.w8(32'h39e5c1a5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80f80e),
	.w1(32'h3a8e1fa6),
	.w2(32'h3a879dc0),
	.w3(32'h398d8115),
	.w4(32'h38df92e5),
	.w5(32'h39e35423),
	.w6(32'h3967b23f),
	.w7(32'hb7e7fd73),
	.w8(32'h3a05326a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8f61),
	.w1(32'h3a400931),
	.w2(32'h39ce27cb),
	.w3(32'h3ac9842e),
	.w4(32'h3a193253),
	.w5(32'h3a03d49b),
	.w6(32'h3b0a8506),
	.w7(32'h3a53c539),
	.w8(32'h399b0b88),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f555b8),
	.w1(32'hbacb0589),
	.w2(32'hb91f3e89),
	.w3(32'hba4f825c),
	.w4(32'hbac64ef9),
	.w5(32'h39c0c82c),
	.w6(32'hba1f9aea),
	.w7(32'hba93b6ae),
	.w8(32'h3a364542),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918c8f9),
	.w1(32'h382ebc27),
	.w2(32'hb6d4e8de),
	.w3(32'h394c5341),
	.w4(32'h38fb61aa),
	.w5(32'h38dfcb60),
	.w6(32'h39360dfa),
	.w7(32'h38815efd),
	.w8(32'h3849fe07),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a90198),
	.w1(32'h37b7e7d4),
	.w2(32'h38252b04),
	.w3(32'h36f0625b),
	.w4(32'h34909d9a),
	.w5(32'hb664d8f9),
	.w6(32'h36891098),
	.w7(32'hb56d011a),
	.w8(32'h37fe96b1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86653f2),
	.w1(32'hb76f69fc),
	.w2(32'hb6f9c758),
	.w3(32'hb757e5ca),
	.w4(32'hb5a8c980),
	.w5(32'hb73268c3),
	.w6(32'hb81871de),
	.w7(32'hb727f41c),
	.w8(32'hb7ae1c34),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393dfd77),
	.w1(32'hb8359300),
	.w2(32'h390bee5e),
	.w3(32'h38bba36e),
	.w4(32'hb8930328),
	.w5(32'h37586231),
	.w6(32'h38061a7b),
	.w7(32'h3742aa5f),
	.w8(32'hb7051c47),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4a77f),
	.w1(32'hbb056b5a),
	.w2(32'hba6cd631),
	.w3(32'hba63bd29),
	.w4(32'hbad5b10e),
	.w5(32'hb824e3eb),
	.w6(32'hbaab0306),
	.w7(32'hbaeb30e1),
	.w8(32'hb9941ead),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941bd1c),
	.w1(32'h39b10367),
	.w2(32'h39bcb0d5),
	.w3(32'h3a081e3c),
	.w4(32'h39b9a07c),
	.w5(32'h39987795),
	.w6(32'h398f633a),
	.w7(32'h39275683),
	.w8(32'h39ba7236),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a967a4a),
	.w1(32'h3b0db72b),
	.w2(32'h3adb3a93),
	.w3(32'h3a8e5961),
	.w4(32'h3afb9b53),
	.w5(32'h3a3dd63f),
	.w6(32'h3b0ac43b),
	.w7(32'h3abd2d7f),
	.w8(32'h3a9b07f6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446376),
	.w1(32'hbb6750a2),
	.w2(32'hba663060),
	.w3(32'hbb1b450f),
	.w4(32'hbb2ee742),
	.w5(32'h3a8fc175),
	.w6(32'hbb60cd62),
	.w7(32'hbb027d18),
	.w8(32'h3a635f8c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923a044),
	.w1(32'hb8ff5aea),
	.w2(32'hb82253b6),
	.w3(32'hb8f4dcaa),
	.w4(32'h375341ac),
	.w5(32'h391385fe),
	.w6(32'hb879ffc5),
	.w7(32'h3841e682),
	.w8(32'h38ebb979),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fdb4ae),
	.w1(32'h38b4a52c),
	.w2(32'h38b3979a),
	.w3(32'h38aa72e5),
	.w4(32'h38ee7fff),
	.w5(32'h38c6e720),
	.w6(32'h38802a07),
	.w7(32'h379e3aec),
	.w8(32'h38d7a532),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82ec7df),
	.w1(32'hb6cc8cfe),
	.w2(32'hb7b2b3b5),
	.w3(32'hb81c2735),
	.w4(32'hb7474bde),
	.w5(32'hb78bfaec),
	.w6(32'hb7c1b1db),
	.w7(32'hb7434224),
	.w8(32'hb7db1bc4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93eb817),
	.w1(32'hba042155),
	.w2(32'hb99865c4),
	.w3(32'hba5fef82),
	.w4(32'hba3cc1b9),
	.w5(32'h38336dd0),
	.w6(32'hba643967),
	.w7(32'hba0ca5fe),
	.w8(32'h3889967c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0787bc),
	.w1(32'h3a1c1e5a),
	.w2(32'h39fb041f),
	.w3(32'h392f43b8),
	.w4(32'h39e267dd),
	.w5(32'h3a994d18),
	.w6(32'h3aba5fe3),
	.w7(32'h3a9c2629),
	.w8(32'h3a911aae),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a00e75),
	.w1(32'hb90cfe81),
	.w2(32'h39c575a8),
	.w3(32'h3a834d7c),
	.w4(32'h3abf3540),
	.w5(32'h3a299f18),
	.w6(32'h3a8e3d6f),
	.w7(32'h3a49d654),
	.w8(32'h399b05cc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984c524),
	.w1(32'h3accb201),
	.w2(32'h3a91bf33),
	.w3(32'h3a330c22),
	.w4(32'h3a993e19),
	.w5(32'h3a07cf50),
	.w6(32'h3a4840cc),
	.w7(32'h3a1baf37),
	.w8(32'h3a084042),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adba121),
	.w1(32'h3a86edd1),
	.w2(32'h392d0158),
	.w3(32'h3a6bf60e),
	.w4(32'h3a13c01f),
	.w5(32'hb970b95b),
	.w6(32'h3a8251a2),
	.w7(32'h389a87ed),
	.w8(32'h3a64f4d5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b37aad),
	.w1(32'hba33ee8c),
	.w2(32'hb8f00e43),
	.w3(32'hba1318fa),
	.w4(32'hba0970f5),
	.w5(32'h36c44222),
	.w6(32'hba2e973b),
	.w7(32'hba0f0f74),
	.w8(32'h382757f6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec1480),
	.w1(32'h363a1e1e),
	.w2(32'hb91eb848),
	.w3(32'h3a4e087a),
	.w4(32'h39c597b2),
	.w5(32'h3805733a),
	.w6(32'h3a5dcb41),
	.w7(32'h39cbb159),
	.w8(32'h39779163),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe07e8),
	.w1(32'hbace9b9e),
	.w2(32'hbb4f5b63),
	.w3(32'h3ad477eb),
	.w4(32'hba514d8c),
	.w5(32'hbb1ddba6),
	.w6(32'h3a0b1582),
	.w7(32'hbab66b11),
	.w8(32'hbb21f08d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52cceb),
	.w1(32'h3b9f9baf),
	.w2(32'h3b4d2d1b),
	.w3(32'h3baf0e0d),
	.w4(32'h3ba876d2),
	.w5(32'h3aefbe6b),
	.w6(32'h3ba2942b),
	.w7(32'h3b5fa0fd),
	.w8(32'h3b1ea990),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba699320),
	.w1(32'hbacb7df7),
	.w2(32'h378d8dbf),
	.w3(32'hbaca5253),
	.w4(32'hba8c47c3),
	.w5(32'h3a3621ff),
	.w6(32'hbaa5469c),
	.w7(32'hbaa65690),
	.w8(32'h38594e82),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37be93),
	.w1(32'h39533285),
	.w2(32'h39c14ebf),
	.w3(32'h395891d9),
	.w4(32'hb991e87b),
	.w5(32'h3a1387c4),
	.w6(32'hb8d021b2),
	.w7(32'h39a5966e),
	.w8(32'h3a3afdec),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75cca4),
	.w1(32'h3b9219a1),
	.w2(32'h3ad22a86),
	.w3(32'h3b954665),
	.w4(32'h3b87f713),
	.w5(32'h3a0ebb68),
	.w6(32'h3b885359),
	.w7(32'h3b063213),
	.w8(32'h3a79da53),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39531840),
	.w1(32'hb9f5ef90),
	.w2(32'hba8ae4d7),
	.w3(32'h3980588b),
	.w4(32'hb891a54a),
	.w5(32'hb97bdc9c),
	.w6(32'h3a7d19b4),
	.w7(32'hb887c225),
	.w8(32'hb7e772a8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11bd83),
	.w1(32'hb867b267),
	.w2(32'h3900f80d),
	.w3(32'h3a19198e),
	.w4(32'hb80e162d),
	.w5(32'h39772472),
	.w6(32'h3a449fde),
	.w7(32'h381cf74b),
	.w8(32'h391b7a95),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5edd6),
	.w1(32'hb8dd4939),
	.w2(32'hb8002daa),
	.w3(32'h39c2b1bf),
	.w4(32'h392a2994),
	.w5(32'h395e6e2a),
	.w6(32'h39d13cbf),
	.w7(32'h389cbc7a),
	.w8(32'h396e386a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933875),
	.w1(32'hbb8ee82c),
	.w2(32'hba3c88f9),
	.w3(32'hbb58f2dd),
	.w4(32'hbb82fdc0),
	.w5(32'h3aa893f3),
	.w6(32'hbb82fac9),
	.w7(32'hbb39e374),
	.w8(32'h3a2cdb4d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ecde9),
	.w1(32'h3a848dcc),
	.w2(32'h3a468c65),
	.w3(32'h3ab4edbe),
	.w4(32'h39b3e3e3),
	.w5(32'hb981b2e1),
	.w6(32'h3aad6c87),
	.w7(32'h38935695),
	.w8(32'hb9dc6155),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f115c7),
	.w1(32'h36ede6ed),
	.w2(32'h3686bbda),
	.w3(32'hb80ecc27),
	.w4(32'h379d10cc),
	.w5(32'h371bb52c),
	.w6(32'hb810bf2d),
	.w7(32'hb6720c1b),
	.w8(32'hb727b71e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d03d12),
	.w1(32'h37b39d2b),
	.w2(32'h3579493b),
	.w3(32'hb80381bb),
	.w4(32'hb6a5d673),
	.w5(32'hb758976c),
	.w6(32'hb7cbda70),
	.w7(32'h359ed21a),
	.w8(32'hb78a4903),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d62a02),
	.w1(32'hb9b71ca5),
	.w2(32'hb90ff006),
	.w3(32'hb921302f),
	.w4(32'hb95fd5a0),
	.w5(32'h3a4c9a24),
	.w6(32'hb938c06d),
	.w7(32'hb98a53e6),
	.w8(32'h3a566e97),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6881d),
	.w1(32'hbb27b958),
	.w2(32'h3983b399),
	.w3(32'hbac1bb34),
	.w4(32'hbad6631e),
	.w5(32'h3730432a),
	.w6(32'hba9e8f50),
	.w7(32'hbaa3939c),
	.w8(32'h37cd2fe4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5967fe),
	.w1(32'hba0d0756),
	.w2(32'h390a9ba9),
	.w3(32'h39e06e97),
	.w4(32'h393c2cb4),
	.w5(32'h3abc8dc3),
	.w6(32'h3911f2c7),
	.w7(32'h394862bf),
	.w8(32'h3ade998b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb58c031f),
	.w1(32'hb70d337c),
	.w2(32'h34a71369),
	.w3(32'h377cfc56),
	.w4(32'hb671f978),
	.w5(32'h3758c565),
	.w6(32'hb7c924d8),
	.w7(32'hb7821309),
	.w8(32'h3453e3fd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fefd8),
	.w1(32'hba7264d8),
	.w2(32'h39077ea5),
	.w3(32'h3a1abc2a),
	.w4(32'hb9f4a4d6),
	.w5(32'h39e09154),
	.w6(32'h3a760a91),
	.w7(32'hb916f927),
	.w8(32'h3a3b5999),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba484442),
	.w1(32'hbac879b2),
	.w2(32'hb96d2fb1),
	.w3(32'hbab2a819),
	.w4(32'hbad4efca),
	.w5(32'h3a2eb1e8),
	.w6(32'hb9ad537e),
	.w7(32'hb9c0f21f),
	.w8(32'h3a49749c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3228ec),
	.w1(32'h3b66bd43),
	.w2(32'h3b43ab40),
	.w3(32'h3b3cddc3),
	.w4(32'h3b62a67f),
	.w5(32'h3b0f3d21),
	.w6(32'h3b3edd8f),
	.w7(32'h3b26f862),
	.w8(32'h3b024cbb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa403de),
	.w1(32'hbb03a455),
	.w2(32'h392cb907),
	.w3(32'hb9cf281f),
	.w4(32'hbb2285c2),
	.w5(32'h3a37ab98),
	.w6(32'hba90d88d),
	.w7(32'hbb11952e),
	.w8(32'hb94a5ba5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2254c7),
	.w1(32'hbaa387a2),
	.w2(32'hba2ae698),
	.w3(32'hba54d2a9),
	.w4(32'hbaa33c44),
	.w5(32'hb636a440),
	.w6(32'hbabc8a9e),
	.w7(32'hba6f27ef),
	.w8(32'hb984a849),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9162b),
	.w1(32'h38badfaa),
	.w2(32'hb9a3b991),
	.w3(32'hb9a99e85),
	.w4(32'hb9c9efbd),
	.w5(32'hba1cc07e),
	.w6(32'hba33b875),
	.w7(32'hbaa1f924),
	.w8(32'hba58ee57),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb837048e),
	.w1(32'hbab5d61f),
	.w2(32'h3889905c),
	.w3(32'hba21141b),
	.w4(32'hba8c32b8),
	.w5(32'h39fbe988),
	.w6(32'h3825b700),
	.w7(32'hba56e5c4),
	.w8(32'h39bbbdb7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd7d11),
	.w1(32'hbadbd2b2),
	.w2(32'hba4bf025),
	.w3(32'hb999b661),
	.w4(32'hbb1ea7e1),
	.w5(32'hba5a0e2b),
	.w6(32'hba87cf7b),
	.w7(32'hba9c85a0),
	.w8(32'hba2fe0ef),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d946a6),
	.w1(32'hba63a9b4),
	.w2(32'hb9bae821),
	.w3(32'hba7f17ed),
	.w4(32'hba8d7bfc),
	.w5(32'hba140f47),
	.w6(32'hba86a822),
	.w7(32'hba7d7897),
	.w8(32'hba0d0034),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5415b2),
	.w1(32'h3b02ff31),
	.w2(32'h3a6fa589),
	.w3(32'h3ac1caeb),
	.w4(32'h3ad4151d),
	.w5(32'h39ba7567),
	.w6(32'h3ade6fbe),
	.w7(32'h3a80f10c),
	.w8(32'h3705bdc1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912f632),
	.w1(32'hb9913d65),
	.w2(32'hb91180bb),
	.w3(32'hb9628c36),
	.w4(32'hb9b4f143),
	.w5(32'hb72aa2d1),
	.w6(32'hb980f820),
	.w7(32'hb98d7800),
	.w8(32'hb8b49e49),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a907a93),
	.w1(32'h3a9f091d),
	.w2(32'h3a4d1bfd),
	.w3(32'h3ab186b0),
	.w4(32'h3a6844d2),
	.w5(32'h398a93fc),
	.w6(32'h3a825ac6),
	.w7(32'h3a4dd21f),
	.w8(32'h39534c78),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906d2f5),
	.w1(32'hb920ea70),
	.w2(32'hb86ee798),
	.w3(32'hb9053046),
	.w4(32'hb90d145a),
	.w5(32'hb6969137),
	.w6(32'hb8e6cfc0),
	.w7(32'hb939e4f9),
	.w8(32'hb83f4d64),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b37fe),
	.w1(32'hba2cb5da),
	.w2(32'hba28f520),
	.w3(32'h39a53c1f),
	.w4(32'hba482543),
	.w5(32'h38438c72),
	.w6(32'h39fc31bb),
	.w7(32'hba11e4f4),
	.w8(32'h3899487e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932b0dc),
	.w1(32'hb9ca7b94),
	.w2(32'hb89c6180),
	.w3(32'hb9a9d1c1),
	.w4(32'hb9bb0cd9),
	.w5(32'hb8db724b),
	.w6(32'hb9035b28),
	.w7(32'hb970a76d),
	.w8(32'hb7f977ac),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71f442),
	.w1(32'hb9ba2171),
	.w2(32'hb9e6a344),
	.w3(32'hb9f86ce8),
	.w4(32'h383c7103),
	.w5(32'hb9a144f0),
	.w6(32'hba37b720),
	.w7(32'hb821fb9e),
	.w8(32'h39939c66),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a87caa),
	.w1(32'hb8a64fb8),
	.w2(32'hb8394347),
	.w3(32'h377b7ea0),
	.w4(32'hb8b9d113),
	.w5(32'hb8344807),
	.w6(32'hb78afb70),
	.w7(32'hb89f1876),
	.w8(32'hb8583fb7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933d8f9),
	.w1(32'h38e4a6a1),
	.w2(32'h39633526),
	.w3(32'hb966d6f9),
	.w4(32'h38dee4e5),
	.w5(32'h393d6662),
	.w6(32'hb64905a4),
	.w7(32'h39440088),
	.w8(32'h395e758f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39821e61),
	.w1(32'hbaa4762a),
	.w2(32'h3a17d741),
	.w3(32'hb8da0d0a),
	.w4(32'hbac05f3e),
	.w5(32'h39031e7a),
	.w6(32'hba3f8078),
	.w7(32'hbab989b8),
	.w8(32'hb9f6e9bf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21b55b),
	.w1(32'h3a8526a3),
	.w2(32'h3ad1123f),
	.w3(32'h3ac57432),
	.w4(32'h3a7f8cbe),
	.w5(32'h39450789),
	.w6(32'h3b97095e),
	.w7(32'h3b0a3ff6),
	.w8(32'h3a14f6a2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abffa2),
	.w1(32'hb9ee3023),
	.w2(32'hb9d74f2c),
	.w3(32'hba204439),
	.w4(32'hb9fa9b5f),
	.w5(32'hb91d345f),
	.w6(32'hba182379),
	.w7(32'hb9f02095),
	.w8(32'h359d4cde),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a9045),
	.w1(32'hbb24c00f),
	.w2(32'hba05566b),
	.w3(32'hbac955de),
	.w4(32'hbb005114),
	.w5(32'h39e106b8),
	.w6(32'hbabfe2e2),
	.w7(32'hbaebefb2),
	.w8(32'h39ac7963),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377232ab),
	.w1(32'hb9b95f17),
	.w2(32'hb9a05fc1),
	.w3(32'hb8e0da67),
	.w4(32'hb9d51242),
	.w5(32'hb9a8e829),
	.w6(32'h38d31b32),
	.w7(32'hb9379890),
	.w8(32'hb9b03d90),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10b7a),
	.w1(32'h3a59eda1),
	.w2(32'h3a928840),
	.w3(32'h3abf1493),
	.w4(32'h3a6701aa),
	.w5(32'h3ac03082),
	.w6(32'h3a59016f),
	.w7(32'h3a1c217a),
	.w8(32'h39ae07f3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac07e31),
	.w1(32'h3a636f2c),
	.w2(32'h3a5a4087),
	.w3(32'h3acb5a27),
	.w4(32'h3a547c66),
	.w5(32'h3a1a5263),
	.w6(32'h3ad7f5af),
	.w7(32'h3a2cba14),
	.w8(32'h3a5429c4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830d86),
	.w1(32'h3b22ad3d),
	.w2(32'h39ddb0ea),
	.w3(32'h3b9ee121),
	.w4(32'h3b41d38a),
	.w5(32'h388442dd),
	.w6(32'h3b82f185),
	.w7(32'h3b0c03fa),
	.w8(32'hb9d25e75),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2da59),
	.w1(32'hb9ec9b62),
	.w2(32'hb904523c),
	.w3(32'hb8f1987c),
	.w4(32'hb9e6ad4a),
	.w5(32'hb9155fb5),
	.w6(32'hb91c8acb),
	.w7(32'hb9b0272a),
	.w8(32'hb9d4e50e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39925b93),
	.w1(32'h38480a8e),
	.w2(32'h3a2f3f4a),
	.w3(32'h3a0afe78),
	.w4(32'h38eb1b7a),
	.w5(32'h39714aed),
	.w6(32'h3a3b3ee0),
	.w7(32'h392c4aa3),
	.w8(32'h392be7bb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d5a5d2),
	.w1(32'h37833df7),
	.w2(32'hb8143399),
	.w3(32'hb6ecb963),
	.w4(32'h379061ad),
	.w5(32'hb7d008c8),
	.w6(32'hb808f749),
	.w7(32'hb7bb070f),
	.w8(32'hb7901cd0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b3f5a),
	.w1(32'h39461bdb),
	.w2(32'hb862e7b0),
	.w3(32'h3a51faf5),
	.w4(32'h38f7a761),
	.w5(32'hb9592e5b),
	.w6(32'h3a31f7b5),
	.w7(32'h39735e22),
	.w8(32'hb97c6589),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9df2a),
	.w1(32'h3987f310),
	.w2(32'hb8d1d121),
	.w3(32'h397b4dd6),
	.w4(32'h39403ef9),
	.w5(32'hb8399eff),
	.w6(32'h39c5d2f2),
	.w7(32'h396f4021),
	.w8(32'hb8e327db),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e3ca),
	.w1(32'h382cfb0e),
	.w2(32'h3a8ed80b),
	.w3(32'h390517c1),
	.w4(32'hb980d599),
	.w5(32'h3a82778d),
	.w6(32'h3a074166),
	.w7(32'h39ee584e),
	.w8(32'h3aae8b80),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb602b7f3),
	.w1(32'h3815ec91),
	.w2(32'hb67e21ee),
	.w3(32'hb74975f1),
	.w4(32'h36263a35),
	.w5(32'hb77b5a19),
	.w6(32'h3809671e),
	.w7(32'h352aed92),
	.w8(32'hb6cf1213),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a064c),
	.w1(32'h391e998f),
	.w2(32'h391fbf6d),
	.w3(32'h392e3ad0),
	.w4(32'h387cfdd4),
	.w5(32'h3815052d),
	.w6(32'h39302dbf),
	.w7(32'h38088d74),
	.w8(32'h38210a96),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ef6dd),
	.w1(32'h3987fde2),
	.w2(32'h382dbb6b),
	.w3(32'hba089d16),
	.w4(32'hb9a0840a),
	.w5(32'h39c7bdab),
	.w6(32'h39e36e0a),
	.w7(32'hb88f7368),
	.w8(32'h3a2ab28d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba357185),
	.w1(32'h3a8154cf),
	.w2(32'h39e23d78),
	.w3(32'hbab3887c),
	.w4(32'hb9a5c63e),
	.w5(32'h3a8eda58),
	.w6(32'hb9296088),
	.w7(32'h3992a489),
	.w8(32'h3aad13c6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2465ed),
	.w1(32'h3a1b5768),
	.w2(32'hb89e7e12),
	.w3(32'h3a2f3182),
	.w4(32'h398c3e20),
	.w5(32'hb9e6520c),
	.w6(32'h3a20c2eb),
	.w7(32'h39a1c945),
	.w8(32'h3907f2d3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f1c8),
	.w1(32'h3a97e89b),
	.w2(32'h38f74fac),
	.w3(32'h3b09ca42),
	.w4(32'h3898e5b6),
	.w5(32'h39e37939),
	.w6(32'h3aabcc9c),
	.w7(32'h39e5faa3),
	.w8(32'hb90ea7d3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2e0a),
	.w1(32'h3ba2c429),
	.w2(32'h3b95138f),
	.w3(32'h3b9ffc63),
	.w4(32'h3bb5996f),
	.w5(32'h3ba17e73),
	.w6(32'h3b8d038e),
	.w7(32'h3b70b67d),
	.w8(32'h3b1d3919),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a975d0e),
	.w1(32'hbb996eb7),
	.w2(32'hbacc46dc),
	.w3(32'hb93d31bc),
	.w4(32'hbba5a6c7),
	.w5(32'hba2f1970),
	.w6(32'hbaa58efd),
	.w7(32'hbb85984c),
	.w8(32'hb9f91752),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967d44f),
	.w1(32'h38cbfc02),
	.w2(32'h3985eb5e),
	.w3(32'hb988bde0),
	.w4(32'h393e5edd),
	.w5(32'h38f64525),
	.w6(32'h36d4bd5a),
	.w7(32'h38ff0620),
	.w8(32'h394600bd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38065359),
	.w1(32'h388a12bc),
	.w2(32'hb7bea2b4),
	.w3(32'h36695a28),
	.w4(32'h37f137b3),
	.w5(32'hb7cdd7b4),
	.w6(32'hb6d03f6f),
	.w7(32'h37802377),
	.w8(32'hb78d0fbb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6b176),
	.w1(32'h398e0131),
	.w2(32'h398f4c1f),
	.w3(32'h38a4bdd4),
	.w4(32'h39242e47),
	.w5(32'h39726e0d),
	.w6(32'h38d27efb),
	.w7(32'h393e42b4),
	.w8(32'h3985fe20),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb728bf84),
	.w1(32'h37553901),
	.w2(32'hb6b2d03d),
	.w3(32'hb8055bb7),
	.w4(32'hb6490740),
	.w5(32'hb6fa46a8),
	.w6(32'hb849870c),
	.w7(32'h36a678cf),
	.w8(32'hb6f92f93),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3654c),
	.w1(32'hb9dfd2e5),
	.w2(32'hb9385803),
	.w3(32'hba08d502),
	.w4(32'hb9d8fb96),
	.w5(32'hb886815b),
	.w6(32'hb9868283),
	.w7(32'hb9653af0),
	.w8(32'h38dfeacd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9ba00),
	.w1(32'h39447543),
	.w2(32'h3a26dac4),
	.w3(32'hb89344bb),
	.w4(32'hba280ff1),
	.w5(32'h38cf6ffa),
	.w6(32'h39e93110),
	.w7(32'h39ae1cc0),
	.w8(32'hb72ec04f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b2f99),
	.w1(32'hbaea8cae),
	.w2(32'h3871f429),
	.w3(32'hba6de942),
	.w4(32'hba3af726),
	.w5(32'h3a490c7c),
	.w6(32'hba6e580f),
	.w7(32'hba6826b6),
	.w8(32'h39fa6899),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c69ef3),
	.w1(32'hb945171b),
	.w2(32'hb952d4c3),
	.w3(32'hb8d0c4c2),
	.w4(32'hb9e94862),
	.w5(32'hb8b784c8),
	.w6(32'h39e56b31),
	.w7(32'hb7a558e5),
	.w8(32'h390b655e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b114fc),
	.w1(32'hbc0ebf11),
	.w2(32'hb990e1e8),
	.w3(32'hb7a60720),
	.w4(32'hbc3604c2),
	.w5(32'hbac29db7),
	.w6(32'h397d3f60),
	.w7(32'hbbc23a9d),
	.w8(32'hbb7924ec),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a0d9d),
	.w1(32'h3bf283ba),
	.w2(32'h3b9d93c7),
	.w3(32'hbb9eda39),
	.w4(32'h3ac89548),
	.w5(32'hbb19be7a),
	.w6(32'hbba836c0),
	.w7(32'hbaecb360),
	.w8(32'hbbab327b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b8059),
	.w1(32'hba8d8880),
	.w2(32'h3c01742b),
	.w3(32'hbc21577e),
	.w4(32'hbb35d7a1),
	.w5(32'hba64ecbf),
	.w6(32'hbc0f0cb5),
	.w7(32'h3b796c8c),
	.w8(32'h3bbe9649),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09038),
	.w1(32'h3bd5e3b6),
	.w2(32'hbc2428ed),
	.w3(32'h3b623a82),
	.w4(32'h3bdd165f),
	.w5(32'hbbf08ef9),
	.w6(32'hbb2add4a),
	.w7(32'h3c70acd6),
	.w8(32'hbc19ae51),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeb6bf),
	.w1(32'h39002a9c),
	.w2(32'h3acede3f),
	.w3(32'h3c1d1ae8),
	.w4(32'h3b18fc7a),
	.w5(32'h3af4f996),
	.w6(32'h3c197800),
	.w7(32'h3abd4059),
	.w8(32'hb84d7697),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f643),
	.w1(32'hbba191f5),
	.w2(32'hbb48149d),
	.w3(32'h3a2753b3),
	.w4(32'hbc1b0de6),
	.w5(32'hbc0543af),
	.w6(32'h3af4b039),
	.w7(32'hbc010900),
	.w8(32'hbc16c174),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb3682),
	.w1(32'hba9175c0),
	.w2(32'hba0d69d0),
	.w3(32'hbb981454),
	.w4(32'hbadf655b),
	.w5(32'hb8b4f712),
	.w6(32'hbb844c3e),
	.w7(32'hba3f42e3),
	.w8(32'h3b23fb8b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a91ed),
	.w1(32'h3bd62225),
	.w2(32'h3c1e3eb9),
	.w3(32'hbb60c255),
	.w4(32'h3beb15a7),
	.w5(32'h3c1bed22),
	.w6(32'hb9baf66b),
	.w7(32'h3b7df1b0),
	.w8(32'h3c611a55),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad02cf6),
	.w1(32'h3a853f9c),
	.w2(32'h3b83a076),
	.w3(32'h3bc59f95),
	.w4(32'hb7b656f5),
	.w5(32'h3c37f085),
	.w6(32'h3bd5fbac),
	.w7(32'hbad1e50a),
	.w8(32'h3c12df6d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa24a67),
	.w1(32'hbc0a9e50),
	.w2(32'hbc09574f),
	.w3(32'hbbc83525),
	.w4(32'hbbaf1b01),
	.w5(32'hbc19ef1c),
	.w6(32'hbc1c9e82),
	.w7(32'hbaf3c10f),
	.w8(32'hbb272aed),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b776a11),
	.w1(32'h3bc0943e),
	.w2(32'hbc0dff37),
	.w3(32'hb9f51d96),
	.w4(32'hba2fd45d),
	.w5(32'h3c1ef0da),
	.w6(32'hbb3e7bfa),
	.w7(32'hba39724d),
	.w8(32'h3c19d04b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43dc01),
	.w1(32'hbbb9df4b),
	.w2(32'hbb15eb6f),
	.w3(32'h3b87959f),
	.w4(32'hba32e6c0),
	.w5(32'hbbfe8b61),
	.w6(32'hbb7dc930),
	.w7(32'h3b4c6e3a),
	.w8(32'hb9e8cb59),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba031999),
	.w1(32'hba8f4678),
	.w2(32'hbba1641f),
	.w3(32'h3a25935c),
	.w4(32'hba9fecdc),
	.w5(32'hbb5a904a),
	.w6(32'h3b55f99d),
	.w7(32'hba9cb1ec),
	.w8(32'hba95f4b6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a0370),
	.w1(32'hb9f8f746),
	.w2(32'h3b28b367),
	.w3(32'hbba420d3),
	.w4(32'hba3beec0),
	.w5(32'hb8f33db2),
	.w6(32'hbb48c27d),
	.w7(32'hba6940c0),
	.w8(32'hbacc87ef),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986a1c8),
	.w1(32'h3b18e21f),
	.w2(32'h3b8af766),
	.w3(32'hbae8a2cf),
	.w4(32'hbb861ad3),
	.w5(32'h3ab5596d),
	.w6(32'h3a62bf3f),
	.w7(32'hba85223b),
	.w8(32'hbb3e2ec8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be631f3),
	.w1(32'h3b21cbce),
	.w2(32'hbb23dd03),
	.w3(32'hb9b2fe37),
	.w4(32'hb9df3975),
	.w5(32'h3b233639),
	.w6(32'h3bebe559),
	.w7(32'h3b5e0013),
	.w8(32'h3b5c5cf1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6dddf),
	.w1(32'hbc24ef1e),
	.w2(32'h3c7d51e2),
	.w3(32'hbbe81f0f),
	.w4(32'hbb5d39ae),
	.w5(32'h3ba65cf9),
	.w6(32'h3aa74f59),
	.w7(32'h3b644cdd),
	.w8(32'hbb1549fd),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06329e),
	.w1(32'h3b972f87),
	.w2(32'hbbbafd9e),
	.w3(32'h3ba07e08),
	.w4(32'hbb93bef5),
	.w5(32'h3cbc95c1),
	.w6(32'hb9935054),
	.w7(32'hbc043e0a),
	.w8(32'h3bc30f22),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951638b),
	.w1(32'h3b1754d6),
	.w2(32'hbc2580c7),
	.w3(32'h3b4df0f2),
	.w4(32'hbabedce6),
	.w5(32'h3895e14b),
	.w6(32'h3aa6a699),
	.w7(32'hbac958e9),
	.w8(32'hba5bbbac),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa6d50),
	.w1(32'h3a999287),
	.w2(32'h3bb2f58f),
	.w3(32'hbbcb8f12),
	.w4(32'h3b8f540a),
	.w5(32'hbb97b0a0),
	.w6(32'hbb8dff7c),
	.w7(32'hb8a7b042),
	.w8(32'h3b7ef46a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0155b),
	.w1(32'h3a8a8bb5),
	.w2(32'hba65060f),
	.w3(32'h3b2b4e2e),
	.w4(32'h3bf21676),
	.w5(32'h3b0c2a5e),
	.w6(32'hbaea9a50),
	.w7(32'hbae109c5),
	.w8(32'h3c0220f1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42b090),
	.w1(32'h3ba9c761),
	.w2(32'hba9fdc9a),
	.w3(32'hba7298e7),
	.w4(32'h3bde2833),
	.w5(32'hba5e8de5),
	.w6(32'h3be2ca99),
	.w7(32'h3aa6dcb4),
	.w8(32'hb98d89eb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcea855),
	.w1(32'h3b41c133),
	.w2(32'h3b3a99f8),
	.w3(32'hbba2c4ec),
	.w4(32'hbb4b5e88),
	.w5(32'hba28256e),
	.w6(32'h3b86766c),
	.w7(32'hbabe2ee2),
	.w8(32'h3ad5f7a9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93ebe7),
	.w1(32'hbb239742),
	.w2(32'hbbac6c32),
	.w3(32'h3b91568b),
	.w4(32'hbaddb977),
	.w5(32'hbbbbfd56),
	.w6(32'hb9afbf01),
	.w7(32'h3b88e136),
	.w8(32'hba73abed),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39885c7e),
	.w1(32'hbb536d52),
	.w2(32'hbb920480),
	.w3(32'h3aabcbed),
	.w4(32'h39c9971b),
	.w5(32'hbb0b597d),
	.w6(32'hbb5431e3),
	.w7(32'h3b732486),
	.w8(32'hba846291),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba864fc9),
	.w1(32'h3bcf618c),
	.w2(32'h38956148),
	.w3(32'h38f9256f),
	.w4(32'hbad4b625),
	.w5(32'h3b0bcf4a),
	.w6(32'h3b6c8e4c),
	.w7(32'h35ad6979),
	.w8(32'h3b9913ed),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f23c6),
	.w1(32'h3b36057e),
	.w2(32'h3bcdd857),
	.w3(32'h3b3450c0),
	.w4(32'hbc12248f),
	.w5(32'h3bbf88c5),
	.w6(32'h3ac8379b),
	.w7(32'hbbdcd7b1),
	.w8(32'h3909da2a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba620667),
	.w1(32'h3b4a0811),
	.w2(32'h3ba391f4),
	.w3(32'hb9d7c494),
	.w4(32'hbae3239c),
	.w5(32'h3b0ee082),
	.w6(32'hbacdc458),
	.w7(32'hbb1b4532),
	.w8(32'h38838a65),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf18cd),
	.w1(32'h3c12a657),
	.w2(32'h3cccd240),
	.w3(32'hba062775),
	.w4(32'h3cbaf63a),
	.w5(32'h3d1572cc),
	.w6(32'hba0d88b9),
	.w7(32'h3c2e2a82),
	.w8(32'h3d1f5251),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa41ba),
	.w1(32'hbbcc761b),
	.w2(32'hbbf6e38d),
	.w3(32'hba6f89d0),
	.w4(32'h3b8cb43a),
	.w5(32'hbc24e40b),
	.w6(32'hba6d399e),
	.w7(32'hbac21f64),
	.w8(32'hbb72610b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a305e3),
	.w1(32'hbabd59f1),
	.w2(32'hbaf0457d),
	.w3(32'h3b071bd1),
	.w4(32'hbaa504f8),
	.w5(32'h3bb6973a),
	.w6(32'h3b0711ec),
	.w7(32'hbbdcb8c0),
	.w8(32'h3c1a3f50),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39532f63),
	.w1(32'h3891c88b),
	.w2(32'hbb4a7c7a),
	.w3(32'h3bc900e9),
	.w4(32'h3b0402a8),
	.w5(32'h3a88a311),
	.w6(32'h3c1882fe),
	.w7(32'hbbb98dc3),
	.w8(32'hbb5ab63e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d8e3c2),
	.w1(32'hba9f54b5),
	.w2(32'hbb8a60d3),
	.w3(32'h3b1d8e57),
	.w4(32'hbba319e1),
	.w5(32'h3c31f4f7),
	.w6(32'h3afb5e50),
	.w7(32'hbb9bab85),
	.w8(32'h3c1b3c2a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba9a6),
	.w1(32'h3c0c3542),
	.w2(32'h3b922c7e),
	.w3(32'h3b3738da),
	.w4(32'h3c29177d),
	.w5(32'h3bd6ebe0),
	.w6(32'h3c1f4bdc),
	.w7(32'h3bb0c8df),
	.w8(32'h3be7a023),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae23e44),
	.w1(32'h3bf834cb),
	.w2(32'h3ba69603),
	.w3(32'hbaf511ab),
	.w4(32'h3b365960),
	.w5(32'h3c7f2efb),
	.w6(32'hbbbf13c6),
	.w7(32'h3a74f5bf),
	.w8(32'h3bde5915),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb438f),
	.w1(32'hba53ee51),
	.w2(32'hbaff85b5),
	.w3(32'hbc27e6be),
	.w4(32'hbad325e3),
	.w5(32'hbbb03bab),
	.w6(32'hbb99f9bb),
	.w7(32'hbb9792b2),
	.w8(32'hbb87fd0d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddaf6d),
	.w1(32'hba62cec8),
	.w2(32'hbbaf5bbc),
	.w3(32'hb9a93e8f),
	.w4(32'hb91bcce4),
	.w5(32'hbb990d54),
	.w6(32'h3b9d6d97),
	.w7(32'hba9f41e7),
	.w8(32'hbaabf7a6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f02f3),
	.w1(32'hbb418b48),
	.w2(32'hbb0394c9),
	.w3(32'hbb391e0d),
	.w4(32'hbafe0083),
	.w5(32'hbad61536),
	.w6(32'hbaef9c4c),
	.w7(32'hbb6695cd),
	.w8(32'hbb13752b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb172b93),
	.w1(32'hb972301d),
	.w2(32'hbba416d3),
	.w3(32'hbbb3d354),
	.w4(32'hbacbfe95),
	.w5(32'hba585619),
	.w6(32'hbad5ff88),
	.w7(32'h39e2f7c4),
	.w8(32'hba94eb73),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51539d),
	.w1(32'h3b00bc94),
	.w2(32'hbb206fef),
	.w3(32'hb96c41b7),
	.w4(32'h3bc373cd),
	.w5(32'hbad081e3),
	.w6(32'h3858b7e9),
	.w7(32'h3a17a3dd),
	.w8(32'h3b089ae1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadad304),
	.w1(32'hb9b66e6e),
	.w2(32'h3b9a86b5),
	.w3(32'hbb29c701),
	.w4(32'hbb52c64c),
	.w5(32'h3c707fa7),
	.w6(32'h3abeb08d),
	.w7(32'hbbfafd7e),
	.w8(32'h3c0e6e82),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09f317),
	.w1(32'hbc0b22cb),
	.w2(32'hbc11c53d),
	.w3(32'h3b3aa8c6),
	.w4(32'h3bbc6740),
	.w5(32'hbc272a61),
	.w6(32'h3bc480e5),
	.w7(32'hbb965be4),
	.w8(32'hbbc8c7a0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8b214),
	.w1(32'hbbcfcf16),
	.w2(32'h3aad0574),
	.w3(32'h3bd50005),
	.w4(32'h3a736991),
	.w5(32'hba70a8d7),
	.w6(32'h3bfaa422),
	.w7(32'h3b25a8ec),
	.w8(32'h3bbe5b2b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2ac8c),
	.w1(32'h3b0b94dc),
	.w2(32'h3ae15e77),
	.w3(32'h3b402339),
	.w4(32'hb9799da9),
	.w5(32'h3aebcc9c),
	.w6(32'h3ac3e644),
	.w7(32'hbb102397),
	.w8(32'h3b370b0f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020ac1),
	.w1(32'hbb7990d2),
	.w2(32'h3c329442),
	.w3(32'h38b3d82a),
	.w4(32'hbb8d6cfb),
	.w5(32'h3b452f59),
	.w6(32'h3b6856e4),
	.w7(32'h3b9cbe00),
	.w8(32'h3b45dfcb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18a286),
	.w1(32'h3a1b3671),
	.w2(32'h3b1bdd62),
	.w3(32'hbb452796),
	.w4(32'hbacb8b09),
	.w5(32'h3b7f084a),
	.w6(32'hbc1d4bab),
	.w7(32'h3b9d47d3),
	.w8(32'h3bc6b8d7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a3b98),
	.w1(32'h3b30ee17),
	.w2(32'hbb31c1d4),
	.w3(32'h3bf2c916),
	.w4(32'h3abbfc69),
	.w5(32'hbb96018d),
	.w6(32'h3bd7d6e7),
	.w7(32'h3a7d3572),
	.w8(32'hbb91d921),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad31261),
	.w1(32'h3b5df687),
	.w2(32'hba98fb51),
	.w3(32'hbbd4da8e),
	.w4(32'h39f23dc2),
	.w5(32'h3ba79dd5),
	.w6(32'hbb857349),
	.w7(32'hbb8adf74),
	.w8(32'h3b971ccf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc8732),
	.w1(32'hba3c07f8),
	.w2(32'h3b7fe30f),
	.w3(32'hbc14c1e3),
	.w4(32'h3b84f472),
	.w5(32'h3b769949),
	.w6(32'hbbe9e122),
	.w7(32'h3c0fb47d),
	.w8(32'h3c0e87f0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14f16d),
	.w1(32'hb9274150),
	.w2(32'h3a8f3d7b),
	.w3(32'h3bcbbc58),
	.w4(32'hbb5f7f39),
	.w5(32'hbada9484),
	.w6(32'h3be8f66f),
	.w7(32'hbb274758),
	.w8(32'hbb870b17),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ae8bf),
	.w1(32'hba733011),
	.w2(32'h3c0fc05e),
	.w3(32'hba8cdb89),
	.w4(32'hb944b9a6),
	.w5(32'h3c12bf40),
	.w6(32'hbb1c0f4d),
	.w7(32'h3b920ba6),
	.w8(32'h3b9f4e36),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0b57f),
	.w1(32'h3a9e9714),
	.w2(32'h3a15c81d),
	.w3(32'hbb2798f5),
	.w4(32'h3acff457),
	.w5(32'hbbbad068),
	.w6(32'hbbcaf143),
	.w7(32'h3a5ca5de),
	.w8(32'hba92ebc0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cf123),
	.w1(32'hbc29778a),
	.w2(32'hbb5463a5),
	.w3(32'h3a8cbef4),
	.w4(32'hbbdd1111),
	.w5(32'hbb8ccb53),
	.w6(32'hb92206c3),
	.w7(32'hbb5901bb),
	.w8(32'hbbf499a4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebec55),
	.w1(32'h3b94fed2),
	.w2(32'h3985a599),
	.w3(32'hbb4935e2),
	.w4(32'h3b947a2f),
	.w5(32'hbb776b19),
	.w6(32'h3b1b8e8c),
	.w7(32'hbac77401),
	.w8(32'hbab77908),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56f3df),
	.w1(32'hbba3d318),
	.w2(32'hbbbbe218),
	.w3(32'hba5c62ab),
	.w4(32'hbb635c06),
	.w5(32'hbb8a751c),
	.w6(32'hbb125376),
	.w7(32'h39c24cb1),
	.w8(32'hbac8da45),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ad19),
	.w1(32'hbb37f2ea),
	.w2(32'h3b1e8a0d),
	.w3(32'h3c2a3bc9),
	.w4(32'h3996e050),
	.w5(32'hba3f6083),
	.w6(32'h3c1d39f9),
	.w7(32'h3b225c82),
	.w8(32'h3bd3544e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38716c),
	.w1(32'h3b78c79a),
	.w2(32'h3c060fb2),
	.w3(32'h3bc5d216),
	.w4(32'hba9ceae8),
	.w5(32'h3b564b24),
	.w6(32'h39a9daa9),
	.w7(32'h3bb8746f),
	.w8(32'h3bb34bba),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fca7a),
	.w1(32'hbb69ec52),
	.w2(32'hbb8054f2),
	.w3(32'hba67ce32),
	.w4(32'hbc67da46),
	.w5(32'hbc013ff8),
	.w6(32'hbb4abbcc),
	.w7(32'hbc48ba58),
	.w8(32'hbb94b971),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17e690),
	.w1(32'hbb9deff0),
	.w2(32'hba588b89),
	.w3(32'h3b54496b),
	.w4(32'hbbf439b4),
	.w5(32'hbb48e8a2),
	.w6(32'hbad3bfe2),
	.w7(32'h38ed64e4),
	.w8(32'hbb675269),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule