module layer_10_featuremap_329(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001cb9),
	.w1(32'h3b8c31a6),
	.w2(32'hbbdcb8b4),
	.w3(32'hbb95e8b3),
	.w4(32'h3af65117),
	.w5(32'h3bce3053),
	.w6(32'h3c66088d),
	.w7(32'h3c047902),
	.w8(32'h3a0bc4c2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb529c04),
	.w1(32'hbad55949),
	.w2(32'h3b9fa84b),
	.w3(32'h39b7e54b),
	.w4(32'h3a577c8c),
	.w5(32'hba7686be),
	.w6(32'hbb9d52ef),
	.w7(32'hbac95a8b),
	.w8(32'hbb6cb41a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e6aa8),
	.w1(32'h3a0aff0a),
	.w2(32'hba0b3e96),
	.w3(32'hbb75906b),
	.w4(32'hbbf75055),
	.w5(32'hba2c3d6a),
	.w6(32'h3abfcaa0),
	.w7(32'h3ba7fd33),
	.w8(32'hba8578f8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2718e),
	.w1(32'hbb20088b),
	.w2(32'hba9f88fe),
	.w3(32'hbae4e257),
	.w4(32'hba27608b),
	.w5(32'hb9b23479),
	.w6(32'hba9723fc),
	.w7(32'hbaef57ac),
	.w8(32'hbc0d184f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7c96),
	.w1(32'hbb5a8c34),
	.w2(32'hbbb38abb),
	.w3(32'h3a1f9855),
	.w4(32'h3a3ed95a),
	.w5(32'hba1dcfad),
	.w6(32'hbb679ef2),
	.w7(32'hbbff9071),
	.w8(32'h3b5fca48),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddee8a),
	.w1(32'hbb497228),
	.w2(32'hbb765a7b),
	.w3(32'hbb00a7b9),
	.w4(32'h3aa4d2a0),
	.w5(32'h3ba60ca7),
	.w6(32'h3ba87609),
	.w7(32'hba87d123),
	.w8(32'hb8f8b1e1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab62e63),
	.w1(32'hbaeffe0c),
	.w2(32'h3aa6f41e),
	.w3(32'hb893871f),
	.w4(32'hbb5155d1),
	.w5(32'hb82adec3),
	.w6(32'hbb303d39),
	.w7(32'hbaffb84b),
	.w8(32'h3b998a4a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47abba),
	.w1(32'h3babbb48),
	.w2(32'hbb25f3fc),
	.w3(32'h387d93b0),
	.w4(32'h3b9aae4c),
	.w5(32'hbac111f8),
	.w6(32'h3bf90fba),
	.w7(32'h3c152c50),
	.w8(32'h3a353e80),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdad696),
	.w1(32'h3a73741a),
	.w2(32'hbb1b7d3e),
	.w3(32'h3b18b79f),
	.w4(32'h3b8e0468),
	.w5(32'hba11600b),
	.w6(32'h3be415f6),
	.w7(32'h3b5bc34c),
	.w8(32'h3ab7c13a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9631),
	.w1(32'hba50b606),
	.w2(32'hbac20012),
	.w3(32'hbb563664),
	.w4(32'h3aff9a8f),
	.w5(32'h3aaec42d),
	.w6(32'hba6fc600),
	.w7(32'hbb4f62e9),
	.w8(32'h3b05d350),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a547433),
	.w1(32'hbb062c3b),
	.w2(32'hbb270706),
	.w3(32'hbb762819),
	.w4(32'hbae9bc64),
	.w5(32'hb9e5d5fb),
	.w6(32'h3be089a1),
	.w7(32'h3b4515e7),
	.w8(32'hba4dbb0f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01fe00),
	.w1(32'h3bb66c2a),
	.w2(32'hbb50a0e5),
	.w3(32'hb9abe489),
	.w4(32'hbb64c7be),
	.w5(32'hbc2238ee),
	.w6(32'hba00e354),
	.w7(32'h3bc466a6),
	.w8(32'hbc23ff1c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b7b6a),
	.w1(32'h3b066a87),
	.w2(32'hba290f25),
	.w3(32'hbbfbdeae),
	.w4(32'hb9d7bd0d),
	.w5(32'h3b8c0a71),
	.w6(32'hba92a99c),
	.w7(32'hbad906e1),
	.w8(32'h3a267bfb),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f26116),
	.w1(32'hbb676f02),
	.w2(32'hbb178ec5),
	.w3(32'h3a9fadaa),
	.w4(32'h3b0e78c0),
	.w5(32'hbbcee9be),
	.w6(32'h39f87598),
	.w7(32'hba211fe8),
	.w8(32'hbb2f859f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b298bed),
	.w1(32'hbb35cc39),
	.w2(32'hbb2202ff),
	.w3(32'hbb8fd86a),
	.w4(32'h3a943bb0),
	.w5(32'h3a61bec3),
	.w6(32'hbb12fbbc),
	.w7(32'hbb37e033),
	.w8(32'hbb6817d6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc178b0),
	.w1(32'hba26996b),
	.w2(32'hb8b32ebd),
	.w3(32'hbbab5a30),
	.w4(32'h39e694a7),
	.w5(32'h3b94bc75),
	.w6(32'hbbde6887),
	.w7(32'hbb7d9ddd),
	.w8(32'hbb4e876c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab01046),
	.w1(32'hb99bb2f7),
	.w2(32'h394e22a0),
	.w3(32'hbb34219b),
	.w4(32'hbb95d109),
	.w5(32'hba331515),
	.w6(32'h39aaab6f),
	.w7(32'h39fd8f1e),
	.w8(32'hb9ca42dc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ccf39),
	.w1(32'hbb305589),
	.w2(32'hbbe38d3d),
	.w3(32'hbb559da6),
	.w4(32'hbbc9d6a6),
	.w5(32'hbbf87475),
	.w6(32'hbbedb0a9),
	.w7(32'hbc3dd3c3),
	.w8(32'hbc7fdfe0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c217),
	.w1(32'hbb650322),
	.w2(32'hbbb93ff8),
	.w3(32'hbb925686),
	.w4(32'hbbf17891),
	.w5(32'h3a2d2740),
	.w6(32'hbc3ad213),
	.w7(32'hbbfbf38c),
	.w8(32'hbb2822b9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ebba4),
	.w1(32'h3b4ec58f),
	.w2(32'h3b06c837),
	.w3(32'h3a4645c3),
	.w4(32'h388c89c7),
	.w5(32'h3af3a9ad),
	.w6(32'hbb15ca04),
	.w7(32'hbb1ec243),
	.w8(32'h3b27b2f2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb160e1d),
	.w1(32'hbaf9dc14),
	.w2(32'h3a0d139a),
	.w3(32'h3aa366d7),
	.w4(32'h3b03480e),
	.w5(32'h3b11a6d9),
	.w6(32'hb9db9c2f),
	.w7(32'hbb4b865c),
	.w8(32'hbad155d1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ce9b),
	.w1(32'h398b37e2),
	.w2(32'h3a53ae18),
	.w3(32'h3b29c515),
	.w4(32'hb8f9d865),
	.w5(32'h3acff214),
	.w6(32'hbb8a1d70),
	.w7(32'hbb20d8ab),
	.w8(32'h3a0faa02),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0e897),
	.w1(32'hbbb5833a),
	.w2(32'hbc0144d6),
	.w3(32'hbbadaf47),
	.w4(32'hbaae6060),
	.w5(32'hbc1d3ce3),
	.w6(32'hbca27818),
	.w7(32'hbc8355e5),
	.w8(32'hbc708010),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f25d8),
	.w1(32'hbb8f3c77),
	.w2(32'h3a5f4c51),
	.w3(32'hbbb57665),
	.w4(32'h3bee872e),
	.w5(32'h3ab25cf8),
	.w6(32'h3b687a1a),
	.w7(32'hbbb493a6),
	.w8(32'hbb88bca7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b871),
	.w1(32'h3b14e3fe),
	.w2(32'h3aa7f639),
	.w3(32'hbb6d49fc),
	.w4(32'hba390696),
	.w5(32'h3a82ce94),
	.w6(32'hbbe81b38),
	.w7(32'hba06e994),
	.w8(32'hbab25604),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818623),
	.w1(32'hbb824fb6),
	.w2(32'hbb4c4c53),
	.w3(32'h3ab1a3b1),
	.w4(32'hbb383aed),
	.w5(32'h3a935641),
	.w6(32'hb9b58585),
	.w7(32'hbb444fd6),
	.w8(32'hb990bb53),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df0f7f),
	.w1(32'hba2f525c),
	.w2(32'hba4020db),
	.w3(32'h3a04fc06),
	.w4(32'h3925f110),
	.w5(32'h39b05e12),
	.w6(32'hb894592e),
	.w7(32'h37e15326),
	.w8(32'h3bcaf676),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed6a41),
	.w1(32'h3aaaf51e),
	.w2(32'hbc1fb767),
	.w3(32'h3ba21b1f),
	.w4(32'h3ba01dda),
	.w5(32'h3b07ec52),
	.w6(32'h3c23b814),
	.w7(32'hbb6c2bc9),
	.w8(32'hbb23398b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949665a),
	.w1(32'h39c34434),
	.w2(32'h3a637dae),
	.w3(32'h3b9c8346),
	.w4(32'h3a31e50f),
	.w5(32'h3b29eac5),
	.w6(32'hbaba83a9),
	.w7(32'hbb5dcc7b),
	.w8(32'hbb46054a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1df48),
	.w1(32'h3b3db6be),
	.w2(32'h3bdc0781),
	.w3(32'hbae19156),
	.w4(32'hb9d220d7),
	.w5(32'hbb9336d0),
	.w6(32'hbae0accc),
	.w7(32'hbaf74ccd),
	.w8(32'h3c57d314),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0404a9),
	.w1(32'hbbb667a8),
	.w2(32'hbbba8ce2),
	.w3(32'h3c205538),
	.w4(32'h3c54b998),
	.w5(32'h3b40f031),
	.w6(32'h3c22b233),
	.w7(32'hbc09c004),
	.w8(32'hbac7b64a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6939b),
	.w1(32'h3b97c0af),
	.w2(32'h3b63c7c9),
	.w3(32'h3951cc9b),
	.w4(32'h3ab0de43),
	.w5(32'h3abfa610),
	.w6(32'hba69c207),
	.w7(32'h3c24723d),
	.w8(32'h3b522531),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaacb1b),
	.w1(32'hba80442d),
	.w2(32'h3a76855d),
	.w3(32'h3b067ebd),
	.w4(32'h399cda9e),
	.w5(32'h3b6b57c4),
	.w6(32'hbb7d70fe),
	.w7(32'h39d53b3d),
	.w8(32'hbaa848c4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba653108),
	.w1(32'h3a8a2d0f),
	.w2(32'h3b04ee94),
	.w3(32'h3b04f583),
	.w4(32'h3aaaf964),
	.w5(32'h3aeb05f4),
	.w6(32'h3979295c),
	.w7(32'hbb2a9e1b),
	.w8(32'h3adf1e3d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba754766),
	.w1(32'h3a395a7a),
	.w2(32'hb9e9349f),
	.w3(32'h3b692058),
	.w4(32'h3ae24f6c),
	.w5(32'hb9f591b8),
	.w6(32'hba07c208),
	.w7(32'hba80041b),
	.w8(32'hba5cb16b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a263a3f),
	.w1(32'h39562546),
	.w2(32'hba866b6e),
	.w3(32'hbb51561a),
	.w4(32'hbb3a036e),
	.w5(32'h3b1959e7),
	.w6(32'hba114005),
	.w7(32'hb99aea94),
	.w8(32'hba825a9e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd45a72),
	.w1(32'h3b54b028),
	.w2(32'h3aefaec6),
	.w3(32'hbb85f40f),
	.w4(32'h3b0f6386),
	.w5(32'hbaef1c44),
	.w6(32'hbc15f608),
	.w7(32'hbaefa8d0),
	.w8(32'hba2ec5e8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b485),
	.w1(32'h3a6be200),
	.w2(32'hbafe0adc),
	.w3(32'hbb9b988c),
	.w4(32'h3b845625),
	.w5(32'hbb72f389),
	.w6(32'hbabca3a9),
	.w7(32'h3aa3a926),
	.w8(32'hbb43ec55),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bf22d),
	.w1(32'h3bbb9013),
	.w2(32'h3ae3abea),
	.w3(32'hbb0f2009),
	.w4(32'h3b79821a),
	.w5(32'h3addc88c),
	.w6(32'h3c0659ab),
	.w7(32'h3ba81189),
	.w8(32'hbbd3198f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6809b1),
	.w1(32'hba0ffeef),
	.w2(32'hbb76bf36),
	.w3(32'h39ad5f3a),
	.w4(32'hbb68198c),
	.w5(32'hbb529985),
	.w6(32'hbb35ce89),
	.w7(32'hbb0e6c72),
	.w8(32'hbb33a6ae),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d83a7),
	.w1(32'hbac48034),
	.w2(32'h39da8674),
	.w3(32'hba8d8d8d),
	.w4(32'hbb68c2af),
	.w5(32'h3b127ef3),
	.w6(32'hbb09046f),
	.w7(32'hba7107a0),
	.w8(32'hbb072e98),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36909b),
	.w1(32'hb9f6a691),
	.w2(32'h3ab787c4),
	.w3(32'hbb194797),
	.w4(32'hbb7db9f4),
	.w5(32'hbb089c74),
	.w6(32'h390d4338),
	.w7(32'hba7cb398),
	.w8(32'h3b0312c8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968b6c1),
	.w1(32'hbb9bd58a),
	.w2(32'hbb67be94),
	.w3(32'hbb7c7c33),
	.w4(32'hbb877312),
	.w5(32'hbadc216e),
	.w6(32'h3aa01696),
	.w7(32'hbac08a8f),
	.w8(32'hb97769d3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb730b0f),
	.w1(32'hbb6db919),
	.w2(32'hbb1dcadd),
	.w3(32'hbbb2ca7e),
	.w4(32'h3aff2bce),
	.w5(32'hb9916373),
	.w6(32'hbc24a6ea),
	.w7(32'hbb517e8a),
	.w8(32'hbb8477fe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea2db8),
	.w1(32'h3b0c150a),
	.w2(32'h3adba098),
	.w3(32'hbbb56742),
	.w4(32'h3a9ac634),
	.w5(32'h3b7dae5d),
	.w6(32'hbb51fd29),
	.w7(32'h3a2c3bf8),
	.w8(32'hbb94f31a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e120),
	.w1(32'h3aaedcc8),
	.w2(32'h3c297bd5),
	.w3(32'hbbb74896),
	.w4(32'hbb0a551f),
	.w5(32'h3b71b140),
	.w6(32'hbc0bc272),
	.w7(32'hba1ca99d),
	.w8(32'h3a9f391b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd2533),
	.w1(32'h3b220809),
	.w2(32'h3afb7138),
	.w3(32'hbb07e042),
	.w4(32'h3a0dae5b),
	.w5(32'hbb23e8ea),
	.w6(32'hbb5b9e2f),
	.w7(32'hbaf686ee),
	.w8(32'hbb885339),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35c14e),
	.w1(32'h3a824d06),
	.w2(32'hbbc89661),
	.w3(32'h3abfb5e1),
	.w4(32'hbb028560),
	.w5(32'hbc74e395),
	.w6(32'hbc085989),
	.w7(32'hbc269e63),
	.w8(32'hbc19cb24),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcb93d),
	.w1(32'hba8a5af3),
	.w2(32'hbb842a98),
	.w3(32'hbb1a2ba6),
	.w4(32'h3b9b1d2b),
	.w5(32'h3b11ef1c),
	.w6(32'h3c676a53),
	.w7(32'h3b00a078),
	.w8(32'hbb17b8c5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13949a),
	.w1(32'hbb19ec4e),
	.w2(32'h39a72185),
	.w3(32'h3b02a103),
	.w4(32'hbb3a52f3),
	.w5(32'hbb94ff5f),
	.w6(32'hbbb72235),
	.w7(32'hbb8dfeac),
	.w8(32'hbb0fa4d0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb110e8a),
	.w1(32'hbad4b206),
	.w2(32'h3adbad0b),
	.w3(32'hbb376a2a),
	.w4(32'hbab159e3),
	.w5(32'h3b3e2696),
	.w6(32'hbb362ce9),
	.w7(32'hbaa8d011),
	.w8(32'h3b8c517b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99bb623),
	.w1(32'hb9c4e7fe),
	.w2(32'h3ae5b8a6),
	.w3(32'h3ac4da7e),
	.w4(32'h3b111e6b),
	.w5(32'hbaa21d71),
	.w6(32'h3a3aed51),
	.w7(32'hba6e7365),
	.w8(32'hbb818402),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9555ca),
	.w1(32'hbb76ee92),
	.w2(32'hbbbf4e3e),
	.w3(32'hbc07a2f2),
	.w4(32'hbbb93f94),
	.w5(32'h3ade37a2),
	.w6(32'hbaf0691b),
	.w7(32'h394c734b),
	.w8(32'hbb7da273),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98f05b),
	.w1(32'h3b81fbac),
	.w2(32'hbaa655d2),
	.w3(32'h3abf5f77),
	.w4(32'hbb85cf12),
	.w5(32'hbb856673),
	.w6(32'hbbb0600a),
	.w7(32'hbb81919e),
	.w8(32'hbb9efc67),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2d13),
	.w1(32'h3a55f09c),
	.w2(32'hba063cbf),
	.w3(32'hbb2f00b5),
	.w4(32'hbb14c4aa),
	.w5(32'hb9a81eb6),
	.w6(32'hbb852704),
	.w7(32'hbb7adcb2),
	.w8(32'hbabb5083),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a0ba8),
	.w1(32'h3adfe3bd),
	.w2(32'h3976548f),
	.w3(32'h3ada22f6),
	.w4(32'h3b551eea),
	.w5(32'hbae5040e),
	.w6(32'hbb0b70e2),
	.w7(32'hba266325),
	.w8(32'hbb0f515b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b7721),
	.w1(32'hbaf04a4b),
	.w2(32'hb9d2e768),
	.w3(32'h3b496ec5),
	.w4(32'h3b845a7e),
	.w5(32'hba8ca46d),
	.w6(32'hbb06ce19),
	.w7(32'h3a57ea4c),
	.w8(32'hbb14a46c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25633e),
	.w1(32'h3acc2aac),
	.w2(32'h39300a41),
	.w3(32'hbb20285d),
	.w4(32'hbb9d5824),
	.w5(32'h3b82e2ba),
	.w6(32'hba82866d),
	.w7(32'hba1c64fe),
	.w8(32'hba76d3c7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7d30d),
	.w1(32'hbb1c3087),
	.w2(32'hb8ec4eb1),
	.w3(32'h3b56104c),
	.w4(32'hbb0bebd5),
	.w5(32'hba98e998),
	.w6(32'hbb58284a),
	.w7(32'hbb3b9e9b),
	.w8(32'hba9b5fab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba169ad),
	.w1(32'h39ff4fbe),
	.w2(32'h3b7d7d54),
	.w3(32'h3bb7a80b),
	.w4(32'hb9ce6947),
	.w5(32'hbb074414),
	.w6(32'hbb7ac4a4),
	.w7(32'h3a9beacb),
	.w8(32'hb9c43a27),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59d89),
	.w1(32'h3b38611d),
	.w2(32'hba44ba73),
	.w3(32'hba744a5f),
	.w4(32'hbac32489),
	.w5(32'h3ae756d8),
	.w6(32'h3b174d97),
	.w7(32'hbb52a27d),
	.w8(32'hbb9eb8f0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb214600),
	.w1(32'hbb8bd24d),
	.w2(32'hba9c79c5),
	.w3(32'hbb0997ef),
	.w4(32'hbab60325),
	.w5(32'hbaa5ce44),
	.w6(32'hbb11b022),
	.w7(32'hbbb20959),
	.w8(32'hbaafeea2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0546de),
	.w1(32'h3aef4b6d),
	.w2(32'h3aae2f96),
	.w3(32'h3b324ce9),
	.w4(32'h3b6bad17),
	.w5(32'h3aa27ab7),
	.w6(32'h3b854535),
	.w7(32'h3b75ed11),
	.w8(32'h3946a181),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e7dd),
	.w1(32'h3ac68ba3),
	.w2(32'hb99d43d0),
	.w3(32'h3b26f060),
	.w4(32'h3b0dfb41),
	.w5(32'h3b888f22),
	.w6(32'hba9ac393),
	.w7(32'hb9533f39),
	.w8(32'h3b77a4cb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ecb71),
	.w1(32'h3b6161e9),
	.w2(32'h3b67256f),
	.w3(32'h3ba17544),
	.w4(32'h3b9d760b),
	.w5(32'hbb48160d),
	.w6(32'h3a1b8df0),
	.w7(32'h3b1264e5),
	.w8(32'hb9bbf29d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad26699),
	.w1(32'hbaaf7a5e),
	.w2(32'hbb19df47),
	.w3(32'hbb65756e),
	.w4(32'hbb0e755e),
	.w5(32'hbab0cf71),
	.w6(32'h3a6d39fd),
	.w7(32'hbaf25804),
	.w8(32'hbb87093b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b041b),
	.w1(32'h3bdd84e4),
	.w2(32'hbb42583f),
	.w3(32'hbbc27d0a),
	.w4(32'h3b01ac67),
	.w5(32'hbbd53962),
	.w6(32'h3b85f75c),
	.w7(32'h3c261fbd),
	.w8(32'hbba4ae7b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7d2d1),
	.w1(32'h3a414e28),
	.w2(32'h3b8a1f7b),
	.w3(32'hbc097758),
	.w4(32'h3b070435),
	.w5(32'hbb0031f8),
	.w6(32'hbbd37225),
	.w7(32'hbb45d12d),
	.w8(32'hb939ecbf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeadd39),
	.w1(32'hbb3db6f1),
	.w2(32'hbb6f8419),
	.w3(32'hbb877bc2),
	.w4(32'hbb3194aa),
	.w5(32'hbc07c87f),
	.w6(32'hbc22a7b4),
	.w7(32'hbbfda5eb),
	.w8(32'hbc44ad3c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a8c0),
	.w1(32'hba08853f),
	.w2(32'h3a016089),
	.w3(32'hbbe726b5),
	.w4(32'h3b0be4e3),
	.w5(32'hba83b0c0),
	.w6(32'hbbd19951),
	.w7(32'hbb270340),
	.w8(32'hbb50478c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992ff7f),
	.w1(32'hba86eb42),
	.w2(32'hb975d2c0),
	.w3(32'hbaa45175),
	.w4(32'hba9e98c1),
	.w5(32'hbaba0ccb),
	.w6(32'h3a652834),
	.w7(32'hbb0edecd),
	.w8(32'hbb9b1a67),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a948fc),
	.w1(32'h3ac96ccc),
	.w2(32'hbb662249),
	.w3(32'hbbac9229),
	.w4(32'hbb1d63fa),
	.w5(32'hbb30089c),
	.w6(32'h3a979824),
	.w7(32'h3aea7aba),
	.w8(32'hbbc7243d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d118f),
	.w1(32'hbafd6ffe),
	.w2(32'hbbb633a4),
	.w3(32'hbb453610),
	.w4(32'hbb20ddac),
	.w5(32'h3ba8ef60),
	.w6(32'h3b6a5bb6),
	.w7(32'h3be89785),
	.w8(32'h3b1d1694),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad21b0f),
	.w1(32'h3b81e97a),
	.w2(32'h3baeba63),
	.w3(32'h3b855732),
	.w4(32'h3b01e4a7),
	.w5(32'hbac1da69),
	.w6(32'h3b105ba3),
	.w7(32'hb9b9604a),
	.w8(32'hbbaa84e8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd3bb6),
	.w1(32'h3b4bd719),
	.w2(32'hbb89321c),
	.w3(32'hbbe9a33d),
	.w4(32'hbba7db73),
	.w5(32'hbbaf6505),
	.w6(32'h3bbddfa3),
	.w7(32'h3bf5e445),
	.w8(32'hba6139e8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b169233),
	.w1(32'h3b6a21ed),
	.w2(32'hbb4c1b65),
	.w3(32'hbac36327),
	.w4(32'hb9c0a4cd),
	.w5(32'hbb69de9e),
	.w6(32'h3a9c8a39),
	.w7(32'hbadfa543),
	.w8(32'hbbeaeafa),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f05b),
	.w1(32'hbb16655e),
	.w2(32'hbbade83c),
	.w3(32'h39a37a7f),
	.w4(32'hbbc27e44),
	.w5(32'hbbb60310),
	.w6(32'hbc1698e5),
	.w7(32'hbc3f82eb),
	.w8(32'hbc342052),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca5033),
	.w1(32'hba1b0bac),
	.w2(32'h3b0cfb99),
	.w3(32'hbaa96f0e),
	.w4(32'h3a75d476),
	.w5(32'h3af8f0af),
	.w6(32'hbb7dd0a5),
	.w7(32'hbac6196d),
	.w8(32'h3a1291eb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a2b15),
	.w1(32'h3a9c5c94),
	.w2(32'hbb876eb4),
	.w3(32'hbb12a107),
	.w4(32'h3bac03a8),
	.w5(32'hb90b895c),
	.w6(32'h3b98bda4),
	.w7(32'h39b88084),
	.w8(32'hbaf54326),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade191d),
	.w1(32'hb983e3a2),
	.w2(32'hbac34003),
	.w3(32'hba905d1a),
	.w4(32'h3b7d5c3a),
	.w5(32'h3aeca58f),
	.w6(32'h3bbc0516),
	.w7(32'hbb0bd6a6),
	.w8(32'h3ba5888e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e0979),
	.w1(32'h3bbab57b),
	.w2(32'h3b3624f6),
	.w3(32'h3bb820b4),
	.w4(32'h3c432ac2),
	.w5(32'hbb03793b),
	.w6(32'h3b9a358e),
	.w7(32'h3c004207),
	.w8(32'h39ed6b1a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a47d6b),
	.w1(32'hbb159427),
	.w2(32'hbbca573d),
	.w3(32'hbb26c480),
	.w4(32'hba538af2),
	.w5(32'hbbb24259),
	.w6(32'h3aa237f3),
	.w7(32'hbbbe6ceb),
	.w8(32'hbbd23ac0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86b2f9),
	.w1(32'hbb8cc90d),
	.w2(32'hbb62c7bf),
	.w3(32'hbb4500ea),
	.w4(32'hba52ee0f),
	.w5(32'hbb9b9915),
	.w6(32'h3a60a01b),
	.w7(32'hbab3c10f),
	.w8(32'hbb4723c0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e0f5b),
	.w1(32'hbb10a534),
	.w2(32'hbb942167),
	.w3(32'hbaa3f520),
	.w4(32'hbabe069d),
	.w5(32'h3b1059ed),
	.w6(32'h3b3340fa),
	.w7(32'h3acba8e0),
	.w8(32'hbaa03e38),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7505b0),
	.w1(32'hba4c7095),
	.w2(32'hbaff3c23),
	.w3(32'h3991b19a),
	.w4(32'hba71229a),
	.w5(32'hbb2687c2),
	.w6(32'hbaa1563f),
	.w7(32'hba2e4185),
	.w8(32'h3b976cf5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4cfc5),
	.w1(32'hbb0528ec),
	.w2(32'hba2e84f3),
	.w3(32'h3aa54a4b),
	.w4(32'h3bb2dcd2),
	.w5(32'hbaf221c8),
	.w6(32'h3c3bcaff),
	.w7(32'h3b919090),
	.w8(32'hbaee1301),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ae7c9),
	.w1(32'h3aa16637),
	.w2(32'h3a5c63d0),
	.w3(32'hbba98d68),
	.w4(32'hbb9f5469),
	.w5(32'h3b060fe0),
	.w6(32'hbb8db7d2),
	.w7(32'hba689483),
	.w8(32'hba0d22c7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeddadc),
	.w1(32'hba7f4c60),
	.w2(32'hb8b9f8d8),
	.w3(32'h3b2ba45d),
	.w4(32'hba1a36b2),
	.w5(32'h3b9f0faf),
	.w6(32'hbb00e200),
	.w7(32'hbbbd1818),
	.w8(32'h3b00c95a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f31c),
	.w1(32'hbb353b2d),
	.w2(32'h3a09298a),
	.w3(32'hbaf55b1b),
	.w4(32'hb9fb1196),
	.w5(32'h3bbc9318),
	.w6(32'hbbb95965),
	.w7(32'hbb93fa6a),
	.w8(32'h3b0bb7db),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9c49),
	.w1(32'hbbce365c),
	.w2(32'hbc0e6c41),
	.w3(32'hbbaa0a3b),
	.w4(32'hbb223d6f),
	.w5(32'hbb135ee9),
	.w6(32'hbc158f53),
	.w7(32'hbc6a274a),
	.w8(32'hbbd74a3d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9433d8),
	.w1(32'h399b6e0b),
	.w2(32'h3a8c8ffb),
	.w3(32'h3b96e4cf),
	.w4(32'h397b970c),
	.w5(32'h3bddc55d),
	.w6(32'hbab23722),
	.w7(32'hbb84f790),
	.w8(32'h3a2a6eae),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6613d),
	.w1(32'hbb55f730),
	.w2(32'hb94ae300),
	.w3(32'hba998d8a),
	.w4(32'hbb12840a),
	.w5(32'h3b410540),
	.w6(32'hbbc136de),
	.w7(32'hbb12796c),
	.w8(32'hbbce74ba),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d5d19),
	.w1(32'hb8c881d8),
	.w2(32'h3b89f95c),
	.w3(32'hb9d1063d),
	.w4(32'h3ac3a76e),
	.w5(32'h3b3c05b0),
	.w6(32'hbbab8f4b),
	.w7(32'hb9efef16),
	.w8(32'h3a85b42e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd4564),
	.w1(32'hbb40739a),
	.w2(32'hbb05f43b),
	.w3(32'hbb1103b6),
	.w4(32'hbb035d6d),
	.w5(32'hbb363dec),
	.w6(32'hbb8b6577),
	.w7(32'hbb275cd2),
	.w8(32'hbb07bf26),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893b10c),
	.w1(32'hba191ba8),
	.w2(32'hbba5a32a),
	.w3(32'hba8ca010),
	.w4(32'h3b51fd11),
	.w5(32'h39931a13),
	.w6(32'h3b1a3e6d),
	.w7(32'h3a9b61a0),
	.w8(32'hbb06d18d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a589993),
	.w1(32'h3a163bc6),
	.w2(32'hbb43282a),
	.w3(32'hbb8a20b3),
	.w4(32'hbb8b62dd),
	.w5(32'h3b84c4a5),
	.w6(32'h3ad90304),
	.w7(32'h3b7bb127),
	.w8(32'h3b1a0d8b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab0ddf),
	.w1(32'h3a9eeb18),
	.w2(32'h3b654f76),
	.w3(32'h3bc6492c),
	.w4(32'h3b8a4b6c),
	.w5(32'hbb10f0af),
	.w6(32'h3b83daab),
	.w7(32'h3b7957e1),
	.w8(32'h3c10c35f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a588),
	.w1(32'hbbb2b31d),
	.w2(32'h3a7f2bf9),
	.w3(32'h3c17508c),
	.w4(32'h3c2c171a),
	.w5(32'h3afdf999),
	.w6(32'hb8f4be2c),
	.w7(32'hbb52553c),
	.w8(32'hb989f74c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca2a56),
	.w1(32'hba511075),
	.w2(32'h3a58ae24),
	.w3(32'hbb0eaeaf),
	.w4(32'h39404fa4),
	.w5(32'hba15e391),
	.w6(32'hbbe4a9a8),
	.w7(32'hbb2052d0),
	.w8(32'hbb718473),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8706),
	.w1(32'hbbe357ae),
	.w2(32'hbbc48006),
	.w3(32'hbb78a225),
	.w4(32'hbb4b7cd2),
	.w5(32'h39ced485),
	.w6(32'hbc7e980d),
	.w7(32'hbc1b5997),
	.w8(32'hbc2ca143),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6b2b),
	.w1(32'hbb48ce1c),
	.w2(32'hbbc4698f),
	.w3(32'hbb99ceb5),
	.w4(32'h3a931c63),
	.w5(32'hbb84e5ff),
	.w6(32'hbc10e9b7),
	.w7(32'h3a6ca8a7),
	.w8(32'hbc18e3ed),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f689),
	.w1(32'h3bf3cc4f),
	.w2(32'h3c723a83),
	.w3(32'hbc090504),
	.w4(32'h3b70cce3),
	.w5(32'hbb840f19),
	.w6(32'hbc58f6ea),
	.w7(32'hbc44efa6),
	.w8(32'hbb946988),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe36d36),
	.w1(32'hbb82febb),
	.w2(32'hbc3af4bf),
	.w3(32'hbc8165cf),
	.w4(32'hbc4162b0),
	.w5(32'hbbb29dd0),
	.w6(32'hbc84623b),
	.w7(32'hbc8c4cb6),
	.w8(32'hbbae6957),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e7a8),
	.w1(32'hbb841e51),
	.w2(32'hba4743f1),
	.w3(32'h3a8d5040),
	.w4(32'h3a867760),
	.w5(32'h3b3ea4d4),
	.w6(32'hba835160),
	.w7(32'h3b8ff56e),
	.w8(32'h3bae0005),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202f6c),
	.w1(32'hbb7ec687),
	.w2(32'hbbe873a1),
	.w3(32'hbb71bbd2),
	.w4(32'hbc30c27a),
	.w5(32'hbbda44a6),
	.w6(32'h3b33fb55),
	.w7(32'hba256057),
	.w8(32'hbc03e4d5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60be0a),
	.w1(32'hbb00754a),
	.w2(32'hbb6aa9b1),
	.w3(32'h3bcfa4dd),
	.w4(32'h3b93227d),
	.w5(32'hbb771260),
	.w6(32'h3b8980db),
	.w7(32'h3a94a717),
	.w8(32'hbb80c02f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8bff),
	.w1(32'hbbab6087),
	.w2(32'hbb542ac8),
	.w3(32'h3ab557d9),
	.w4(32'h3b6c5216),
	.w5(32'h3940ec9d),
	.w6(32'h3954a58d),
	.w7(32'hb9593ff7),
	.w8(32'hba750a9e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9cbbb),
	.w1(32'hbba276c1),
	.w2(32'hbac9d113),
	.w3(32'hbb28acf5),
	.w4(32'h3a98bdd8),
	.w5(32'h3acde8e5),
	.w6(32'hbb499466),
	.w7(32'hb9a4626b),
	.w8(32'h3b0db10c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba26a3),
	.w1(32'h3ae06e7f),
	.w2(32'h3b3a1ff3),
	.w3(32'hba7d7f54),
	.w4(32'h3bc0336f),
	.w5(32'hb7feb764),
	.w6(32'hbbf1b89a),
	.w7(32'h3b0e0ee2),
	.w8(32'h384e52b0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f7d53),
	.w1(32'h3b27607d),
	.w2(32'h3b777113),
	.w3(32'hbb52bb28),
	.w4(32'h3b65d151),
	.w5(32'hbaaee3ce),
	.w6(32'hbb8a22d2),
	.w7(32'hba52c4eb),
	.w8(32'hba9a272e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d2cbb),
	.w1(32'hbb632dd9),
	.w2(32'hbb01900e),
	.w3(32'hbb2d01dc),
	.w4(32'hbaafd489),
	.w5(32'hbc721c82),
	.w6(32'hbb238c5c),
	.w7(32'h3a7c5ed1),
	.w8(32'hbc1b71ef),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da074),
	.w1(32'hbc5a3441),
	.w2(32'hbc131cda),
	.w3(32'hbc1da5c0),
	.w4(32'hbbee96c4),
	.w5(32'h3b9ac1f7),
	.w6(32'hbc0380ce),
	.w7(32'hbc007a15),
	.w8(32'h3b47ac54),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89a64f),
	.w1(32'h3b0336e6),
	.w2(32'hb809c05a),
	.w3(32'h3a9c6951),
	.w4(32'h3ac9d573),
	.w5(32'h3b9da318),
	.w6(32'hba2ec525),
	.w7(32'h3accc4f3),
	.w8(32'hbab83889),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33e0c9),
	.w1(32'hbba1e49f),
	.w2(32'hbb11acb9),
	.w3(32'h3a2161f5),
	.w4(32'h3c12f73f),
	.w5(32'h3bc4a12d),
	.w6(32'h3bbb410f),
	.w7(32'h3be74b04),
	.w8(32'h3ba87948),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b404244),
	.w1(32'h39deaf4c),
	.w2(32'h3aae9c13),
	.w3(32'h3aa08f95),
	.w4(32'h3bb8fcd4),
	.w5(32'hbc6ab835),
	.w6(32'hbb8d1305),
	.w7(32'h39fba394),
	.w8(32'hbc19dcde),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc427329),
	.w1(32'hbc87c637),
	.w2(32'hbc594537),
	.w3(32'hbbebb761),
	.w4(32'hbc2fbc91),
	.w5(32'h3abac1d9),
	.w6(32'hbc511373),
	.w7(32'hbc29dc5e),
	.w8(32'h3b1a919d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad13613),
	.w1(32'hbae31a3c),
	.w2(32'hbb18ba2d),
	.w3(32'h3a0dfce5),
	.w4(32'h3b48917c),
	.w5(32'hbb25d90a),
	.w6(32'h398a5427),
	.w7(32'hb9dc4a14),
	.w8(32'hba9f8a95),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2fb37),
	.w1(32'hbb8573f1),
	.w2(32'hb975a5f4),
	.w3(32'hbbe5b9d4),
	.w4(32'hbb7c8052),
	.w5(32'hbaa02dac),
	.w6(32'h3bcd12f5),
	.w7(32'hbb5a3231),
	.w8(32'h3b4f9863),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c4b7),
	.w1(32'h3aad3500),
	.w2(32'hbab3fb72),
	.w3(32'hbb2665c9),
	.w4(32'hbb6cf969),
	.w5(32'hba97f11d),
	.w6(32'h3adb509a),
	.w7(32'h3a04e7e2),
	.w8(32'h3b8d99bc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1b9b),
	.w1(32'h3b30565c),
	.w2(32'h3bb93dc9),
	.w3(32'hbba7ec18),
	.w4(32'hbb881cac),
	.w5(32'hbbcc6eeb),
	.w6(32'hbb1fa7bd),
	.w7(32'h3b31fdae),
	.w8(32'hba7c7eed),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c423318),
	.w1(32'h3b871341),
	.w2(32'h3b1694c3),
	.w3(32'hbc01dff9),
	.w4(32'hbc02a97b),
	.w5(32'hba81195e),
	.w6(32'hbbf87a5c),
	.w7(32'hbb7b53b7),
	.w8(32'h3a28fa90),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac73595),
	.w1(32'hbaa91533),
	.w2(32'hba7ac4db),
	.w3(32'hb8ed1a4c),
	.w4(32'hbc003010),
	.w5(32'hbb24c455),
	.w6(32'hba0911d5),
	.w7(32'hbb4272ef),
	.w8(32'h3a4ae8fd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953fa37),
	.w1(32'h3ab1ff87),
	.w2(32'h3b4b9808),
	.w3(32'hbb168d46),
	.w4(32'h3b786170),
	.w5(32'h3b8dd31f),
	.w6(32'h3bdb44a8),
	.w7(32'h3940906b),
	.w8(32'h39f8327f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1474f9),
	.w1(32'h3a39165c),
	.w2(32'hb681f010),
	.w3(32'h3b0dde54),
	.w4(32'h3a646ea5),
	.w5(32'h3b0c429b),
	.w6(32'h3b3ffd80),
	.w7(32'h3b20df7a),
	.w8(32'h3b066d3d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395cf31d),
	.w1(32'h3bdf01e6),
	.w2(32'h3b992104),
	.w3(32'hba5ce293),
	.w4(32'h3a5f3989),
	.w5(32'hbbce5a88),
	.w6(32'h3b32f342),
	.w7(32'hbab4094e),
	.w8(32'hbc821339),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5bd84),
	.w1(32'hbc00f262),
	.w2(32'hb9678634),
	.w3(32'hbc6c3da1),
	.w4(32'hbb0d8fe0),
	.w5(32'hbad094b3),
	.w6(32'hbc1abae1),
	.w7(32'hbc24a8e3),
	.w8(32'hbacd061b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5acde9),
	.w1(32'hbab0050d),
	.w2(32'hbade98e2),
	.w3(32'hbab881a6),
	.w4(32'h3acc162d),
	.w5(32'h3b4be910),
	.w6(32'hbb0c968b),
	.w7(32'hba51006e),
	.w8(32'h3afc4f69),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d6482),
	.w1(32'h3ad6ce78),
	.w2(32'h39e63adc),
	.w3(32'hbb017bb4),
	.w4(32'hbb029865),
	.w5(32'hbb4496e3),
	.w6(32'hbab4fbbd),
	.w7(32'hbb88cbb4),
	.w8(32'hbbbb94b1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf07e8f),
	.w1(32'h3a697fb0),
	.w2(32'h3a54ae2f),
	.w3(32'hbbec2afe),
	.w4(32'hbaea2d79),
	.w5(32'h3b0819b2),
	.w6(32'hbc1037b6),
	.w7(32'hbb811108),
	.w8(32'h3ba2319f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad62019),
	.w1(32'h3a72d336),
	.w2(32'hbbac7b51),
	.w3(32'hbb895d35),
	.w4(32'hbb1abd0b),
	.w5(32'hbb713cb7),
	.w6(32'hba9fdfba),
	.w7(32'hbbb03335),
	.w8(32'hbbd88afb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8d14d),
	.w1(32'hbbae6be4),
	.w2(32'hbb2e7451),
	.w3(32'h3b4df2cc),
	.w4(32'hbb5ffcfa),
	.w5(32'hbadf524f),
	.w6(32'hbb9cdfa2),
	.w7(32'hbb61ccb6),
	.w8(32'hbb24061d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb495d67),
	.w1(32'hba4b1b46),
	.w2(32'h3a655daa),
	.w3(32'h3a410afe),
	.w4(32'h3b3e5907),
	.w5(32'hbad7d669),
	.w6(32'h38a1159a),
	.w7(32'h38ef19c5),
	.w8(32'h3c9bfa47),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a230230),
	.w1(32'hbbb44dea),
	.w2(32'hbc1d53fc),
	.w3(32'hbc5d796b),
	.w4(32'hbc3ba01f),
	.w5(32'hba9a752c),
	.w6(32'h3c306641),
	.w7(32'h3be397e2),
	.w8(32'hba4478eb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978ae28),
	.w1(32'h3b5d7a55),
	.w2(32'h3b691d59),
	.w3(32'hbb1f399f),
	.w4(32'h3b483b49),
	.w5(32'h3b29c155),
	.w6(32'h3ab6fd0d),
	.w7(32'h3b655d9c),
	.w8(32'h394aa1fa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dba11),
	.w1(32'hbb89b9a0),
	.w2(32'hbba5e375),
	.w3(32'hbab09996),
	.w4(32'h3a12399d),
	.w5(32'hbbe43f06),
	.w6(32'hbb8311a4),
	.w7(32'hbba28025),
	.w8(32'hbc0ac9b4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba12cac),
	.w1(32'hbb88e31f),
	.w2(32'h394d9458),
	.w3(32'hbb83df98),
	.w4(32'h3a83105d),
	.w5(32'h3a9af113),
	.w6(32'hbae969e7),
	.w7(32'h386e1204),
	.w8(32'h3a7b5c81),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bfdf6),
	.w1(32'hbb0fee57),
	.w2(32'hbb375b61),
	.w3(32'hbab5f05c),
	.w4(32'h3b83a2cb),
	.w5(32'hbb645343),
	.w6(32'hbb97722c),
	.w7(32'h3a52ef7d),
	.w8(32'hbb13cf41),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72ba9),
	.w1(32'hbac40ad8),
	.w2(32'hbb07799c),
	.w3(32'hbb8b1832),
	.w4(32'hbacb1390),
	.w5(32'hbb49f220),
	.w6(32'hbbd20530),
	.w7(32'hbb90f480),
	.w8(32'hbb1426a7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab27860),
	.w1(32'h3b780fcd),
	.w2(32'h3bd96549),
	.w3(32'hbb8483b9),
	.w4(32'h337880ce),
	.w5(32'hb989e5e1),
	.w6(32'h3b2c1a7e),
	.w7(32'h3a60ac99),
	.w8(32'h3bedbf7a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e921c),
	.w1(32'h3c0edf63),
	.w2(32'h3c3ef89e),
	.w3(32'hba5f9c9b),
	.w4(32'h3c28fa77),
	.w5(32'hba169217),
	.w6(32'h3b8a5d5d),
	.w7(32'h3c3c88d6),
	.w8(32'h3ab8c670),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3a4b),
	.w1(32'hbc36d6a6),
	.w2(32'hbc1a812c),
	.w3(32'hb9dc14b3),
	.w4(32'hbb6070c5),
	.w5(32'hbbc44151),
	.w6(32'h3ae26e84),
	.w7(32'h3bd1c57e),
	.w8(32'h3b882664),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0fe67),
	.w1(32'hbbea3bfa),
	.w2(32'hba4c6759),
	.w3(32'hbc8c401c),
	.w4(32'h3ba23254),
	.w5(32'h3b22af37),
	.w6(32'hbb4d3d4d),
	.w7(32'h3bbb00f8),
	.w8(32'h3a3e5506),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969dd35),
	.w1(32'hb955e9e4),
	.w2(32'h3ab4ae24),
	.w3(32'h3a9370f2),
	.w4(32'h3ab14e7b),
	.w5(32'hbbcb383b),
	.w6(32'h39a7281b),
	.w7(32'h3ab638d3),
	.w8(32'hbbf9a311),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35d1b2),
	.w1(32'hbb691469),
	.w2(32'hbb3e696d),
	.w3(32'hbba6a6ca),
	.w4(32'hbbbb80cb),
	.w5(32'h3b4aa9be),
	.w6(32'h39f67ca6),
	.w7(32'hba7373a3),
	.w8(32'h3b38cb0a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b5e3),
	.w1(32'h3b086da1),
	.w2(32'h3af11aa7),
	.w3(32'h3aed70d4),
	.w4(32'h3b73f41f),
	.w5(32'hbb1129e7),
	.w6(32'h3b32d77f),
	.w7(32'h3b96003b),
	.w8(32'h3b2f6dd1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aab6e4),
	.w1(32'hb901a12f),
	.w2(32'hbaa0a99e),
	.w3(32'h39ce9648),
	.w4(32'hb9cfb1b1),
	.w5(32'hbb8feb06),
	.w6(32'h3ad95405),
	.w7(32'h3ac83376),
	.w8(32'h3ac2e2f6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c71f39),
	.w1(32'hb9e1c9f7),
	.w2(32'h3ab857ad),
	.w3(32'hbb15a55d),
	.w4(32'hbaa7c7b9),
	.w5(32'h3ade42a8),
	.w6(32'h3afd5c20),
	.w7(32'h3bcfaccc),
	.w8(32'hbb9999e8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc158168),
	.w1(32'hbacfc32c),
	.w2(32'h3b7d5511),
	.w3(32'h3b1e4497),
	.w4(32'hbc1ba495),
	.w5(32'h3a924c47),
	.w6(32'h3c442a38),
	.w7(32'hbb8110c8),
	.w8(32'hbb80df74),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29c8ce),
	.w1(32'h3a6f8836),
	.w2(32'hb939b4e4),
	.w3(32'h3ae1dbb6),
	.w4(32'hbabaaf86),
	.w5(32'h3a98caf8),
	.w6(32'h3b505dcd),
	.w7(32'h3912e06c),
	.w8(32'h3aac9388),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988ff33),
	.w1(32'h3a981fe6),
	.w2(32'h3b7047f9),
	.w3(32'h3a20d472),
	.w4(32'h3bdd28d4),
	.w5(32'hbb375063),
	.w6(32'hbb9c4469),
	.w7(32'hb97e36d7),
	.w8(32'hbba58fc3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178cd7),
	.w1(32'hbbd7931d),
	.w2(32'hbc221d03),
	.w3(32'hbb49210d),
	.w4(32'h3b90ce0f),
	.w5(32'hbaf42799),
	.w6(32'hbbd902d4),
	.w7(32'hbb900ed7),
	.w8(32'hbb736c3e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc563725),
	.w1(32'hbbbe67fd),
	.w2(32'hbc18f3eb),
	.w3(32'hbbe0b3d3),
	.w4(32'hbbc4163d),
	.w5(32'hbc4d3600),
	.w6(32'hbb3b5d38),
	.w7(32'hbbada0cd),
	.w8(32'hbc579291),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7ddf3),
	.w1(32'hbac9f276),
	.w2(32'hbb1f8bfd),
	.w3(32'hbbbb8a3b),
	.w4(32'h3b277989),
	.w5(32'h3ab85ae4),
	.w6(32'hbc3c095f),
	.w7(32'hbc767992),
	.w8(32'hbb7c49e2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec527),
	.w1(32'hbbc05085),
	.w2(32'hbaedb1fd),
	.w3(32'hbb058196),
	.w4(32'hbad570da),
	.w5(32'h3b2ae17a),
	.w6(32'hbbd4a139),
	.w7(32'h39bee262),
	.w8(32'h3aa1b357),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437e94),
	.w1(32'hbb74d666),
	.w2(32'hb9984c7b),
	.w3(32'hba317de8),
	.w4(32'hbabc2dca),
	.w5(32'hbaf24262),
	.w6(32'hba88f118),
	.w7(32'h3abf7e97),
	.w8(32'hb98e3d39),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a5fc),
	.w1(32'h3aabaafe),
	.w2(32'hb9761b8b),
	.w3(32'hbb5ccedc),
	.w4(32'h3b546c7f),
	.w5(32'hbc0dc1f4),
	.w6(32'hbbc0f56e),
	.w7(32'hba6aa84a),
	.w8(32'hbc606aca),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab406f),
	.w1(32'h3a34cdc5),
	.w2(32'h3ae93b00),
	.w3(32'hbc76b8ed),
	.w4(32'h3c9149a8),
	.w5(32'hbb0057af),
	.w6(32'hbc847c37),
	.w7(32'hbc151162),
	.w8(32'hbba5a55b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2778d6),
	.w1(32'hbb26d2a8),
	.w2(32'hb974e90a),
	.w3(32'h3b19ac23),
	.w4(32'hbba4bd6a),
	.w5(32'h3b428ed7),
	.w6(32'h3a82bd22),
	.w7(32'h3a00e1cd),
	.w8(32'hbc0228d3),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5d996),
	.w1(32'hbbdc9f09),
	.w2(32'hbc121e58),
	.w3(32'h3b29c603),
	.w4(32'h3bee552d),
	.w5(32'h3b9daa42),
	.w6(32'h3a81f06f),
	.w7(32'hbacef480),
	.w8(32'h3bbe455e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58806c),
	.w1(32'h3bb6673d),
	.w2(32'hb9de3eb6),
	.w3(32'h390f1432),
	.w4(32'hb9d98c6f),
	.w5(32'hbb45e6f8),
	.w6(32'h3bd03b3b),
	.w7(32'hb93c2929),
	.w8(32'hbbcf1212),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e3f5),
	.w1(32'hbbbd581b),
	.w2(32'hbadf0d83),
	.w3(32'hbba19e05),
	.w4(32'hbb61479c),
	.w5(32'hbb2dbbb2),
	.w6(32'hbbd8dcc0),
	.w7(32'h3b3e9c50),
	.w8(32'h3a52d09e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf06bc),
	.w1(32'hbb60388d),
	.w2(32'hbb5846f0),
	.w3(32'hbb851ceb),
	.w4(32'h3b0a632c),
	.w5(32'hbb826b63),
	.w6(32'hba4ffdeb),
	.w7(32'h386525e0),
	.w8(32'h3a125184),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b84d0),
	.w1(32'h39e2e362),
	.w2(32'hbb25b683),
	.w3(32'h39805a74),
	.w4(32'hbbd6813d),
	.w5(32'hb9be9844),
	.w6(32'h3c4a3a8d),
	.w7(32'h39b6513c),
	.w8(32'hbb607d4f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06197c),
	.w1(32'h3b39b770),
	.w2(32'h3b7054cd),
	.w3(32'h3c06c81e),
	.w4(32'h3c0a662e),
	.w5(32'h3b5bff2e),
	.w6(32'hbb2bd8f5),
	.w7(32'h3a55333f),
	.w8(32'hbabccd57),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc70651),
	.w1(32'hbbd2ee0c),
	.w2(32'hba87a41b),
	.w3(32'h3ba66d0c),
	.w4(32'h3b72c594),
	.w5(32'h3b787f89),
	.w6(32'h3aece2a4),
	.w7(32'h3bb04d29),
	.w8(32'h3a6c8807),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf9b5b),
	.w1(32'h3a532284),
	.w2(32'h3b932876),
	.w3(32'hbb28c0f4),
	.w4(32'hbb4793aa),
	.w5(32'hbaa22448),
	.w6(32'hbabe4f34),
	.w7(32'hbaa68ca1),
	.w8(32'hba0b897d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe49f82),
	.w1(32'hbb289323),
	.w2(32'hba978036),
	.w3(32'hb9f78691),
	.w4(32'hbb2a0d11),
	.w5(32'h3b0c4500),
	.w6(32'hba86b9e8),
	.w7(32'hb98978a0),
	.w8(32'hbaafffdb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca695),
	.w1(32'hbb9586dd),
	.w2(32'hbb492038),
	.w3(32'hbacf4659),
	.w4(32'h3bdfa78c),
	.w5(32'hbbf231ac),
	.w6(32'hbbe02070),
	.w7(32'h3b250f34),
	.w8(32'h3ad7d86e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ad1e),
	.w1(32'h3c1f931e),
	.w2(32'h3ba4b9f7),
	.w3(32'hbc259c6a),
	.w4(32'h3c720e49),
	.w5(32'h3b7e6835),
	.w6(32'hbc0e6b3f),
	.w7(32'h3b230041),
	.w8(32'hbb96de9c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6185),
	.w1(32'hbba67518),
	.w2(32'hb9bb1022),
	.w3(32'h3aa28611),
	.w4(32'hbad7175c),
	.w5(32'hbb57a357),
	.w6(32'hbb7d77ab),
	.w7(32'h393fb6fc),
	.w8(32'h3b58ad9d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40b25d),
	.w1(32'h39e61c82),
	.w2(32'hba1fb4bd),
	.w3(32'hbb6c391c),
	.w4(32'hba27bc3d),
	.w5(32'hb902e046),
	.w6(32'hbad72615),
	.w7(32'hb9e8dc26),
	.w8(32'h3accb6a8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cf591),
	.w1(32'h3b3d9321),
	.w2(32'h3b679920),
	.w3(32'hbc1daa16),
	.w4(32'hba9c8b65),
	.w5(32'hba0c41e7),
	.w6(32'hba31f4b9),
	.w7(32'h3aaaec52),
	.w8(32'hbb422bca),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9278cb0),
	.w1(32'hba9a1e95),
	.w2(32'h3a5ad535),
	.w3(32'hb91a4efb),
	.w4(32'h39af80d7),
	.w5(32'h3acf4bc1),
	.w6(32'hbbb3f789),
	.w7(32'hbabd5529),
	.w8(32'hbbeea652),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf4d6a),
	.w1(32'hbbabfc80),
	.w2(32'hbba844c9),
	.w3(32'hbb35a110),
	.w4(32'hbb84c33e),
	.w5(32'h3a8466d2),
	.w6(32'hbc261680),
	.w7(32'hbc189452),
	.w8(32'hbac8cb7a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9a7e2),
	.w1(32'hba43e712),
	.w2(32'h3b34c045),
	.w3(32'h3a8640ae),
	.w4(32'hbaa6cb36),
	.w5(32'h3b81f2cc),
	.w6(32'hbb9e44df),
	.w7(32'hbb014e4f),
	.w8(32'h3b36e83a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bfccc),
	.w1(32'h3aa66ee3),
	.w2(32'hb99c374b),
	.w3(32'h3a7e895a),
	.w4(32'h3b829ee9),
	.w5(32'h3b1dfab6),
	.w6(32'h3a5ed5ab),
	.w7(32'h3b5293f3),
	.w8(32'h3a0f98c9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11065f),
	.w1(32'hb8b4588b),
	.w2(32'h3a821ff7),
	.w3(32'h3b1c44f8),
	.w4(32'h3bd994b1),
	.w5(32'h3b070b70),
	.w6(32'hba8114d3),
	.w7(32'h3ba5824b),
	.w8(32'h3a354169),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb262d6b),
	.w1(32'hbb588fd8),
	.w2(32'hba712b49),
	.w3(32'h3a816740),
	.w4(32'h3aa6a8a2),
	.w5(32'hb9bac4c3),
	.w6(32'hbb34649c),
	.w7(32'h39ff049f),
	.w8(32'hb9d4aa8b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf8fb1),
	.w1(32'hbc673439),
	.w2(32'hbbaf64a3),
	.w3(32'hbbb27d41),
	.w4(32'h3a95c53c),
	.w5(32'hba76961d),
	.w6(32'hbc152c80),
	.w7(32'h396fac49),
	.w8(32'h3bfa51d3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85049e),
	.w1(32'h3b83e897),
	.w2(32'h3aa35e47),
	.w3(32'hbbc7f59d),
	.w4(32'hba7c5d4b),
	.w5(32'hbc27cb14),
	.w6(32'h3bc27a0f),
	.w7(32'hb9bf77ff),
	.w8(32'h3c03d00a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac9c35),
	.w1(32'h3c7a2b7e),
	.w2(32'h3c483bd0),
	.w3(32'hbc24d53e),
	.w4(32'h3b5397c8),
	.w5(32'h3b105395),
	.w6(32'h3b1c2ede),
	.w7(32'h3beee9b5),
	.w8(32'h3a371b10),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4a82),
	.w1(32'hbb469a82),
	.w2(32'h3943ba33),
	.w3(32'h3adcd461),
	.w4(32'hbb282236),
	.w5(32'h3c217115),
	.w6(32'h3ac32912),
	.w7(32'h3b36256c),
	.w8(32'h3c28c7cf),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50206e),
	.w1(32'h3ca56f1e),
	.w2(32'h3c83c42b),
	.w3(32'h3c5e0068),
	.w4(32'h3b6d4d96),
	.w5(32'hbb9851a5),
	.w6(32'h3ce4d6d6),
	.w7(32'h3c522a2d),
	.w8(32'h3b17e1f5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf22899),
	.w1(32'hbacdc6be),
	.w2(32'hbb957322),
	.w3(32'hbc1dee3e),
	.w4(32'hbc18f7d5),
	.w5(32'hbc16d7a0),
	.w6(32'h3bfb6ba8),
	.w7(32'hbbdd5167),
	.w8(32'hbbcf31dc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba941d1d),
	.w1(32'h3a511e1e),
	.w2(32'hbba22412),
	.w3(32'hbbec7791),
	.w4(32'h39f254b3),
	.w5(32'hbbf97645),
	.w6(32'hbc27999a),
	.w7(32'hbc01cb7f),
	.w8(32'hbbc518f8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f776c),
	.w1(32'h3b523666),
	.w2(32'h3baaa538),
	.w3(32'hbb914380),
	.w4(32'hbbd4f4c4),
	.w5(32'h3afcec7d),
	.w6(32'h3b5e6a94),
	.w7(32'hba9db1c9),
	.w8(32'h37ec5fcb),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae28d81),
	.w1(32'hbbe8714c),
	.w2(32'hbb4a1918),
	.w3(32'hbb12948b),
	.w4(32'hbad95232),
	.w5(32'hb9e92f34),
	.w6(32'hbbc2796f),
	.w7(32'hbb2bfd0e),
	.w8(32'hbb3d947a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d4ecc),
	.w1(32'h3acfc4e1),
	.w2(32'h3b8a6178),
	.w3(32'h39672197),
	.w4(32'hbbe7fa18),
	.w5(32'h3acb4641),
	.w6(32'hbc0e6275),
	.w7(32'hbc078f09),
	.w8(32'hbb84b89f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc07e9),
	.w1(32'hba83ad59),
	.w2(32'hba45143c),
	.w3(32'h3a9fc3b4),
	.w4(32'h3a6132d6),
	.w5(32'h3b275246),
	.w6(32'h3ae18b6e),
	.w7(32'h3b88cb46),
	.w8(32'hbb22b61f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb663f09),
	.w1(32'hbb67c538),
	.w2(32'hbb86084f),
	.w3(32'h3b2e4002),
	.w4(32'h3aab0bf2),
	.w5(32'h3acb7cbe),
	.w6(32'hba41ad1f),
	.w7(32'hbb19c811),
	.w8(32'h3c9a1cab),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643aa1),
	.w1(32'hbb957613),
	.w2(32'hbbc2761f),
	.w3(32'h3b4c1b93),
	.w4(32'hb9355587),
	.w5(32'hbc461648),
	.w6(32'h3cf158b2),
	.w7(32'h3cbdca1b),
	.w8(32'hbc0ff016),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cc0ff),
	.w1(32'hbbc4c7ee),
	.w2(32'hbc0b0f49),
	.w3(32'hbc2f55f7),
	.w4(32'hbc210525),
	.w5(32'h3c83e279),
	.w6(32'hbb30f9ac),
	.w7(32'hbc0dc713),
	.w8(32'h3c3d78d3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ff70f),
	.w1(32'h3cfd11f8),
	.w2(32'h3cef3283),
	.w3(32'h3c5f5b91),
	.w4(32'hb9eb7216),
	.w5(32'h3b8628c7),
	.w6(32'h3d12df27),
	.w7(32'h3c93ff43),
	.w8(32'h3cb4d87f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf6537),
	.w1(32'h3cbc79e9),
	.w2(32'h3c953557),
	.w3(32'h3b667afd),
	.w4(32'h3c12f0d6),
	.w5(32'hbb5fa850),
	.w6(32'h3cb5425e),
	.w7(32'h3c8a1934),
	.w8(32'h398409dd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb84c28),
	.w1(32'hbb8085e5),
	.w2(32'h39b49447),
	.w3(32'hbb5a180c),
	.w4(32'hbb1be125),
	.w5(32'h3b09ae83),
	.w6(32'hbb0ffd9a),
	.w7(32'hba273449),
	.w8(32'h3abfc650),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aa742),
	.w1(32'h3aa86432),
	.w2(32'h3b55ca42),
	.w3(32'hbb571793),
	.w4(32'h3a8ecd40),
	.w5(32'h3aa3685b),
	.w6(32'hbbb91838),
	.w7(32'hb9aad980),
	.w8(32'h3b9fab3c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c26da),
	.w1(32'h3ca96cab),
	.w2(32'h3cb1adf6),
	.w3(32'hbb5f57f0),
	.w4(32'hba7fb108),
	.w5(32'hbb4327ca),
	.w6(32'h3c07436f),
	.w7(32'h3be1b37f),
	.w8(32'h3b2e00e9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a865222),
	.w1(32'h3aac2f84),
	.w2(32'hb9110a40),
	.w3(32'hbbbd395e),
	.w4(32'hba37406c),
	.w5(32'h3ab5e48b),
	.w6(32'hbc5404de),
	.w7(32'hbb8cabb2),
	.w8(32'hb9891cbc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40f008),
	.w1(32'hbb43edb6),
	.w2(32'hbb05207f),
	.w3(32'hb9c1bbdd),
	.w4(32'h3a3ad1a5),
	.w5(32'h39e5038d),
	.w6(32'hbacc6dda),
	.w7(32'h3b6f1c21),
	.w8(32'hbb38ec2f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7fcf6),
	.w1(32'hbb5f8dc4),
	.w2(32'hbb1e14ad),
	.w3(32'hbb08bc70),
	.w4(32'hb8a5fcc3),
	.w5(32'h3a8d77c3),
	.w6(32'hbbb4592d),
	.w7(32'hbad54284),
	.w8(32'hbb373be1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f70947),
	.w1(32'h3b03ea29),
	.w2(32'hbad8435c),
	.w3(32'hb9413366),
	.w4(32'h3a91eb52),
	.w5(32'hbb4293db),
	.w6(32'hbb9cff98),
	.w7(32'hbba955e7),
	.w8(32'hba068874),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac2fb3),
	.w1(32'hbb483a00),
	.w2(32'hbb219883),
	.w3(32'h3ae661f6),
	.w4(32'h3b89486f),
	.w5(32'hbaf06c5f),
	.w6(32'h3b1f3cc5),
	.w7(32'h3931b8ef),
	.w8(32'h3991f04f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b082a88),
	.w1(32'h3b81eae7),
	.w2(32'h3b9e8638),
	.w3(32'hb723a24c),
	.w4(32'h3ac14add),
	.w5(32'hbb317f0b),
	.w6(32'h3b04729e),
	.w7(32'hb972cb0c),
	.w8(32'h3a04399b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5aadeb),
	.w1(32'h3905f872),
	.w2(32'hbac366dd),
	.w3(32'hbb45a8ab),
	.w4(32'h3b7f40a1),
	.w5(32'hbc2a8b93),
	.w6(32'h3a25b7b9),
	.w7(32'h3bab6b09),
	.w8(32'hbb69ef4a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb901366),
	.w1(32'hbafcc770),
	.w2(32'hbbdc1de4),
	.w3(32'hbc4b7b3e),
	.w4(32'hbafe9fb9),
	.w5(32'h3a31069f),
	.w6(32'hbb774c3e),
	.w7(32'hba929fa6),
	.w8(32'h3afea74b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bab4d),
	.w1(32'hba5c480e),
	.w2(32'hba892ef8),
	.w3(32'h39f7935c),
	.w4(32'h3b034126),
	.w5(32'hbb589676),
	.w6(32'h3b126e37),
	.w7(32'h3a4f7e8d),
	.w8(32'hba53eb8c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d654a),
	.w1(32'h3a9860f0),
	.w2(32'h3ba374d0),
	.w3(32'hbb4898b9),
	.w4(32'h3b9816ea),
	.w5(32'h39f3be3c),
	.w6(32'hbbaab376),
	.w7(32'h3b2fe3dc),
	.w8(32'h38bd12a8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc453),
	.w1(32'h38bcfe1f),
	.w2(32'h3a95e7c1),
	.w3(32'h3a0beb0d),
	.w4(32'h3bc682dc),
	.w5(32'hbb0be273),
	.w6(32'h38abcad3),
	.w7(32'h3b6238c6),
	.w8(32'h3a8a7dac),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9b91),
	.w1(32'hba89970a),
	.w2(32'h3ac977dd),
	.w3(32'hbb96d5d2),
	.w4(32'hbb678dc2),
	.w5(32'h3b752660),
	.w6(32'hbba2299d),
	.w7(32'hbb179dc8),
	.w8(32'h362bbabd),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869b9ae),
	.w1(32'hbb5e4694),
	.w2(32'hba216e76),
	.w3(32'h3b463f81),
	.w4(32'h3b7b25f8),
	.w5(32'h3aae1721),
	.w6(32'hbb30ebc0),
	.w7(32'h3a33ca7a),
	.w8(32'hbbb95ce5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b336485),
	.w1(32'h3bcff98a),
	.w2(32'h3bd7b5a1),
	.w3(32'hbaa831a5),
	.w4(32'hbb2008d8),
	.w5(32'hbb2f1ca9),
	.w6(32'hbc18394f),
	.w7(32'hbc1969a9),
	.w8(32'h3ad7bd68),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0afe3b),
	.w1(32'hba3cab7e),
	.w2(32'h3a87fee3),
	.w3(32'hbb5b861d),
	.w4(32'hbb8bdff7),
	.w5(32'h3c238c9b),
	.w6(32'hbb8d5e6e),
	.w7(32'hbb8b1a3e),
	.w8(32'hba7f5a8d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b175aa3),
	.w1(32'h3c1263b2),
	.w2(32'h3c13fc2f),
	.w3(32'h3babe061),
	.w4(32'h3c549034),
	.w5(32'hbb9967e9),
	.w6(32'hbc23e254),
	.w7(32'hbb95a8e9),
	.w8(32'hbc08a61d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8c4cb),
	.w1(32'h3b866b6e),
	.w2(32'h3b9e4cfc),
	.w3(32'h39e549e4),
	.w4(32'h3badbc46),
	.w5(32'h3b3b30a4),
	.w6(32'hbafc46a8),
	.w7(32'hbb8085ba),
	.w8(32'hba49b16c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e85ca),
	.w1(32'hbb987457),
	.w2(32'h3ac245be),
	.w3(32'h3b188640),
	.w4(32'hbb9cc70a),
	.w5(32'hbc323cd5),
	.w6(32'h3a2a37e6),
	.w7(32'h3a61ec56),
	.w8(32'hbc14d3a3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81642b),
	.w1(32'hb979e2f6),
	.w2(32'hba54e93b),
	.w3(32'hbc303587),
	.w4(32'hbc2afb60),
	.w5(32'hb7ab9794),
	.w6(32'hbb000888),
	.w7(32'hbbdb94a6),
	.w8(32'h3ab72a11),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adca911),
	.w1(32'hba1969ce),
	.w2(32'hba6dadbb),
	.w3(32'h3a43f043),
	.w4(32'h3b8f69cb),
	.w5(32'hbba08f61),
	.w6(32'h398da620),
	.w7(32'h3b50b58a),
	.w8(32'h39c72752),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367247),
	.w1(32'hbc0a9eb1),
	.w2(32'hba9e7319),
	.w3(32'hbb8dce49),
	.w4(32'h3b69882c),
	.w5(32'h3b5ba907),
	.w6(32'hbba2a147),
	.w7(32'h3b864f9a),
	.w8(32'h3b821991),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6302),
	.w1(32'hbaf7c891),
	.w2(32'hbb8a99f7),
	.w3(32'hbb220f76),
	.w4(32'hbbb4baea),
	.w5(32'hbbca2db7),
	.w6(32'hbbbb6bcd),
	.w7(32'hbbe56b19),
	.w8(32'hbc2302a7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc3900),
	.w1(32'hbb85ce15),
	.w2(32'hbbd87332),
	.w3(32'hbb8eb5e6),
	.w4(32'hbbe554fc),
	.w5(32'h3b63a6e3),
	.w6(32'hbbf65ef9),
	.w7(32'hbc2f93b6),
	.w8(32'hbb2ffa86),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7883b5),
	.w1(32'hbb96895f),
	.w2(32'hbbe7288b),
	.w3(32'hbbdfcada),
	.w4(32'hbbb87c6a),
	.w5(32'hbb672b45),
	.w6(32'h3b55750f),
	.w7(32'h3b53d434),
	.w8(32'h3af1f56f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b469a46),
	.w1(32'h3b7fe205),
	.w2(32'h3bc939b3),
	.w3(32'hb9ae9312),
	.w4(32'h3a3a6752),
	.w5(32'h3a2302a2),
	.w6(32'h3b9b04a1),
	.w7(32'h3ba31099),
	.w8(32'hbad79042),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a17bf),
	.w1(32'hbacc789e),
	.w2(32'hbb0481a6),
	.w3(32'hbae35890),
	.w4(32'hbae0a68f),
	.w5(32'h3b9d0fcd),
	.w6(32'hbb2119bd),
	.w7(32'hbb0de30f),
	.w8(32'h3ad45c76),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab2c55),
	.w1(32'h3b469487),
	.w2(32'h3b76d080),
	.w3(32'h3b48b24f),
	.w4(32'h3b1ac2dd),
	.w5(32'hbad4d2c2),
	.w6(32'h3ac99269),
	.w7(32'h3aafdfcb),
	.w8(32'h3a14e81b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65fb62),
	.w1(32'hba597cca),
	.w2(32'hba70da47),
	.w3(32'hbb2c055a),
	.w4(32'h3b6d25ea),
	.w5(32'hbb239be0),
	.w6(32'hbbdfdcec),
	.w7(32'hba39886b),
	.w8(32'hb8f938ae),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad087c1),
	.w1(32'hbc370091),
	.w2(32'hbc466c36),
	.w3(32'hbbb16753),
	.w4(32'h3b0a4989),
	.w5(32'hbb4d5e96),
	.w6(32'h3ad2b3d5),
	.w7(32'h3b363d17),
	.w8(32'hbb8db060),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e9e8c),
	.w1(32'hbb174fbc),
	.w2(32'hbb2c3036),
	.w3(32'hbb232e2b),
	.w4(32'h393a0119),
	.w5(32'hbb14b451),
	.w6(32'hbb8e8420),
	.w7(32'hbb26a14f),
	.w8(32'hbb978684),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54239e),
	.w1(32'hbb9e7f33),
	.w2(32'hbba2e729),
	.w3(32'hbc409ef2),
	.w4(32'hbbdb5608),
	.w5(32'hbb20137a),
	.w6(32'hbc20c365),
	.w7(32'hbc126301),
	.w8(32'hbbb0015d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb322aa2),
	.w1(32'hba922d1c),
	.w2(32'hbb3f629b),
	.w3(32'hba653247),
	.w4(32'h3b776cb5),
	.w5(32'h3b8318f8),
	.w6(32'hbb479fd6),
	.w7(32'h3986efe8),
	.w8(32'h3ac93511),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b297a49),
	.w1(32'hbb83e98e),
	.w2(32'hbb4fee52),
	.w3(32'hba86e88d),
	.w4(32'h3b6b4452),
	.w5(32'hb9304bdc),
	.w6(32'hbb563c88),
	.w7(32'h3a655e11),
	.w8(32'hbae59288),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb303a4),
	.w1(32'hbaf1a2df),
	.w2(32'hbb7541d5),
	.w3(32'hbbfea473),
	.w4(32'hbacf8924),
	.w5(32'h3b7c546d),
	.w6(32'hbc6f159f),
	.w7(32'hbbf669d0),
	.w8(32'hbb93836a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ed537),
	.w1(32'hb9d69fe1),
	.w2(32'h3aeca194),
	.w3(32'h3b647db1),
	.w4(32'h3bdcdd02),
	.w5(32'hbb6ada7e),
	.w6(32'h3ab3de99),
	.w7(32'h3b88bea5),
	.w8(32'h3893a4b7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6115af),
	.w1(32'h3a5ce5a3),
	.w2(32'h3acdd710),
	.w3(32'hbb222470),
	.w4(32'hbb79b5b4),
	.w5(32'hbaca6594),
	.w6(32'hbbfe7a3b),
	.w7(32'h3a847974),
	.w8(32'hba97fce4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba435eb),
	.w1(32'hba20a3f1),
	.w2(32'hba2732ba),
	.w3(32'hbb15628e),
	.w4(32'hbb0872fc),
	.w5(32'hbaece8bf),
	.w6(32'h3bfa1b8e),
	.w7(32'hbb9231b7),
	.w8(32'hbba4fa94),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6636f0),
	.w1(32'h3bdcf9b2),
	.w2(32'h3a036311),
	.w3(32'hbbad3ea3),
	.w4(32'h3b28bd6c),
	.w5(32'h3992d7b2),
	.w6(32'h3b2af941),
	.w7(32'h3ac2c584),
	.w8(32'h3b8a931c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817fad),
	.w1(32'h3c0e47c3),
	.w2(32'h37734bcd),
	.w3(32'h3b1f26ce),
	.w4(32'hbaa1daec),
	.w5(32'hbb15127e),
	.w6(32'h3ae11b96),
	.w7(32'hb8f31707),
	.w8(32'hbb761bed),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca412d),
	.w1(32'h39df1e20),
	.w2(32'hbaec8e17),
	.w3(32'h3a416d80),
	.w4(32'hbb04c93f),
	.w5(32'hbafa3915),
	.w6(32'hbb15cff0),
	.w7(32'hbba7f6e0),
	.w8(32'hbb75fa0a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78d245),
	.w1(32'h3ba2cc4f),
	.w2(32'hb911a971),
	.w3(32'h3b9502fd),
	.w4(32'h3b23f87f),
	.w5(32'hbac9ab67),
	.w6(32'h3c4648f4),
	.w7(32'h3b7d4ae2),
	.w8(32'hbb7c22af),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdb336),
	.w1(32'h3bb2c7a8),
	.w2(32'hbaab3be5),
	.w3(32'h3a1d2923),
	.w4(32'h3b4a9c03),
	.w5(32'hb98c9bad),
	.w6(32'hbaa9db1a),
	.w7(32'hbafde48a),
	.w8(32'h3ab10ea4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd1d61),
	.w1(32'h3abba34e),
	.w2(32'hba875581),
	.w3(32'hbc025b0c),
	.w4(32'hba5107aa),
	.w5(32'hbac8454a),
	.w6(32'hbbeddbae),
	.w7(32'hbbce5a05),
	.w8(32'hbbe162c3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19f859),
	.w1(32'h3b0204d9),
	.w2(32'h3c098dcb),
	.w3(32'hba168b46),
	.w4(32'h3b805a1a),
	.w5(32'h3b990bba),
	.w6(32'h3bca8803),
	.w7(32'h3c22b4b6),
	.w8(32'h3be11160),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba632966),
	.w1(32'hba6bc14e),
	.w2(32'h3b0a936f),
	.w3(32'h3b8a2d79),
	.w4(32'h3bd97d17),
	.w5(32'hbbb58642),
	.w6(32'hbba19af2),
	.w7(32'hb98b956c),
	.w8(32'hbabf77a1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53f35),
	.w1(32'hbb356657),
	.w2(32'hbbb07c58),
	.w3(32'hbc1624f7),
	.w4(32'hb9753e1a),
	.w5(32'h3b9c5ab9),
	.w6(32'hbab444b0),
	.w7(32'hbb731914),
	.w8(32'h3babf939),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd21a60),
	.w1(32'h3b7cf3b7),
	.w2(32'h3a97593b),
	.w3(32'hbab498ae),
	.w4(32'h3a98a152),
	.w5(32'h3baa2578),
	.w6(32'hba9324ba),
	.w7(32'h3b4e4c27),
	.w8(32'h3afc4341),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c7d5),
	.w1(32'hbb7d825d),
	.w2(32'hba3f98dd),
	.w3(32'h3aff9aad),
	.w4(32'h3a09db37),
	.w5(32'hbbd8e6c6),
	.w6(32'hbbad935e),
	.w7(32'hbb1778b6),
	.w8(32'hbb80af65),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a0054),
	.w1(32'hbbefed5e),
	.w2(32'hbaeb39ce),
	.w3(32'hbb47def6),
	.w4(32'hbb934491),
	.w5(32'h3b132fe8),
	.w6(32'hbc0138a7),
	.w7(32'hbac7a306),
	.w8(32'h3ae72adc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e8882),
	.w1(32'hbb08c869),
	.w2(32'h388f31ff),
	.w3(32'hbb472f49),
	.w4(32'h3a2499c9),
	.w5(32'hbad8926a),
	.w6(32'hbb87a469),
	.w7(32'hbae45986),
	.w8(32'hbbceb517),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c000),
	.w1(32'h3adb79f6),
	.w2(32'h3a742614),
	.w3(32'hbaa9e4d9),
	.w4(32'h3aca8ce9),
	.w5(32'hbb4bc2d8),
	.w6(32'hbb3496f4),
	.w7(32'h39d0e3ca),
	.w8(32'hb735618f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcfb2a),
	.w1(32'hbb7c52b1),
	.w2(32'hba8ec6b3),
	.w3(32'h39036a0a),
	.w4(32'hb90f68ac),
	.w5(32'hba81625d),
	.w6(32'h3a3eaec0),
	.w7(32'h3b02803e),
	.w8(32'h3b2960cc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b757170),
	.w1(32'hbb0a8387),
	.w2(32'hbaac058d),
	.w3(32'h3a36d208),
	.w4(32'hbba6c7cb),
	.w5(32'h3b71f0af),
	.w6(32'h3b57ebcb),
	.w7(32'h3a1a7c39),
	.w8(32'hbb30f4c8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332211),
	.w1(32'h3bdc3802),
	.w2(32'hba026374),
	.w3(32'hbc47c5ba),
	.w4(32'hb9ded2a2),
	.w5(32'h3a4737d9),
	.w6(32'hba5b579e),
	.w7(32'hbb49f8aa),
	.w8(32'hbbd421cf),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86dfd2),
	.w1(32'hba136dee),
	.w2(32'h3a148b7a),
	.w3(32'h3b99c8a8),
	.w4(32'hbc0d20b5),
	.w5(32'h3aadee28),
	.w6(32'h3c8421ee),
	.w7(32'h3a6a2155),
	.w8(32'h3b19e4aa),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5295fa),
	.w1(32'h3bf8815b),
	.w2(32'hbc03cc57),
	.w3(32'hbb1706c8),
	.w4(32'h3aa74738),
	.w5(32'h3a7d9764),
	.w6(32'hbc3b821e),
	.w7(32'hbab96ba4),
	.w8(32'h3b55f532),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375272),
	.w1(32'hbb53dcd3),
	.w2(32'hbb1bddab),
	.w3(32'hbb9ae45b),
	.w4(32'h3a39280b),
	.w5(32'h3ae62afc),
	.w6(32'hbbc94fe1),
	.w7(32'hbb7103a2),
	.w8(32'hba93eebd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a909254),
	.w1(32'h3bc4a902),
	.w2(32'h3a42a5a6),
	.w3(32'h3b1cbac5),
	.w4(32'h389546ad),
	.w5(32'hb9a14d73),
	.w6(32'h3bdaf965),
	.w7(32'hba2e8e3a),
	.w8(32'h3b27e3fa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c9f30),
	.w1(32'hbb0dcafa),
	.w2(32'hbb9300d7),
	.w3(32'hbbb347e1),
	.w4(32'hbb6f68b0),
	.w5(32'hbbe58f67),
	.w6(32'hbbb26cb9),
	.w7(32'hbbc52f44),
	.w8(32'hbc133e3b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule