module layer_8_featuremap_175(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedb216),
	.w1(32'hbbce476d),
	.w2(32'hbb7e50bd),
	.w3(32'hbb2931cc),
	.w4(32'hbb93eceb),
	.w5(32'hbbd24536),
	.w6(32'hbc1f39ec),
	.w7(32'hbc5cae16),
	.w8(32'hbb08ae11),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7adf1e),
	.w1(32'h3b829a34),
	.w2(32'hba994ed3),
	.w3(32'hbaae5c43),
	.w4(32'h3b22e747),
	.w5(32'hba7c0fa0),
	.w6(32'h3b996df2),
	.w7(32'h399d82c5),
	.w8(32'h36fea541),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f2206),
	.w1(32'hbb4dcb3f),
	.w2(32'hbc345208),
	.w3(32'hba82bb34),
	.w4(32'hbc13bde0),
	.w5(32'hbb7e199d),
	.w6(32'h39dee6dc),
	.w7(32'hbb898d24),
	.w8(32'h3b288a92),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4f88),
	.w1(32'h3ba86f30),
	.w2(32'hbb0ce10a),
	.w3(32'h3a657633),
	.w4(32'h3aa78cb6),
	.w5(32'hbaf8f414),
	.w6(32'hbb1dfa87),
	.w7(32'h3abec392),
	.w8(32'h3c000d99),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0192b5),
	.w1(32'h3c03c0cf),
	.w2(32'hbac42fdf),
	.w3(32'h3b05386c),
	.w4(32'h3a8b7ae9),
	.w5(32'hbbdb695f),
	.w6(32'h3c226161),
	.w7(32'h3bc3b668),
	.w8(32'hba271e96),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c137a),
	.w1(32'h3bbeba7f),
	.w2(32'h3c95716b),
	.w3(32'hbb7af761),
	.w4(32'h3c33a49d),
	.w5(32'h3be7ebaf),
	.w6(32'hbb6c44c1),
	.w7(32'h3b86e281),
	.w8(32'h3c4d1a0d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab231ba),
	.w1(32'h3a281aba),
	.w2(32'h3b0c144a),
	.w3(32'hbbb09ce2),
	.w4(32'h3a66058b),
	.w5(32'h39b56135),
	.w6(32'h3a5b5b0e),
	.w7(32'h3ab4fffe),
	.w8(32'h3a0cab30),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79b4a2),
	.w1(32'hbc081562),
	.w2(32'h3b9b4f35),
	.w3(32'h3b2ddffa),
	.w4(32'hb95655d4),
	.w5(32'h3c97a043),
	.w6(32'hba9037f9),
	.w7(32'hbb507c51),
	.w8(32'h3be383d7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c555b21),
	.w1(32'hb90e1717),
	.w2(32'hbc2ab825),
	.w3(32'h3bf5d3f0),
	.w4(32'hbbc8d24f),
	.w5(32'hbc56e27c),
	.w6(32'h3b9594c8),
	.w7(32'hbb3f79d7),
	.w8(32'hbc0bffda),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d361f),
	.w1(32'hba5a7c0b),
	.w2(32'hbbb2c165),
	.w3(32'hbb9e3953),
	.w4(32'hbb2598aa),
	.w5(32'hbb23f9c6),
	.w6(32'h3946fbd7),
	.w7(32'hbbc6d0b3),
	.w8(32'h39e37e9c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08a05d),
	.w1(32'hb9a29c91),
	.w2(32'h37ca12eb),
	.w3(32'hbaa0e4b1),
	.w4(32'h3ba84012),
	.w5(32'h3ad7465a),
	.w6(32'hba29876a),
	.w7(32'h3b330743),
	.w8(32'h3b5eb4df),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d134d8),
	.w1(32'hbaf65f22),
	.w2(32'hbb13f28e),
	.w3(32'hbb857272),
	.w4(32'h3a7b386c),
	.w5(32'hbb06f06b),
	.w6(32'hb9ac86c9),
	.w7(32'hbb22024e),
	.w8(32'h3a9ac2ac),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a03ec7),
	.w1(32'h3b0b2dae),
	.w2(32'hbae321a5),
	.w3(32'hbb418c9a),
	.w4(32'hba8fb44f),
	.w5(32'hb998ad3a),
	.w6(32'hbb7ffffa),
	.w7(32'h3b82895d),
	.w8(32'h3a96ede4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893f3ac),
	.w1(32'hb8346e60),
	.w2(32'h3a1c475c),
	.w3(32'h3ad4379e),
	.w4(32'hba06f6f1),
	.w5(32'h3b954cb0),
	.w6(32'h3b735e0b),
	.w7(32'h39ec5ff5),
	.w8(32'h3a0aaa4d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395f64),
	.w1(32'hbafe849c),
	.w2(32'h3afa4844),
	.w3(32'h3c13463f),
	.w4(32'hbb07103d),
	.w5(32'h3b34d4cf),
	.w6(32'hbb143d8e),
	.w7(32'h39e588a6),
	.w8(32'h3a226b00),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7be7bf),
	.w1(32'h3bf2c74f),
	.w2(32'h3ac6eb79),
	.w3(32'h3bab1890),
	.w4(32'h3b6fd6be),
	.w5(32'hbc1729f5),
	.w6(32'hbb194a45),
	.w7(32'h3a97dca3),
	.w8(32'h3a436a50),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb925),
	.w1(32'h3b8790c1),
	.w2(32'hbbc7041a),
	.w3(32'hbaf12d63),
	.w4(32'hbbb23bbe),
	.w5(32'hbc0233e0),
	.w6(32'hb9d9afbc),
	.w7(32'hbb1020a4),
	.w8(32'hbbf0d836),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0d66),
	.w1(32'h3a41f208),
	.w2(32'hbc173785),
	.w3(32'hbba1a3b8),
	.w4(32'hbb337dda),
	.w5(32'hbb8faabd),
	.w6(32'h3c08ad38),
	.w7(32'hbb55067b),
	.w8(32'hb9d52175),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e1147),
	.w1(32'h3af89f0b),
	.w2(32'h3b0e6f3f),
	.w3(32'h3c3a9a84),
	.w4(32'hbb25cf9e),
	.w5(32'h371f2b43),
	.w6(32'h39ed8c10),
	.w7(32'hb9bfcc2d),
	.w8(32'h39e7b4ff),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97e396),
	.w1(32'hba83eb50),
	.w2(32'h3b315970),
	.w3(32'h3c16dcc0),
	.w4(32'hbb5210c9),
	.w5(32'hba42da8b),
	.w6(32'hbbbf6e4d),
	.w7(32'hbb485a18),
	.w8(32'hbae15098),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaaa6a),
	.w1(32'h3bdf2c69),
	.w2(32'h3b643382),
	.w3(32'hba3d8af6),
	.w4(32'hbbe760d8),
	.w5(32'hbc4cbed5),
	.w6(32'h3b0f38ae),
	.w7(32'h3b9bc126),
	.w8(32'hba8df2ce),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a31c),
	.w1(32'h3bbdf1e9),
	.w2(32'h3c160641),
	.w3(32'hbc2f82f5),
	.w4(32'h3c0e3ca6),
	.w5(32'h3c06891f),
	.w6(32'h3b6c2b5b),
	.w7(32'h3c5e46ad),
	.w8(32'hbb186cbf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a5739),
	.w1(32'hbb563536),
	.w2(32'h3b2b1b86),
	.w3(32'h39575a45),
	.w4(32'h3a4121ed),
	.w5(32'h3c6852ea),
	.w6(32'hbbceb51e),
	.w7(32'hbc5356cb),
	.w8(32'hbb86e016),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed4978),
	.w1(32'h3b62daae),
	.w2(32'h3b2d7997),
	.w3(32'h3a9190cc),
	.w4(32'h3bc01ba3),
	.w5(32'h3c21a803),
	.w6(32'h3b396968),
	.w7(32'h3c0fa40c),
	.w8(32'hbb84e10d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c1506),
	.w1(32'h3b4f45d5),
	.w2(32'h3be972ef),
	.w3(32'h3aeecc1c),
	.w4(32'hbaaa6975),
	.w5(32'h3bbe9b1c),
	.w6(32'h3b68624d),
	.w7(32'h3b913cf8),
	.w8(32'h3b1f39c7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2dd48),
	.w1(32'hbc282155),
	.w2(32'hba8df3c4),
	.w3(32'h3b9ca514),
	.w4(32'h3a8803e9),
	.w5(32'h3b92926d),
	.w6(32'hba643e71),
	.w7(32'hbbf5f382),
	.w8(32'hbaaffa50),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be921cc),
	.w1(32'hbb9a7828),
	.w2(32'hbae30cad),
	.w3(32'hbb838e04),
	.w4(32'h3bbf5591),
	.w5(32'h3a370bca),
	.w6(32'hbb016d60),
	.w7(32'hbadb2c7b),
	.w8(32'h3c042fa7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7772c),
	.w1(32'h39e39b8e),
	.w2(32'hbba7560b),
	.w3(32'hbaac6954),
	.w4(32'hbb86da9d),
	.w5(32'h3b78ca82),
	.w6(32'h3bc419dd),
	.w7(32'hbbe06072),
	.w8(32'hbb77e3f6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5cf9f),
	.w1(32'h3baaf0fd),
	.w2(32'h3bf3129f),
	.w3(32'h3b03ee7e),
	.w4(32'h3bf193ec),
	.w5(32'hbb2ff418),
	.w6(32'hbbac72fa),
	.w7(32'h3b098dd6),
	.w8(32'h3c1e0a96),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07401d),
	.w1(32'hb87816b2),
	.w2(32'h3b514af6),
	.w3(32'hbc1952bf),
	.w4(32'hbb591288),
	.w5(32'hbb5d31a3),
	.w6(32'h3abe0b12),
	.w7(32'h3b47f41d),
	.w8(32'h39de3ebc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2385cb),
	.w1(32'h3c288ad5),
	.w2(32'h3c592982),
	.w3(32'hbb672622),
	.w4(32'h3c126770),
	.w5(32'hba931017),
	.w6(32'hbadebd94),
	.w7(32'h3c2295dd),
	.w8(32'h3bd35410),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb744f74),
	.w1(32'hbb665567),
	.w2(32'hbc10cb98),
	.w3(32'hbc1d42a5),
	.w4(32'hbbfac5d0),
	.w5(32'hbbdf00c0),
	.w6(32'hbba300fe),
	.w7(32'hbbc2f3c6),
	.w8(32'hbc1a1497),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53ec3),
	.w1(32'hbbf27f92),
	.w2(32'hbc1a384e),
	.w3(32'hbae53c75),
	.w4(32'hbbef3bb1),
	.w5(32'h3b9b01bb),
	.w6(32'h3aae9183),
	.w7(32'hbb3b6179),
	.w8(32'hbb84ca3a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8a317),
	.w1(32'hbba98a67),
	.w2(32'hbc187fd0),
	.w3(32'h3b4e0141),
	.w4(32'hbbc36b9c),
	.w5(32'hbb98502a),
	.w6(32'hbc17194d),
	.w7(32'hbc3aa5b5),
	.w8(32'hbbaf6344),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdd7e2),
	.w1(32'h3af9087a),
	.w2(32'h3aacdcba),
	.w3(32'hbbdba2e1),
	.w4(32'hba698334),
	.w5(32'hbac77a68),
	.w6(32'hba49b7fb),
	.w7(32'h3aa6e9da),
	.w8(32'h3a4e7ee1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaf569),
	.w1(32'hbae97a57),
	.w2(32'hbb83a3c1),
	.w3(32'hbb1914be),
	.w4(32'h3a8f96e9),
	.w5(32'hba246a1d),
	.w6(32'h3ac248ad),
	.w7(32'hba29edcc),
	.w8(32'h3b993ebc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a515fd7),
	.w1(32'hb9cb2738),
	.w2(32'hba3085c8),
	.w3(32'h3b8aba08),
	.w4(32'hb9d873d7),
	.w5(32'hbadbc993),
	.w6(32'hba243fa4),
	.w7(32'hbaff430b),
	.w8(32'h3ab20932),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3ca2e),
	.w1(32'h3a08cf89),
	.w2(32'hbaf77bad),
	.w3(32'h38f35c16),
	.w4(32'hbacf888a),
	.w5(32'hba909440),
	.w6(32'h3ab831f6),
	.w7(32'h3a37a11b),
	.w8(32'hb985f542),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c48b4),
	.w1(32'h3b446464),
	.w2(32'hbb0c9b78),
	.w3(32'h3b46e609),
	.w4(32'hbac23128),
	.w5(32'h3b9b68a8),
	.w6(32'hbaf1372e),
	.w7(32'hbb23e678),
	.w8(32'hbaa4a83f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5fc05),
	.w1(32'h3b0542a1),
	.w2(32'h3b9e96b7),
	.w3(32'h3be31d4e),
	.w4(32'h3a662646),
	.w5(32'hb9b3a094),
	.w6(32'hbb0db6a4),
	.w7(32'hbb9f7500),
	.w8(32'h39ace27a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485699),
	.w1(32'h3b2b372c),
	.w2(32'h3a05df58),
	.w3(32'hbb6385b1),
	.w4(32'h3ab3240a),
	.w5(32'hbab50020),
	.w6(32'h3aec60d7),
	.w7(32'hb9a26f82),
	.w8(32'h3af70049),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277c1f),
	.w1(32'hbc0a430b),
	.w2(32'hbbc607a2),
	.w3(32'hba5f277c),
	.w4(32'hbab8c25b),
	.w5(32'h3b738386),
	.w6(32'hbbc79539),
	.w7(32'hbc5a4ac0),
	.w8(32'hbb9d5838),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e8c2ff),
	.w1(32'hba3ae81d),
	.w2(32'hb96d663f),
	.w3(32'hba875f41),
	.w4(32'hb84ecbe7),
	.w5(32'hbb1a0608),
	.w6(32'hbb7b7bcc),
	.w7(32'hbb285f05),
	.w8(32'h3aadaaa0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af28e2a),
	.w1(32'h3b197f1e),
	.w2(32'hbbc2ad6b),
	.w3(32'hba8d643c),
	.w4(32'hbab4be3e),
	.w5(32'hbb891760),
	.w6(32'h3ba0fd83),
	.w7(32'hb962e21f),
	.w8(32'h3ab9fb99),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3bb71),
	.w1(32'h38b975bd),
	.w2(32'hbb88f2d5),
	.w3(32'h3c4da9d6),
	.w4(32'hb82cb576),
	.w5(32'hbb3ba216),
	.w6(32'hbb75ff06),
	.w7(32'hbbe4fe9c),
	.w8(32'hbc0a6c6c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb38bc),
	.w1(32'hba98c673),
	.w2(32'h3b349553),
	.w3(32'hbba648d4),
	.w4(32'h3aeae1a9),
	.w5(32'h3bb23c34),
	.w6(32'hbab14725),
	.w7(32'hba96d05d),
	.w8(32'h3b22baaf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1aa8),
	.w1(32'h3b165f65),
	.w2(32'h3b9c108d),
	.w3(32'h3b60b9d2),
	.w4(32'hbad2a13d),
	.w5(32'h3a733e2f),
	.w6(32'h3b2e7d18),
	.w7(32'h3b837ea5),
	.w8(32'hba00df99),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec8e90),
	.w1(32'h3b3c181e),
	.w2(32'h3b7db947),
	.w3(32'h3996cccc),
	.w4(32'hbb56f208),
	.w5(32'h3b86ed1d),
	.w6(32'hbbc8a196),
	.w7(32'h3b047d57),
	.w8(32'h3bb1609b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1844c9),
	.w1(32'h3ba6142b),
	.w2(32'h3ba3a97f),
	.w3(32'h3a9fbeac),
	.w4(32'hbbe9fc8d),
	.w5(32'h3b7237fd),
	.w6(32'h3b8ce1fc),
	.w7(32'h3c0a9045),
	.w8(32'h3b24b221),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117e75),
	.w1(32'h3aea88e6),
	.w2(32'hbb657d8f),
	.w3(32'h3ae3efc6),
	.w4(32'hbb6323c4),
	.w5(32'hbbf47a17),
	.w6(32'h3c19b640),
	.w7(32'h3aafacc5),
	.w8(32'h3a11cef0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba173dd8),
	.w1(32'h3acd9cdc),
	.w2(32'h3b3ea56c),
	.w3(32'hba980e95),
	.w4(32'h3a289fd7),
	.w5(32'hba99292b),
	.w6(32'hb93cc78d),
	.w7(32'hbb791b19),
	.w8(32'h3b1d206d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b759f17),
	.w1(32'h3b8a36dd),
	.w2(32'h3bd350e0),
	.w3(32'hb926e9dc),
	.w4(32'h3b865df5),
	.w5(32'h3b3fbcb4),
	.w6(32'h371dfca6),
	.w7(32'hb9057ffb),
	.w8(32'h3bd5e640),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa1ec),
	.w1(32'h3a461c26),
	.w2(32'h39ac0dc2),
	.w3(32'h393088eb),
	.w4(32'hbaad720d),
	.w5(32'h3a219aef),
	.w6(32'hba4aa088),
	.w7(32'hba4c301b),
	.w8(32'hb8c8c506),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2d818),
	.w1(32'hbc144662),
	.w2(32'hba07bf59),
	.w3(32'hbaaf59d2),
	.w4(32'hbb552021),
	.w5(32'h3c2e2d20),
	.w6(32'h3aaf970d),
	.w7(32'h391ff8cb),
	.w8(32'h3a70cb21),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac29c55),
	.w1(32'hbbea84b4),
	.w2(32'hbbd32e05),
	.w3(32'hba97f2ea),
	.w4(32'hbbf330ea),
	.w5(32'h38b8c6db),
	.w6(32'hba479eee),
	.w7(32'hbb891848),
	.w8(32'hbaabed62),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762744),
	.w1(32'h3bddef80),
	.w2(32'hbaa9ef0e),
	.w3(32'h3c460d14),
	.w4(32'h3aff5b8f),
	.w5(32'h3b7aa214),
	.w6(32'hba8b9d46),
	.w7(32'h3b1cc714),
	.w8(32'h3b3bba45),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63ff2f),
	.w1(32'hba6e2865),
	.w2(32'h3b6a2fb3),
	.w3(32'h3ba95377),
	.w4(32'h3b867943),
	.w5(32'h39bed1db),
	.w6(32'h3ba7a19c),
	.w7(32'h3ace1982),
	.w8(32'h3abf959d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62dd67),
	.w1(32'h3b93447b),
	.w2(32'h3aba1b85),
	.w3(32'h3ad884de),
	.w4(32'h3b4db274),
	.w5(32'hbbc16ff3),
	.w6(32'h3b28e5f9),
	.w7(32'h3b50625d),
	.w8(32'h3bb9f2f2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b8fd2),
	.w1(32'hbb561852),
	.w2(32'hbb2723ce),
	.w3(32'hbaf63744),
	.w4(32'hbafcd668),
	.w5(32'hbb56c99b),
	.w6(32'hbb3801bf),
	.w7(32'hbb726dce),
	.w8(32'hbb40c3ab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb869545),
	.w1(32'h3b620494),
	.w2(32'h3c488c9e),
	.w3(32'hbb850d01),
	.w4(32'h3c2df6df),
	.w5(32'h3bdebe52),
	.w6(32'hbb7584f3),
	.w7(32'h3b0aa4fb),
	.w8(32'hbaf5a290),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08ecf),
	.w1(32'h3b16e0b7),
	.w2(32'h3aa2cd29),
	.w3(32'hbbaec874),
	.w4(32'hb7475b06),
	.w5(32'h3bee247d),
	.w6(32'h3bf34684),
	.w7(32'h3ba6452a),
	.w8(32'h3beff0c2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41c38),
	.w1(32'hbbc800f9),
	.w2(32'hbbeb1759),
	.w3(32'h3b5c512f),
	.w4(32'hbc1c3092),
	.w5(32'hbb4f3cb9),
	.w6(32'h39b2e45e),
	.w7(32'hbbd91044),
	.w8(32'hbbf7d207),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5c3c),
	.w1(32'hbc1622f0),
	.w2(32'hbb8cceaf),
	.w3(32'h3ba7eed6),
	.w4(32'hba8deede),
	.w5(32'hbb9afe3d),
	.w6(32'hbc076100),
	.w7(32'hbc2b7dd4),
	.w8(32'hbb9a72d2),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e2397),
	.w1(32'hbba6afd9),
	.w2(32'hbbd86168),
	.w3(32'hbbee31d9),
	.w4(32'hbb2e8221),
	.w5(32'hbb911efc),
	.w6(32'hbace3a32),
	.w7(32'hbb842373),
	.w8(32'hbb5c6c4d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9a09),
	.w1(32'hbb7b6448),
	.w2(32'h3b2fcf8f),
	.w3(32'hbb8c988f),
	.w4(32'h3abad83b),
	.w5(32'h3bacc185),
	.w6(32'hbb8cac8d),
	.w7(32'hbb0f629e),
	.w8(32'h3add8a48),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dbc7a),
	.w1(32'hbb771e29),
	.w2(32'h3ac37bdf),
	.w3(32'h3aebf5ef),
	.w4(32'hb93e6236),
	.w5(32'h3b579167),
	.w6(32'hbb022e94),
	.w7(32'h3a80505d),
	.w8(32'hbb5835f4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7814),
	.w1(32'h3c2bd6de),
	.w2(32'hba7cf811),
	.w3(32'hbb6d255f),
	.w4(32'h3a08466f),
	.w5(32'hbb200044),
	.w6(32'hba1bad65),
	.w7(32'h3c10398f),
	.w8(32'hbb40c4c4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fda40),
	.w1(32'h3bc1a3f9),
	.w2(32'hba1706ad),
	.w3(32'hb9575fe3),
	.w4(32'hbba0730c),
	.w5(32'h3ab2d4d4),
	.w6(32'h3bbf0b04),
	.w7(32'hbb498a07),
	.w8(32'hbc043633),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba361cd),
	.w1(32'hb89fa65c),
	.w2(32'hbb18791c),
	.w3(32'hbb71d095),
	.w4(32'hba15f27f),
	.w5(32'h39c40e7a),
	.w6(32'h3b753139),
	.w7(32'hbbfa3af4),
	.w8(32'hbc0d0179),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f4963),
	.w1(32'h3c3894d3),
	.w2(32'h3c0d7d96),
	.w3(32'hbaab76f8),
	.w4(32'h3b1fcecb),
	.w5(32'hbb6a900d),
	.w6(32'hbb4ce89e),
	.w7(32'h3c82b6cc),
	.w8(32'h3bf3db3f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b7545),
	.w1(32'hbc2d7cab),
	.w2(32'hbc23f555),
	.w3(32'hba4012df),
	.w4(32'hbc14f9da),
	.w5(32'hbb7aa184),
	.w6(32'hbc08ba93),
	.w7(32'hbc163cc6),
	.w8(32'hbc3b0790),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda0da0),
	.w1(32'hb9a93f1a),
	.w2(32'hbc2d1919),
	.w3(32'hbb2ed522),
	.w4(32'h3aa0ca2d),
	.w5(32'hbb251aaa),
	.w6(32'h3adc1e2b),
	.w7(32'hbba8d621),
	.w8(32'h3aec24e8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f826),
	.w1(32'hba8fed4a),
	.w2(32'hbc0c066d),
	.w3(32'h3bab1b79),
	.w4(32'hba9dc170),
	.w5(32'h3b3b8b46),
	.w6(32'hbab9139f),
	.w7(32'hbbbc5a85),
	.w8(32'hb7098994),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4be40e),
	.w1(32'h3bb78339),
	.w2(32'h3b926424),
	.w3(32'h3be5b01c),
	.w4(32'hbb8d0f34),
	.w5(32'hbc427f66),
	.w6(32'hbb7240db),
	.w7(32'h3b0dc0a1),
	.w8(32'hba9861b9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd6617),
	.w1(32'h3b3f4387),
	.w2(32'h3bc31da7),
	.w3(32'hbbf8d4d2),
	.w4(32'h3b673792),
	.w5(32'h3bcf385d),
	.w6(32'hb93d200b),
	.w7(32'h3b2aa28d),
	.w8(32'h3b7a1c98),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370547),
	.w1(32'hbbf7dc7b),
	.w2(32'hb9b7eac6),
	.w3(32'h3bc72e10),
	.w4(32'hbc20add3),
	.w5(32'hba58df70),
	.w6(32'hba27bc99),
	.w7(32'hbb4adae2),
	.w8(32'hbbb7b8bf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35689f),
	.w1(32'h3bcc146f),
	.w2(32'h3bc6e7fc),
	.w3(32'hbb184f45),
	.w4(32'h3b9e2071),
	.w5(32'hbb57e5ba),
	.w6(32'h390e9e6d),
	.w7(32'h3b49ae9b),
	.w8(32'h3bc10004),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70c664),
	.w1(32'h3bdef301),
	.w2(32'h3b3978ee),
	.w3(32'hbbec657b),
	.w4(32'h3bbccf77),
	.w5(32'hbabdd900),
	.w6(32'h3ab7ab5d),
	.w7(32'h38b1f391),
	.w8(32'h3bab0358),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd452),
	.w1(32'hbb7e8e02),
	.w2(32'hbbd97e44),
	.w3(32'hb95bda85),
	.w4(32'hbc00c08a),
	.w5(32'hbb2e9ba0),
	.w6(32'hbbbb019f),
	.w7(32'hbc0c5f2b),
	.w8(32'hbac1f7e0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa00ffe),
	.w1(32'hba18399e),
	.w2(32'h3a20fbf4),
	.w3(32'h3b2377f7),
	.w4(32'hbbf016e5),
	.w5(32'h3a2f4ff4),
	.w6(32'h3addbdc1),
	.w7(32'hbb865dc6),
	.w8(32'hb980394d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12fc98),
	.w1(32'h3a9f7127),
	.w2(32'hbc14bdd4),
	.w3(32'h3b2c1e72),
	.w4(32'hbbaf7f25),
	.w5(32'hbc234778),
	.w6(32'hbad0537d),
	.w7(32'hbb6a9d2a),
	.w8(32'hbb87f7ab),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931f1f),
	.w1(32'hbb189ec4),
	.w2(32'hbbe2c1a8),
	.w3(32'hb9881865),
	.w4(32'h3b0a873f),
	.w5(32'h3b1b9493),
	.w6(32'hbbe937c2),
	.w7(32'hbbb95873),
	.w8(32'hbb9e172e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3952d9),
	.w1(32'hba60891f),
	.w2(32'hbc16aeaa),
	.w3(32'hbb82cf4e),
	.w4(32'hbc0e69e2),
	.w5(32'hbbe3c017),
	.w6(32'h3ba82274),
	.w7(32'hbc0e883b),
	.w8(32'hbb446f9d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2265b),
	.w1(32'hba7f0dd4),
	.w2(32'hbba65267),
	.w3(32'h3abf7ba7),
	.w4(32'hbac92072),
	.w5(32'h3bc1cc2a),
	.w6(32'hbbbb200e),
	.w7(32'hbb2d3bf5),
	.w8(32'hbbd6e85e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a541b),
	.w1(32'h3ba34c41),
	.w2(32'hbb743845),
	.w3(32'h3bcdc742),
	.w4(32'hbb90dcff),
	.w5(32'hbbc1e039),
	.w6(32'h3b157db2),
	.w7(32'hbb57bbb8),
	.w8(32'hbb660b93),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2fc5a),
	.w1(32'h3b199cdf),
	.w2(32'h3b02a70c),
	.w3(32'h3bd47835),
	.w4(32'h3c26868c),
	.w5(32'hbabcc5c6),
	.w6(32'hbc1ef544),
	.w7(32'h3b0e606f),
	.w8(32'h3c1ba7bb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818c50),
	.w1(32'h3b37508b),
	.w2(32'h3b417cf2),
	.w3(32'hbc0c6420),
	.w4(32'h3afbbcaf),
	.w5(32'h3aad285e),
	.w6(32'hba7c8489),
	.w7(32'h3b929b92),
	.w8(32'h3b1d6379),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a171766),
	.w1(32'hbc456314),
	.w2(32'hbbacc59e),
	.w3(32'hbb4a2192),
	.w4(32'hbc0528fc),
	.w5(32'h3b05be48),
	.w6(32'hbb2f2743),
	.w7(32'hbc20d7b5),
	.w8(32'hbbeb8242),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b495dcd),
	.w1(32'h3bd0f017),
	.w2(32'h3b8b02d4),
	.w3(32'h3bd03357),
	.w4(32'h3ba06aea),
	.w5(32'h3ab4a490),
	.w6(32'hbabb1737),
	.w7(32'h3ba6a454),
	.w8(32'h3ba473ce),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84daf1),
	.w1(32'h3a2a9994),
	.w2(32'h3bb8ec65),
	.w3(32'hba7782f6),
	.w4(32'hbb420b28),
	.w5(32'hbba03113),
	.w6(32'hbbb0d86a),
	.w7(32'hb87fa6e7),
	.w8(32'h3a69b2d5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6b8a3),
	.w1(32'h39b8ca51),
	.w2(32'hbc0c8655),
	.w3(32'hbc08864a),
	.w4(32'h3a3a2854),
	.w5(32'hba46ee77),
	.w6(32'hbaf0fa47),
	.w7(32'hbb144c57),
	.w8(32'hb92eac95),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9013),
	.w1(32'hbb05efe8),
	.w2(32'hbbc98dca),
	.w3(32'h3b589f33),
	.w4(32'hbb4aeb07),
	.w5(32'hbb23c19a),
	.w6(32'hbb386d44),
	.w7(32'hba63cb58),
	.w8(32'hbc096b64),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04c430),
	.w1(32'hbb1f4d2c),
	.w2(32'hbbaeabc7),
	.w3(32'hbbea8623),
	.w4(32'hbaecd45b),
	.w5(32'hbbc6a057),
	.w6(32'hbabf8e26),
	.w7(32'hbb3535c3),
	.w8(32'hbba8310e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb921555),
	.w1(32'h3b615637),
	.w2(32'h3aabefa7),
	.w3(32'hbbbef9ff),
	.w4(32'h3ac73022),
	.w5(32'h39da28b7),
	.w6(32'h3af44081),
	.w7(32'hba703e1b),
	.w8(32'hbaca9ae6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d323cb),
	.w1(32'h3badaf26),
	.w2(32'h3c3b063b),
	.w3(32'hb9aa1216),
	.w4(32'h3b4b3213),
	.w5(32'hbc0bcda1),
	.w6(32'hba429a59),
	.w7(32'h3c71b4de),
	.w8(32'h3c0d1925),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6659e2),
	.w1(32'h3b61d8d5),
	.w2(32'hbad432eb),
	.w3(32'hbbc6aba4),
	.w4(32'h38b1cb60),
	.w5(32'hbbd5b15b),
	.w6(32'h3993f5ef),
	.w7(32'h39c150ed),
	.w8(32'h3a2c66c0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f72e1),
	.w1(32'h3b94d3f9),
	.w2(32'h3c13b1ba),
	.w3(32'hbbb543b4),
	.w4(32'h3b11e39a),
	.w5(32'h3b8422f4),
	.w6(32'h3aa69c01),
	.w7(32'h3b2c4ecb),
	.w8(32'h3bb563b8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b318b2c),
	.w1(32'hbbe20752),
	.w2(32'hbadc2afb),
	.w3(32'hbbded777),
	.w4(32'hbafd9f26),
	.w5(32'h3a3065be),
	.w6(32'h3ad2f3e0),
	.w7(32'h3a8a4f7f),
	.w8(32'hbb9b8e47),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4b119),
	.w1(32'hbc1048a9),
	.w2(32'hbba414c7),
	.w3(32'h3b8ed1fe),
	.w4(32'hbc2663f8),
	.w5(32'hbbaf508b),
	.w6(32'hbb9dae22),
	.w7(32'hbbc8a2b1),
	.w8(32'h39bdb857),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d48d),
	.w1(32'hbc0e776a),
	.w2(32'hbbfd581e),
	.w3(32'h3b88ad8f),
	.w4(32'hbbb782b4),
	.w5(32'h3c47531d),
	.w6(32'hbbce117a),
	.w7(32'hbbb032f8),
	.w8(32'hbb0ae88e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eca38),
	.w1(32'hbb8bb29f),
	.w2(32'hbc161de5),
	.w3(32'h3c00f5c0),
	.w4(32'hbba36a9f),
	.w5(32'hbbec2a95),
	.w6(32'h3bc2779c),
	.w7(32'hba95ab67),
	.w8(32'hbb51f78f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74f9bb),
	.w1(32'hbbac8b9e),
	.w2(32'h39020d49),
	.w3(32'hbbd5c9c6),
	.w4(32'h3bbe90c0),
	.w5(32'hbb769f6a),
	.w6(32'hbaa97b8b),
	.w7(32'hbbbae508),
	.w8(32'h3b8549e9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e3f7),
	.w1(32'h3b950043),
	.w2(32'h3adb34e8),
	.w3(32'hbb7b2405),
	.w4(32'h3b8e9220),
	.w5(32'h3b9a16d7),
	.w6(32'h3bd5a387),
	.w7(32'hb9d71f98),
	.w8(32'hbb4326e5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0cac),
	.w1(32'hbb3e933e),
	.w2(32'hbb133f8b),
	.w3(32'h3ae5a7d6),
	.w4(32'hbb1870bb),
	.w5(32'hbb703482),
	.w6(32'h3b936543),
	.w7(32'h3a30d061),
	.w8(32'hbb2ae9ce),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e4ca8),
	.w1(32'hbb9b5bcf),
	.w2(32'hbbe5a361),
	.w3(32'hbbd9e08d),
	.w4(32'hbb7a2552),
	.w5(32'h3b53fd3c),
	.w6(32'hbac4c8e1),
	.w7(32'hbc175f38),
	.w8(32'hbaeb4e49),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc376),
	.w1(32'hbb882bf7),
	.w2(32'h3a7c710f),
	.w3(32'hbaabd009),
	.w4(32'hbb3b49e5),
	.w5(32'h3b21edbd),
	.w6(32'hbbf7afe6),
	.w7(32'hbbe165d2),
	.w8(32'hb7e4364d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c3235),
	.w1(32'h3c352931),
	.w2(32'h3c6a6f9f),
	.w3(32'h39e6f8ba),
	.w4(32'h3baf56b7),
	.w5(32'hbaab1e5d),
	.w6(32'hbbbf632e),
	.w7(32'h3c42f1ae),
	.w8(32'h3bdefa90),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcc8d8),
	.w1(32'hbbf44938),
	.w2(32'hbbfed3d6),
	.w3(32'hbb5c4afe),
	.w4(32'hbc1cb584),
	.w5(32'hbc1c07b5),
	.w6(32'hbbb1152a),
	.w7(32'hbc140a3e),
	.w8(32'hbb3e531f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39735d9d),
	.w1(32'hb9a210b3),
	.w2(32'hba2639f3),
	.w3(32'h3b519fd7),
	.w4(32'h3b01cd27),
	.w5(32'h3bb19f63),
	.w6(32'h37393bb4),
	.w7(32'hbb9087b1),
	.w8(32'h3931ce73),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc13888),
	.w1(32'h3a59f39f),
	.w2(32'hbac5f085),
	.w3(32'h3b7d4e7a),
	.w4(32'h3a409796),
	.w5(32'hb8903d53),
	.w6(32'h39da8df0),
	.w7(32'hbb4d19f2),
	.w8(32'hbb1570ed),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a32e),
	.w1(32'h3b56f697),
	.w2(32'hbb1b9be6),
	.w3(32'hba576abe),
	.w4(32'h3b23f7b1),
	.w5(32'h3b194cda),
	.w6(32'h3b0f6824),
	.w7(32'hbaa29818),
	.w8(32'h3a73e141),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae79d14),
	.w1(32'hbb93c918),
	.w2(32'hbacdf0f3),
	.w3(32'h3b3b5fca),
	.w4(32'hbb3d107b),
	.w5(32'hba5ced50),
	.w6(32'hbb6ad0fb),
	.w7(32'hbb683cde),
	.w8(32'hbb4c1b05),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1481d4),
	.w1(32'hbb43ddf8),
	.w2(32'hbb01a933),
	.w3(32'hbb5e2ac8),
	.w4(32'h39405ac6),
	.w5(32'hba949405),
	.w6(32'hbba4580a),
	.w7(32'hbbafa9dd),
	.w8(32'hbb5e2774),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe38463),
	.w1(32'hbbf4f968),
	.w2(32'hbb4b2d19),
	.w3(32'hbbc50e46),
	.w4(32'hbbad9b83),
	.w5(32'h3b8cb73b),
	.w6(32'hbb6b7b48),
	.w7(32'hbbc8c62e),
	.w8(32'hbb9d4918),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4da5be),
	.w1(32'hba003f7b),
	.w2(32'hbad7ed77),
	.w3(32'h3aa62547),
	.w4(32'hb9579481),
	.w5(32'h38ae096b),
	.w6(32'hbb00dcac),
	.w7(32'h39368cef),
	.w8(32'h3b23128c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb216911),
	.w1(32'h38abbc2b),
	.w2(32'h3aa5dd24),
	.w3(32'hba5e5dec),
	.w4(32'h3b00566c),
	.w5(32'h3b3e1494),
	.w6(32'hb99ec755),
	.w7(32'hba961d0f),
	.w8(32'h3a0cfe3f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbaba3),
	.w1(32'hba7a7077),
	.w2(32'h39e7c8e5),
	.w3(32'h3a55c0f1),
	.w4(32'hbb4c4631),
	.w5(32'hb9cd7d4d),
	.w6(32'h3afb98e8),
	.w7(32'hba985194),
	.w8(32'h39d086a5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e64b),
	.w1(32'hbba272c8),
	.w2(32'hbbbe3e85),
	.w3(32'h3acfa6cf),
	.w4(32'hbb17d84d),
	.w5(32'hbb99482b),
	.w6(32'hba1d7ec3),
	.w7(32'hbbd00f08),
	.w8(32'hbba4b669),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e5f0),
	.w1(32'hbb0f51e3),
	.w2(32'hba5c6e3a),
	.w3(32'hbb902a07),
	.w4(32'h3bcd8d8d),
	.w5(32'h3be9de62),
	.w6(32'hbaa4bd66),
	.w7(32'hbbbcb4f3),
	.w8(32'hbb443994),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a456),
	.w1(32'h3af65dc5),
	.w2(32'h389e9b28),
	.w3(32'h3bb7c140),
	.w4(32'h399e1aa8),
	.w5(32'hba399e14),
	.w6(32'h3b2f6c48),
	.w7(32'h3ad4ca8b),
	.w8(32'h3b00bedf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ba570),
	.w1(32'hbb37f321),
	.w2(32'hbac1327b),
	.w3(32'hb814d03d),
	.w4(32'hbb7c5f5b),
	.w5(32'hbb1043a6),
	.w6(32'h3af644ff),
	.w7(32'hbbc11ea9),
	.w8(32'hbba01ba4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6b77),
	.w1(32'hba9ea7ea),
	.w2(32'hbb34cb6c),
	.w3(32'hbb70e396),
	.w4(32'hbbd084a3),
	.w5(32'h3b641ca9),
	.w6(32'hba3d316a),
	.w7(32'hbb1c9ab5),
	.w8(32'hba95a9f0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1af8a),
	.w1(32'hbb191844),
	.w2(32'hbbdf3370),
	.w3(32'h3c13a016),
	.w4(32'hbaea786b),
	.w5(32'hbba13109),
	.w6(32'h39ebd77e),
	.w7(32'hbb537d7a),
	.w8(32'hbb8868bc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef11a6),
	.w1(32'hbb62b2aa),
	.w2(32'hbb8de5bb),
	.w3(32'hbba558a8),
	.w4(32'h3a61a39d),
	.w5(32'h3b37b8cd),
	.w6(32'hba4e1529),
	.w7(32'hbba18b78),
	.w8(32'hbb5911b5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29367b),
	.w1(32'hb98fe666),
	.w2(32'hbbc1b67b),
	.w3(32'hbb0895be),
	.w4(32'hbb9528f9),
	.w5(32'h3bae44b3),
	.w6(32'h3ae0cdaa),
	.w7(32'hbb96f594),
	.w8(32'hbb4aa5c9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ee2e9),
	.w1(32'hbb68e1de),
	.w2(32'h3b85ecdd),
	.w3(32'h3c51bc80),
	.w4(32'hbb6de8e5),
	.w5(32'hbb941fe1),
	.w6(32'hbbddf2d2),
	.w7(32'h3b5755d9),
	.w8(32'h3a3d6156),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81a924),
	.w1(32'hbc15cbf7),
	.w2(32'hbcc1ffbe),
	.w3(32'hbb65c40f),
	.w4(32'hbc147423),
	.w5(32'hbc863512),
	.w6(32'hbb7c9302),
	.w7(32'hbbf09714),
	.w8(32'h3a18cdc6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f7af),
	.w1(32'hbb482a76),
	.w2(32'hbbee723c),
	.w3(32'hbb5c7308),
	.w4(32'hbb6fe2df),
	.w5(32'hbc4a13a2),
	.w6(32'h3ba3d96d),
	.w7(32'hbbf6aacd),
	.w8(32'hbb1ff35b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule