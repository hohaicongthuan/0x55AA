module layer_6_featuremap_38(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eba95),
	.w1(32'hbc1b6b49),
	.w2(32'h398eabe4),
	.w3(32'hba892e09),
	.w4(32'hbbb00b0a),
	.w5(32'hbc093d13),
	.w6(32'hbc0a3afb),
	.w7(32'hbb872f4a),
	.w8(32'hba74038f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85378a),
	.w1(32'hbc091e10),
	.w2(32'hba6bf7ad),
	.w3(32'hbc57d47e),
	.w4(32'hbc3e325d),
	.w5(32'hbbd5e4a2),
	.w6(32'hbc86dd8b),
	.w7(32'hbc242364),
	.w8(32'hbc18abe3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca0aa7),
	.w1(32'h3b39ba79),
	.w2(32'hbcb5c4ff),
	.w3(32'h3c87ee5a),
	.w4(32'h3bdd8e76),
	.w5(32'hbbf464cd),
	.w6(32'h3c695ea5),
	.w7(32'h3aecebac),
	.w8(32'hbc209bad),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bb37f),
	.w1(32'hbb5d6db4),
	.w2(32'hbb80c232),
	.w3(32'hbbce6e41),
	.w4(32'hba513a5d),
	.w5(32'h3978bba7),
	.w6(32'hbb9f1277),
	.w7(32'hbad912c0),
	.w8(32'hbad03500),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993aac),
	.w1(32'h3c1c9ee9),
	.w2(32'h3cb69b16),
	.w3(32'hbac6e3fa),
	.w4(32'hbb8392ba),
	.w5(32'hbc0274e8),
	.w6(32'hbc37ddf1),
	.w7(32'h3a91600e),
	.w8(32'h3c1f1710),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f790a),
	.w1(32'hbaf71eaf),
	.w2(32'hbae5bca7),
	.w3(32'h3c20b72c),
	.w4(32'h3a81176e),
	.w5(32'hbb302873),
	.w6(32'h3a4675c1),
	.w7(32'hbacd22c0),
	.w8(32'hba833242),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147cf6),
	.w1(32'hba0cccff),
	.w2(32'h3b54a735),
	.w3(32'hb9069e2f),
	.w4(32'h3bc00a6c),
	.w5(32'h3c44914c),
	.w6(32'h36e3e935),
	.w7(32'hb6a6e327),
	.w8(32'h3a2229dc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85bf8b),
	.w1(32'h3c128cc0),
	.w2(32'hbc2e0920),
	.w3(32'h3c1227d2),
	.w4(32'h3c173213),
	.w5(32'h3bfea177),
	.w6(32'h3c25160e),
	.w7(32'h3c643269),
	.w8(32'h3bf7ca7a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad7682),
	.w1(32'h3b9b5286),
	.w2(32'h3ce10cca),
	.w3(32'hbbb090b4),
	.w4(32'h3c22ade2),
	.w5(32'h3c124db2),
	.w6(32'hbb190625),
	.w7(32'h3cc33730),
	.w8(32'h3c8823d2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22ea58),
	.w1(32'h3a9009ae),
	.w2(32'hbb107ab9),
	.w3(32'h3c16909d),
	.w4(32'h3bb52699),
	.w5(32'h3b4002e1),
	.w6(32'h3af2d56d),
	.w7(32'h3b01d7a5),
	.w8(32'hba5c568c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79b164),
	.w1(32'h3ca4f5ea),
	.w2(32'h39bb1603),
	.w3(32'h3bc03f09),
	.w4(32'h3cab234f),
	.w5(32'hbbaeac6a),
	.w6(32'h3c96a647),
	.w7(32'h3cd840f4),
	.w8(32'h3a96f9f5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bb52b),
	.w1(32'hbc508344),
	.w2(32'hbc88d2e0),
	.w3(32'hbbaf922d),
	.w4(32'h3ab6b26d),
	.w5(32'h3706c6f5),
	.w6(32'hbc41f722),
	.w7(32'hbc0c7b60),
	.w8(32'h3af91306),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0607c7),
	.w1(32'h3b6d26a5),
	.w2(32'h3b952bb8),
	.w3(32'hbb336077),
	.w4(32'hbb39c242),
	.w5(32'h39f55a94),
	.w6(32'hbbb2ce9f),
	.w7(32'hbb949bce),
	.w8(32'hbba044be),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1b4c5),
	.w1(32'hbc024874),
	.w2(32'h3ac7ab1e),
	.w3(32'hbb7e88f9),
	.w4(32'hbc0afded),
	.w5(32'hba7848b5),
	.w6(32'hbc5796c1),
	.w7(32'h3aa88690),
	.w8(32'h3c9d2ba9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c646fca),
	.w1(32'hbc4aaec7),
	.w2(32'h3bac028a),
	.w3(32'h39bfff25),
	.w4(32'h3b3a1da4),
	.w5(32'h3a0d2d08),
	.w6(32'hba208910),
	.w7(32'h3c8e0f6c),
	.w8(32'h3beff6c5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ed79d),
	.w1(32'hbb2385de),
	.w2(32'hbbea7f2c),
	.w3(32'h3853524f),
	.w4(32'hbb474cf6),
	.w5(32'hbba522d5),
	.w6(32'hb9c440ad),
	.w7(32'hbb3a68b1),
	.w8(32'hbbe1b07d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0e930),
	.w1(32'h3c62be45),
	.w2(32'h3c95ca50),
	.w3(32'hbc964c0d),
	.w4(32'hbc1fb5a9),
	.w5(32'hbcf38aba),
	.w6(32'h3cbb5149),
	.w7(32'h3c0adced),
	.w8(32'hbc3c4f55),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b52c),
	.w1(32'hbb01da07),
	.w2(32'hba2fa85e),
	.w3(32'h3aac2d6f),
	.w4(32'h3ad50770),
	.w5(32'h3a9dfdac),
	.w6(32'hbb445b82),
	.w7(32'hbb690de3),
	.w8(32'hbb8e4f55),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44caad),
	.w1(32'h3afec493),
	.w2(32'hbbaabe55),
	.w3(32'h3bd9e57b),
	.w4(32'h3bab1082),
	.w5(32'h3af173c0),
	.w6(32'h3b441177),
	.w7(32'hbab1a0dc),
	.w8(32'hbb77dc72),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb98f1),
	.w1(32'h3cd2e48d),
	.w2(32'h3b6c20f2),
	.w3(32'hbb677f25),
	.w4(32'hbcb83f2f),
	.w5(32'hbcb94955),
	.w6(32'h3bee0899),
	.w7(32'hbc1f062a),
	.w8(32'h39cc9ce0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8646d5),
	.w1(32'hbb72d671),
	.w2(32'hbb806d98),
	.w3(32'h38f243a1),
	.w4(32'hbb25aa4c),
	.w5(32'hb93090c8),
	.w6(32'hbaa8bc2f),
	.w7(32'hbb27ca62),
	.w8(32'hbb089489),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99650),
	.w1(32'hbb8168e2),
	.w2(32'hbc430510),
	.w3(32'hbbfa1fa0),
	.w4(32'hbb2bbba6),
	.w5(32'hbb8c47bb),
	.w6(32'hbbb98c9c),
	.w7(32'hba7b0a0f),
	.w8(32'h3a4751fe),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a9b26),
	.w1(32'h3cd7b22d),
	.w2(32'h3ca1a7a5),
	.w3(32'hbba04a16),
	.w4(32'hbcb78442),
	.w5(32'hbc9cb9cd),
	.w6(32'h3c3282dd),
	.w7(32'h3c472bd8),
	.w8(32'hbbe9eb8d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d7255),
	.w1(32'hbb80e89b),
	.w2(32'hba32e574),
	.w3(32'hbc0da6fa),
	.w4(32'hbc95d48c),
	.w5(32'hbc495cab),
	.w6(32'hbcc1f6f7),
	.w7(32'hbd42a75f),
	.w8(32'hbcc490eb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b381e),
	.w1(32'hbcd63d76),
	.w2(32'hbbb9076a),
	.w3(32'hbc113d41),
	.w4(32'h3a402a3f),
	.w5(32'h3cd73fd1),
	.w6(32'hbc8ac4fc),
	.w7(32'hbc73829a),
	.w8(32'h3cecaa31),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c003499),
	.w1(32'h3b04c057),
	.w2(32'hbc06a2e7),
	.w3(32'h3b81d973),
	.w4(32'hbca4fd72),
	.w5(32'hbcbe1423),
	.w6(32'h3b3c03ea),
	.w7(32'hbc8384f1),
	.w8(32'hbc630631),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca9f30),
	.w1(32'hbbb96d6c),
	.w2(32'hbb852b2a),
	.w3(32'h3c040de5),
	.w4(32'h3d00af9a),
	.w5(32'h3c8ab11a),
	.w6(32'h3c7372e1),
	.w7(32'h3cbdd541),
	.w8(32'h3ca2daae),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf0eb),
	.w1(32'hb8e18483),
	.w2(32'hbb1ce77f),
	.w3(32'h3b5975bb),
	.w4(32'h3b9866e7),
	.w5(32'h3bc085b0),
	.w6(32'h3a559cf1),
	.w7(32'hba0514de),
	.w8(32'h3a6fbf29),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab65abf),
	.w1(32'h3a077f08),
	.w2(32'hb9f25481),
	.w3(32'h3a9f543a),
	.w4(32'h3b53bf5a),
	.w5(32'h3b1b239b),
	.w6(32'h3b56706a),
	.w7(32'h3b45322e),
	.w8(32'h3a3059da),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5c12),
	.w1(32'hbbd9dfc5),
	.w2(32'h3c64ed94),
	.w3(32'hbce14a5e),
	.w4(32'hbccde915),
	.w5(32'h3a3ba2e2),
	.w6(32'hbcd50c09),
	.w7(32'hbc8b0642),
	.w8(32'hbb901ce6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b989a23),
	.w1(32'hbc36f1e1),
	.w2(32'hbceafa95),
	.w3(32'h3cad595a),
	.w4(32'h3c506921),
	.w5(32'h3ace73ad),
	.w6(32'h3c9dfbd8),
	.w7(32'h3c182e4c),
	.w8(32'hbb39487a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0234e2),
	.w1(32'hbc584fa5),
	.w2(32'h3b933f60),
	.w3(32'h3bcd8ff0),
	.w4(32'hbca560f8),
	.w5(32'hbc46cde1),
	.w6(32'hbcb64b7f),
	.w7(32'hbd03fcf5),
	.w8(32'hbc834dd3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2b0865),
	.w1(32'h3d148877),
	.w2(32'h3cb833f0),
	.w3(32'hbbc8474b),
	.w4(32'hbcc9b5df),
	.w5(32'hbd1a3a96),
	.w6(32'h3bbee2c9),
	.w7(32'hbad4c9b5),
	.w8(32'hbcac462e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82403c),
	.w1(32'h3c1ce860),
	.w2(32'h3bfc306d),
	.w3(32'hbc8e0aef),
	.w4(32'hbcae330f),
	.w5(32'hbc472376),
	.w6(32'hbbbc9d5d),
	.w7(32'hbc08e041),
	.w8(32'hb969250b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4285),
	.w1(32'hbb3ec816),
	.w2(32'hbad102b3),
	.w3(32'h3ab1d27d),
	.w4(32'hba0e50de),
	.w5(32'hbbb7c24b),
	.w6(32'h3b0519d1),
	.w7(32'h3bb1ea46),
	.w8(32'hbb7284ec),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40799f),
	.w1(32'hba909202),
	.w2(32'hbb16f48a),
	.w3(32'hb9feac09),
	.w4(32'hbbb84dd0),
	.w5(32'hbc539793),
	.w6(32'hbc6e22f9),
	.w7(32'hbc5408eb),
	.w8(32'hba616ad2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c362a),
	.w1(32'hbbede616),
	.w2(32'hb94c7f7f),
	.w3(32'h3a785d25),
	.w4(32'hbb76adfc),
	.w5(32'hbb8e85a2),
	.w6(32'hbb3bd5bd),
	.w7(32'hbb254470),
	.w8(32'hbb2b3041),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae38f19),
	.w1(32'hbb499987),
	.w2(32'hbb1ff023),
	.w3(32'hbb83306e),
	.w4(32'hbb19686f),
	.w5(32'hbb032938),
	.w6(32'hbb1613dc),
	.w7(32'hbb5002e3),
	.w8(32'hbaced050),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3c3c),
	.w1(32'hbc5d01bd),
	.w2(32'hbcc02d15),
	.w3(32'h3aa51aa2),
	.w4(32'h3cd74d3c),
	.w5(32'h3cb398c7),
	.w6(32'h3c7e7a09),
	.w7(32'h3d035167),
	.w8(32'h3c53192f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeef993),
	.w1(32'hbc271eaa),
	.w2(32'hbc73a44e),
	.w3(32'h3c527a3b),
	.w4(32'hbbe8bfdd),
	.w5(32'hba3f8635),
	.w6(32'hbba771b4),
	.w7(32'hbc61e4c8),
	.w8(32'h3c285d71),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb132d),
	.w1(32'h3c0e15d6),
	.w2(32'hbc2d6dbe),
	.w3(32'h3c84e679),
	.w4(32'h3c1ff211),
	.w5(32'h3aca7f5d),
	.w6(32'h3c1386bb),
	.w7(32'h3aaf38a0),
	.w8(32'hbc9249ec),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23da97),
	.w1(32'hbb651ec1),
	.w2(32'hbb8b4806),
	.w3(32'hbb98dc96),
	.w4(32'hbb0421e9),
	.w5(32'hbac98084),
	.w6(32'hbb55a314),
	.w7(32'hbb4c2bc2),
	.w8(32'hbb8a9305),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaacd5e),
	.w1(32'hbaeeb613),
	.w2(32'h3b130a8e),
	.w3(32'hbb5c74fc),
	.w4(32'hbc1e96cf),
	.w5(32'hbbd9cc44),
	.w6(32'h3b0cfdbe),
	.w7(32'h3bcb5513),
	.w8(32'h39cf6001),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90356e3),
	.w1(32'hbafe4c56),
	.w2(32'hbc12a6a0),
	.w3(32'h3bbfdac6),
	.w4(32'h3a930ef9),
	.w5(32'h3af76b11),
	.w6(32'h3b054d2a),
	.w7(32'hbb264c46),
	.w8(32'hbbed9c6c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba47202),
	.w1(32'hbbb74bfa),
	.w2(32'hbb95b2a4),
	.w3(32'hbb33df85),
	.w4(32'hbb5bed40),
	.w5(32'hbb34bedb),
	.w6(32'hbb678f9d),
	.w7(32'hb9d83e90),
	.w8(32'hba65a802),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7658d5),
	.w1(32'hbc9f1aaf),
	.w2(32'hbca9969d),
	.w3(32'h3ce80ba8),
	.w4(32'h3d045fc4),
	.w5(32'h3c21609f),
	.w6(32'h3ce4cff6),
	.w7(32'h3d0d69b6),
	.w8(32'h3c17b493),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc688272),
	.w1(32'h3ad994c1),
	.w2(32'hba892673),
	.w3(32'h3b622a77),
	.w4(32'hbb272357),
	.w5(32'h3b87186b),
	.w6(32'hbc260d3e),
	.w7(32'hbc87237e),
	.w8(32'hbc02f0b5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d2fbc),
	.w1(32'h3ce7b44d),
	.w2(32'h3c7b6959),
	.w3(32'hbca5fd92),
	.w4(32'hbd4ca74d),
	.w5(32'hbd3e4995),
	.w6(32'hbbf06b8c),
	.w7(32'h3b8705c5),
	.w8(32'h3b9532ce),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b808eb3),
	.w1(32'h3b185163),
	.w2(32'h3ba5df57),
	.w3(32'h3b6e315d),
	.w4(32'h3aa73273),
	.w5(32'h398ac3da),
	.w6(32'h3b380cdc),
	.w7(32'h3b149392),
	.w8(32'h3a216604),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445ddd),
	.w1(32'h3b2949db),
	.w2(32'hbb6492e0),
	.w3(32'hbb4de860),
	.w4(32'hbb321a83),
	.w5(32'h3bb16368),
	.w6(32'hbc89a654),
	.w7(32'hbcf52a8f),
	.w8(32'h3b091228),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c72a),
	.w1(32'hbb329409),
	.w2(32'hbb83e46e),
	.w3(32'hbba4fa98),
	.w4(32'hba784d72),
	.w5(32'h3a5195a6),
	.w6(32'hbbbe757c),
	.w7(32'hbb654c47),
	.w8(32'hbb3ca58d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77ff87),
	.w1(32'hbba0e81c),
	.w2(32'hbc0c4bc8),
	.w3(32'h3b3e4dba),
	.w4(32'hbbae474e),
	.w5(32'hbc0b3c35),
	.w6(32'hbae96154),
	.w7(32'hbc099846),
	.w8(32'hbc375ae7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e13a7),
	.w1(32'hbae7bb73),
	.w2(32'hbbed8956),
	.w3(32'hba429c6c),
	.w4(32'hbb2678d7),
	.w5(32'h3a647a8c),
	.w6(32'hbb27ea98),
	.w7(32'hbb919694),
	.w8(32'hbba2b687),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a00b),
	.w1(32'hbbf27eab),
	.w2(32'hbb8519dd),
	.w3(32'hbb6d4923),
	.w4(32'hbb85ad78),
	.w5(32'h3b86801c),
	.w6(32'hbbc2b8fe),
	.w7(32'hbb052092),
	.w8(32'h3ba2e5d8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0044e1),
	.w1(32'hbae0dec4),
	.w2(32'hbb339751),
	.w3(32'hbc2c5f71),
	.w4(32'hbc0caffe),
	.w5(32'hbbb55623),
	.w6(32'hbc465b2e),
	.w7(32'hbc0d51fb),
	.w8(32'hbc035366),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9e8f),
	.w1(32'hbc4023ac),
	.w2(32'hbc66a31e),
	.w3(32'hbbaf2f3b),
	.w4(32'hbc0ddbf0),
	.w5(32'hbbe10e98),
	.w6(32'hbc04bed9),
	.w7(32'hbc235d67),
	.w8(32'hbc044383),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e4bc8),
	.w1(32'h3934e44f),
	.w2(32'h3bc096ad),
	.w3(32'hbb3524bb),
	.w4(32'h3c07b4fb),
	.w5(32'h3b38c971),
	.w6(32'h3bd10952),
	.w7(32'h3c89a2bd),
	.w8(32'h3c044882),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc329),
	.w1(32'h3b1c30af),
	.w2(32'h3ae1a83c),
	.w3(32'hbbad85a2),
	.w4(32'hbb3ffd2f),
	.w5(32'hbb0226b7),
	.w6(32'hb9c3df51),
	.w7(32'hbab5660e),
	.w8(32'hbbcf4af3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8721a),
	.w1(32'h3c55add2),
	.w2(32'h3c95f9a3),
	.w3(32'h3bfcd6df),
	.w4(32'h3c5813ac),
	.w5(32'h3c72697b),
	.w6(32'h3c628864),
	.w7(32'h3c9558d0),
	.w8(32'h3c963cc8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a9b1c),
	.w1(32'h3b0fb906),
	.w2(32'h3c7fff1e),
	.w3(32'hbb019cdf),
	.w4(32'h3b52fb5c),
	.w5(32'h3c55c982),
	.w6(32'hbb9a15ec),
	.w7(32'h3bccb7c8),
	.w8(32'h3c6ba805),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c724378),
	.w1(32'h3c5e2e28),
	.w2(32'h3cb6988d),
	.w3(32'h3c09575b),
	.w4(32'h3c2a5b0b),
	.w5(32'h3c4f7c8b),
	.w6(32'h3c893a38),
	.w7(32'h3cab4cc7),
	.w8(32'h3c8fbb2b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89d21a),
	.w1(32'h3b4d59a9),
	.w2(32'hbb684fcd),
	.w3(32'h3bb3cf74),
	.w4(32'h3b3ef7ab),
	.w5(32'h3a4a1997),
	.w6(32'hbaf2cdef),
	.w7(32'hbbd97c3f),
	.w8(32'hbaef2e62),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba584487),
	.w1(32'hbb4aa003),
	.w2(32'hbb885dff),
	.w3(32'h3b877279),
	.w4(32'h3c801866),
	.w5(32'h3c397146),
	.w6(32'hb9ca702b),
	.w7(32'h3a949d86),
	.w8(32'h3bbaddd1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9b2a),
	.w1(32'h3dbaa48b),
	.w2(32'h3e327032),
	.w3(32'h3d94e326),
	.w4(32'h3e0c6eb4),
	.w5(32'h3dc82449),
	.w6(32'h3e0447c4),
	.w7(32'h3e63e461),
	.w8(32'h3e339217),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule