module layer_10_featuremap_286(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c276806),
	.w1(32'h3c1e5160),
	.w2(32'h3c3061e0),
	.w3(32'h3c0cbf48),
	.w4(32'h3c167300),
	.w5(32'h3a9a0a27),
	.w6(32'h3c18100e),
	.w7(32'h3c2ed103),
	.w8(32'hb97420b3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbac80),
	.w1(32'h394a7fb3),
	.w2(32'h3aea709a),
	.w3(32'h39061fd0),
	.w4(32'hbab392ed),
	.w5(32'hbb8f8a8d),
	.w6(32'h39926aa6),
	.w7(32'h39874940),
	.w8(32'hb9acca7a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad00345),
	.w1(32'hba1e7ee8),
	.w2(32'h36a2e796),
	.w3(32'hbb1ce500),
	.w4(32'hbab90208),
	.w5(32'hbaf3a91a),
	.w6(32'hbaab1998),
	.w7(32'h3b5d1da9),
	.w8(32'hbb289621),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76adcc),
	.w1(32'hbb4a6988),
	.w2(32'hbb38df7d),
	.w3(32'hbae7af35),
	.w4(32'hbaabd294),
	.w5(32'h3ab5fa99),
	.w6(32'hba811142),
	.w7(32'hbb30e04e),
	.w8(32'h3a8c296a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c976f),
	.w1(32'hbad8f92e),
	.w2(32'h39bae220),
	.w3(32'h395736ff),
	.w4(32'h3b276927),
	.w5(32'hbaaaadaa),
	.w6(32'hbb0b6726),
	.w7(32'h38a02cfc),
	.w8(32'hbb2da437),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29992d),
	.w1(32'hbafdbbbb),
	.w2(32'hba6eaf5d),
	.w3(32'hba442f97),
	.w4(32'hba683bed),
	.w5(32'hbaf9a03c),
	.w6(32'hbaafff82),
	.w7(32'hbaf0025c),
	.w8(32'hbb243746),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368d16),
	.w1(32'h39d55075),
	.w2(32'hba048e49),
	.w3(32'hbb0a81ca),
	.w4(32'h3b6bafe1),
	.w5(32'h3acc689b),
	.w6(32'hbaffcf5a),
	.w7(32'h3b1d428f),
	.w8(32'h3b062450),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1afde1),
	.w1(32'h3ba891f4),
	.w2(32'hbadbe8a8),
	.w3(32'h3c054ea9),
	.w4(32'h3c33fb80),
	.w5(32'hbb2aa060),
	.w6(32'h3c02e162),
	.w7(32'h3b81ca40),
	.w8(32'hba3176bf),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c91f),
	.w1(32'h3b4a48c0),
	.w2(32'h3bb9d3d1),
	.w3(32'h394a3af5),
	.w4(32'h3b240660),
	.w5(32'h3a422d5f),
	.w6(32'h3b056ff2),
	.w7(32'h3b92af03),
	.w8(32'hba7ca864),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb814d3f),
	.w1(32'hbbaead9a),
	.w2(32'hbbf841e6),
	.w3(32'hbaa07eda),
	.w4(32'h37e24c46),
	.w5(32'hbb935875),
	.w6(32'h39a66d75),
	.w7(32'hb89e09e7),
	.w8(32'hbba1c2ee),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4be794),
	.w1(32'hbb4b1859),
	.w2(32'hbb859ba2),
	.w3(32'hbae65bec),
	.w4(32'hbb23fbfb),
	.w5(32'h3b2e4bf5),
	.w6(32'hbacaa2ca),
	.w7(32'hbb8014be),
	.w8(32'hb910404e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06e299),
	.w1(32'h3b19af03),
	.w2(32'h3b511031),
	.w3(32'h3b03143b),
	.w4(32'h3bf3b99a),
	.w5(32'h3be77d58),
	.w6(32'h3a962694),
	.w7(32'h3baa3588),
	.w8(32'h3baf2693),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43041f),
	.w1(32'hbb0f172a),
	.w2(32'hbb964383),
	.w3(32'h3a2ecbe6),
	.w4(32'h3b46b2f1),
	.w5(32'hbad5944f),
	.w6(32'h3b38cef2),
	.w7(32'h3b9218aa),
	.w8(32'h3af5bb0e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56767),
	.w1(32'hba9ef123),
	.w2(32'h39f5be9b),
	.w3(32'hba798a26),
	.w4(32'h3b12588e),
	.w5(32'hbb3e97f6),
	.w6(32'hbaf7b4fc),
	.w7(32'h3a0496b6),
	.w8(32'hbb18b993),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8452d4),
	.w1(32'hbb47e20b),
	.w2(32'hbb0423b5),
	.w3(32'hba5977f6),
	.w4(32'hba092aef),
	.w5(32'h3baf31af),
	.w6(32'h3998e3af),
	.w7(32'h3a7796cb),
	.w8(32'h3b83e5c3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de0a3),
	.w1(32'hbaa883ee),
	.w2(32'hbb37d11c),
	.w3(32'h3bab1426),
	.w4(32'hba13bb60),
	.w5(32'hba94bc25),
	.w6(32'h3bd277b7),
	.w7(32'h3a073754),
	.w8(32'hbb7b0174),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab28b14),
	.w1(32'h3af868b1),
	.w2(32'h3b8aafb0),
	.w3(32'h3b08669d),
	.w4(32'h3b06cc4f),
	.w5(32'hba89f7e7),
	.w6(32'h3aafb2cb),
	.w7(32'h3b803ffd),
	.w8(32'hba34ec1f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fd52e0),
	.w1(32'hba855a07),
	.w2(32'hbb9b44bb),
	.w3(32'h3b104779),
	.w4(32'h3b37c6b4),
	.w5(32'hbbe3da3c),
	.w6(32'h3b0d4726),
	.w7(32'h38dd8516),
	.w8(32'hbc17d268),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6bcae),
	.w1(32'hbba43b16),
	.w2(32'hbbcbd2d0),
	.w3(32'hbaa1816e),
	.w4(32'hb9ff067c),
	.w5(32'hb842174e),
	.w6(32'hbb151cf8),
	.w7(32'hbb31628b),
	.w8(32'h3aecb41f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbab801),
	.w1(32'h3b490e2e),
	.w2(32'h3b4d4bee),
	.w3(32'h3b6ab444),
	.w4(32'h3c1a15cd),
	.w5(32'h3b4897cf),
	.w6(32'h37e0f5af),
	.w7(32'h3c0cfc5b),
	.w8(32'h3b6a620f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215f4d),
	.w1(32'h3aca09ce),
	.w2(32'h38e2356c),
	.w3(32'h3abbd943),
	.w4(32'hb9c5a698),
	.w5(32'h3ab07326),
	.w6(32'h3b59217b),
	.w7(32'h3a0bf6b9),
	.w8(32'h3b06ff31),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abab48c),
	.w1(32'h3b726cff),
	.w2(32'h3b8e4832),
	.w3(32'h3adab7ec),
	.w4(32'h3b64276b),
	.w5(32'h3b79a449),
	.w6(32'h3b3df600),
	.w7(32'h3b5a024d),
	.w8(32'h3b377229),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04dbf8),
	.w1(32'h3ab78da1),
	.w2(32'hbb401a73),
	.w3(32'h3c7836d3),
	.w4(32'h3c05c917),
	.w5(32'h3a83f907),
	.w6(32'h3c1d6e56),
	.w7(32'h3a72b8e0),
	.w8(32'hbba0eeca),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4270dc),
	.w1(32'hbb8394f7),
	.w2(32'hbbe7bbdb),
	.w3(32'hb98760b1),
	.w4(32'hbad90316),
	.w5(32'h3b179044),
	.w6(32'h3b14991e),
	.w7(32'hbb2423a1),
	.w8(32'h3bf02a96),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a7f71),
	.w1(32'h3c2c6313),
	.w2(32'h3c467be5),
	.w3(32'h3a05bcd5),
	.w4(32'hb9d588da),
	.w5(32'hba81c20d),
	.w6(32'h3c2dd87e),
	.w7(32'h3c2fa49d),
	.w8(32'hbaae6445),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77c8d8),
	.w1(32'hbb3d13d1),
	.w2(32'hbad4d599),
	.w3(32'h39246393),
	.w4(32'h39c5b3b6),
	.w5(32'h3ba825da),
	.w6(32'hb9ee23b2),
	.w7(32'hb9fd4216),
	.w8(32'h3bda597d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95fd7c),
	.w1(32'h3bc424d7),
	.w2(32'h3c088569),
	.w3(32'h3ba83009),
	.w4(32'h3be16b3d),
	.w5(32'h3bdcce21),
	.w6(32'h3be629ba),
	.w7(32'h3c1683d7),
	.w8(32'h3bbf592b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79c8b2),
	.w1(32'h3b7ea7cc),
	.w2(32'h3c0b3398),
	.w3(32'h3b88ea3c),
	.w4(32'h3c123c2e),
	.w5(32'h3b8a1e74),
	.w6(32'h3a7279ed),
	.w7(32'h3bd06b60),
	.w8(32'h3b43d2d1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecc4d2),
	.w1(32'h3abc244a),
	.w2(32'h3b204409),
	.w3(32'hbb56a1f2),
	.w4(32'h3b10f1ac),
	.w5(32'hbba7941f),
	.w6(32'h38ca80ae),
	.w7(32'h37bf8b78),
	.w8(32'hbb73be1b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe181f9),
	.w1(32'hbbf1ed7e),
	.w2(32'hbbac8163),
	.w3(32'hbb467122),
	.w4(32'hbaaf6982),
	.w5(32'h398fb651),
	.w6(32'hbbd13c99),
	.w7(32'h3957d5f8),
	.w8(32'h3b3ced1b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3f58),
	.w1(32'hbb42764b),
	.w2(32'hba988c0b),
	.w3(32'h3bb241ae),
	.w4(32'h3be50ae7),
	.w5(32'h3a86ec78),
	.w6(32'hbb07ddd9),
	.w7(32'hb96ffa38),
	.w8(32'h39aadf52),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308c64),
	.w1(32'hbaa093fa),
	.w2(32'h394671f3),
	.w3(32'hbb0d5eed),
	.w4(32'hbafbe497),
	.w5(32'h39cda9f6),
	.w6(32'hbb1b193c),
	.w7(32'hbb55a051),
	.w8(32'h3a219cab),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a6e3a),
	.w1(32'hba3dcf5e),
	.w2(32'hba18f608),
	.w3(32'hb91fa182),
	.w4(32'h3b107353),
	.w5(32'h3a6a3642),
	.w6(32'hbaea07ea),
	.w7(32'h3b57865a),
	.w8(32'h3a7fe14e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b62fb),
	.w1(32'h39f65100),
	.w2(32'h3a5b9460),
	.w3(32'h39db20ea),
	.w4(32'hba7916f7),
	.w5(32'h3ba89624),
	.w6(32'h3b49c89c),
	.w7(32'hba5492e6),
	.w8(32'h3b8e0a98),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9048ed),
	.w1(32'h3be18969),
	.w2(32'h3bcddbd7),
	.w3(32'h3b6eba6a),
	.w4(32'hbaa0764b),
	.w5(32'hbb14e000),
	.w6(32'h3c290326),
	.w7(32'h3b41dee5),
	.w8(32'h3a160578),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc4cd1),
	.w1(32'hbabd5eba),
	.w2(32'hba46f37f),
	.w3(32'hbaffa6e6),
	.w4(32'h3ad7e1b6),
	.w5(32'h3b8e689a),
	.w6(32'hba2daf1d),
	.w7(32'h3b1f93f6),
	.w8(32'h3b556925),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa4ee2),
	.w1(32'h3c1c4e03),
	.w2(32'h3bfe6ba5),
	.w3(32'hbb773235),
	.w4(32'hbb1220ef),
	.w5(32'h3bce19f5),
	.w6(32'hb99f6bf9),
	.w7(32'h3ab36ba4),
	.w8(32'h3b797a70),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b3bb5),
	.w1(32'h3b381d14),
	.w2(32'h3bf17d59),
	.w3(32'hbb3e3c46),
	.w4(32'hbad84986),
	.w5(32'hba4c7cda),
	.w6(32'hba20b64b),
	.w7(32'h3b25cf24),
	.w8(32'hbb02f111),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8b58),
	.w1(32'hbb3fbd96),
	.w2(32'h3aba22ca),
	.w3(32'hbb575b95),
	.w4(32'hbb20908f),
	.w5(32'hbb54cb55),
	.w6(32'hbbcf35b6),
	.w7(32'h3929b804),
	.w8(32'hbb87275b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc194),
	.w1(32'hbbca7ccf),
	.w2(32'hbb984c7a),
	.w3(32'hbb9104b4),
	.w4(32'hbb23858d),
	.w5(32'h3b9e558a),
	.w6(32'hbbb2c3a0),
	.w7(32'hbb5560e0),
	.w8(32'h3ac752a6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f1957),
	.w1(32'h3b2d2b66),
	.w2(32'h3b68bb35),
	.w3(32'h3b944a04),
	.w4(32'h3bab07fb),
	.w5(32'hba0c7bdb),
	.w6(32'h3c0ac961),
	.w7(32'h3a64ec2a),
	.w8(32'hbaebc7ec),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27d5e4),
	.w1(32'hbad7ab1c),
	.w2(32'hb9f4c65c),
	.w3(32'hba72fe5f),
	.w4(32'h3a1f1400),
	.w5(32'hbb4ab793),
	.w6(32'hba5b9882),
	.w7(32'hba38f03c),
	.w8(32'hbb1b6698),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bb06),
	.w1(32'hba3400fd),
	.w2(32'hbab2aaf2),
	.w3(32'hbb806dba),
	.w4(32'hbb144d51),
	.w5(32'h3b0fbceb),
	.w6(32'hbb0b8ce2),
	.w7(32'hbb250768),
	.w8(32'h3941246e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd7ad),
	.w1(32'hbb4560e4),
	.w2(32'hbbd81ce3),
	.w3(32'h3a7d62d5),
	.w4(32'h3a4c6211),
	.w5(32'hbba7c3cc),
	.w6(32'hba6ce349),
	.w7(32'h3a0b3e22),
	.w8(32'hbc224225),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863e9d),
	.w1(32'hbb979af8),
	.w2(32'hbbdf23ec),
	.w3(32'hba270ea4),
	.w4(32'hbb1d6403),
	.w5(32'h3b97cbef),
	.w6(32'hbae616fd),
	.w7(32'hbb894519),
	.w8(32'h3b86ba1d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18d11),
	.w1(32'h3a597d20),
	.w2(32'h390e42ff),
	.w3(32'h3b463ff3),
	.w4(32'h3b62232c),
	.w5(32'h3af71ee0),
	.w6(32'h3a84425a),
	.w7(32'h3b334d66),
	.w8(32'h3b26bdd3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349528),
	.w1(32'h3a59ac11),
	.w2(32'h3a4b7ece),
	.w3(32'h3b796e7a),
	.w4(32'h3b0cc5ad),
	.w5(32'h39381291),
	.w6(32'h3b5d77cc),
	.w7(32'h3b3fca78),
	.w8(32'h3ac6b17f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e1aea),
	.w1(32'h3ac6a143),
	.w2(32'h3abf8c2b),
	.w3(32'h3ab6d241),
	.w4(32'h3ba2326a),
	.w5(32'hbb43ad63),
	.w6(32'h3bc5e90b),
	.w7(32'h3bde5e6c),
	.w8(32'hbb50ac8f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec2cbd),
	.w1(32'h386ad65b),
	.w2(32'h395f2e3a),
	.w3(32'hba0b6a0f),
	.w4(32'hba0529f1),
	.w5(32'h381c2f62),
	.w6(32'h3a861eaf),
	.w7(32'h39db084c),
	.w8(32'h39633638),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f01991),
	.w1(32'h3add17c0),
	.w2(32'h3b6820cc),
	.w3(32'h3a459f2a),
	.w4(32'h3b510487),
	.w5(32'h3b9dff95),
	.w6(32'h3849d5ca),
	.w7(32'h3b1642aa),
	.w8(32'h3bbdce5f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b65243),
	.w1(32'hbb05c950),
	.w2(32'h39c32c7a),
	.w3(32'hbabe7e66),
	.w4(32'hb9a41169),
	.w5(32'hba63837d),
	.w6(32'hbb2a5da1),
	.w7(32'h3aa2475b),
	.w8(32'hbadf4fb4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c77fc),
	.w1(32'hbb720878),
	.w2(32'hbbc6cd23),
	.w3(32'hbabbb7fd),
	.w4(32'hbacd498a),
	.w5(32'hba75fada),
	.w6(32'hbb46da40),
	.w7(32'hbb567a37),
	.w8(32'hbb1392ab),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae32628),
	.w1(32'hbb066b67),
	.w2(32'hbb77f70a),
	.w3(32'h3aa8c0bb),
	.w4(32'h3a5d2e8e),
	.w5(32'h39efbff3),
	.w6(32'hb9838f4f),
	.w7(32'hbafec0ad),
	.w8(32'hb8096f8f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d77aa),
	.w1(32'h3a1c8658),
	.w2(32'hbb838513),
	.w3(32'h3bc049a5),
	.w4(32'h3b950ae7),
	.w5(32'hba13e3fd),
	.w6(32'h3b944e59),
	.w7(32'h3b36d071),
	.w8(32'hbb7c7c80),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e904b),
	.w1(32'h3ae9ec25),
	.w2(32'h3abd0ff1),
	.w3(32'h3bb6aeea),
	.w4(32'h3bf59295),
	.w5(32'h3b2bd476),
	.w6(32'hba35d735),
	.w7(32'h3b7ee1b5),
	.w8(32'h3b5b96e6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d304a),
	.w1(32'h3b619e8e),
	.w2(32'h3b172f62),
	.w3(32'hba3b9775),
	.w4(32'hbb950a2d),
	.w5(32'h3beb5937),
	.w6(32'h3bbd717c),
	.w7(32'hbb3e90ae),
	.w8(32'h3baa26cd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaa7db),
	.w1(32'h3bd3aea4),
	.w2(32'h3bd3729d),
	.w3(32'h3b9f7c1c),
	.w4(32'h3b2fd89b),
	.w5(32'h3b4cad71),
	.w6(32'h3c356670),
	.w7(32'h3ad686dd),
	.w8(32'h3b78e12f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f0f48),
	.w1(32'h3b1cd488),
	.w2(32'hb99d292b),
	.w3(32'h3b9cd65e),
	.w4(32'h3b93fe7e),
	.w5(32'hbaf6ca80),
	.w6(32'h3b0a0e82),
	.w7(32'h3b27a6d7),
	.w8(32'hbabf628f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4861e),
	.w1(32'h3a3a3c94),
	.w2(32'h3b22ac7e),
	.w3(32'hbaada7ed),
	.w4(32'h3ac771c8),
	.w5(32'h3bc8139b),
	.w6(32'hbad2fe6d),
	.w7(32'h3a070622),
	.w8(32'h3bf5dbb1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09eb16),
	.w1(32'h3c309886),
	.w2(32'h3be27ea7),
	.w3(32'h3bd25247),
	.w4(32'h3bb4684b),
	.w5(32'hba0c8752),
	.w6(32'h3bf5ddac),
	.w7(32'h3bda42e6),
	.w8(32'hba9bb326),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80276e),
	.w1(32'hba9379fb),
	.w2(32'hb9a3573a),
	.w3(32'h3b47e6f8),
	.w4(32'h3ba39edb),
	.w5(32'h3b606155),
	.w6(32'h3aad1245),
	.w7(32'h3b8b8c1d),
	.w8(32'hba4287c9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f7f5d),
	.w1(32'h3a12afdd),
	.w2(32'h3b4d50d2),
	.w3(32'h3bac53b5),
	.w4(32'h3baec180),
	.w5(32'hbab710dd),
	.w6(32'h3ac3f1e3),
	.w7(32'h3b0cf5c9),
	.w8(32'hbb86eb8e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12fcbc),
	.w1(32'h3b0ec6ec),
	.w2(32'h3a78be8c),
	.w3(32'h39281b19),
	.w4(32'hba75150c),
	.w5(32'h3b2c0025),
	.w6(32'hba116d15),
	.w7(32'hba4eff9b),
	.w8(32'h3b14822d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa911),
	.w1(32'h3a94e6ff),
	.w2(32'hb912d449),
	.w3(32'h3b35177e),
	.w4(32'hbaa76ae4),
	.w5(32'h3b237099),
	.w6(32'h3bf3313a),
	.w7(32'hbafbac7c),
	.w8(32'h3a7048ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9daafea),
	.w1(32'h38814bec),
	.w2(32'hb8804f0f),
	.w3(32'h3b3be074),
	.w4(32'hbad6e4e6),
	.w5(32'h3bacd66d),
	.w6(32'h3a339af9),
	.w7(32'hba59247e),
	.w8(32'hba6dc772),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a881f93),
	.w1(32'h3a81ecca),
	.w2(32'h37d95582),
	.w3(32'h3bd5f800),
	.w4(32'h3bcb10dc),
	.w5(32'hbb4648e3),
	.w6(32'h39a06dfa),
	.w7(32'hba1df568),
	.w8(32'hbb66be43),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca370e),
	.w1(32'hbb95408e),
	.w2(32'hbbe6433a),
	.w3(32'hbae61b71),
	.w4(32'hb9946c7c),
	.w5(32'hbc42bf63),
	.w6(32'h3b833cc3),
	.w7(32'h3ba7fea9),
	.w8(32'hbc1d7b5b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d4974),
	.w1(32'h3b1aae50),
	.w2(32'hbb0a7a7e),
	.w3(32'hbb0bbe9f),
	.w4(32'hbb8d0785),
	.w5(32'hbb73b4ce),
	.w6(32'h3bc09372),
	.w7(32'h3b1d0f1c),
	.w8(32'hbb59b7cc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ba4f1),
	.w1(32'h3b0e7876),
	.w2(32'h3b9cfd34),
	.w3(32'h3b94e90c),
	.w4(32'h3bedb6c5),
	.w5(32'hbbbcb083),
	.w6(32'h3aa0a000),
	.w7(32'h3c076c8f),
	.w8(32'hbbd53943),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e8a61),
	.w1(32'hbb1c576c),
	.w2(32'hbb066b93),
	.w3(32'hbb84fbe3),
	.w4(32'hba50a7cd),
	.w5(32'h39bfa640),
	.w6(32'hbb4b0d4a),
	.w7(32'hba33eac6),
	.w8(32'hb7f9d2c0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90451d),
	.w1(32'h3b189f65),
	.w2(32'h3adca1ff),
	.w3(32'h3a007dab),
	.w4(32'h3aa16951),
	.w5(32'hb9fdbdc3),
	.w6(32'h3b060a82),
	.w7(32'h3a918616),
	.w8(32'hba90209b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2d8d4),
	.w1(32'hba562c3a),
	.w2(32'hba2f330b),
	.w3(32'hb794d787),
	.w4(32'h3a98066a),
	.w5(32'hbb3bd370),
	.w6(32'h3a6a558f),
	.w7(32'h3ac74837),
	.w8(32'hbb21a12e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9880c0c),
	.w1(32'hb98595ac),
	.w2(32'hb9eaae98),
	.w3(32'hbb25fff7),
	.w4(32'hbb305596),
	.w5(32'h39ca5c23),
	.w6(32'hb9dd1cdc),
	.w7(32'hbae5d73e),
	.w8(32'h3a8d6e19),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b306bbe),
	.w1(32'h3a4c065b),
	.w2(32'hba2a87c8),
	.w3(32'hb844fe26),
	.w4(32'hb8746022),
	.w5(32'hb9490a32),
	.w6(32'h37e4e27d),
	.w7(32'h384cb2d7),
	.w8(32'hbae6424f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8492),
	.w1(32'h3a77e410),
	.w2(32'h3a66c353),
	.w3(32'h3b1902f7),
	.w4(32'h3a281578),
	.w5(32'h3afe6d70),
	.w6(32'h3b39a553),
	.w7(32'h3b085685),
	.w8(32'h3b4ffe17),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f94af),
	.w1(32'h3ae1a3d5),
	.w2(32'hba52803e),
	.w3(32'h3afb7803),
	.w4(32'h3a7ad6ec),
	.w5(32'h3be0e0ba),
	.w6(32'h3ba1a153),
	.w7(32'h3b1df25f),
	.w8(32'h3b7eaecd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc184e1),
	.w1(32'h3b70030c),
	.w2(32'hb98d373e),
	.w3(32'h3c2e7990),
	.w4(32'h3c020aec),
	.w5(32'hba543dfe),
	.w6(32'h3c2061b2),
	.w7(32'h3a151dac),
	.w8(32'hbb68b260),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc171cdd),
	.w1(32'hbc2d4fdd),
	.w2(32'hbc079762),
	.w3(32'hbbf085dc),
	.w4(32'hbbc31f6e),
	.w5(32'hbaccada6),
	.w6(32'hbbb3052e),
	.w7(32'hbbbc4ce2),
	.w8(32'hb816e94d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f455e),
	.w1(32'h39db31ef),
	.w2(32'hbac09614),
	.w3(32'h3b3c655a),
	.w4(32'h3b3d89d4),
	.w5(32'hb97fac05),
	.w6(32'h3b21f9e1),
	.w7(32'h3a396492),
	.w8(32'hbb182939),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9da34),
	.w1(32'h3a74de83),
	.w2(32'h3a8bc5bd),
	.w3(32'hb89c9732),
	.w4(32'h3a62a7d8),
	.w5(32'hbaf6da94),
	.w6(32'h3b5e9c4f),
	.w7(32'h3bbcecb5),
	.w8(32'h3ac67af9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d83d3),
	.w1(32'h3b4003ea),
	.w2(32'h3b0e9cfd),
	.w3(32'h3b0320d6),
	.w4(32'h3b87b888),
	.w5(32'h3a817cfa),
	.w6(32'h3b915060),
	.w7(32'h3b53acb6),
	.w8(32'h3ae08e9d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba478b),
	.w1(32'hbab5faf3),
	.w2(32'hbb222efa),
	.w3(32'h3a87e568),
	.w4(32'h3aa608d0),
	.w5(32'hb9a0eef6),
	.w6(32'h3b514b85),
	.w7(32'h3abdb34f),
	.w8(32'hbaaf9ae1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba6475),
	.w1(32'hba499719),
	.w2(32'hb96ec16c),
	.w3(32'h3b0f415f),
	.w4(32'h39057c78),
	.w5(32'hbb8816ff),
	.w6(32'hb92f0a88),
	.w7(32'hb88bff1a),
	.w8(32'hbb9b4180),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16223),
	.w1(32'hbb90dc1d),
	.w2(32'hbb88e4e0),
	.w3(32'hbba46299),
	.w4(32'hbb8c654b),
	.w5(32'h3b0198b9),
	.w6(32'hbb6c1443),
	.w7(32'hbb5fbf57),
	.w8(32'h3aa68b5a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a407529),
	.w1(32'hb8900cbc),
	.w2(32'h38a39cd9),
	.w3(32'h3b3554fb),
	.w4(32'h3a1fdfb2),
	.w5(32'h3b7ddd06),
	.w6(32'hba78a7cf),
	.w7(32'hb85c6350),
	.w8(32'h3ad89643),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47869d),
	.w1(32'h3b11253d),
	.w2(32'hb9fb0e3a),
	.w3(32'h3b82ce69),
	.w4(32'h3b4301d2),
	.w5(32'hbb2eb589),
	.w6(32'h3a50f921),
	.w7(32'hba0cb5d3),
	.w8(32'hbac0b0a7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1da156),
	.w1(32'hbb2eabb0),
	.w2(32'h3ac4a3f1),
	.w3(32'h38c7e8cd),
	.w4(32'hba478dec),
	.w5(32'h3b949b9f),
	.w6(32'hbad66fe4),
	.w7(32'h3afd7e87),
	.w8(32'h3b106c6a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c3d24),
	.w1(32'hb6b8ac99),
	.w2(32'hba563c22),
	.w3(32'h3b879b37),
	.w4(32'h3b908bff),
	.w5(32'h3a6c5912),
	.w6(32'hbaccac6e),
	.w7(32'hb9fed612),
	.w8(32'h3a1b1d70),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a291636),
	.w1(32'h3958d1cc),
	.w2(32'h3ac98af6),
	.w3(32'hb9670583),
	.w4(32'h3a09e57d),
	.w5(32'hbb08fe15),
	.w6(32'hb8d5445c),
	.w7(32'h39f7c5ab),
	.w8(32'hbb4eb7a2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4e1c),
	.w1(32'hbbb29625),
	.w2(32'hbb2097fb),
	.w3(32'h3b17cf39),
	.w4(32'hbb21225b),
	.w5(32'h3aa1e329),
	.w6(32'h3b6979f7),
	.w7(32'hbb753919),
	.w8(32'hba6d4dfc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a158a),
	.w1(32'hba728a1d),
	.w2(32'h3b128e51),
	.w3(32'hbab82a97),
	.w4(32'h3b36f0b7),
	.w5(32'hb9bc88e7),
	.w6(32'hbafd2e21),
	.w7(32'h3b13c2e6),
	.w8(32'hb9452dc5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae69c71),
	.w1(32'hbbbcaa6a),
	.w2(32'hbc04c3c3),
	.w3(32'hbb63f1d7),
	.w4(32'hbaf77979),
	.w5(32'h3b145730),
	.w6(32'hbb5cc25d),
	.w7(32'hbb0834f6),
	.w8(32'h3a8e898c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99c687),
	.w1(32'h38ecd574),
	.w2(32'h3adc2c9c),
	.w3(32'hbacbe54a),
	.w4(32'hba06033d),
	.w5(32'h3930a02e),
	.w6(32'hb9b22d4b),
	.w7(32'hba4de92e),
	.w8(32'h3b5b109c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65e015),
	.w1(32'h3b1b7092),
	.w2(32'hbaf42ea4),
	.w3(32'h3b3da595),
	.w4(32'hb999c9e4),
	.w5(32'h397ffec5),
	.w6(32'h3b9f875f),
	.w7(32'h3b0fda7c),
	.w8(32'hbb44dee6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a903a),
	.w1(32'h39756860),
	.w2(32'h39a64b0e),
	.w3(32'h3b9dc2da),
	.w4(32'h3b36f6ef),
	.w5(32'hbb869c18),
	.w6(32'h3b83591c),
	.w7(32'h3b36b598),
	.w8(32'hbb8aaa7a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea95f),
	.w1(32'hbb96145f),
	.w2(32'hbb92d66c),
	.w3(32'hbb3e9cd8),
	.w4(32'hbb514236),
	.w5(32'hbb15ccc3),
	.w6(32'hbb1adf3b),
	.w7(32'hbad6568e),
	.w8(32'hb91abfb0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83d47e),
	.w1(32'hba4e8092),
	.w2(32'hba8013c3),
	.w3(32'hbb0c64f1),
	.w4(32'hbae8351e),
	.w5(32'h3a4d7a73),
	.w6(32'hbb1db00a),
	.w7(32'hbb629d62),
	.w8(32'hba7d3a19),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f9464),
	.w1(32'hbbe3ed71),
	.w2(32'hbc19384a),
	.w3(32'hbacbfc7e),
	.w4(32'h394f3c9a),
	.w5(32'hbb0cea9d),
	.w6(32'hbb01df85),
	.w7(32'hbbc2657f),
	.w8(32'hbb7b0a3a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b165e7a),
	.w1(32'hbb00159c),
	.w2(32'hbb2f33c4),
	.w3(32'hbb0fff0c),
	.w4(32'hba222a7a),
	.w5(32'hbb21905f),
	.w6(32'hbab5afa6),
	.w7(32'h3a99a171),
	.w8(32'hbb31f6c2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f489f),
	.w1(32'h3b82a1e5),
	.w2(32'h3bf367d1),
	.w3(32'h3b395768),
	.w4(32'h3ae18fca),
	.w5(32'h3c02763b),
	.w6(32'h3b3ee9f4),
	.w7(32'hba3a6299),
	.w8(32'hbb202555),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bf0812),
	.w1(32'h3b482d2f),
	.w2(32'h3ac9fa3a),
	.w3(32'h3b612d3b),
	.w4(32'h3b8403e7),
	.w5(32'h3b23d407),
	.w6(32'hb82764fb),
	.w7(32'h3acf5ce2),
	.w8(32'h3b4b3da2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6db0b),
	.w1(32'hbb02a3d7),
	.w2(32'hba1bcd9b),
	.w3(32'hba9f52c9),
	.w4(32'hbad3437f),
	.w5(32'hbadb46eb),
	.w6(32'hb89675f2),
	.w7(32'h39862776),
	.w8(32'hbaab76f9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b042b),
	.w1(32'h3aec4bdc),
	.w2(32'hb8b28d0b),
	.w3(32'hbad42bd5),
	.w4(32'hb9bb034b),
	.w5(32'h3ba6c833),
	.w6(32'h3a12647a),
	.w7(32'h3a754864),
	.w8(32'h3b1693ee),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3dff6),
	.w1(32'h3b4e6f76),
	.w2(32'h3adfbb33),
	.w3(32'h3b9d1a3e),
	.w4(32'h3ba4c47b),
	.w5(32'hbafd29ad),
	.w6(32'h3b0e3995),
	.w7(32'h3b9b5a7b),
	.w8(32'hbb193c82),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80699),
	.w1(32'h3bbfd23d),
	.w2(32'h3b957a4f),
	.w3(32'h3a29bc42),
	.w4(32'h3aab541b),
	.w5(32'h3c1a6fda),
	.w6(32'h3a9c771b),
	.w7(32'h3b0b7788),
	.w8(32'h3b84b98c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18bce6),
	.w1(32'hbb710298),
	.w2(32'hbb259436),
	.w3(32'hbb2f8872),
	.w4(32'hbb1050e6),
	.w5(32'h3bb7f134),
	.w6(32'hbb1b5e5f),
	.w7(32'hba535005),
	.w8(32'h3b5772f3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01d6e9),
	.w1(32'h39d136c7),
	.w2(32'h3aee4762),
	.w3(32'hba49e9ee),
	.w4(32'hbab45a8f),
	.w5(32'h3a46d633),
	.w6(32'h3a93bff8),
	.w7(32'h39d2cd17),
	.w8(32'hb92aeff6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393fdc77),
	.w1(32'hbaa9a5bd),
	.w2(32'h3a81a447),
	.w3(32'h3a01be9c),
	.w4(32'hba8ed4ca),
	.w5(32'h3a457cc8),
	.w6(32'h384d7331),
	.w7(32'h365a284e),
	.w8(32'hba931f67),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad00289),
	.w1(32'hbbab6fcb),
	.w2(32'hbb9a0514),
	.w3(32'hbb4b3692),
	.w4(32'hba7ae703),
	.w5(32'hbb4a9d2b),
	.w6(32'hbb9ff74d),
	.w7(32'hba775693),
	.w8(32'hbb3d3f7f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f73c),
	.w1(32'hbb41a157),
	.w2(32'hbb0397d4),
	.w3(32'hbb038fc2),
	.w4(32'hba7acf82),
	.w5(32'hba0e1952),
	.w6(32'hbb339848),
	.w7(32'hbacdace8),
	.w8(32'hba8c8da3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c6fe4),
	.w1(32'hbb26b492),
	.w2(32'hba5650cb),
	.w3(32'h3abff1db),
	.w4(32'h3adfe137),
	.w5(32'hb8670938),
	.w6(32'hbac8da97),
	.w7(32'h3a8dd2ea),
	.w8(32'hb9b36094),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04d120),
	.w1(32'hbac93638),
	.w2(32'hbacf463d),
	.w3(32'h3903380c),
	.w4(32'hbb1cbba9),
	.w5(32'hbb7df2e6),
	.w6(32'h3ad44b18),
	.w7(32'hbb15d67d),
	.w8(32'hbb7eb087),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb40f),
	.w1(32'hba7ff50f),
	.w2(32'hba18ff3d),
	.w3(32'hbb8f8370),
	.w4(32'hbb0c318b),
	.w5(32'hb87d7902),
	.w6(32'hbb188cbe),
	.w7(32'hbb83a435),
	.w8(32'hbb15efed),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa8b0),
	.w1(32'hba2e902f),
	.w2(32'hba52f208),
	.w3(32'h3a80f179),
	.w4(32'hba984d07),
	.w5(32'hbb657bfa),
	.w6(32'h3b087a83),
	.w7(32'h3a7c9679),
	.w8(32'hbb8cb611),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be089a),
	.w1(32'hbb1d6c1a),
	.w2(32'hbb98d7e5),
	.w3(32'hbb31d87c),
	.w4(32'hbb437c56),
	.w5(32'hbb431d4e),
	.w6(32'hbb425765),
	.w7(32'hbb8a1076),
	.w8(32'hbabafc03),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ad191),
	.w1(32'h399e8c17),
	.w2(32'h3ae9719a),
	.w3(32'h3a8fa7ed),
	.w4(32'h39acc9f5),
	.w5(32'hb91ca33c),
	.w6(32'h3b1fdffb),
	.w7(32'h3a0e523e),
	.w8(32'h3a1164cb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98aff3),
	.w1(32'h39f1e7d7),
	.w2(32'hba9d1062),
	.w3(32'hba499125),
	.w4(32'hba866def),
	.w5(32'hbb412c91),
	.w6(32'hb9bb5555),
	.w7(32'hba68c43b),
	.w8(32'hbb1916e9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e12b1),
	.w1(32'hbaec3931),
	.w2(32'hb9906929),
	.w3(32'hbb2ab7fd),
	.w4(32'hbb300103),
	.w5(32'hb883bab8),
	.w6(32'hbb376475),
	.w7(32'hbae76a7f),
	.w8(32'hba6fa8f1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399de2d4),
	.w1(32'hba8c4047),
	.w2(32'hba979569),
	.w3(32'hba5744a3),
	.w4(32'hba41390c),
	.w5(32'h3ab563d8),
	.w6(32'hbaf79d1a),
	.w7(32'hba0897dc),
	.w8(32'hbae86a0b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cb59a),
	.w1(32'hbb85229a),
	.w2(32'hbb533011),
	.w3(32'hba2e92e8),
	.w4(32'hb89933ff),
	.w5(32'hba819ce1),
	.w6(32'hbb86d933),
	.w7(32'hba6d70b2),
	.w8(32'h3a84dc9b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c6fc3),
	.w1(32'h3ac66714),
	.w2(32'h3984dee2),
	.w3(32'h3afa5e1f),
	.w4(32'h3ad6371d),
	.w5(32'h39e252ad),
	.w6(32'h3b99567c),
	.w7(32'h3b29739a),
	.w8(32'h3981e995),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3ffa1),
	.w1(32'hbabf965d),
	.w2(32'hba81c054),
	.w3(32'hba2e80ce),
	.w4(32'h3b04fcb2),
	.w5(32'hbadd729a),
	.w6(32'h3ab17a22),
	.w7(32'h3a928712),
	.w8(32'hbab2961b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab26d3e),
	.w1(32'hbb580cc1),
	.w2(32'hba172f6a),
	.w3(32'hbb6dd612),
	.w4(32'hbba653de),
	.w5(32'hbb895802),
	.w6(32'hbaf89976),
	.w7(32'hbae615a2),
	.w8(32'hbb57662d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb196d37),
	.w1(32'hbaff68f6),
	.w2(32'hbab7f1cf),
	.w3(32'hbb14c78c),
	.w4(32'hbb162546),
	.w5(32'hba641cee),
	.w6(32'hbb01c57b),
	.w7(32'hbaa00e77),
	.w8(32'hba3aedf4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bea5b),
	.w1(32'hba380c4e),
	.w2(32'hba9786b5),
	.w3(32'hba60edfa),
	.w4(32'hbaac481f),
	.w5(32'hb9b681e8),
	.w6(32'hba9433b5),
	.w7(32'hbab86573),
	.w8(32'hb9539a39),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d5e3b),
	.w1(32'h3afc422a),
	.w2(32'h3a7dcd19),
	.w3(32'hba60b17e),
	.w4(32'h3987a3cc),
	.w5(32'h39e7ee89),
	.w6(32'hb9bba4c4),
	.w7(32'h3a1f1692),
	.w8(32'h3a15af84),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8898b2f),
	.w1(32'hbb11a0b9),
	.w2(32'hba8c2e79),
	.w3(32'hbb08da2a),
	.w4(32'hbb0a9787),
	.w5(32'h3a2066d2),
	.w6(32'hbb120ea9),
	.w7(32'hba4ffc27),
	.w8(32'h3a0f3897),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e0c42),
	.w1(32'h3b20ce95),
	.w2(32'hb98a1f92),
	.w3(32'hbb8ebc70),
	.w4(32'h3b13a13f),
	.w5(32'hbaeb1d2d),
	.w6(32'hba6e434e),
	.w7(32'hbb0c2541),
	.w8(32'hbb9c59d9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30293f),
	.w1(32'hbb956b37),
	.w2(32'hbbfbdc46),
	.w3(32'hba1421a0),
	.w4(32'hba912a10),
	.w5(32'hbbbfa8dc),
	.w6(32'h3aef943c),
	.w7(32'hba0ea4f2),
	.w8(32'hbb8f869f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987114d),
	.w1(32'hba52d046),
	.w2(32'hba326926),
	.w3(32'hba8f0f12),
	.w4(32'hbaaf756f),
	.w5(32'hba53dfc9),
	.w6(32'h3ace7186),
	.w7(32'hb9aa5ad6),
	.w8(32'hba852abe),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62fee1),
	.w1(32'hb673739f),
	.w2(32'h3ab96998),
	.w3(32'hba2b5a81),
	.w4(32'hb9e36453),
	.w5(32'hba2d5602),
	.w6(32'h3a499533),
	.w7(32'hb9f17ed3),
	.w8(32'hba4fe1c2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb6682),
	.w1(32'hb9ddaefd),
	.w2(32'h392524fa),
	.w3(32'hba6a1b04),
	.w4(32'hb9dcdbe4),
	.w5(32'hbb41ea4f),
	.w6(32'hbae5ac1a),
	.w7(32'h39102a50),
	.w8(32'hbb6258fa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99eb630),
	.w1(32'hb99db054),
	.w2(32'hba0067b3),
	.w3(32'hbb504782),
	.w4(32'hbadcc8c6),
	.w5(32'hbacb17a6),
	.w6(32'hbb923ab3),
	.w7(32'hbb085ddf),
	.w8(32'hbaf5a801),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6848),
	.w1(32'hba8b84d3),
	.w2(32'hba2a3b91),
	.w3(32'h3a48c2fa),
	.w4(32'hba983c0f),
	.w5(32'hbb0da2fc),
	.w6(32'h3a0445ca),
	.w7(32'hbaa8d6ae),
	.w8(32'hbb44a081),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f539e),
	.w1(32'hbaf22616),
	.w2(32'hbb8bf814),
	.w3(32'hba28a6da),
	.w4(32'h3ace29f6),
	.w5(32'hbb2da9d9),
	.w6(32'h3b091fe1),
	.w7(32'h3b080c5b),
	.w8(32'hbb52c8a8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10a676),
	.w1(32'hba8ea8dc),
	.w2(32'hbae8ff25),
	.w3(32'hb96535fe),
	.w4(32'hbade0cb9),
	.w5(32'hbab7eb42),
	.w6(32'hba81ac29),
	.w7(32'hbb0073ec),
	.w8(32'hbac0bbbb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f70d8),
	.w1(32'hbb2c43cd),
	.w2(32'hbb82f9fe),
	.w3(32'hb9fd2cba),
	.w4(32'hbab3208d),
	.w5(32'hba813b29),
	.w6(32'h394509cf),
	.w7(32'hbac5e9c7),
	.w8(32'hb9accf6e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ca8e6),
	.w1(32'h3aaf6f09),
	.w2(32'hbaffd50f),
	.w3(32'h3ae21929),
	.w4(32'h3b14c74a),
	.w5(32'hba0f08b2),
	.w6(32'h3a8ea9b6),
	.w7(32'h3b0b478a),
	.w8(32'hbb0703fc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98871df),
	.w1(32'hba6aa891),
	.w2(32'hb9aafa7c),
	.w3(32'hbb028460),
	.w4(32'hbb3dcc44),
	.w5(32'hba2908b7),
	.w6(32'hbacb546b),
	.w7(32'hbb328475),
	.w8(32'hba958fea),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7fe5c),
	.w1(32'hbadf1f02),
	.w2(32'hbafaa013),
	.w3(32'h37a980d6),
	.w4(32'hb9ff8331),
	.w5(32'hbaf249ab),
	.w6(32'h3adf2069),
	.w7(32'h3a40a409),
	.w8(32'hbb5162bc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae44811),
	.w1(32'hba88ad6a),
	.w2(32'hbb2fc6e9),
	.w3(32'hb9e02a5b),
	.w4(32'hba85b1b9),
	.w5(32'h3a48c73f),
	.w6(32'hb9ff7df2),
	.w7(32'hbb0705fa),
	.w8(32'h3ab78e8a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d22e0d),
	.w1(32'hba0eb85b),
	.w2(32'hbb6a64e6),
	.w3(32'hba30da23),
	.w4(32'h396520fc),
	.w5(32'hbaacee23),
	.w6(32'h39a9f55e),
	.w7(32'hb778ab04),
	.w8(32'hb9dcfb00),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abae7a8),
	.w1(32'hb9908543),
	.w2(32'h39d21ce0),
	.w3(32'h3ad86be1),
	.w4(32'h3b064c2e),
	.w5(32'hba0528e3),
	.w6(32'hbadeb1e4),
	.w7(32'hb5b3fda2),
	.w8(32'hba53a4c0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b26a11),
	.w1(32'hb90d985d),
	.w2(32'h3aa1d093),
	.w3(32'hb8d06d6a),
	.w4(32'h3aa5fec6),
	.w5(32'hba6f5d51),
	.w6(32'h3a7bfbda),
	.w7(32'h3af6c302),
	.w8(32'hbaee2bdb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9f038),
	.w1(32'hbaef76be),
	.w2(32'hb9f9a7aa),
	.w3(32'hba8ea0a7),
	.w4(32'hbac122af),
	.w5(32'hba7f3f90),
	.w6(32'hbad1734b),
	.w7(32'hba971dc8),
	.w8(32'hba2a88a6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98c724),
	.w1(32'hbab7c85b),
	.w2(32'hba66f8ef),
	.w3(32'hba757db0),
	.w4(32'hba26340a),
	.w5(32'h3ad80144),
	.w6(32'hba043be2),
	.w7(32'hb9928a35),
	.w8(32'h3a4ab53c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f8c571),
	.w1(32'hbb0f212c),
	.w2(32'hba052387),
	.w3(32'h39d9a4e1),
	.w4(32'h39cd1bad),
	.w5(32'hba8c3df3),
	.w6(32'h39cf9ea2),
	.w7(32'h3b150416),
	.w8(32'h398c3048),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e50b),
	.w1(32'hbbabcd80),
	.w2(32'hbbe8759b),
	.w3(32'hbb5ca312),
	.w4(32'hba88d4a4),
	.w5(32'hbb06412b),
	.w6(32'hbb0c143f),
	.w7(32'hba9b52d3),
	.w8(32'h38a76439),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac81fc0),
	.w1(32'h3a482145),
	.w2(32'h39eb0c1b),
	.w3(32'hb9c8da0e),
	.w4(32'hb9e6b63d),
	.w5(32'h3aaebbd4),
	.w6(32'h39d10594),
	.w7(32'h3a9eb1a3),
	.w8(32'h3ab41297),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9618a2),
	.w1(32'hbacda13b),
	.w2(32'hbbad43c7),
	.w3(32'h3a4a02dc),
	.w4(32'h3ada73e4),
	.w5(32'hbb16efc5),
	.w6(32'hb9558e89),
	.w7(32'h3a8c00fc),
	.w8(32'hbaf44c15),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21a855),
	.w1(32'hbaec1b9c),
	.w2(32'hbb1a89e6),
	.w3(32'hba9e208a),
	.w4(32'hbb427d39),
	.w5(32'hba77a4a3),
	.w6(32'h3a1f1b9b),
	.w7(32'hba2ca367),
	.w8(32'hba31e727),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e7f0a),
	.w1(32'hbb265663),
	.w2(32'hbb6367b3),
	.w3(32'hbb07df07),
	.w4(32'h3adabcca),
	.w5(32'hba6241db),
	.w6(32'h3a99fce6),
	.w7(32'h3b09e5b9),
	.w8(32'hba38fc08),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15aa75),
	.w1(32'hbb2df0b6),
	.w2(32'h389212ef),
	.w3(32'h394bee07),
	.w4(32'hbad7600d),
	.w5(32'hbac32596),
	.w6(32'hbacca44b),
	.w7(32'h3aa89265),
	.w8(32'hbaf04768),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4865d2),
	.w1(32'h39bc2c1f),
	.w2(32'h3a6445d4),
	.w3(32'h3a5cf75a),
	.w4(32'hba6f87d7),
	.w5(32'hb9692696),
	.w6(32'hba658278),
	.w7(32'hba554d8c),
	.w8(32'hba8a509c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba523351),
	.w1(32'hba5ebd78),
	.w2(32'h391c8784),
	.w3(32'hbad6d463),
	.w4(32'hba925234),
	.w5(32'hbaff579b),
	.w6(32'hba7c06a1),
	.w7(32'hbaaa94e9),
	.w8(32'hbad6ee7a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf59ff5),
	.w1(32'hbaf67bb1),
	.w2(32'hbaf21847),
	.w3(32'hbac66c67),
	.w4(32'hba8a7d36),
	.w5(32'h3b17153c),
	.w6(32'hbae5d4b5),
	.w7(32'hbab6c41a),
	.w8(32'h3b4aef98),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afce5f7),
	.w1(32'h3aec4a96),
	.w2(32'h3b3d7ae8),
	.w3(32'h3a2a92d2),
	.w4(32'hbac84a3a),
	.w5(32'hb9b2c17e),
	.w6(32'h3a9536e9),
	.w7(32'h3ac2d818),
	.w8(32'h3a301af1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d404c),
	.w1(32'hba260694),
	.w2(32'h3abf3905),
	.w3(32'hba334919),
	.w4(32'hb8ee01bd),
	.w5(32'hb9cbaaf4),
	.w6(32'hba81a7fa),
	.w7(32'h3a01109a),
	.w8(32'hb579bb2e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5711c),
	.w1(32'hbad48b99),
	.w2(32'hbaa677b9),
	.w3(32'hb9e88e3c),
	.w4(32'h392e9689),
	.w5(32'hbab872d6),
	.w6(32'hb9c7d640),
	.w7(32'h390b74c6),
	.w8(32'h3a2a8d2c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d93d21),
	.w1(32'hb9b5272e),
	.w2(32'h39ed64c7),
	.w3(32'hbb26ab83),
	.w4(32'hbb42a0d3),
	.w5(32'h3b038a06),
	.w6(32'hba95a9aa),
	.w7(32'hba922a52),
	.w8(32'h3a7d0d69),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e5c721),
	.w1(32'hbaa18d52),
	.w2(32'hbaa8ce45),
	.w3(32'h3b4c2b2e),
	.w4(32'h3b38a099),
	.w5(32'hbac81d12),
	.w6(32'h3b0feb4f),
	.w7(32'h3a3504f8),
	.w8(32'hbb3acaf2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae7630),
	.w1(32'hba49206a),
	.w2(32'hbb6d2af2),
	.w3(32'hba04776a),
	.w4(32'hbb176b56),
	.w5(32'hba8497f7),
	.w6(32'hb6d30a08),
	.w7(32'hbb2e9ff5),
	.w8(32'hb9b181ce),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a785c50),
	.w1(32'hb9b5cee2),
	.w2(32'hba4da037),
	.w3(32'hba40b667),
	.w4(32'hba83e7ad),
	.w5(32'hbaf91985),
	.w6(32'hb9a41c3e),
	.w7(32'h3a2cec87),
	.w8(32'h39d5ceef),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08eaed),
	.w1(32'hbad807c8),
	.w2(32'hbb17df0a),
	.w3(32'hba55c1f8),
	.w4(32'hbac19178),
	.w5(32'hbab142a3),
	.w6(32'h395992a0),
	.w7(32'hbb1ad020),
	.w8(32'hbada1bae),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90b296),
	.w1(32'hbad68a08),
	.w2(32'hbb165b1a),
	.w3(32'hb9907b27),
	.w4(32'h3b2dd866),
	.w5(32'hb9e3df31),
	.w6(32'hbb268f1b),
	.w7(32'h3b0bd7fa),
	.w8(32'hba74db97),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925aa77),
	.w1(32'h39bdb5e4),
	.w2(32'hb95ab080),
	.w3(32'hb9fdbe9b),
	.w4(32'hba94e836),
	.w5(32'hbac6e2c0),
	.w6(32'h3ab210c5),
	.w7(32'hba0ed392),
	.w8(32'hbb086c83),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aa362),
	.w1(32'hba801671),
	.w2(32'hba5f2fe6),
	.w3(32'hbb098f8e),
	.w4(32'hbb070d91),
	.w5(32'h3b701db5),
	.w6(32'hbabcf504),
	.w7(32'hbaaf7b6f),
	.w8(32'h3b5af45a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5636e),
	.w1(32'h3b901312),
	.w2(32'h3b219f1a),
	.w3(32'h3baa6546),
	.w4(32'h3bba3f51),
	.w5(32'h37f9d258),
	.w6(32'h3b28521f),
	.w7(32'h3b8da66c),
	.w8(32'hb5fbde02),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f2348),
	.w1(32'h3a37290e),
	.w2(32'hbb1bcb43),
	.w3(32'h3b4ea27c),
	.w4(32'h3b486c38),
	.w5(32'h3aa54c45),
	.w6(32'h3bacde1d),
	.w7(32'h3b622f93),
	.w8(32'h38b24eb7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec458),
	.w1(32'hba137722),
	.w2(32'hb905bf19),
	.w3(32'hbae12fea),
	.w4(32'hba64fd21),
	.w5(32'hbb56f135),
	.w6(32'hbb2d88b6),
	.w7(32'hb99f63cc),
	.w8(32'hbb10d9e3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ca59c),
	.w1(32'hbb838ad5),
	.w2(32'hbb307231),
	.w3(32'hbb1652b9),
	.w4(32'hba82ba4c),
	.w5(32'hbb85d8d1),
	.w6(32'hba904727),
	.w7(32'hb93f7808),
	.w8(32'hbb70e00a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf06f24),
	.w1(32'hbb8be7d1),
	.w2(32'hba3968b4),
	.w3(32'hbb1de942),
	.w4(32'hbb0aeb99),
	.w5(32'h3a66dffc),
	.w6(32'hba873540),
	.w7(32'hbb0095b3),
	.w8(32'hbab03eb7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb701b53),
	.w1(32'hbb9972c6),
	.w2(32'hbbb25c30),
	.w3(32'h3ac2d796),
	.w4(32'h3b2201be),
	.w5(32'hbb62e074),
	.w6(32'hba6ee321),
	.w7(32'h3b2ac193),
	.w8(32'hbb8436af),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecda58),
	.w1(32'hba9b024b),
	.w2(32'hbaf7cb8a),
	.w3(32'hba0c2e56),
	.w4(32'h393e9bda),
	.w5(32'h3acba547),
	.w6(32'hbb1fb0c5),
	.w7(32'hbad7f278),
	.w8(32'hbaabfb91),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b582119),
	.w1(32'hbac5dcca),
	.w2(32'hbb858047),
	.w3(32'h3b5d9b6b),
	.w4(32'h3b4e6220),
	.w5(32'hba8d8d3a),
	.w6(32'h3ab2c463),
	.w7(32'h3b092652),
	.w8(32'hbb0ca20b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3058f),
	.w1(32'hb8a67e81),
	.w2(32'hb8a42c6d),
	.w3(32'hbab4db9a),
	.w4(32'hb9f8e7c7),
	.w5(32'hbac7c018),
	.w6(32'hba84a6df),
	.w7(32'hba0c1346),
	.w8(32'hbb0b87b8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a5f6),
	.w1(32'hbb630f83),
	.w2(32'hbbb4ff5f),
	.w3(32'hb9fd310c),
	.w4(32'hbabbbe9a),
	.w5(32'hba9348a2),
	.w6(32'h38d1b305),
	.w7(32'hbacb77d9),
	.w8(32'hba195ad8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a907a67),
	.w1(32'h3a2cb60a),
	.w2(32'h39a20c5c),
	.w3(32'hb8c31de9),
	.w4(32'h3a2d43fa),
	.w5(32'hbb6101d3),
	.w6(32'hba01fdad),
	.w7(32'hb80cae91),
	.w8(32'hbb44adcd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab90a75),
	.w1(32'h397007dc),
	.w2(32'hb9071271),
	.w3(32'h3b103bd1),
	.w4(32'h39aae6dd),
	.w5(32'hbb0a911e),
	.w6(32'h3b6f335c),
	.w7(32'h38e0e116),
	.w8(32'hbb11a2a9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27e734),
	.w1(32'hba1caea0),
	.w2(32'hb9adea37),
	.w3(32'hbb199bf8),
	.w4(32'hbaaf254e),
	.w5(32'h39844988),
	.w6(32'hbb0737e6),
	.w7(32'hbac3a8dc),
	.w8(32'h3a1ffe3d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a644c13),
	.w1(32'hbb554fb9),
	.w2(32'hbb54d67c),
	.w3(32'hba34aaf6),
	.w4(32'hbb041578),
	.w5(32'hbb90db7a),
	.w6(32'h3b189d98),
	.w7(32'h3a3a5aa4),
	.w8(32'hbb6fa082),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaa6c8),
	.w1(32'hba36509d),
	.w2(32'h3b2aff0d),
	.w3(32'hb8130e88),
	.w4(32'h3ae8eadc),
	.w5(32'h39c84896),
	.w6(32'hb8b71f8f),
	.w7(32'h3af49a07),
	.w8(32'h3a0ccbc8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6efd6e),
	.w1(32'h3a303975),
	.w2(32'hb94ddf4b),
	.w3(32'hba3bb54a),
	.w4(32'h39c24204),
	.w5(32'hbaf347b9),
	.w6(32'hba8e085e),
	.w7(32'hba063487),
	.w8(32'hba73ec54),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89ce4e),
	.w1(32'hbab4ddee),
	.w2(32'hba8a7258),
	.w3(32'hbb34eef9),
	.w4(32'hbb5cd1ef),
	.w5(32'hbb03f6f7),
	.w6(32'hbaaf206c),
	.w7(32'hbabbf437),
	.w8(32'hba0e5f69),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8f28b),
	.w1(32'hba97d6f5),
	.w2(32'hbac6e689),
	.w3(32'hbb273e87),
	.w4(32'hbb0c1f0f),
	.w5(32'hbb238076),
	.w6(32'hba0da060),
	.w7(32'hba1874f6),
	.w8(32'hba8de14e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb8550),
	.w1(32'h39eba689),
	.w2(32'h3b07d24e),
	.w3(32'hbaccc925),
	.w4(32'hbab221b5),
	.w5(32'h3bb7f44c),
	.w6(32'h393fd6d6),
	.w7(32'h39f0e793),
	.w8(32'h3ba6ab9a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46e619),
	.w1(32'hb91db4b6),
	.w2(32'hba443a01),
	.w3(32'h3833b228),
	.w4(32'hb942ae64),
	.w5(32'hba676d7f),
	.w6(32'hb6800481),
	.w7(32'hb9deea7a),
	.w8(32'hbb2d6187),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd3621),
	.w1(32'hbbc902dc),
	.w2(32'hbbc0a990),
	.w3(32'hba975ba7),
	.w4(32'h3bd395f2),
	.w5(32'h3a36de76),
	.w6(32'hbb3a77b9),
	.w7(32'h3b5f183b),
	.w8(32'h39dcf051),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fca0c),
	.w1(32'hbbc5baf0),
	.w2(32'hbb00109a),
	.w3(32'hb914a4f1),
	.w4(32'hbb64d1b9),
	.w5(32'hbb37a3e7),
	.w6(32'hbb17b8e6),
	.w7(32'hbb16a9f3),
	.w8(32'hbb9706e0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d052a8),
	.w1(32'hbac16aeb),
	.w2(32'hba88628c),
	.w3(32'hbb40d45d),
	.w4(32'hba381524),
	.w5(32'h39a40bfa),
	.w6(32'hbb22c1cf),
	.w7(32'hba38a920),
	.w8(32'hba2c3808),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c0bf77),
	.w1(32'h3a023d38),
	.w2(32'h3a3663ae),
	.w3(32'hbabace34),
	.w4(32'h38089375),
	.w5(32'h37d5e40d),
	.w6(32'hba7d8281),
	.w7(32'hb91626bf),
	.w8(32'h39f0ff65),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f0ba4),
	.w1(32'h3a49e316),
	.w2(32'h39b05a85),
	.w3(32'h3a857c74),
	.w4(32'hba425057),
	.w5(32'h39543db4),
	.w6(32'h3aea5282),
	.w7(32'h39ba4f39),
	.w8(32'h3a8e84c1),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbe836),
	.w1(32'h3a9a7037),
	.w2(32'h39ba1d02),
	.w3(32'hba7ab26f),
	.w4(32'h39350bbd),
	.w5(32'hbadf7a68),
	.w6(32'hb98ba540),
	.w7(32'h39b58526),
	.w8(32'hbaeb14f5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1f764),
	.w1(32'hb96e1153),
	.w2(32'h3a137d1c),
	.w3(32'hbb1ec8b2),
	.w4(32'h3af1b351),
	.w5(32'h3affd559),
	.w6(32'hbb0fb609),
	.w7(32'h39c60b1d),
	.w8(32'hb929d345),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad77e82),
	.w1(32'hba930286),
	.w2(32'hba31c447),
	.w3(32'h3aa940d2),
	.w4(32'h3a27e58c),
	.w5(32'hbb1adaf0),
	.w6(32'h39dee94f),
	.w7(32'hba8b4198),
	.w8(32'hbb9b9702),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a0f5),
	.w1(32'hbb45b0df),
	.w2(32'hba1e72d0),
	.w3(32'hbb2457e4),
	.w4(32'hbaaaa891),
	.w5(32'hba2ebdd1),
	.w6(32'hbb470fbe),
	.w7(32'hbb108878),
	.w8(32'hbab9ac15),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba072f0e),
	.w1(32'h3a06c02b),
	.w2(32'h3a96d595),
	.w3(32'h3a134e0c),
	.w4(32'h3a2cd9e3),
	.w5(32'hbadfbcf2),
	.w6(32'h3a3eb24a),
	.w7(32'hb90534a0),
	.w8(32'hba88e3b1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4831ac),
	.w1(32'hbbc956e5),
	.w2(32'hbbe640f3),
	.w3(32'hbb4a1b74),
	.w4(32'hbaeb8ed7),
	.w5(32'hbb3ddbec),
	.w6(32'hbb103073),
	.w7(32'hbb013b14),
	.w8(32'hbb0c9935),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09523e),
	.w1(32'hbaba5f2c),
	.w2(32'h39c6792d),
	.w3(32'hbaeb51c0),
	.w4(32'hb96d283d),
	.w5(32'h3b563dc8),
	.w6(32'hbaf69dab),
	.w7(32'hbaa2c325),
	.w8(32'h3b73d41f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b547baa),
	.w1(32'h3a97dd92),
	.w2(32'h3afe6671),
	.w3(32'h3b85fe4f),
	.w4(32'h3a04b9ad),
	.w5(32'hbac70b4a),
	.w6(32'h3b5ef4dd),
	.w7(32'h3acb5e10),
	.w8(32'h3a10f107),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9add82),
	.w1(32'h3ad09bd3),
	.w2(32'h3a19faa9),
	.w3(32'h391205d1),
	.w4(32'h39bfe197),
	.w5(32'hba847b30),
	.w6(32'h3afd9fdb),
	.w7(32'hba2e77d7),
	.w8(32'hbaa075ad),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9507bbf),
	.w1(32'hb99cb2c3),
	.w2(32'hbb038465),
	.w3(32'hb892a820),
	.w4(32'hba822191),
	.w5(32'h399d9fee),
	.w6(32'h3a11df66),
	.w7(32'hb93c5f5a),
	.w8(32'h397b11f4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a704af),
	.w1(32'hbb224de6),
	.w2(32'h39dd6a9e),
	.w3(32'hbb07371b),
	.w4(32'hb9778e5a),
	.w5(32'hb9803260),
	.w6(32'hba8ca4c5),
	.w7(32'h3a91b46d),
	.w8(32'hb9c77f86),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971a16c),
	.w1(32'h39e5fc74),
	.w2(32'h3a70216a),
	.w3(32'hb82f67d4),
	.w4(32'hbb438f65),
	.w5(32'h3a585b69),
	.w6(32'h3afe4f25),
	.w7(32'hb98a3902),
	.w8(32'hb873ff66),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4738fd),
	.w1(32'hba762663),
	.w2(32'hba04bc04),
	.w3(32'hbaa26a32),
	.w4(32'hbaac2951),
	.w5(32'hba2ea0a5),
	.w6(32'h38cb9fcf),
	.w7(32'hba0120b1),
	.w8(32'hbb3b4200),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8dc4d),
	.w1(32'hb98b5dd7),
	.w2(32'hb91ad777),
	.w3(32'hbaf84956),
	.w4(32'hba190f08),
	.w5(32'h38d9c56c),
	.w6(32'hbb4c2556),
	.w7(32'hba58e3c5),
	.w8(32'hb99b4776),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ea9e3),
	.w1(32'hbaa7e15f),
	.w2(32'hbad7097f),
	.w3(32'hb8b49918),
	.w4(32'hb8bfd3b3),
	.w5(32'hbb76becf),
	.w6(32'hb9de656a),
	.w7(32'h39a5080b),
	.w8(32'hbb8ec489),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084a27),
	.w1(32'hbb67f987),
	.w2(32'hbb82007c),
	.w3(32'hbb0af410),
	.w4(32'hba960faf),
	.w5(32'h39b5fea1),
	.w6(32'hbb1b24f7),
	.w7(32'hba4f99e1),
	.w8(32'hb8e7c9e5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb924a39),
	.w1(32'hbb5420b4),
	.w2(32'hbb947937),
	.w3(32'h3af0281d),
	.w4(32'h3b5b9c12),
	.w5(32'hbb7c93a5),
	.w6(32'h3b57f23f),
	.w7(32'h3a8ccc1f),
	.w8(32'hba9881e8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9ceb3),
	.w1(32'hba993344),
	.w2(32'hbb1824c6),
	.w3(32'h3a66698b),
	.w4(32'hb96fb073),
	.w5(32'h39484e64),
	.w6(32'h3a62017d),
	.w7(32'hb99e5cb8),
	.w8(32'h399ab699),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79b314),
	.w1(32'h3a4ff80c),
	.w2(32'h3b36a48d),
	.w3(32'h3adec70e),
	.w4(32'h38c06dbd),
	.w5(32'h3b1448eb),
	.w6(32'h3b17f2b9),
	.w7(32'h3ab15cc7),
	.w8(32'h3ae6c907),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66f5ae),
	.w1(32'h3ae6e8b2),
	.w2(32'h3afc1237),
	.w3(32'hbb716943),
	.w4(32'hbad1453d),
	.w5(32'hbae92f65),
	.w6(32'hb9c8d61e),
	.w7(32'hb8fb66e6),
	.w8(32'hbac9ecb7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bddd7),
	.w1(32'h3ab7d8c4),
	.w2(32'hb9fdc73f),
	.w3(32'h3b836e14),
	.w4(32'h3b03d8eb),
	.w5(32'hba8e1acc),
	.w6(32'h3ba943d3),
	.w7(32'h3b117bc7),
	.w8(32'hbaedbeb2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080baa),
	.w1(32'hbb58f548),
	.w2(32'hbb87a836),
	.w3(32'hbb359bce),
	.w4(32'hbb64079d),
	.w5(32'hbb6007fd),
	.w6(32'hbb203db1),
	.w7(32'hbafa9552),
	.w8(32'hbb2919e4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb196e21),
	.w1(32'hbb537073),
	.w2(32'hbb27a7f8),
	.w3(32'hbbc86959),
	.w4(32'hbb22fc79),
	.w5(32'hbadebc34),
	.w6(32'h39e7ad6c),
	.w7(32'h3ae12e67),
	.w8(32'hbb6ef1c3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27b45b),
	.w1(32'hb9203314),
	.w2(32'hb910c3de),
	.w3(32'hba44da5c),
	.w4(32'h38f5bae8),
	.w5(32'hbac09e82),
	.w6(32'hba598fa8),
	.w7(32'hb972008e),
	.w8(32'hbb163057),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884ba7),
	.w1(32'hbad80479),
	.w2(32'hbae356a7),
	.w3(32'hbaa50416),
	.w4(32'hbae2e328),
	.w5(32'hbaa2a467),
	.w6(32'hbaffb884),
	.w7(32'hbae5c08c),
	.w8(32'hb9646fff),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7949f7),
	.w1(32'h3b88d026),
	.w2(32'h3bd41b38),
	.w3(32'h3b3eeec6),
	.w4(32'h3b950cba),
	.w5(32'h3c20cdc2),
	.w6(32'h3ad55e2b),
	.w7(32'h3bbdbe84),
	.w8(32'h3baed725),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ec288),
	.w1(32'hb9b5797c),
	.w2(32'hbb5ea331),
	.w3(32'hba0ba737),
	.w4(32'h3bda5bc4),
	.w5(32'hbb6c5dd0),
	.w6(32'h3ac11566),
	.w7(32'h3ab3729f),
	.w8(32'hbba08233),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ea5cc),
	.w1(32'hba3f5f63),
	.w2(32'hba6403ba),
	.w3(32'hb99d4f26),
	.w4(32'h3a2a38aa),
	.w5(32'hbb1e28d0),
	.w6(32'h3a792564),
	.w7(32'h3a38b7d0),
	.w8(32'hbb8c1082),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b873b),
	.w1(32'hbb87ff69),
	.w2(32'hbb46d205),
	.w3(32'hbb888db6),
	.w4(32'hbb8618b4),
	.w5(32'h3947c37d),
	.w6(32'hbba8f39b),
	.w7(32'hbb65fbd3),
	.w8(32'h3a820b46),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e2d38),
	.w1(32'hba984fa2),
	.w2(32'h3abea722),
	.w3(32'h391c91b4),
	.w4(32'hbac08467),
	.w5(32'hb99b62a0),
	.w6(32'h3a674e51),
	.w7(32'h3a56927d),
	.w8(32'h3ac17d97),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9582311),
	.w1(32'h3aaeca36),
	.w2(32'hb8e41d02),
	.w3(32'h39d00ec8),
	.w4(32'hb9834704),
	.w5(32'hbb1e0981),
	.w6(32'h3b1c4f94),
	.w7(32'h3a1c60a0),
	.w8(32'hbad39fa4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab549da),
	.w1(32'h394f4b82),
	.w2(32'h3b3860a9),
	.w3(32'hba8dda44),
	.w4(32'h3929b3cf),
	.w5(32'h3a5506da),
	.w6(32'h39dcfe6d),
	.w7(32'h3ad0c767),
	.w8(32'h3adbac00),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199f5e),
	.w1(32'h3b04bbf5),
	.w2(32'h3a624734),
	.w3(32'h399f99d6),
	.w4(32'h3b3b16fb),
	.w5(32'h393a4529),
	.w6(32'h3a3a55de),
	.w7(32'h3b37e33a),
	.w8(32'hbb1b27d9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01df6a),
	.w1(32'h38804489),
	.w2(32'hbaa13968),
	.w3(32'hba9e0826),
	.w4(32'h3a0e908d),
	.w5(32'hba09bbed),
	.w6(32'h3a7c806d),
	.w7(32'h3a4cf085),
	.w8(32'hba260ea4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10eebb),
	.w1(32'hb98af91d),
	.w2(32'h3aa142c0),
	.w3(32'hba2884a1),
	.w4(32'h3a5c0321),
	.w5(32'h3aa4506b),
	.w6(32'hba516a16),
	.w7(32'h3a3e5080),
	.w8(32'h3a078ad0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da600e),
	.w1(32'hb87f6d2e),
	.w2(32'hbab3b7b7),
	.w3(32'h3915533a),
	.w4(32'h3abb7ca6),
	.w5(32'hbacfedfe),
	.w6(32'h38d689c6),
	.w7(32'h3a0c3550),
	.w8(32'hbb2e0cee),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbc044),
	.w1(32'hbb0f902b),
	.w2(32'hbadb936b),
	.w3(32'hba61e33a),
	.w4(32'hba5e1fc3),
	.w5(32'h3a03b187),
	.w6(32'hbae8b81a),
	.w7(32'hbaa2c509),
	.w8(32'h3a1567d3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab966cc),
	.w1(32'h3ab17a5a),
	.w2(32'h3a58f49e),
	.w3(32'h3a82a5bf),
	.w4(32'h3a45f5d6),
	.w5(32'h39d3d787),
	.w6(32'h3a30568e),
	.w7(32'h3a2b0715),
	.w8(32'h39b5ed48),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a6c5b),
	.w1(32'h3af92c0e),
	.w2(32'h3b0475b6),
	.w3(32'hbaece704),
	.w4(32'h3b20410d),
	.w5(32'h3b2f4f77),
	.w6(32'h3a285529),
	.w7(32'h3b78c133),
	.w8(32'h38fae47d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba122069),
	.w1(32'hba6b0e3f),
	.w2(32'hbb175661),
	.w3(32'h38e84698),
	.w4(32'h3a1650d3),
	.w5(32'h3850cee0),
	.w6(32'h3a435cb9),
	.w7(32'h3954f508),
	.w8(32'hbacf3372),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815dc72),
	.w1(32'h38e05547),
	.w2(32'h385b9208),
	.w3(32'hb8e7f4bd),
	.w4(32'hb9be3f7d),
	.w5(32'h395480de),
	.w6(32'hb977d5b4),
	.w7(32'hba0b4f8a),
	.w8(32'h3a283fdd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a527e3f),
	.w1(32'h39a9eb9f),
	.w2(32'hba9aba81),
	.w3(32'hb99d4bc1),
	.w4(32'h39ed815d),
	.w5(32'hba77c11e),
	.w6(32'h3a20c6d7),
	.w7(32'h3a8808a8),
	.w8(32'hbab45dd6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2ae4f),
	.w1(32'hb9d8fb5c),
	.w2(32'h39968fc6),
	.w3(32'hba88fd95),
	.w4(32'hba0ab8b1),
	.w5(32'h396ab93e),
	.w6(32'hba95a356),
	.w7(32'hb99759d6),
	.w8(32'h39c9c8de),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f34666),
	.w1(32'hb9987890),
	.w2(32'hb9db3f6e),
	.w3(32'hb8f74c82),
	.w4(32'hb9c3935f),
	.w5(32'hba1b6abd),
	.w6(32'h391338c1),
	.w7(32'hb88aca87),
	.w8(32'hba500009),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f97673),
	.w1(32'hb9f2bbd9),
	.w2(32'h3997f6ea),
	.w3(32'hb93f771d),
	.w4(32'h399fac95),
	.w5(32'h3996cd53),
	.w6(32'hb9f8be97),
	.w7(32'hb8221c12),
	.w8(32'h39f2cd7c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a018b83),
	.w1(32'h39a15806),
	.w2(32'h3a2e7b0a),
	.w3(32'hb7f62f2c),
	.w4(32'h39251a4a),
	.w5(32'h3951bce5),
	.w6(32'hb82fa1cc),
	.w7(32'h399baefd),
	.w8(32'hb826f0dd),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9866f2),
	.w1(32'hba271c27),
	.w2(32'hb966d5ec),
	.w3(32'hba0c2338),
	.w4(32'hba4b4e55),
	.w5(32'h3a8023c3),
	.w6(32'hba410564),
	.w7(32'hba10fe14),
	.w8(32'h3ab01eb4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ef830),
	.w1(32'hbb7d93d6),
	.w2(32'hbbc7d54b),
	.w3(32'h3ab107d4),
	.w4(32'h3ab049a6),
	.w5(32'hbb5e477f),
	.w6(32'h3b266b76),
	.w7(32'h3afbcbd2),
	.w8(32'hbb5bf585),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29de7c),
	.w1(32'h3b0f765c),
	.w2(32'hba8906ae),
	.w3(32'h3b23e4df),
	.w4(32'h3b71c721),
	.w5(32'hba598901),
	.w6(32'h3ae98e47),
	.w7(32'h3b201ab2),
	.w8(32'hba05fc8c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69e5fc),
	.w1(32'hb9fc603a),
	.w2(32'hbb0e636e),
	.w3(32'h37111695),
	.w4(32'h3ad0d2e2),
	.w5(32'hbb4266c8),
	.w6(32'h3ae1850d),
	.w7(32'h3b605e76),
	.w8(32'hbb1c08bd),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8636e3),
	.w1(32'h39e0af94),
	.w2(32'hb9bb58b7),
	.w3(32'hba72b418),
	.w4(32'hbaccfa21),
	.w5(32'h3b030ab9),
	.w6(32'hb993983e),
	.w7(32'hba91aa2e),
	.w8(32'h3ac46f1a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a958675),
	.w1(32'h3a1bea26),
	.w2(32'h38a297a0),
	.w3(32'h3af2bf2a),
	.w4(32'h3a91bd0a),
	.w5(32'h396562f1),
	.w6(32'h3adb0767),
	.w7(32'h3a239504),
	.w8(32'h39d724c7),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03d17f),
	.w1(32'h3958313e),
	.w2(32'hb8e5e93a),
	.w3(32'hb867785a),
	.w4(32'hb9de3cbb),
	.w5(32'h36b2332c),
	.w6(32'hb7f296fa),
	.w7(32'hb9d9ff63),
	.w8(32'hb988b9e6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9857db3),
	.w1(32'hba21d15f),
	.w2(32'hb9562b6a),
	.w3(32'hb9a7ec29),
	.w4(32'h39053c47),
	.w5(32'hba11aeb8),
	.w6(32'hb98a8cab),
	.w7(32'h3863635e),
	.w8(32'hb99e382e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb1dc8),
	.w1(32'hb9bf4b69),
	.w2(32'hbab0a50b),
	.w3(32'h3b0bb3fb),
	.w4(32'h3a7027a6),
	.w5(32'hbb9f76b6),
	.w6(32'h3b0039b4),
	.w7(32'h3a7fc02c),
	.w8(32'hbbb40f07),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2543a),
	.w1(32'hbab5a281),
	.w2(32'hb9fc69f2),
	.w3(32'hbaa3c948),
	.w4(32'hba0cf6fb),
	.w5(32'h39f39b89),
	.w6(32'hbab32f63),
	.w7(32'hba23c3bd),
	.w8(32'hb78ead82),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cbab0),
	.w1(32'hbadbed8b),
	.w2(32'hbad6d529),
	.w3(32'hb953209b),
	.w4(32'hba9e3a47),
	.w5(32'hb902f8cf),
	.w6(32'h38b0aaa1),
	.w7(32'hbafdc45a),
	.w8(32'hb99086f0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afae51a),
	.w1(32'h3b11e4cb),
	.w2(32'h3ab23159),
	.w3(32'h3b105176),
	.w4(32'h3a970107),
	.w5(32'h3a9263f2),
	.w6(32'h3b250d32),
	.w7(32'h39ddf56e),
	.w8(32'h39d76811),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9271f4d),
	.w1(32'hba04a342),
	.w2(32'hba1f0d2f),
	.w3(32'h3a973e9d),
	.w4(32'h3a4b2768),
	.w5(32'h3927ceb7),
	.w6(32'h397e3d7e),
	.w7(32'h395864a1),
	.w8(32'h39c4b82c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ac6ed),
	.w1(32'h394a7e6e),
	.w2(32'hb98f6cdf),
	.w3(32'hb9d71379),
	.w4(32'h39059bab),
	.w5(32'hb9f7d481),
	.w6(32'h399d0310),
	.w7(32'h38cebf3f),
	.w8(32'h38b0f97c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dca897),
	.w1(32'hb9b3c703),
	.w2(32'hb833e528),
	.w3(32'h3a97e225),
	.w4(32'h3a4e9c71),
	.w5(32'hb86ac15b),
	.w6(32'h3ad5d008),
	.w7(32'h3abfc273),
	.w8(32'h396d55a8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7e521),
	.w1(32'hba857127),
	.w2(32'hbb29b27f),
	.w3(32'h3ad85bed),
	.w4(32'hbabe5007),
	.w5(32'hbbc72fc4),
	.w6(32'h3b11a02a),
	.w7(32'h39f4481e),
	.w8(32'hbc1da9a5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942eeb9),
	.w1(32'h39cb9776),
	.w2(32'h3a3d4c73),
	.w3(32'h3858b598),
	.w4(32'h39be8dea),
	.w5(32'hba041a01),
	.w6(32'hb816cc9d),
	.w7(32'h3a21e636),
	.w8(32'h39bd1026),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9852d1),
	.w1(32'h3b5433d3),
	.w2(32'h3a6736ae),
	.w3(32'hb9c96f95),
	.w4(32'hbada8c4d),
	.w5(32'h39144c10),
	.w6(32'h358aebaa),
	.w7(32'hbb05b162),
	.w8(32'h3986f6d5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule