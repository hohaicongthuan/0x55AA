module layer_8_featuremap_213(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b2fa4),
	.w1(32'h3ba0b760),
	.w2(32'h3a1f402d),
	.w3(32'h3c07155a),
	.w4(32'h3aa40e0e),
	.w5(32'h3c419b16),
	.w6(32'h3b1a3ed9),
	.w7(32'h3c48f09d),
	.w8(32'hbb623e83),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94fde8),
	.w1(32'h3bc5a605),
	.w2(32'h3b27a204),
	.w3(32'h3c3a2504),
	.w4(32'h3bb91ec3),
	.w5(32'h3aeed77f),
	.w6(32'h3b5558c2),
	.w7(32'h3a2707cb),
	.w8(32'hbba14691),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42e979),
	.w1(32'h3a0cf199),
	.w2(32'hbc06246f),
	.w3(32'hbc004ca2),
	.w4(32'h3c1255e9),
	.w5(32'h3b195776),
	.w6(32'h3af58552),
	.w7(32'hbba3ec6f),
	.w8(32'h39113e0f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27f6aa),
	.w1(32'hbcbc0aa1),
	.w2(32'hbc1bd56c),
	.w3(32'h3bb55a33),
	.w4(32'hbbaa253a),
	.w5(32'hbb4d90d3),
	.w6(32'hbba1d50d),
	.w7(32'h3933a0b2),
	.w8(32'h3be4c9cd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d217),
	.w1(32'hbc452a5f),
	.w2(32'hbb511a9a),
	.w3(32'h3bee67b5),
	.w4(32'hbc0d7fb9),
	.w5(32'hbb41e7d4),
	.w6(32'hbb8f78df),
	.w7(32'hbb894889),
	.w8(32'hbb5303d4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55742c),
	.w1(32'h3d50ca6e),
	.w2(32'h3c14c741),
	.w3(32'h3c1b0877),
	.w4(32'h3cd3a0d9),
	.w5(32'hbc95ed65),
	.w6(32'h3cdb20cc),
	.w7(32'h3c8603fd),
	.w8(32'hbac74dcd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb18be7),
	.w1(32'hbc0121ad),
	.w2(32'hba140978),
	.w3(32'hbc302e6f),
	.w4(32'hbbb635c9),
	.w5(32'hba8c6733),
	.w6(32'hbb79ca32),
	.w7(32'hbb31ab8f),
	.w8(32'h3aa4ea14),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095b3d),
	.w1(32'hbc0e4e27),
	.w2(32'h3ac8e1a3),
	.w3(32'h3b88b5be),
	.w4(32'hbc8c62ed),
	.w5(32'h3afbff45),
	.w6(32'hbb2ff746),
	.w7(32'hbbee6888),
	.w8(32'hbc228e5c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc043e9),
	.w1(32'hbc48a89c),
	.w2(32'h3b014a38),
	.w3(32'h3bbcddbc),
	.w4(32'hbc110d24),
	.w5(32'h39f920f4),
	.w6(32'hbb337cc6),
	.w7(32'hba628e9b),
	.w8(32'h3c3bcce0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3bbcf),
	.w1(32'hbc042d6b),
	.w2(32'hbb23ab36),
	.w3(32'h3c93b09f),
	.w4(32'hbbcf8675),
	.w5(32'hbb987acf),
	.w6(32'h3bcfa2fb),
	.w7(32'h3b694f08),
	.w8(32'hbc2df323),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf48dac),
	.w1(32'h3c80e596),
	.w2(32'hbb130e71),
	.w3(32'hb8f2deec),
	.w4(32'h3c82fe4c),
	.w5(32'h3bf0f72b),
	.w6(32'h3c01cab5),
	.w7(32'hba7653ae),
	.w8(32'hbc50c415),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc85332),
	.w1(32'h3bba92e1),
	.w2(32'hbb1b7f41),
	.w3(32'hbc39a6aa),
	.w4(32'h3be9a613),
	.w5(32'hb95fa6ca),
	.w6(32'h3b8e6258),
	.w7(32'hbbc4c3a3),
	.w8(32'hb98ef5ae),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd211e),
	.w1(32'hbc0c8a1b),
	.w2(32'hbbeb3e46),
	.w3(32'h3be347fe),
	.w4(32'h3bab65cb),
	.w5(32'hba9210df),
	.w6(32'h3ab29f8e),
	.w7(32'h3b3c7df2),
	.w8(32'hba228520),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084b1f),
	.w1(32'h3b1ed23c),
	.w2(32'hbbfc87b0),
	.w3(32'hba64d0f7),
	.w4(32'h391d0419),
	.w5(32'hb72c79dd),
	.w6(32'hbb3b58d0),
	.w7(32'hbbc27f9e),
	.w8(32'hbc22f923),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92591b),
	.w1(32'hbb807c59),
	.w2(32'hbaa089ec),
	.w3(32'h3b8f45a3),
	.w4(32'hbade821c),
	.w5(32'hb9af0b94),
	.w6(32'h3a897209),
	.w7(32'hbac1eb7b),
	.w8(32'h3c5a8fb6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafb575),
	.w1(32'h3c8d2c5c),
	.w2(32'hbc75196b),
	.w3(32'h3c725c95),
	.w4(32'h3c2cdeed),
	.w5(32'hbbcf6dd9),
	.w6(32'h3c09a77c),
	.w7(32'hbbc07991),
	.w8(32'hbb5ea368),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede076),
	.w1(32'hbb601c8e),
	.w2(32'hbac37726),
	.w3(32'h39cd37f3),
	.w4(32'h39cb7cf5),
	.w5(32'h3b412bfe),
	.w6(32'h3ba035ff),
	.w7(32'hbb660752),
	.w8(32'h3c30581d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e59a5),
	.w1(32'h3a7faf6a),
	.w2(32'hbc906b04),
	.w3(32'h39fc5847),
	.w4(32'hba95bfaa),
	.w5(32'hbc67fabf),
	.w6(32'hbb31e845),
	.w7(32'hbc9c35ec),
	.w8(32'hbc2e0538),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce36d0b),
	.w1(32'hbb33fee6),
	.w2(32'h3c78ec3e),
	.w3(32'hbc57edd3),
	.w4(32'h3c471291),
	.w5(32'h3ca966d8),
	.w6(32'hbad4e0f8),
	.w7(32'h3c0d3d6e),
	.w8(32'h3a58896c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c450154),
	.w1(32'h389732b3),
	.w2(32'h392f4931),
	.w3(32'hbb89b1c9),
	.w4(32'hbabf5ab1),
	.w5(32'hbb3f1a74),
	.w6(32'h3ba39e58),
	.w7(32'h3a0dbf6d),
	.w8(32'h3b8c519a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c247184),
	.w1(32'h3b8e136f),
	.w2(32'hbc6c2e24),
	.w3(32'h3b764063),
	.w4(32'hbc0c8f13),
	.w5(32'hbc79c9d0),
	.w6(32'hba14186d),
	.w7(32'h3bf9a5e9),
	.w8(32'hbba2e88a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc546c8c),
	.w1(32'hbab754b5),
	.w2(32'hbbc03dc8),
	.w3(32'hbbf7aeac),
	.w4(32'h382e8b9c),
	.w5(32'hbba500f4),
	.w6(32'h3922d137),
	.w7(32'hbb1f8adc),
	.w8(32'hbbc9cb84),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb381241),
	.w1(32'hbc2f2c37),
	.w2(32'hbaa9f548),
	.w3(32'hbc3d175e),
	.w4(32'hbc0b5457),
	.w5(32'hbbbdfb5a),
	.w6(32'hbc0aea17),
	.w7(32'h3c500edd),
	.w8(32'hbb9b3cdb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ca4b1),
	.w1(32'h3baaba00),
	.w2(32'hbbe0c0aa),
	.w3(32'hbc4fc9f3),
	.w4(32'hbc5ff843),
	.w5(32'hbc22a706),
	.w6(32'h3a23e12a),
	.w7(32'hbc16a0a7),
	.w8(32'hbc451687),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a929),
	.w1(32'hbc580062),
	.w2(32'hbbfab941),
	.w3(32'h3b0d9f45),
	.w4(32'h3bad3c55),
	.w5(32'hba1581a3),
	.w6(32'hbc428ae2),
	.w7(32'h3a1aae30),
	.w8(32'h3bb1af49),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5c8f8),
	.w1(32'h3b950eb2),
	.w2(32'hbac4c016),
	.w3(32'hbb2069ff),
	.w4(32'h3c2e4258),
	.w5(32'h3c6a1db5),
	.w6(32'h3c161829),
	.w7(32'h3b02f4f6),
	.w8(32'h3a78724d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07204d),
	.w1(32'h3b89e146),
	.w2(32'hba0f21bc),
	.w3(32'h3a3983c9),
	.w4(32'h3acba133),
	.w5(32'hbc0f0d4c),
	.w6(32'h3bfe5546),
	.w7(32'h3a91b6f3),
	.w8(32'h3bd6d477),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd218b45),
	.w1(32'hbd24bf8f),
	.w2(32'hbd6d069e),
	.w3(32'hbd092b51),
	.w4(32'hbd7c62f3),
	.w5(32'hbcfa30b7),
	.w6(32'hbce2c8e2),
	.w7(32'h3c6e2bfc),
	.w8(32'h3d83435f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa8b34),
	.w1(32'h3c957ee6),
	.w2(32'hbd0158c5),
	.w3(32'h3c9d4a3c),
	.w4(32'h3c3ae55c),
	.w5(32'hbcc11a33),
	.w6(32'h3ca1129d),
	.w7(32'hbc1a8242),
	.w8(32'hbbdb135d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc508fcc),
	.w1(32'h3ae61918),
	.w2(32'hba691685),
	.w3(32'hbb123df5),
	.w4(32'h3af0cab6),
	.w5(32'hb9ef3e48),
	.w6(32'h3ab47bc6),
	.w7(32'h3970b089),
	.w8(32'h3b48081b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c146a61),
	.w1(32'h3a35db3e),
	.w2(32'hbc9468c5),
	.w3(32'h3c124cc2),
	.w4(32'hbc412237),
	.w5(32'hbbfc06b2),
	.w6(32'h3c14e726),
	.w7(32'hbb539da8),
	.w8(32'hbc9632e1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc139bcf),
	.w1(32'h3c21e188),
	.w2(32'hb99781ee),
	.w3(32'h3c2f9a5b),
	.w4(32'h3bc85db0),
	.w5(32'h3a906e49),
	.w6(32'h3bbb2acd),
	.w7(32'hbaf27215),
	.w8(32'hbb3dfa4b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc525141),
	.w1(32'hba4ab6e2),
	.w2(32'h3b86aa57),
	.w3(32'hbc3a2d48),
	.w4(32'hba7d3603),
	.w5(32'h3adc16ff),
	.w6(32'hbb9aea35),
	.w7(32'h3a536cf5),
	.w8(32'h394c939b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c694049),
	.w1(32'hbb526149),
	.w2(32'hbae30628),
	.w3(32'h3bb06bb3),
	.w4(32'hb901aa5a),
	.w5(32'hbb320d85),
	.w6(32'hbb8f0a14),
	.w7(32'hbb76d610),
	.w8(32'hba308665),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae01ff3),
	.w1(32'hbc04a3e7),
	.w2(32'hbbded30c),
	.w3(32'h39611d3d),
	.w4(32'h3aee65bd),
	.w5(32'h3b1eea0c),
	.w6(32'hbb614b4b),
	.w7(32'hbbe087bf),
	.w8(32'hba4e4fe8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dadbe),
	.w1(32'hbc1ce286),
	.w2(32'hbc1b062f),
	.w3(32'h3be89ebc),
	.w4(32'hbb64ef6f),
	.w5(32'h3878f03b),
	.w6(32'hbb030a21),
	.w7(32'hb94119e1),
	.w8(32'h3b2d9fdb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba181b8e),
	.w1(32'hbbf30daa),
	.w2(32'hbc9cfcc6),
	.w3(32'hb9c11806),
	.w4(32'hbb98cd35),
	.w5(32'hbc9c13c2),
	.w6(32'hbb5feee6),
	.w7(32'hbc4ccf33),
	.w8(32'h3a8562c8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb668d1b),
	.w1(32'hbbf87b08),
	.w2(32'hbb629e7b),
	.w3(32'hbbead778),
	.w4(32'hbbbde7cb),
	.w5(32'hbb55af7e),
	.w6(32'hbad7770c),
	.w7(32'hbb260489),
	.w8(32'h3c3b3b99),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97ad0d),
	.w1(32'h38c92dc7),
	.w2(32'hbc20eaf9),
	.w3(32'h3c430d83),
	.w4(32'hbaa735a9),
	.w5(32'hbbe1982b),
	.w6(32'h39617cdc),
	.w7(32'hbc19f662),
	.w8(32'hbc252072),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc454381),
	.w1(32'hbb13a22e),
	.w2(32'hbaedccdd),
	.w3(32'hbc5f16f7),
	.w4(32'hbb8cedea),
	.w5(32'hbc138624),
	.w6(32'hbc1c3b71),
	.w7(32'hbb47cbd9),
	.w8(32'h3a3ab88e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc1822),
	.w1(32'h3bd253e0),
	.w2(32'hba38f5a3),
	.w3(32'hbb694c8a),
	.w4(32'h3c07ebf3),
	.w5(32'hbbbd66bd),
	.w6(32'h3c584193),
	.w7(32'h3b86522c),
	.w8(32'hbb46c919),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bec13),
	.w1(32'h3c337f8e),
	.w2(32'h3d454ac2),
	.w3(32'hba4696bc),
	.w4(32'h3bc0fa83),
	.w5(32'h3d005623),
	.w6(32'hbaf7751a),
	.w7(32'h3cc64cee),
	.w8(32'h3b66d26f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba545de9),
	.w1(32'hbbe9a269),
	.w2(32'hbcf5f880),
	.w3(32'hbb02d226),
	.w4(32'h3b6f57ae),
	.w5(32'hbc732fa7),
	.w6(32'hbb287349),
	.w7(32'hbc8ce3dc),
	.w8(32'hba812f46),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb0c02),
	.w1(32'h3aea9f07),
	.w2(32'hbc78fc01),
	.w3(32'hba6d3641),
	.w4(32'h3b2caaf4),
	.w5(32'hbc2f2227),
	.w6(32'h3b5eb525),
	.w7(32'hbb78f13e),
	.w8(32'hbbd0f316),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4a68),
	.w1(32'hbc81824c),
	.w2(32'hbbdf0a48),
	.w3(32'hbbcd7084),
	.w4(32'hbc4d191e),
	.w5(32'hbc00e912),
	.w6(32'hbbb63ca7),
	.w7(32'hba7a0cb4),
	.w8(32'h3c9e1525),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1a958),
	.w1(32'hbc17dba9),
	.w2(32'h39d3722e),
	.w3(32'h3ad9d57c),
	.w4(32'hba4f7628),
	.w5(32'h3bc3ba98),
	.w6(32'hbbcf2924),
	.w7(32'h3a212407),
	.w8(32'h3a869bee),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1356cb),
	.w1(32'hba7c449c),
	.w2(32'hbc87f683),
	.w3(32'hb88c5166),
	.w4(32'h3b5875c5),
	.w5(32'hbc465f30),
	.w6(32'hbb46da5a),
	.w7(32'hbc13d6fc),
	.w8(32'hbb3c1d77),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff4a6),
	.w1(32'h3bf405e6),
	.w2(32'hbbdfb93a),
	.w3(32'h3b6bb619),
	.w4(32'hbbdafa3a),
	.w5(32'hbbb3c140),
	.w6(32'h3b6f70f1),
	.w7(32'h3bdaca63),
	.w8(32'h3c0256ba),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb264d53),
	.w1(32'hbb8086df),
	.w2(32'hbc8ff8c0),
	.w3(32'hbb083e6a),
	.w4(32'hbc1ff2db),
	.w5(32'hbc616a3d),
	.w6(32'h3bb6fe34),
	.w7(32'hbb8e34cb),
	.w8(32'h3a25f8d6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cbdbe),
	.w1(32'h3cfac16b),
	.w2(32'hbbc9d805),
	.w3(32'h3ba9d837),
	.w4(32'h3cc16806),
	.w5(32'h3b50d11c),
	.w6(32'h3cad6815),
	.w7(32'hbc276145),
	.w8(32'h3b2eaa8c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e37a1),
	.w1(32'hba1072e0),
	.w2(32'hbb50c856),
	.w3(32'hbb099dc1),
	.w4(32'h3b5baa63),
	.w5(32'h3b432877),
	.w6(32'h3b512e0d),
	.w7(32'h3b1214b7),
	.w8(32'h3b9173c9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf8f4a),
	.w1(32'h3b96c302),
	.w2(32'h3ca44070),
	.w3(32'hbbccca32),
	.w4(32'hbc27c6e1),
	.w5(32'h391980bf),
	.w6(32'h3acc0f79),
	.w7(32'h3c171ee4),
	.w8(32'hbbc12047),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34acf),
	.w1(32'hb9825b6e),
	.w2(32'hbbc807b8),
	.w3(32'hbadab0e9),
	.w4(32'hbba3ac0a),
	.w5(32'hbbee8250),
	.w6(32'h3b274442),
	.w7(32'hbbac046a),
	.w8(32'hbb34836d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e335a),
	.w1(32'h3b83d1db),
	.w2(32'h3b63e565),
	.w3(32'hbb913a93),
	.w4(32'h3a1ae0a5),
	.w5(32'h3b16fa88),
	.w6(32'h3bf93beb),
	.w7(32'h3bded9d4),
	.w8(32'h39d3266e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9285eb),
	.w1(32'hbcbd65e0),
	.w2(32'h393ff71e),
	.w3(32'hbb1ea923),
	.w4(32'hbc959a00),
	.w5(32'hbbab8cd6),
	.w6(32'hbc769437),
	.w7(32'h3b30beeb),
	.w8(32'hbbb1d28c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc259651),
	.w1(32'hbb4aebcf),
	.w2(32'hbc055496),
	.w3(32'h3a0ae242),
	.w4(32'h39f5611e),
	.w5(32'hbc1bce62),
	.w6(32'hbad86590),
	.w7(32'hbc0f2a12),
	.w8(32'hbb99c0c0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2480e0),
	.w1(32'hbbac9807),
	.w2(32'hbc3824c7),
	.w3(32'hbbf8b196),
	.w4(32'hbb69a5eb),
	.w5(32'h3bfbc776),
	.w6(32'h3b8246a2),
	.w7(32'hbc4cfc37),
	.w8(32'h3ca9d0f7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4246a3),
	.w1(32'hbc0017cb),
	.w2(32'hbcfda3cf),
	.w3(32'h3d15989a),
	.w4(32'hbb9f9afc),
	.w5(32'hbcec1a73),
	.w6(32'h3a7df3d3),
	.w7(32'hbc983a91),
	.w8(32'h3af69ed7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af012f5),
	.w1(32'hbbafaed3),
	.w2(32'hbbf582e3),
	.w3(32'h3b238605),
	.w4(32'hbbfefc13),
	.w5(32'hbc0507c6),
	.w6(32'hbb861766),
	.w7(32'hbac3e9aa),
	.w8(32'hbb405ebb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7495fc),
	.w1(32'h3b2a08b9),
	.w2(32'hbc5f21e7),
	.w3(32'hbbcc3183),
	.w4(32'hbad8aa78),
	.w5(32'hbc47beab),
	.w6(32'hba7399a2),
	.w7(32'hbae64b13),
	.w8(32'hbc14685e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbdd89),
	.w1(32'hba8f5573),
	.w2(32'hba82db81),
	.w3(32'hbb0e685a),
	.w4(32'hbb8f264e),
	.w5(32'hbbda1747),
	.w6(32'h3b6d3904),
	.w7(32'h3b89cefb),
	.w8(32'h3c6dcd14),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ebc80),
	.w1(32'hbbd90f99),
	.w2(32'h3baebdf4),
	.w3(32'h3b204ed5),
	.w4(32'h3aa9b768),
	.w5(32'h3b594e04),
	.w6(32'hbbfb35e7),
	.w7(32'h3acfc9b8),
	.w8(32'h3c4115be),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f4a95),
	.w1(32'h3c81a545),
	.w2(32'h3a5bf3a9),
	.w3(32'hbc0c40e7),
	.w4(32'h3c521a45),
	.w5(32'hbb54eeb1),
	.w6(32'h3c55b281),
	.w7(32'hbaf4beda),
	.w8(32'hbc9c4f24),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf1302),
	.w1(32'hbb072d44),
	.w2(32'hbb961764),
	.w3(32'hbc8dedc4),
	.w4(32'h3a94784d),
	.w5(32'hb9cf0e3e),
	.w6(32'h3ae8fb2e),
	.w7(32'hbb27ea03),
	.w8(32'hbae1051f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4333f),
	.w1(32'h3c6aed6a),
	.w2(32'hba381abb),
	.w3(32'h3b1b3516),
	.w4(32'h3c306ba5),
	.w5(32'hba71fa56),
	.w6(32'h3c138843),
	.w7(32'h3b11eb4c),
	.w8(32'hbbbcc3b7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35b68d),
	.w1(32'hbb01b6a0),
	.w2(32'hb9baf110),
	.w3(32'hbbbcb278),
	.w4(32'hbac0d665),
	.w5(32'hbbcadf42),
	.w6(32'hba45ea84),
	.w7(32'hbb107e68),
	.w8(32'hbad95591),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba461354),
	.w1(32'hbb136557),
	.w2(32'h3c178f4c),
	.w3(32'hbb8b93a2),
	.w4(32'h3b425930),
	.w5(32'h3b69f7ec),
	.w6(32'h3b8b93ac),
	.w7(32'h3c1c442e),
	.w8(32'h3c67c9b7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63b93a),
	.w1(32'hbc35a4b9),
	.w2(32'hbb37ed11),
	.w3(32'h3c099e73),
	.w4(32'hbbfff3f8),
	.w5(32'hbb8299d6),
	.w6(32'h38628c9b),
	.w7(32'hbba48015),
	.w8(32'hbb66da0a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3a125),
	.w1(32'h3c0aacb1),
	.w2(32'hbbb06454),
	.w3(32'hbc057a56),
	.w4(32'h3b5877c8),
	.w5(32'h394c3f08),
	.w6(32'h3b54183c),
	.w7(32'h3ba95505),
	.w8(32'hbb4da934),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bf77a),
	.w1(32'hbb564a7e),
	.w2(32'hbcab0195),
	.w3(32'hbb42b9c7),
	.w4(32'hbbd0dc4c),
	.w5(32'hbc1711e1),
	.w6(32'h3babcf88),
	.w7(32'h3b9a3a9a),
	.w8(32'h3c64dc4a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd91e7a),
	.w1(32'hb8c7f9d9),
	.w2(32'h3cf0b96f),
	.w3(32'h3c14d462),
	.w4(32'h3adcb623),
	.w5(32'h3ccb67f1),
	.w6(32'h388555a4),
	.w7(32'h3c05b942),
	.w8(32'hbb11ef82),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf341fb),
	.w1(32'hbba50d99),
	.w2(32'hbb271e35),
	.w3(32'h3b83737e),
	.w4(32'hbc5c7dfa),
	.w5(32'hbc230706),
	.w6(32'hbb5d40ab),
	.w7(32'hbb90d9ec),
	.w8(32'hba897f5f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c105be8),
	.w1(32'h38834674),
	.w2(32'hbb711f0c),
	.w3(32'hbaa59eb8),
	.w4(32'hba92ad1e),
	.w5(32'h39860928),
	.w6(32'h3b6221dd),
	.w7(32'hbafd92f7),
	.w8(32'h3b187a72),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb7ac),
	.w1(32'hbb9a232c),
	.w2(32'hbd16bc8f),
	.w3(32'h3bd7d5a5),
	.w4(32'hbb0b3740),
	.w5(32'hbca91cfb),
	.w6(32'h3b14c289),
	.w7(32'hbc8b9ab5),
	.w8(32'hbbbb3ebc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc140215),
	.w1(32'h3aa9a0fc),
	.w2(32'h3c119487),
	.w3(32'h3ba5366e),
	.w4(32'hba1e6d37),
	.w5(32'h3c596bbf),
	.w6(32'h3b0be7f7),
	.w7(32'h3b427201),
	.w8(32'hbb759bd0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe829),
	.w1(32'hbc43c374),
	.w2(32'hbc8d11c8),
	.w3(32'hbb611095),
	.w4(32'hbc8470e9),
	.w5(32'hbc6ccfa9),
	.w6(32'hbb2dc31c),
	.w7(32'hbc210127),
	.w8(32'hbb828187),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cf107),
	.w1(32'hbbfe89fb),
	.w2(32'hbcd8d988),
	.w3(32'hbbdc9ed3),
	.w4(32'hbc5df2b3),
	.w5(32'hbc845868),
	.w6(32'hbbcd0b4a),
	.w7(32'hbc776ce0),
	.w8(32'h3a857e4d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0276a8),
	.w1(32'hbc5159b4),
	.w2(32'hbcc4e92d),
	.w3(32'h3b8793c1),
	.w4(32'hbc4a2e1b),
	.w5(32'hbc9fe59b),
	.w6(32'hbbf4fff2),
	.w7(32'hbc4a1208),
	.w8(32'hb9f3c703),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1ef82),
	.w1(32'hbb551a0c),
	.w2(32'h3c68640b),
	.w3(32'hbb1cdd23),
	.w4(32'hba1ff01a),
	.w5(32'h3c165b5e),
	.w6(32'hbbb22396),
	.w7(32'h3c239588),
	.w8(32'h3b47c2cb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe11e2),
	.w1(32'hbc863593),
	.w2(32'hbbb498f1),
	.w3(32'h3b5a35f3),
	.w4(32'hbc556381),
	.w5(32'hbc1a9035),
	.w6(32'hbc334ac8),
	.w7(32'hbb208bcc),
	.w8(32'hbbf5986f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb714),
	.w1(32'hba84b090),
	.w2(32'hbb970890),
	.w3(32'h3b1e8826),
	.w4(32'hba9e672e),
	.w5(32'hbb7870ba),
	.w6(32'hbb595a74),
	.w7(32'h3add3287),
	.w8(32'h3b878d62),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb019a),
	.w1(32'hb98633f3),
	.w2(32'h3be68ebc),
	.w3(32'hbb4e74ec),
	.w4(32'h3b9db963),
	.w5(32'hbb818913),
	.w6(32'hbba3464f),
	.w7(32'hbadbef6e),
	.w8(32'hbb107171),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37b712),
	.w1(32'h3c706a84),
	.w2(32'h3a99ca54),
	.w3(32'h3b29f658),
	.w4(32'h3c130d76),
	.w5(32'hbc37e1a0),
	.w6(32'h3c2f7c97),
	.w7(32'h3b955115),
	.w8(32'h3a9abd8c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1709b),
	.w1(32'hbacbfe90),
	.w2(32'h3c6dd4bf),
	.w3(32'h3bacdbbc),
	.w4(32'h3ae84f86),
	.w5(32'h3c0d6795),
	.w6(32'h3b3fb510),
	.w7(32'h3c34fa49),
	.w8(32'h3a7f3dac),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1394db),
	.w1(32'hbc026ade),
	.w2(32'hbbc568c3),
	.w3(32'h3b737013),
	.w4(32'h3b1703e2),
	.w5(32'h3c0aa6b9),
	.w6(32'h3b7df346),
	.w7(32'h3c27c7e7),
	.w8(32'h3ad8e799),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b4de3),
	.w1(32'h3c54a0f5),
	.w2(32'hbaf1b76e),
	.w3(32'h3c118c42),
	.w4(32'hbb6b7d03),
	.w5(32'hbceed5e1),
	.w6(32'h3c93b03d),
	.w7(32'h3cac68b4),
	.w8(32'h38d22277),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc953704),
	.w1(32'h3a352abe),
	.w2(32'h3ba9f47d),
	.w3(32'hb7ae9aef),
	.w4(32'h3a3957aa),
	.w5(32'h3bb0e3d9),
	.w6(32'h3a66d576),
	.w7(32'h3bb37c57),
	.w8(32'hbc00c1b3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefc738),
	.w1(32'h3c19c345),
	.w2(32'hb9a5d1b4),
	.w3(32'hbb0dfefb),
	.w4(32'h3cb0ef79),
	.w5(32'hbb03f949),
	.w6(32'hb96e88c4),
	.w7(32'h3bd15ce4),
	.w8(32'h3c08b39a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d96f8),
	.w1(32'hbbb6f845),
	.w2(32'hbc1cade8),
	.w3(32'hbc9ff7cd),
	.w4(32'hba0eea27),
	.w5(32'hb93d0a39),
	.w6(32'h3b1726db),
	.w7(32'hb9873ca3),
	.w8(32'hbbabbfaa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3855b),
	.w1(32'h3c809d6a),
	.w2(32'hbba8cedc),
	.w3(32'h3be5bd38),
	.w4(32'hbbd3d258),
	.w5(32'hbb491de0),
	.w6(32'h3a975723),
	.w7(32'hbba14989),
	.w8(32'h3bb11340),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22393e),
	.w1(32'hba9aea75),
	.w2(32'h3b7aa4a6),
	.w3(32'h3c0a1271),
	.w4(32'hbbc4b176),
	.w5(32'hbaff241d),
	.w6(32'hba9c153a),
	.w7(32'hba38827d),
	.w8(32'hbab10925),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe94cf),
	.w1(32'hbaa2ca4a),
	.w2(32'hbb627e2a),
	.w3(32'h3a8565d6),
	.w4(32'hbbb853ba),
	.w5(32'hbb5aba90),
	.w6(32'hba12d82d),
	.w7(32'hba8e8e1e),
	.w8(32'hbb32a4bb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b887),
	.w1(32'h3b8be81e),
	.w2(32'h3bfa8889),
	.w3(32'hb8cb5fe2),
	.w4(32'hbac669d6),
	.w5(32'h3b0daed5),
	.w6(32'h3a89f4c1),
	.w7(32'h3b5f7d54),
	.w8(32'h3a19907e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5281f),
	.w1(32'h3c1fa780),
	.w2(32'h3bad8349),
	.w3(32'h39e00002),
	.w4(32'h3c000fbc),
	.w5(32'h3b11e8b2),
	.w6(32'h3b9b8453),
	.w7(32'h3b38b81b),
	.w8(32'hbb1292cb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9c4e5),
	.w1(32'h3d320d5e),
	.w2(32'hbccefb96),
	.w3(32'h3ace83ea),
	.w4(32'h3d0fb9f4),
	.w5(32'hbc92e826),
	.w6(32'h3cc2e0a7),
	.w7(32'hbb931cda),
	.w8(32'hbc90fb08),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce97b6a),
	.w1(32'hbc398813),
	.w2(32'hbcc7484e),
	.w3(32'hbc55775d),
	.w4(32'hbbbd113a),
	.w5(32'hbc579414),
	.w6(32'hbb8a6b93),
	.w7(32'hbc473c89),
	.w8(32'h3b2ee03a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7337f3),
	.w1(32'hbaa6e0ff),
	.w2(32'hbb8b3fca),
	.w3(32'h3ba933d1),
	.w4(32'hbb4fbe7a),
	.w5(32'hbbeb003f),
	.w6(32'h3a03bd80),
	.w7(32'hbb8ad5cf),
	.w8(32'hbbc55c1d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc864939),
	.w1(32'h3ac8d4df),
	.w2(32'hbc54fc17),
	.w3(32'hbbbf2ac5),
	.w4(32'hbaec387a),
	.w5(32'hbbc6ecb1),
	.w6(32'hb9b18b31),
	.w7(32'hbc56e704),
	.w8(32'hbc1e7aa9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3a1f),
	.w1(32'h3bd80382),
	.w2(32'hbc6e79c0),
	.w3(32'hbc57dcf5),
	.w4(32'h3b7ea554),
	.w5(32'hbc34e41c),
	.w6(32'h3b2479d5),
	.w7(32'hbc09226e),
	.w8(32'hbb887673),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ad1fc),
	.w1(32'hbbff3dec),
	.w2(32'hbc06aa68),
	.w3(32'h3b91ef62),
	.w4(32'hbc57fc4b),
	.w5(32'hbbd3c5ba),
	.w6(32'h3aa8d2e0),
	.w7(32'h3ba65912),
	.w8(32'h3c3f98e9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89a60d),
	.w1(32'hbb8335f4),
	.w2(32'h3c2acd5e),
	.w3(32'h3c95092f),
	.w4(32'hbb997777),
	.w5(32'h392fb198),
	.w6(32'hb9d91706),
	.w7(32'h3c46dc31),
	.w8(32'hbb27d38e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d89f7),
	.w1(32'hbc35fcb3),
	.w2(32'h3b8927a4),
	.w3(32'h3b026842),
	.w4(32'h3bd02d7b),
	.w5(32'h3bf44aaf),
	.w6(32'hb8a9ad5b),
	.w7(32'hbc470519),
	.w8(32'h3bef2913),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6538a3),
	.w1(32'h3b58f05e),
	.w2(32'h3bae92e3),
	.w3(32'h3b341b62),
	.w4(32'h3b6efafe),
	.w5(32'h3c111635),
	.w6(32'hbb4312cc),
	.w7(32'hb9dc8343),
	.w8(32'hbb815791),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78b018),
	.w1(32'hbc19be96),
	.w2(32'hbb3cdd86),
	.w3(32'hbb5bd6d2),
	.w4(32'hbc8b80ec),
	.w5(32'h3b0dcf88),
	.w6(32'h3b51a671),
	.w7(32'hbca69f5f),
	.w8(32'h3c194273),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc39ef1),
	.w1(32'h3ca5ed07),
	.w2(32'h3ca4d27c),
	.w3(32'h3caaefda),
	.w4(32'h3c77b9f5),
	.w5(32'h3c9802ac),
	.w6(32'h3c5a45fe),
	.w7(32'h3c4d5acf),
	.w8(32'hb9ab10e7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45445a),
	.w1(32'hb87086b6),
	.w2(32'hb624fab6),
	.w3(32'hbbede9e0),
	.w4(32'hb990bfda),
	.w5(32'h3af7efb5),
	.w6(32'h37dbe0eb),
	.w7(32'h3b7d14af),
	.w8(32'h3bf73d5b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15700f),
	.w1(32'hbc072fa6),
	.w2(32'hbcef47c9),
	.w3(32'h3c0baa71),
	.w4(32'hbc36eb1b),
	.w5(32'hbc6ec7fd),
	.w6(32'h3c15edd9),
	.w7(32'hba9b738a),
	.w8(32'hbc7b4d05),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7ecf),
	.w1(32'hbc6373a2),
	.w2(32'hbce4d71e),
	.w3(32'h3a4227f2),
	.w4(32'h3a72c1f1),
	.w5(32'hbc9fa519),
	.w6(32'hbc0ace02),
	.w7(32'hbc7f00aa),
	.w8(32'h3aebe959),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd455b4),
	.w1(32'hbb6df39e),
	.w2(32'h3bd22241),
	.w3(32'hbbb60f4a),
	.w4(32'hbbd66d89),
	.w5(32'h3b7b76d2),
	.w6(32'hbbd0e742),
	.w7(32'hba8f3bb0),
	.w8(32'h3b79204d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc183b0),
	.w1(32'h3b90fa8a),
	.w2(32'h3b8934e5),
	.w3(32'h3bbc7e32),
	.w4(32'h3b098ef2),
	.w5(32'h3b265d0a),
	.w6(32'hba3749fa),
	.w7(32'h3aaf7e09),
	.w8(32'hbbbcf691),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1609f0),
	.w1(32'h3b963538),
	.w2(32'h3bc8532a),
	.w3(32'hbba78398),
	.w4(32'h3c0a7db4),
	.w5(32'h3c1d0bda),
	.w6(32'h387db1ca),
	.w7(32'hba34eee1),
	.w8(32'hb8071684),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f409),
	.w1(32'h3c3650b0),
	.w2(32'h3c076590),
	.w3(32'hbb644241),
	.w4(32'h3c552c30),
	.w5(32'h3c1f05b6),
	.w6(32'h3c635acd),
	.w7(32'h3c3a9cb7),
	.w8(32'h3bceb783),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad779de),
	.w1(32'h3bd69efa),
	.w2(32'h3a4b2704),
	.w3(32'h3bc4788f),
	.w4(32'h3bb19a5b),
	.w5(32'h3b9821da),
	.w6(32'h3b403ce7),
	.w7(32'h3a337f94),
	.w8(32'hba016d8c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38242fed),
	.w1(32'hba05fee8),
	.w2(32'hbb549fc1),
	.w3(32'h3a5314c6),
	.w4(32'h3bd003d8),
	.w5(32'hbaae3a40),
	.w6(32'hbc1e242b),
	.w7(32'hbacc6dad),
	.w8(32'h3c825470),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a41863),
	.w1(32'hbb22ba89),
	.w2(32'h3c7f9f31),
	.w3(32'hbb45bf92),
	.w4(32'hbb8dd6f2),
	.w5(32'h3c55546d),
	.w6(32'hbb5a9033),
	.w7(32'h3bbb6d3c),
	.w8(32'hbb4626a7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb492ed),
	.w1(32'h3bc1af54),
	.w2(32'hbb97d3b8),
	.w3(32'h3c1ea571),
	.w4(32'h3b93e2a4),
	.w5(32'hbba20347),
	.w6(32'h3b478881),
	.w7(32'hbaccaa4a),
	.w8(32'hbc1bebeb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc527b2d),
	.w1(32'hbac8820d),
	.w2(32'hbb03703a),
	.w3(32'hbc40cac8),
	.w4(32'hbc0d7418),
	.w5(32'hbb831fe0),
	.w6(32'hbb710c26),
	.w7(32'hbbbb7e96),
	.w8(32'hbbcfbd0c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2412),
	.w1(32'hba9690f7),
	.w2(32'h3ac22b9b),
	.w3(32'hbc56bb25),
	.w4(32'hbb076441),
	.w5(32'h3b6c077e),
	.w6(32'hbb013c2c),
	.w7(32'hbadff877),
	.w8(32'h3b1a1f82),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09a47e),
	.w1(32'h3bcf5b24),
	.w2(32'hbbde9244),
	.w3(32'hbb8cae2b),
	.w4(32'h3c84ef4f),
	.w5(32'hbb205587),
	.w6(32'hbbb7dd71),
	.w7(32'hbc903c99),
	.w8(32'h3b0402c6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c56c9),
	.w1(32'hbb1a130c),
	.w2(32'h3c77d646),
	.w3(32'hbb2826da),
	.w4(32'hbb0fdc3e),
	.w5(32'h3c409620),
	.w6(32'hbbb2150a),
	.w7(32'h3b4ea236),
	.w8(32'h3b93d4e4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca22dde),
	.w1(32'h3c2c34b8),
	.w2(32'h3a4e628f),
	.w3(32'h3bab05f5),
	.w4(32'h3b5dfb9b),
	.w5(32'hbaf95ec0),
	.w6(32'h3ba0de24),
	.w7(32'h3b428354),
	.w8(32'h3bd3c8c0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7d0b6),
	.w1(32'hbc1a9bba),
	.w2(32'hbbd848cc),
	.w3(32'h3b06b661),
	.w4(32'hba7ac394),
	.w5(32'hbb0d96f3),
	.w6(32'h3b9ac89e),
	.w7(32'hbaad8e29),
	.w8(32'h3b083213),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39249f7d),
	.w1(32'h3b8c0171),
	.w2(32'h3bb1bf0e),
	.w3(32'hbb1172c1),
	.w4(32'h3bba4d33),
	.w5(32'h3b4c8f01),
	.w6(32'h3ac61cbc),
	.w7(32'h3aa6f025),
	.w8(32'hbac962e0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba702b24),
	.w1(32'h3c27b046),
	.w2(32'h3b1c9234),
	.w3(32'h3b241d5c),
	.w4(32'h3b9dfa2c),
	.w5(32'h3b8be78d),
	.w6(32'h3c18cbf4),
	.w7(32'hba8436d5),
	.w8(32'hb882c7ca),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a11b0d),
	.w1(32'hba553ad2),
	.w2(32'hbc74d58f),
	.w3(32'hba2a6d7c),
	.w4(32'h3b71929f),
	.w5(32'hbba4ae07),
	.w6(32'hbc131d63),
	.w7(32'hbc0c58d9),
	.w8(32'h3c28ccc4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f9f9b),
	.w1(32'h3a8842cd),
	.w2(32'hbbe6a894),
	.w3(32'h3bc279cd),
	.w4(32'hbc059482),
	.w5(32'h3b26509c),
	.w6(32'hb9ba72bc),
	.w7(32'h3c190fb9),
	.w8(32'h3bf649e1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29d062),
	.w1(32'hbb311db6),
	.w2(32'h3b3173fe),
	.w3(32'h3b56703e),
	.w4(32'h39db6d8e),
	.w5(32'h3b95834e),
	.w6(32'h3a980f17),
	.w7(32'h3bbfe530),
	.w8(32'h39e00b18),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b368a),
	.w1(32'hbba5f9e5),
	.w2(32'hbb696583),
	.w3(32'hbb14399c),
	.w4(32'hb9ee88b0),
	.w5(32'h3c113ece),
	.w6(32'hbb0f8023),
	.w7(32'hbb864deb),
	.w8(32'h3b44d7ce),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule