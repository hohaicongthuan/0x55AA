module layer_10_featuremap_426(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada26d6),
	.w1(32'hbb447d68),
	.w2(32'hbb82c86b),
	.w3(32'hbba3f88f),
	.w4(32'hbb9243bc),
	.w5(32'hbc3d62b3),
	.w6(32'hbc058d23),
	.w7(32'hbb94e054),
	.w8(32'hbbc1a6b9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a59e),
	.w1(32'h3b3f4c07),
	.w2(32'h3ba6856d),
	.w3(32'hbb3bd648),
	.w4(32'h39009c4d),
	.w5(32'hbb49c201),
	.w6(32'hbaef030c),
	.w7(32'h3a83d93f),
	.w8(32'hbaa8f81e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdae698),
	.w1(32'h3a56f0e5),
	.w2(32'hbb67c10a),
	.w3(32'h3c1e3892),
	.w4(32'hbb4cf973),
	.w5(32'hbbab3909),
	.w6(32'h3c33662e),
	.w7(32'hbc12e7a8),
	.w8(32'hbba9b399),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e28dd),
	.w1(32'hbc2d92d6),
	.w2(32'h39c302b6),
	.w3(32'h3b870932),
	.w4(32'hbbd6d314),
	.w5(32'h3af03e8c),
	.w6(32'hbb6acc93),
	.w7(32'hbbaf0f92),
	.w8(32'hbab344f5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25c706),
	.w1(32'hbad1de71),
	.w2(32'h3a83c7ee),
	.w3(32'hbbc904e5),
	.w4(32'h3ac74c23),
	.w5(32'h3c26f7ea),
	.w6(32'hbb35d1d0),
	.w7(32'hbbc47dc3),
	.w8(32'hb9349087),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d495c6),
	.w1(32'h3b53b80c),
	.w2(32'h3b8704be),
	.w3(32'h3c182dfb),
	.w4(32'h3c138f05),
	.w5(32'hbba3a1db),
	.w6(32'h3b9e6c14),
	.w7(32'h3adf2914),
	.w8(32'hbbf3b680),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf657e),
	.w1(32'h3c191ad7),
	.w2(32'h3c403fc4),
	.w3(32'h3b3ee29b),
	.w4(32'h3bedaa4d),
	.w5(32'h3c40f4d5),
	.w6(32'hbb4e9f64),
	.w7(32'h3c5c371b),
	.w8(32'h3c31b81f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be53731),
	.w1(32'h3b306977),
	.w2(32'h394cd106),
	.w3(32'h3bea9677),
	.w4(32'h3bb784b9),
	.w5(32'hbb1421f8),
	.w6(32'h3b9f0ad9),
	.w7(32'h39df0ad7),
	.w8(32'hbb5164c4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b052c),
	.w1(32'hbb39ce48),
	.w2(32'h3980bc78),
	.w3(32'hbc0ef04e),
	.w4(32'hbbd40665),
	.w5(32'h3b40df52),
	.w6(32'hbc46cec8),
	.w7(32'hbad72f1f),
	.w8(32'hba9694e6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3827d5),
	.w1(32'hb9bc77ba),
	.w2(32'h3bb92802),
	.w3(32'h3b6cd807),
	.w4(32'hbb1292d6),
	.w5(32'h3bb96de0),
	.w6(32'h3b739188),
	.w7(32'hb91eb812),
	.w8(32'h3bdae287),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9956cc3),
	.w1(32'h3bf0e15e),
	.w2(32'h3bd569c2),
	.w3(32'h3a1fa875),
	.w4(32'h3aeaf8b4),
	.w5(32'h3b71fc0d),
	.w6(32'hba5f465c),
	.w7(32'h3b0bd0b0),
	.w8(32'h3b5c9408),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4a2f7),
	.w1(32'h3c19eb82),
	.w2(32'h3b51ffab),
	.w3(32'h3bd19e4b),
	.w4(32'h3c419ee0),
	.w5(32'h3bf18c49),
	.w6(32'h3bb9f598),
	.w7(32'h3b8c083f),
	.w8(32'h3b1f3197),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdb315),
	.w1(32'hbb45c8ff),
	.w2(32'hbb9a8366),
	.w3(32'h3c646eb0),
	.w4(32'hbaf126e9),
	.w5(32'hbb9df313),
	.w6(32'h3b91c078),
	.w7(32'hbb9257f1),
	.w8(32'hbaed3be1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb956eb8),
	.w1(32'h3a26148f),
	.w2(32'hbb45f4bf),
	.w3(32'h3c347550),
	.w4(32'hb98fca65),
	.w5(32'hbad9a896),
	.w6(32'h3aa3dcd7),
	.w7(32'hbba218cd),
	.w8(32'hbb405496),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55c9cd),
	.w1(32'hbb03e3b1),
	.w2(32'hbbec74e7),
	.w3(32'hbbbc79fa),
	.w4(32'h3b94d4a3),
	.w5(32'h3b93da43),
	.w6(32'hba9a9020),
	.w7(32'h39141963),
	.w8(32'h3b863e91),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2244a),
	.w1(32'h3ba36895),
	.w2(32'h3b8c80d9),
	.w3(32'h3b5d17a0),
	.w4(32'h3ba5ca5e),
	.w5(32'h3b98db6d),
	.w6(32'h3baffbd1),
	.w7(32'h3b48791f),
	.w8(32'h3b8e2c2a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38123e8b),
	.w1(32'hbc08f003),
	.w2(32'hbc2043b7),
	.w3(32'h3b319f6b),
	.w4(32'hbc2799b1),
	.w5(32'hbc044210),
	.w6(32'hbb3ad3d6),
	.w7(32'hbb94074f),
	.w8(32'hb98b21f2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ed59f),
	.w1(32'hbbe01080),
	.w2(32'hbb90ad1c),
	.w3(32'h3aa85a31),
	.w4(32'hbc59b211),
	.w5(32'hbc699ef2),
	.w6(32'h3bc22040),
	.w7(32'hbbe1e9c9),
	.w8(32'hbbe7068f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad488c1),
	.w1(32'h3a9a323a),
	.w2(32'hbb2f6660),
	.w3(32'hbbdee3fb),
	.w4(32'h3aab9af8),
	.w5(32'h3c2f243a),
	.w6(32'hbb33b52a),
	.w7(32'hbae8ef5e),
	.w8(32'h3b0eb575),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9030798),
	.w1(32'hbb093f5e),
	.w2(32'hbbd4dbfa),
	.w3(32'h3c2e1ee5),
	.w4(32'hbb10aa68),
	.w5(32'hbb03d815),
	.w6(32'h3bfc8700),
	.w7(32'h3b2eef46),
	.w8(32'hba23700e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78d923),
	.w1(32'h3c6dce22),
	.w2(32'h3c1b286c),
	.w3(32'h3b90890e),
	.w4(32'h3caf8482),
	.w5(32'h3c4212d4),
	.w6(32'h3bc35f31),
	.w7(32'h3c6b540a),
	.w8(32'h3c5f1976),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7edec4),
	.w1(32'h3bb7969f),
	.w2(32'hbae79f0a),
	.w3(32'h3c479e84),
	.w4(32'h3c4906bb),
	.w5(32'hbbc5ffe7),
	.w6(32'h3c0ee7fe),
	.w7(32'h3bcd9f13),
	.w8(32'hbba17060),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb790b),
	.w1(32'h3bbfe9a0),
	.w2(32'h3c204474),
	.w3(32'h3b4041d0),
	.w4(32'h3bbd9635),
	.w5(32'h3c17a3d2),
	.w6(32'hbb387979),
	.w7(32'h3b011b7b),
	.w8(32'h3ac393fb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b717bcf),
	.w1(32'hbc17e33c),
	.w2(32'h3bce6088),
	.w3(32'h3b33dce5),
	.w4(32'hb8bacf2a),
	.w5(32'h3c8fde06),
	.w6(32'h3a225eda),
	.w7(32'hbbece5f2),
	.w8(32'h3c18b015),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b1ce5),
	.w1(32'h3a4a960b),
	.w2(32'h3c15e24e),
	.w3(32'h3ce4fd5f),
	.w4(32'hbafe3a74),
	.w5(32'h3b7c9091),
	.w6(32'h3c63d1e0),
	.w7(32'hbb50725c),
	.w8(32'hbb4636de),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b781eaf),
	.w1(32'h3baae5e4),
	.w2(32'h3b9941d3),
	.w3(32'hbb9214ad),
	.w4(32'h3b97e94a),
	.w5(32'h3a3ffbc3),
	.w6(32'hba96a740),
	.w7(32'h3c2ab4b1),
	.w8(32'h3ac06280),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109ea5),
	.w1(32'hbaf00b25),
	.w2(32'hbc0817fb),
	.w3(32'hbbb9c2f9),
	.w4(32'hbb533299),
	.w5(32'hbbaca8c2),
	.w6(32'h3ad62ae5),
	.w7(32'hbb36b24f),
	.w8(32'hbbd6eb6a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bcfea),
	.w1(32'hb994e704),
	.w2(32'h3bd1883c),
	.w3(32'hbbb33da1),
	.w4(32'hba920a55),
	.w5(32'h3babb85c),
	.w6(32'hbc0d8a47),
	.w7(32'h3a9c74f2),
	.w8(32'h3ada00bd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba151014),
	.w1(32'h3ae9c298),
	.w2(32'h3b0ced71),
	.w3(32'hbae07ea6),
	.w4(32'hb9ccc77d),
	.w5(32'hb9d5da17),
	.w6(32'h39232d45),
	.w7(32'h3ba55639),
	.w8(32'h3b352e49),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38907d33),
	.w1(32'h3b84649d),
	.w2(32'h3b5da630),
	.w3(32'h3ac2699f),
	.w4(32'h3b87c27b),
	.w5(32'h3bdff7d7),
	.w6(32'h3c0983dd),
	.w7(32'hbb4b01b5),
	.w8(32'hb925bd3b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6bbea),
	.w1(32'h3ba1bdc3),
	.w2(32'h3b64f9e7),
	.w3(32'h3bc83f21),
	.w4(32'hbbdb1c70),
	.w5(32'hbbd94af4),
	.w6(32'h3a10f230),
	.w7(32'h3a35b3b7),
	.w8(32'h3aebf6e6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e5f09),
	.w1(32'h3b367428),
	.w2(32'h3a96bfb7),
	.w3(32'hbb8214f5),
	.w4(32'h3ba86f2c),
	.w5(32'hbb38665b),
	.w6(32'h3bdab91b),
	.w7(32'h3b9e284a),
	.w8(32'h3a8b136a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15dddd),
	.w1(32'h3aed8a3a),
	.w2(32'h3af8e533),
	.w3(32'h3b370634),
	.w4(32'hbb87ac39),
	.w5(32'h3b9d24ef),
	.w6(32'h3ae682ec),
	.w7(32'h39e12247),
	.w8(32'h3b881010),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8322),
	.w1(32'h3abf2555),
	.w2(32'h3a49630c),
	.w3(32'h3a4e8e0b),
	.w4(32'hb9a325e9),
	.w5(32'h3b48f7fc),
	.w6(32'h399c511c),
	.w7(32'h3b95df73),
	.w8(32'hbba2db6b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44e5e7),
	.w1(32'hb99b769b),
	.w2(32'hbab7f2c5),
	.w3(32'hbb57d82c),
	.w4(32'hbb02369b),
	.w5(32'hba3cccec),
	.w6(32'hbbf57cad),
	.w7(32'hbaf42f3b),
	.w8(32'h3b5c7cd8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b12b),
	.w1(32'h3953e9bf),
	.w2(32'h3b8a6772),
	.w3(32'hbb8f90af),
	.w4(32'h3b13c669),
	.w5(32'hbb388d96),
	.w6(32'hbb453a95),
	.w7(32'h3b9dc792),
	.w8(32'h3ad059a6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb660e6),
	.w1(32'h3b813b58),
	.w2(32'h3c03a07a),
	.w3(32'hbb90c600),
	.w4(32'hbbf80d02),
	.w5(32'hbb816a46),
	.w6(32'hbbbe9374),
	.w7(32'hbc09a88d),
	.w8(32'hbbb8fc5a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c599777),
	.w1(32'hbbc7de63),
	.w2(32'hb965e629),
	.w3(32'h3b88f507),
	.w4(32'hbc5132ec),
	.w5(32'hbc0d2af1),
	.w6(32'h3b4e0d80),
	.w7(32'hbc2cd283),
	.w8(32'hbc059136),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e14c4),
	.w1(32'hbb80c8ac),
	.w2(32'h39b3643a),
	.w3(32'h3c295020),
	.w4(32'hbb9c470f),
	.w5(32'hbb288103),
	.w6(32'h3b5f82b2),
	.w7(32'hbbfda140),
	.w8(32'hbb9a23e0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f4c0c),
	.w1(32'hbbd48c1c),
	.w2(32'h3bb8f92e),
	.w3(32'hbc762326),
	.w4(32'hbbac4cdd),
	.w5(32'h3b065da0),
	.w6(32'hbc269c77),
	.w7(32'hbb0950a0),
	.w8(32'h3b34917b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2fd36),
	.w1(32'hbb950b53),
	.w2(32'hba19f8cb),
	.w3(32'h3855baec),
	.w4(32'hbb34937e),
	.w5(32'h3b303202),
	.w6(32'h3af585e7),
	.w7(32'hbc0407f3),
	.w8(32'hbb403ee3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af914),
	.w1(32'hbb92f2d5),
	.w2(32'hbb951bff),
	.w3(32'hbc040bb1),
	.w4(32'hb9f58533),
	.w5(32'h393dede5),
	.w6(32'hbba9a205),
	.w7(32'hbb0a8de0),
	.w8(32'hbabff0e6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e89ba6),
	.w1(32'h39baae81),
	.w2(32'h3ad6d148),
	.w3(32'h3b594e34),
	.w4(32'hbaa0dc49),
	.w5(32'hbb636c95),
	.w6(32'hbadb30e0),
	.w7(32'hbba22d5f),
	.w8(32'hbbbef6a9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873eda),
	.w1(32'hbb18a671),
	.w2(32'h3b5652f5),
	.w3(32'hbba5b08e),
	.w4(32'hbb1e09a8),
	.w5(32'hbac1738a),
	.w6(32'h39a614a1),
	.w7(32'hbb13f470),
	.w8(32'h3aa4dd06),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfe71c),
	.w1(32'hbb92cb4b),
	.w2(32'hbabe2ae2),
	.w3(32'hbb96eb25),
	.w4(32'hbbe8aadb),
	.w5(32'hba8263e3),
	.w6(32'hbb07a588),
	.w7(32'hbc23702d),
	.w8(32'hbbee81f8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8f6a5),
	.w1(32'h3b420b36),
	.w2(32'h3c07b009),
	.w3(32'hbaa99769),
	.w4(32'hbb0df524),
	.w5(32'h3bdaa192),
	.w6(32'hba0f42ba),
	.w7(32'hbb2bf2cd),
	.w8(32'h3c0e2d35),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7efb25),
	.w1(32'h3ab86235),
	.w2(32'hbaceba5e),
	.w3(32'h3ba1d21f),
	.w4(32'hbaf0b81c),
	.w5(32'hba8ab080),
	.w6(32'h3a13fa49),
	.w7(32'hbaa39280),
	.w8(32'h3be9267a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93021f),
	.w1(32'h3b8f2dcf),
	.w2(32'h3bc6f0b4),
	.w3(32'h3c110c8f),
	.w4(32'h3bfeda47),
	.w5(32'h3bc4242c),
	.w6(32'h3ba9502c),
	.w7(32'h3bcbe3fa),
	.w8(32'h3bfd04c4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2fae),
	.w1(32'h3b9ff8a2),
	.w2(32'h3b81f5b4),
	.w3(32'hbb1dda4e),
	.w4(32'h3c286a9e),
	.w5(32'h3bddf8de),
	.w6(32'hbaf13aa6),
	.w7(32'h3c00b900),
	.w8(32'h3a841d9b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40ca9c),
	.w1(32'h3bff5b45),
	.w2(32'h3b62aebe),
	.w3(32'hbbb44030),
	.w4(32'h3c6f9941),
	.w5(32'hbb60860a),
	.w6(32'hba0889ce),
	.w7(32'h3c460d19),
	.w8(32'h3b099d86),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7f046),
	.w1(32'hbb4fe14c),
	.w2(32'hbbad532d),
	.w3(32'hbb2d80e6),
	.w4(32'h3b0d645e),
	.w5(32'hbb2ad5bb),
	.w6(32'h3a9c1588),
	.w7(32'hbb5455f4),
	.w8(32'hbad94d81),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab90329),
	.w1(32'hbb9bdeb2),
	.w2(32'hb93b3146),
	.w3(32'h3c78e037),
	.w4(32'hbbe42a15),
	.w5(32'hbae41a4e),
	.w6(32'h3c0da458),
	.w7(32'hbb9d1c31),
	.w8(32'hbb05dfc0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2b7f),
	.w1(32'h3c16cb3b),
	.w2(32'h3c44a6e7),
	.w3(32'hbbb9a501),
	.w4(32'h3c39bc56),
	.w5(32'h3b53037a),
	.w6(32'hbb3b41b5),
	.w7(32'h3c28cf68),
	.w8(32'hbb10676e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2152f4),
	.w1(32'h3c0a558f),
	.w2(32'h3c57b0ef),
	.w3(32'h3a0bf7cf),
	.w4(32'h3aae84c3),
	.w5(32'h3b81607e),
	.w6(32'hbb2d5102),
	.w7(32'h3bc2223f),
	.w8(32'h3aa0ff71),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdfcbf),
	.w1(32'hbbdcc3c4),
	.w2(32'h3a3eb523),
	.w3(32'h3b2de095),
	.w4(32'hbc203f12),
	.w5(32'hbb1fcd46),
	.w6(32'hbc291464),
	.w7(32'hbbed7ca7),
	.w8(32'hbb101c7a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dfd993),
	.w1(32'hbb2baf6e),
	.w2(32'h3c085dc4),
	.w3(32'hbb3c3501),
	.w4(32'hbb91fb44),
	.w5(32'hbad6c1bc),
	.w6(32'hbabc756e),
	.w7(32'hba96db06),
	.w8(32'h39836fe2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4c2e9),
	.w1(32'h3b8faa7d),
	.w2(32'h3a174810),
	.w3(32'h3b7526fd),
	.w4(32'h3b09ea08),
	.w5(32'h3c1de309),
	.w6(32'h3b661dce),
	.w7(32'hbaa83065),
	.w8(32'h3b696e49),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0942e),
	.w1(32'hbb6348e6),
	.w2(32'h3b548028),
	.w3(32'h3c32ea47),
	.w4(32'hbaede9ee),
	.w5(32'h3b83ecf7),
	.w6(32'h3bd64971),
	.w7(32'hbb295ec1),
	.w8(32'hbb94a323),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0ba5),
	.w1(32'hba39bf4f),
	.w2(32'hb9483a72),
	.w3(32'h3ae2e2d9),
	.w4(32'h3a157785),
	.w5(32'hbaa7c088),
	.w6(32'hbb317e27),
	.w7(32'hbace237e),
	.w8(32'hbb074e94),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38fa0d),
	.w1(32'hbb2635e3),
	.w2(32'h3b4f86f7),
	.w3(32'hba5e554e),
	.w4(32'h3b36808d),
	.w5(32'h3bd283d8),
	.w6(32'hba25d8a8),
	.w7(32'h3b92c722),
	.w8(32'h3b98583c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fba41),
	.w1(32'hba8d9194),
	.w2(32'hbab582be),
	.w3(32'h3b5a8c39),
	.w4(32'hbad5f803),
	.w5(32'hb8e25049),
	.w6(32'h3ac525e1),
	.w7(32'hbb6e46d2),
	.w8(32'h3a57ce81),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e39e6),
	.w1(32'h3b0f11f1),
	.w2(32'hbb155c50),
	.w3(32'h3b30511d),
	.w4(32'h3b95acc3),
	.w5(32'h3b93c37f),
	.w6(32'hbb220384),
	.w7(32'hb9b2b6b2),
	.w8(32'hba19a925),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983d3b1),
	.w1(32'hbbf264be),
	.w2(32'hbaac3b86),
	.w3(32'h3ad28302),
	.w4(32'hbc010706),
	.w5(32'hbc007068),
	.w6(32'h3b041687),
	.w7(32'hbbe4306b),
	.w8(32'hbbd3c85c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78acc),
	.w1(32'h39cc2721),
	.w2(32'hbb8478a6),
	.w3(32'hbc5011d2),
	.w4(32'hba39aa06),
	.w5(32'hba8362db),
	.w6(32'hbbbb4746),
	.w7(32'hb8c98c1d),
	.w8(32'hbb5019f6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27719b),
	.w1(32'h3b4956f6),
	.w2(32'h3a96c161),
	.w3(32'h3ba430f7),
	.w4(32'h3b93bdfd),
	.w5(32'h3a6ff6f6),
	.w6(32'hba7a6072),
	.w7(32'h3ae91440),
	.w8(32'hbabae5e0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd4fe4),
	.w1(32'h3c5f7f57),
	.w2(32'h3c2609ca),
	.w3(32'hbbadc125),
	.w4(32'h3c872fbf),
	.w5(32'h3c782212),
	.w6(32'hbc078540),
	.w7(32'h3c355b69),
	.w8(32'h3c11ae00),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b112745),
	.w1(32'h3c29cce2),
	.w2(32'h3c044eb9),
	.w3(32'hbb4354de),
	.w4(32'h3c34234e),
	.w5(32'h3a170c02),
	.w6(32'hbb4f35da),
	.w7(32'h3c14d937),
	.w8(32'h3b754766),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137d60),
	.w1(32'h3ad318c2),
	.w2(32'h3c314325),
	.w3(32'h3a3e366b),
	.w4(32'hbb78c2e7),
	.w5(32'h3b3b9ba4),
	.w6(32'h3a854da6),
	.w7(32'hbb4ea995),
	.w8(32'h3bad6503),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf68ef9),
	.w1(32'h3b6d747a),
	.w2(32'h3bfb50fa),
	.w3(32'h3b3a3d27),
	.w4(32'h3a4be7cf),
	.w5(32'hb9985c7f),
	.w6(32'h3ba648d8),
	.w7(32'h3b04a40a),
	.w8(32'h3b217851),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb674f2),
	.w1(32'hbbb58139),
	.w2(32'h3bcd755a),
	.w3(32'h3c8db6bd),
	.w4(32'hbb9d6dc3),
	.w5(32'h3b042fcf),
	.w6(32'h3cb65208),
	.w7(32'hbc0a6ea6),
	.w8(32'h3a1a51a2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9caf58),
	.w1(32'h38f4f5d6),
	.w2(32'hbad3d978),
	.w3(32'h3af041e9),
	.w4(32'hbba2c528),
	.w5(32'h3b53cdb7),
	.w6(32'h3aabb202),
	.w7(32'h3a908956),
	.w8(32'h3aec1370),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48d87e),
	.w1(32'h3b9dc43d),
	.w2(32'h3bc3c6e0),
	.w3(32'h3a95bb95),
	.w4(32'hba913b3b),
	.w5(32'h3b6409d0),
	.w6(32'h3b8275a0),
	.w7(32'hbb66591a),
	.w8(32'hbb626286),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2755d),
	.w1(32'h3b588b42),
	.w2(32'hb8851ee0),
	.w3(32'hbaf88f83),
	.w4(32'h3c3a15af),
	.w5(32'h3b36959a),
	.w6(32'hbb271678),
	.w7(32'h3b1c2a14),
	.w8(32'h3b13038c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc5901),
	.w1(32'hba80f5b4),
	.w2(32'h391aa68c),
	.w3(32'h3b0f034a),
	.w4(32'h3b0128a4),
	.w5(32'h3b095530),
	.w6(32'h3c0565b2),
	.w7(32'h3ad995f6),
	.w8(32'h39e5dd3d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d9806),
	.w1(32'hbb867e8a),
	.w2(32'h3abd2647),
	.w3(32'hba3d6042),
	.w4(32'h38bcc473),
	.w5(32'hbb49fab1),
	.w6(32'h3b1d22d4),
	.w7(32'hba320604),
	.w8(32'h3b6e3356),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cb704),
	.w1(32'hbac16225),
	.w2(32'hba4f7e8c),
	.w3(32'h3aa49094),
	.w4(32'h3b050474),
	.w5(32'hbaa8b7eb),
	.w6(32'h3ab7211d),
	.w7(32'h38fdda35),
	.w8(32'hba2c5b8c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e4880),
	.w1(32'h3b914159),
	.w2(32'h3b2e732f),
	.w3(32'hba8b78e5),
	.w4(32'h3b5f162e),
	.w5(32'h3be64b13),
	.w6(32'h3aeac912),
	.w7(32'h3a91c936),
	.w8(32'hba3f092e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0294f4),
	.w1(32'hbaf32f38),
	.w2(32'h3c18ebe8),
	.w3(32'h3b891aa9),
	.w4(32'h3b8af607),
	.w5(32'h3c3f0260),
	.w6(32'h3bb8ee3c),
	.w7(32'hbb6dfbcb),
	.w8(32'hbaadea93),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e293),
	.w1(32'h39873478),
	.w2(32'hba564eef),
	.w3(32'h3bbee40c),
	.w4(32'h3a7900b9),
	.w5(32'h3a3c89f4),
	.w6(32'hbb23edb5),
	.w7(32'h3b50607f),
	.w8(32'h3b5e05c0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ddc5f),
	.w1(32'hbb23d19b),
	.w2(32'hba0acbf2),
	.w3(32'h3b53ceca),
	.w4(32'hbacc01e6),
	.w5(32'h3bb6a7db),
	.w6(32'h3b762f01),
	.w7(32'h3b3a38dc),
	.w8(32'hbbbea713),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b5fc1),
	.w1(32'h3c11be11),
	.w2(32'h3ab0b8df),
	.w3(32'hbba4d60a),
	.w4(32'h3bb7fce7),
	.w5(32'hbbb07826),
	.w6(32'hbaa475c3),
	.w7(32'h3b971141),
	.w8(32'h3ae409cb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc32beb),
	.w1(32'hb9c7c063),
	.w2(32'hba7a4009),
	.w3(32'h3b668223),
	.w4(32'hbaba14d9),
	.w5(32'h3b18dab2),
	.w6(32'h3b3c6d89),
	.w7(32'hba933839),
	.w8(32'hba9003d9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e92fc),
	.w1(32'hbb4f1ffa),
	.w2(32'hbb6e8187),
	.w3(32'h3b3efd3f),
	.w4(32'hbb128550),
	.w5(32'hbb3b32d9),
	.w6(32'hbb238255),
	.w7(32'h3afdc4a8),
	.w8(32'h3bd74b9d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb658922),
	.w1(32'hbaca68cb),
	.w2(32'h3b0e9c58),
	.w3(32'h3b487f8b),
	.w4(32'hba2f1420),
	.w5(32'h3a4b1a15),
	.w6(32'h3b84e368),
	.w7(32'hba2ab7f4),
	.w8(32'hbb3bb1e8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba893f98),
	.w1(32'h3b07f576),
	.w2(32'hb972713a),
	.w3(32'h3b2e10f2),
	.w4(32'h39cdb0cf),
	.w5(32'hb93e3e2d),
	.w6(32'hbb35e0b5),
	.w7(32'hbadd3eef),
	.w8(32'h3b16596c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ff481),
	.w1(32'h3ae1e3f3),
	.w2(32'h3a63d0b9),
	.w3(32'h3b19cf36),
	.w4(32'h3b0f3842),
	.w5(32'hbb2ef4b1),
	.w6(32'h39c19ee4),
	.w7(32'h39d6fcae),
	.w8(32'hba0cdd65),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b684934),
	.w1(32'h3b661011),
	.w2(32'h3b3206da),
	.w3(32'h3af13567),
	.w4(32'h3ae6c99b),
	.w5(32'hbb50a552),
	.w6(32'hbad8f7e9),
	.w7(32'h3a7e6b8c),
	.w8(32'h3b990600),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3bb4a),
	.w1(32'hbaba1913),
	.w2(32'hbadd1dc5),
	.w3(32'hbb862ee1),
	.w4(32'h3a82c787),
	.w5(32'h3ac20661),
	.w6(32'h3b5b9074),
	.w7(32'h3b60ba09),
	.w8(32'h3bd79419),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9533f2),
	.w1(32'h3b2dc815),
	.w2(32'h3b8869a0),
	.w3(32'h3b7aa9b8),
	.w4(32'h3a196c5f),
	.w5(32'h3b454680),
	.w6(32'h3bc0a092),
	.w7(32'hbaa13019),
	.w8(32'h3a4997de),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840581),
	.w1(32'h39d3aa1f),
	.w2(32'h3c0fdd63),
	.w3(32'h38466387),
	.w4(32'h3bd39b5a),
	.w5(32'h3c9868d5),
	.w6(32'h3ae7dfd7),
	.w7(32'h3b580abf),
	.w8(32'h3bc7c745),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d9df2),
	.w1(32'hbb2e8c89),
	.w2(32'h3b97b3ed),
	.w3(32'h3be73d27),
	.w4(32'hbb59a7c2),
	.w5(32'h3bc48cfa),
	.w6(32'h3b9beb2f),
	.w7(32'hbb41eed3),
	.w8(32'hbb4b43f6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08f030),
	.w1(32'h39ae2244),
	.w2(32'h3ba31465),
	.w3(32'h39bcbe2d),
	.w4(32'h3b366f27),
	.w5(32'h3ca9ca4d),
	.w6(32'hbbbb78ed),
	.w7(32'hbb1f6cbb),
	.w8(32'h3b539fd0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0db65),
	.w1(32'h3a6d8d8a),
	.w2(32'h3af98a73),
	.w3(32'h3c21955d),
	.w4(32'hba273082),
	.w5(32'hbb31c74b),
	.w6(32'hba885951),
	.w7(32'hb997f345),
	.w8(32'hbaae6d19),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2f73),
	.w1(32'h3b89a830),
	.w2(32'h3b6fac83),
	.w3(32'h3a90a881),
	.w4(32'h3b07c81f),
	.w5(32'hb9b99429),
	.w6(32'h3aba3fbf),
	.w7(32'h3b8c66df),
	.w8(32'h3b941c6d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add5e4b),
	.w1(32'hb92ba034),
	.w2(32'h39891500),
	.w3(32'h3bca8a97),
	.w4(32'h3a71ccf6),
	.w5(32'h3c1dfccf),
	.w6(32'h3aaf1b02),
	.w7(32'hbb33eb4f),
	.w8(32'h3ae8c2b2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947f7dc),
	.w1(32'hbb99cd3c),
	.w2(32'h3b075d1f),
	.w3(32'h3aeeaa7c),
	.w4(32'hbbf9f4fe),
	.w5(32'h3b6f9a13),
	.w6(32'h3bdabd1f),
	.w7(32'hbbd460b3),
	.w8(32'hbba33774),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5159b0),
	.w1(32'h3a901143),
	.w2(32'hb9a94ef0),
	.w3(32'hbb9a62d9),
	.w4(32'h3abef1bf),
	.w5(32'h3b51f629),
	.w6(32'hb9fc5608),
	.w7(32'h3b8d5e96),
	.w8(32'h3b82ee1c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c282fb0),
	.w1(32'h3c47e053),
	.w2(32'h3c6cdf4c),
	.w3(32'h3c2a2abc),
	.w4(32'h3c075356),
	.w5(32'h3c26a499),
	.w6(32'h3c2a9d45),
	.w7(32'h3c34a4e4),
	.w8(32'h3c1124f7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3b1ab),
	.w1(32'h3c25208f),
	.w2(32'h3c9f1a24),
	.w3(32'h3bbacd92),
	.w4(32'h3c3f28ca),
	.w5(32'h3ceeb875),
	.w6(32'h3baecc6f),
	.w7(32'h3bf6fbfb),
	.w8(32'h3940af1d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b8530),
	.w1(32'hbb79d91a),
	.w2(32'h3c264382),
	.w3(32'h3c9b5e2e),
	.w4(32'h3b7d16a8),
	.w5(32'h3c802ee1),
	.w6(32'h3bd7e579),
	.w7(32'hbbd04f59),
	.w8(32'h3c1481e1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb37215),
	.w1(32'hbb34f6ad),
	.w2(32'h3b07d14c),
	.w3(32'h3c996460),
	.w4(32'hbbf38266),
	.w5(32'hbaabef95),
	.w6(32'h3c2712e8),
	.w7(32'hbbd18359),
	.w8(32'hbb2ee3a0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b279343),
	.w1(32'h3a8a0abd),
	.w2(32'h3bd7abe2),
	.w3(32'h3b95c8de),
	.w4(32'hbc19c5b2),
	.w5(32'h3b97f03f),
	.w6(32'h3be40073),
	.w7(32'hbbd3fb52),
	.w8(32'h3b098a3e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5885cb),
	.w1(32'hbb54ff65),
	.w2(32'hba866f07),
	.w3(32'h3b67c9cf),
	.w4(32'hbaa67a65),
	.w5(32'hb991bed1),
	.w6(32'hbb7361b1),
	.w7(32'hbb7e8bf1),
	.w8(32'h3b9dac8e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1f219),
	.w1(32'hb956a257),
	.w2(32'hba2cdf30),
	.w3(32'hbb4d1168),
	.w4(32'hbb492f61),
	.w5(32'hbb927585),
	.w6(32'hbb18c048),
	.w7(32'hb91b44c3),
	.w8(32'hba13dd72),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c5aea),
	.w1(32'h3ab9cba1),
	.w2(32'h3bd396b0),
	.w3(32'h3ba08afe),
	.w4(32'hbad2f692),
	.w5(32'h3bc3847e),
	.w6(32'hbb370ab5),
	.w7(32'hbbf9b598),
	.w8(32'h3bde3fff),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74724b),
	.w1(32'hba612b59),
	.w2(32'h39eb9056),
	.w3(32'h3bb4e24e),
	.w4(32'h39aa9bf9),
	.w5(32'h3b934867),
	.w6(32'h3c195e60),
	.w7(32'hba34facf),
	.w8(32'h3ad8d68f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa35bb),
	.w1(32'hb9e5306a),
	.w2(32'hbabf7869),
	.w3(32'h39ff4c49),
	.w4(32'hbb6dcbe3),
	.w5(32'h3b1bfe12),
	.w6(32'hba1bb025),
	.w7(32'hbafd0100),
	.w8(32'h3a7316da),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147b7e),
	.w1(32'h3aa88e4d),
	.w2(32'hbb62d4e5),
	.w3(32'h3c038200),
	.w4(32'hba1064fc),
	.w5(32'h3c0e3112),
	.w6(32'h3b9e0ada),
	.w7(32'hba255a9d),
	.w8(32'h3b003579),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba26c6),
	.w1(32'h3b689d02),
	.w2(32'h3be5dd69),
	.w3(32'h3bd48193),
	.w4(32'h3c2308ef),
	.w5(32'h3ba0f238),
	.w6(32'h3c1c4ae0),
	.w7(32'h3a7f6b14),
	.w8(32'hb778fa0c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee222),
	.w1(32'hbbc708b6),
	.w2(32'h3af4fbee),
	.w3(32'h3b1dce98),
	.w4(32'hbb70a342),
	.w5(32'h3c0276b7),
	.w6(32'hbb25a140),
	.w7(32'hbb127a42),
	.w8(32'h3baf143e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3572d),
	.w1(32'hbb25f173),
	.w2(32'h3b83f3f2),
	.w3(32'h3a914f01),
	.w4(32'h3adb6e67),
	.w5(32'h3c4a6059),
	.w6(32'h3b9a8c88),
	.w7(32'hbae28f09),
	.w8(32'hbb06b39a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53e772),
	.w1(32'h3bd7d300),
	.w2(32'h3c0df25e),
	.w3(32'h3bbeaa7a),
	.w4(32'hbaf92f39),
	.w5(32'h3b0cbfce),
	.w6(32'hbb9db17b),
	.w7(32'hbb25800d),
	.w8(32'h3a9e607d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa63875),
	.w1(32'hb9f5c8ad),
	.w2(32'h3a1f7c4a),
	.w3(32'hbabfb24a),
	.w4(32'h3b62d135),
	.w5(32'h3aee6491),
	.w6(32'h3a8fd4a6),
	.w7(32'hba92d8f1),
	.w8(32'hbb01ffdd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b1824),
	.w1(32'hba0c4ac1),
	.w2(32'hbb7c8b47),
	.w3(32'h3bec6d34),
	.w4(32'hbbfa3073),
	.w5(32'hbc2e1dff),
	.w6(32'h3bbc59f3),
	.w7(32'hbc0716ee),
	.w8(32'hba91e1ca),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4ca27),
	.w1(32'h3ad8216d),
	.w2(32'h3c07e1cd),
	.w3(32'h3a80dcda),
	.w4(32'h3ba306ac),
	.w5(32'h3958410f),
	.w6(32'h3b3c58e9),
	.w7(32'hb988d2b4),
	.w8(32'h3b0cd541),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af017c4),
	.w1(32'h3a604142),
	.w2(32'hb92ad117),
	.w3(32'h3b3632a2),
	.w4(32'hbb0f11ef),
	.w5(32'h3aadd6bf),
	.w6(32'hbacb7758),
	.w7(32'h384df35f),
	.w8(32'h3adaa640),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390756c1),
	.w1(32'h3944f608),
	.w2(32'h3a5c6d97),
	.w3(32'h3af95d24),
	.w4(32'h3b633ec4),
	.w5(32'hbaf0de70),
	.w6(32'h3ba51d1d),
	.w7(32'hba8bcf1b),
	.w8(32'h3a92ce7b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0959a1),
	.w1(32'h3bb0f951),
	.w2(32'h3b7a7109),
	.w3(32'h3bd5bacd),
	.w4(32'h3b20736d),
	.w5(32'h3a42181d),
	.w6(32'h3b64387b),
	.w7(32'h3a4ebfc8),
	.w8(32'hbab8bc09),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1123ff),
	.w1(32'h3b0e4563),
	.w2(32'h3aa6917b),
	.w3(32'hba279647),
	.w4(32'h3a63a99b),
	.w5(32'h3bad64bb),
	.w6(32'hba54ca08),
	.w7(32'hb8dad33a),
	.w8(32'hbb4e99cc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba583de),
	.w1(32'hbb063e11),
	.w2(32'h3b190e39),
	.w3(32'h3b18c4be),
	.w4(32'hbb583c3c),
	.w5(32'hba75862e),
	.w6(32'hb88888e8),
	.w7(32'hbb25aa11),
	.w8(32'hba8cb0b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f246),
	.w1(32'h3a9cee7d),
	.w2(32'h3b59f7cd),
	.w3(32'hbb53d11e),
	.w4(32'h38fd83e4),
	.w5(32'hbb65d5ef),
	.w6(32'h3b85fd92),
	.w7(32'h392e582b),
	.w8(32'hbabc6921),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1418b2),
	.w1(32'hbb6ed25a),
	.w2(32'h3bf739c5),
	.w3(32'h3ac7d012),
	.w4(32'h3c1bf8cd),
	.w5(32'h3b90724a),
	.w6(32'h3a648592),
	.w7(32'h3af4bd87),
	.w8(32'hbb2a2646),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bfc34),
	.w1(32'h39b17d11),
	.w2(32'h3b19bd30),
	.w3(32'h3b9da16c),
	.w4(32'hbbb499f3),
	.w5(32'h3b7b7607),
	.w6(32'h3a06cf9e),
	.w7(32'hbb594a59),
	.w8(32'h3b58a7b5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987317),
	.w1(32'h3b1a9ed7),
	.w2(32'hbaf38237),
	.w3(32'h3aed7e22),
	.w4(32'h3ae1f5b8),
	.w5(32'hbbaf08fe),
	.w6(32'h3b86df4b),
	.w7(32'h3b8492eb),
	.w8(32'hbb2b67ba),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4c7de),
	.w1(32'h3c03b334),
	.w2(32'h3c47a9d8),
	.w3(32'hbaacdca4),
	.w4(32'h3b4d2aa1),
	.w5(32'h3bb02883),
	.w6(32'hbb0558fe),
	.w7(32'hbb0fbf61),
	.w8(32'hbb36a049),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b264a),
	.w1(32'hb99a8ff2),
	.w2(32'h39ce3f0e),
	.w3(32'h3a64df8f),
	.w4(32'hbb2e987f),
	.w5(32'hb9dcd194),
	.w6(32'hb7dffbcf),
	.w7(32'hbb00fa6a),
	.w8(32'h3b62a687),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8733ab),
	.w1(32'hb990d055),
	.w2(32'hbbaa404d),
	.w3(32'h3afd55ec),
	.w4(32'hbbf9dfab),
	.w5(32'hba8171a2),
	.w6(32'h3aa5f402),
	.w7(32'hbb6849d7),
	.w8(32'hbc060394),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d55a),
	.w1(32'h3b0f950b),
	.w2(32'h3b6991f6),
	.w3(32'hbbc76745),
	.w4(32'h3b800339),
	.w5(32'h3bd5b876),
	.w6(32'hbad848d9),
	.w7(32'h3be64cdb),
	.w8(32'h3c51fd65),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42dc96),
	.w1(32'h3beac709),
	.w2(32'h3bc20025),
	.w3(32'h3b96b84e),
	.w4(32'h3bb09330),
	.w5(32'h3bdda66b),
	.w6(32'h3ade8327),
	.w7(32'h3af62fa9),
	.w8(32'h3b7e7e5b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fa70c),
	.w1(32'hba026d84),
	.w2(32'h3ba53931),
	.w3(32'h3a6c4a62),
	.w4(32'hbbaab642),
	.w5(32'hb9902c1c),
	.w6(32'hbb29ebea),
	.w7(32'hbb350198),
	.w8(32'hba857f1a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390409),
	.w1(32'h3a73a587),
	.w2(32'h3b034540),
	.w3(32'h3b96eae5),
	.w4(32'hba909662),
	.w5(32'hb7d2937b),
	.w6(32'h3b8ffc19),
	.w7(32'hbad39fc0),
	.w8(32'hbb55be10),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8aa4f),
	.w1(32'h3b1ee902),
	.w2(32'h3b903a56),
	.w3(32'hb96ca53d),
	.w4(32'h3a80a43d),
	.w5(32'h3a876b1b),
	.w6(32'h3acdc99a),
	.w7(32'h39c23370),
	.w8(32'h3b29568f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedd5bb),
	.w1(32'hba5603ae),
	.w2(32'h3a3aa62f),
	.w3(32'hb971dc9a),
	.w4(32'hbaf4ae34),
	.w5(32'hbb76c561),
	.w6(32'h3b84bea4),
	.w7(32'hbb68ad62),
	.w8(32'hbb212523),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3d0c8),
	.w1(32'h3b030f37),
	.w2(32'h3b98f7fd),
	.w3(32'hba941781),
	.w4(32'hbaf07356),
	.w5(32'hbb4a7f5f),
	.w6(32'hbae935d1),
	.w7(32'hbadf1bde),
	.w8(32'h3b6b3827),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aef3e),
	.w1(32'h398ae9be),
	.w2(32'h3ae45b80),
	.w3(32'h3b89f976),
	.w4(32'h3be276e7),
	.w5(32'h3c4121e4),
	.w6(32'h3b0466ca),
	.w7(32'h3b8035c3),
	.w8(32'h3be0f1f3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14881f),
	.w1(32'h3a7ba756),
	.w2(32'h3812abcc),
	.w3(32'h3babbc7d),
	.w4(32'hba9e9cbe),
	.w5(32'hba2455e9),
	.w6(32'h3bc9b892),
	.w7(32'hbb082aa5),
	.w8(32'hbbe24c3c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe3f83),
	.w1(32'h3b333366),
	.w2(32'h3bb04b8f),
	.w3(32'h3b8ee8d2),
	.w4(32'h3b9e3d02),
	.w5(32'h3b4a5dd3),
	.w6(32'hbbdba073),
	.w7(32'hbac70de1),
	.w8(32'h3b48db50),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2b316),
	.w1(32'hbb28847f),
	.w2(32'h3bc22001),
	.w3(32'h3983beac),
	.w4(32'h3b13b517),
	.w5(32'h3ad77d2b),
	.w6(32'h3bbfd749),
	.w7(32'hba997a08),
	.w8(32'h3a724909),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83793f),
	.w1(32'hbaee0702),
	.w2(32'h393f3894),
	.w3(32'h3af222e6),
	.w4(32'hbbb66de9),
	.w5(32'hbb2848af),
	.w6(32'hb999681c),
	.w7(32'hbbf4644a),
	.w8(32'hbb7887eb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4bcd8),
	.w1(32'h3adc93c4),
	.w2(32'h3a2cd417),
	.w3(32'hba9dd74b),
	.w4(32'hba0384a0),
	.w5(32'h3b0659c1),
	.w6(32'hb94d47be),
	.w7(32'h398dc16b),
	.w8(32'h3b3252e2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967f23e),
	.w1(32'h3a904a7f),
	.w2(32'h399a8a9f),
	.w3(32'hb96bda30),
	.w4(32'hbb2804ae),
	.w5(32'hba1a7c36),
	.w6(32'h3abcffbf),
	.w7(32'h3ae52502),
	.w8(32'h3b517cd1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a8664),
	.w1(32'hbb6bdbed),
	.w2(32'h3aa1e36b),
	.w3(32'h3be442aa),
	.w4(32'hbb1a4a07),
	.w5(32'h3b3b8f4c),
	.w6(32'h3a8be937),
	.w7(32'hbb914a93),
	.w8(32'h3c01bffe),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba055c2),
	.w1(32'h3ba69bc4),
	.w2(32'h3bb33172),
	.w3(32'h3be9fa22),
	.w4(32'hba91ff46),
	.w5(32'h3b8ba296),
	.w6(32'h3c0bcfef),
	.w7(32'hba5a35a1),
	.w8(32'h38a6b822),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6469c5),
	.w1(32'h39c05ee9),
	.w2(32'hbb402f63),
	.w3(32'h3c18ef7e),
	.w4(32'hbb06fc5a),
	.w5(32'h3c08b6d7),
	.w6(32'hbaa20927),
	.w7(32'h3a3fc6f7),
	.w8(32'hb961522b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ecf7),
	.w1(32'hbb2b4ea5),
	.w2(32'hbb288521),
	.w3(32'h3badb781),
	.w4(32'hba84cde5),
	.w5(32'h3b8d82d8),
	.w6(32'h3b9a7ba8),
	.w7(32'hbb8a8476),
	.w8(32'hb9360617),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba04b4d),
	.w1(32'h3a839610),
	.w2(32'h3af1e3d7),
	.w3(32'h3b1c2f1b),
	.w4(32'h39583095),
	.w5(32'h3b517a30),
	.w6(32'h3b31b111),
	.w7(32'h3a423a0a),
	.w8(32'h39fd146c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc46e97),
	.w1(32'h3bd91958),
	.w2(32'h3bc87085),
	.w3(32'h3bc7995c),
	.w4(32'hba864b1c),
	.w5(32'hbb8bd01f),
	.w6(32'h3ba2251e),
	.w7(32'hb9f5cb17),
	.w8(32'h3b8d18f5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa62a7),
	.w1(32'h3be3e239),
	.w2(32'h3c00a244),
	.w3(32'h3b9f06fe),
	.w4(32'h3b00bf4e),
	.w5(32'h3af39345),
	.w6(32'h3c17ebca),
	.w7(32'h3a74c805),
	.w8(32'h3c006d7d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b513ebe),
	.w1(32'h3b581c82),
	.w2(32'hba5baabd),
	.w3(32'hbaa645a5),
	.w4(32'hba8e550a),
	.w5(32'hbbbe7e68),
	.w6(32'hbad77e94),
	.w7(32'hb9d04fd8),
	.w8(32'hbacdb3e8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dba7a),
	.w1(32'h3b50b187),
	.w2(32'h3bb64344),
	.w3(32'h3bc2bfc5),
	.w4(32'h3b508a6a),
	.w5(32'hb91a458b),
	.w6(32'hbb844cb3),
	.w7(32'h39442e15),
	.w8(32'h3bbd157c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8018a0d),
	.w1(32'h3bb20fc3),
	.w2(32'h3be06536),
	.w3(32'h3c15c080),
	.w4(32'h3ba24d6f),
	.w5(32'h3b9bb66b),
	.w6(32'hba741721),
	.w7(32'h3b80ae3f),
	.w8(32'h3c071955),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a062f2b),
	.w1(32'h3c0c82a2),
	.w2(32'h3c5a9435),
	.w3(32'h3bf4ac7b),
	.w4(32'h3b8a8b43),
	.w5(32'h3bbf5e46),
	.w6(32'h3c32f1fb),
	.w7(32'h3ae9bb4e),
	.w8(32'h3ba3017d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f760),
	.w1(32'hbc0802e7),
	.w2(32'h3bcaed64),
	.w3(32'h3b271962),
	.w4(32'hbc1343f6),
	.w5(32'hbb934dc0),
	.w6(32'h3b38702f),
	.w7(32'hbc049da5),
	.w8(32'h3b9d79b2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818308),
	.w1(32'hbaa60f60),
	.w2(32'hba42a495),
	.w3(32'h3b8ca43d),
	.w4(32'h3ace91fa),
	.w5(32'hbb3c782c),
	.w6(32'h3c0d61e9),
	.w7(32'h3b5856ce),
	.w8(32'h3a8ecc06),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af163de),
	.w1(32'h3ba4ae64),
	.w2(32'hbb13a4a5),
	.w3(32'h3b606683),
	.w4(32'h3734f990),
	.w5(32'hbb840abe),
	.w6(32'h3bd25ae0),
	.w7(32'h3a999b1c),
	.w8(32'h3be9e340),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9b3dc),
	.w1(32'hb7cfd7e9),
	.w2(32'h3c0552d0),
	.w3(32'h3b0b2d17),
	.w4(32'h3bb13068),
	.w5(32'h3bca24fd),
	.w6(32'h3aadb7d8),
	.w7(32'hb77a75a2),
	.w8(32'hbaef4cc1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08f8b6),
	.w1(32'h3af0e7c8),
	.w2(32'h3bc6dcc4),
	.w3(32'h3b080643),
	.w4(32'hbb8062ef),
	.w5(32'h3ac1f1fe),
	.w6(32'h3b5bf02a),
	.w7(32'hbb6a1477),
	.w8(32'hbbc73ee5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10941a),
	.w1(32'hbba9f3ff),
	.w2(32'hbbe61d9b),
	.w3(32'hbbd64840),
	.w4(32'hbc112a86),
	.w5(32'hbc077656),
	.w6(32'hbb4ef480),
	.w7(32'hbbc2a22d),
	.w8(32'hbbb135e9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc34f21),
	.w1(32'h3ae00148),
	.w2(32'h3b29f6e4),
	.w3(32'hba0f45c1),
	.w4(32'h3b90bb93),
	.w5(32'h3bb69a82),
	.w6(32'hba5fbfc6),
	.w7(32'hbb8ab957),
	.w8(32'hbaf1c8ef),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb0ee9),
	.w1(32'h3a3eca49),
	.w2(32'h3b24a479),
	.w3(32'h3b60d05a),
	.w4(32'hbb4f51b0),
	.w5(32'h3acac277),
	.w6(32'hb80cb0a0),
	.w7(32'hbb9101a6),
	.w8(32'hbb19b156),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d424),
	.w1(32'h3a555b67),
	.w2(32'h3ad3f851),
	.w3(32'h39df34e7),
	.w4(32'h3ad22753),
	.w5(32'hbb0d5ddf),
	.w6(32'h39cd4870),
	.w7(32'hbaa36452),
	.w8(32'h3a1e098c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af85feb),
	.w1(32'h3b48c1f7),
	.w2(32'h3c821f7f),
	.w3(32'hbabed5d3),
	.w4(32'h3c37ff2c),
	.w5(32'h3c63234c),
	.w6(32'h3a1194b3),
	.w7(32'hb68dac58),
	.w8(32'hbae77e56),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c232c5f),
	.w1(32'hba8ef90a),
	.w2(32'hbab696ac),
	.w3(32'h3bbb7ada),
	.w4(32'hbb12df41),
	.w5(32'hbbda332b),
	.w6(32'h3b3b614b),
	.w7(32'hbb598dc1),
	.w8(32'h3a7ad53a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0154cd),
	.w1(32'h3b6e4438),
	.w2(32'h3b3b4dab),
	.w3(32'hbad63bcb),
	.w4(32'h3aa39bfc),
	.w5(32'h3b9801f4),
	.w6(32'h3b55c540),
	.w7(32'h3bac8e21),
	.w8(32'h38e268ff),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96cd3e),
	.w1(32'hb87d29e3),
	.w2(32'hbb086c0d),
	.w3(32'hba8e4ae6),
	.w4(32'hbb05a8d5),
	.w5(32'hbad10ce5),
	.w6(32'h3a12ff9f),
	.w7(32'hbb712d38),
	.w8(32'hbb5d3d48),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb896e),
	.w1(32'hbad6736a),
	.w2(32'hba0c2cb4),
	.w3(32'hbb22cb8b),
	.w4(32'hbaee7c6c),
	.w5(32'hb8590426),
	.w6(32'hbbac59e1),
	.w7(32'hbac1837a),
	.w8(32'hbb73d27b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dc801),
	.w1(32'h3b33a800),
	.w2(32'hb9d5d50f),
	.w3(32'hb703b144),
	.w4(32'h3bd5d808),
	.w5(32'h3bf21530),
	.w6(32'hbb5ac101),
	.w7(32'h3a7197d1),
	.w8(32'hbb19ad6c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b288e94),
	.w1(32'hba8fd036),
	.w2(32'h3b54bb3a),
	.w3(32'hba626bf6),
	.w4(32'h3a1cd32e),
	.w5(32'hbb5a2b7f),
	.w6(32'h3b0615a2),
	.w7(32'h3a2b11fd),
	.w8(32'h3b443ed7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd79528),
	.w1(32'h3b1b77c6),
	.w2(32'h3b0c76b2),
	.w3(32'h3b75e034),
	.w4(32'hbb5c79b8),
	.w5(32'hbb1e7204),
	.w6(32'h3bc495ca),
	.w7(32'h3b2e1700),
	.w8(32'h3c4caa78),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c3deba),
	.w1(32'hbb07bcce),
	.w2(32'hbb263b8a),
	.w3(32'h3985b151),
	.w4(32'hbb7b5b2a),
	.w5(32'hbb22764b),
	.w6(32'h3a55a72b),
	.w7(32'hbac1b1cc),
	.w8(32'h3955d8f5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fe9ae),
	.w1(32'h3bd19844),
	.w2(32'h3c17e925),
	.w3(32'h3bd7f203),
	.w4(32'h3b8234ca),
	.w5(32'h3c0b778b),
	.w6(32'h3a88623d),
	.w7(32'h3b978adb),
	.w8(32'h3bff89e7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38661f),
	.w1(32'hbb87f014),
	.w2(32'hbb88222b),
	.w3(32'h3a398bce),
	.w4(32'hbb80a3e2),
	.w5(32'hbc58a408),
	.w6(32'hba10ef4f),
	.w7(32'hbb959404),
	.w8(32'hbb469024),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d9457),
	.w1(32'h3b862dad),
	.w2(32'h3b9fa13a),
	.w3(32'h3a20b249),
	.w4(32'h3b6d009f),
	.w5(32'h3979fc6d),
	.w6(32'h3afe029a),
	.w7(32'h3bc9020e),
	.w8(32'h3b8e7765),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f396a),
	.w1(32'hba3ec8d0),
	.w2(32'h3b63e0c9),
	.w3(32'hba08a5da),
	.w4(32'hbb0caecc),
	.w5(32'h3ca5c562),
	.w6(32'h3bb0fc2a),
	.w7(32'hbb2b6557),
	.w8(32'h3a9d6622),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c225874),
	.w1(32'hb995e2ad),
	.w2(32'h39741c63),
	.w3(32'h3c00c6ef),
	.w4(32'h3b891870),
	.w5(32'h3c80e137),
	.w6(32'h3b73f12a),
	.w7(32'h3b9bcc2e),
	.w8(32'h3c4d6e8d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae7873),
	.w1(32'h3b822f95),
	.w2(32'h3b39ad84),
	.w3(32'h3bdea083),
	.w4(32'h3baa7f12),
	.w5(32'h3c48fd00),
	.w6(32'h3a036945),
	.w7(32'hb94c90d4),
	.w8(32'hba7e6195),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6cae),
	.w1(32'h3b025119),
	.w2(32'hb8f0dba4),
	.w3(32'h3a823e73),
	.w4(32'h3b19f65f),
	.w5(32'h3b0f5128),
	.w6(32'h398a6ad3),
	.w7(32'h3a4144fa),
	.w8(32'h3b23127f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8576a13),
	.w1(32'hb9c1c724),
	.w2(32'hbb8c1cf4),
	.w3(32'hb793964b),
	.w4(32'h3881c2d0),
	.w5(32'h3b147420),
	.w6(32'h39c709e3),
	.w7(32'hbaecd242),
	.w8(32'hbb719ab4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14d61c),
	.w1(32'h3ae6372a),
	.w2(32'h3ae243c2),
	.w3(32'h3b321a50),
	.w4(32'h3a04367d),
	.w5(32'hbbc34753),
	.w6(32'h3a0a246d),
	.w7(32'hbb185f50),
	.w8(32'h39e5fc74),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83a486),
	.w1(32'h3b90f49c),
	.w2(32'h3a9ee01d),
	.w3(32'h3b128852),
	.w4(32'h3a06397d),
	.w5(32'hbaca5ca3),
	.w6(32'h3ba494f7),
	.w7(32'h3b62f5e0),
	.w8(32'hba54975d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc9add),
	.w1(32'h3a133237),
	.w2(32'h3b313d6e),
	.w3(32'h3bf0c691),
	.w4(32'h3b8117e6),
	.w5(32'h3b7dc5b2),
	.w6(32'h3ba06828),
	.w7(32'h3b019f92),
	.w8(32'h3929de24),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ded73),
	.w1(32'h3b85af03),
	.w2(32'h3b4c932a),
	.w3(32'h3a31b7ee),
	.w4(32'h3b7696d0),
	.w5(32'hbb141043),
	.w6(32'h383ac102),
	.w7(32'h3b625664),
	.w8(32'hb988cbd2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae895ca),
	.w1(32'hbaddd104),
	.w2(32'hbaa6b5b1),
	.w3(32'h3af2016c),
	.w4(32'hbb361ad4),
	.w5(32'h3b654eba),
	.w6(32'hbb5b0321),
	.w7(32'hbaa68d19),
	.w8(32'h3a06ead7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a200866),
	.w1(32'hbaca5b41),
	.w2(32'h3abca383),
	.w3(32'h3a76acbe),
	.w4(32'hbbb05c40),
	.w5(32'hba848dd0),
	.w6(32'hbaa1d2ab),
	.w7(32'hbb2de237),
	.w8(32'h3a624fff),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61e0c7),
	.w1(32'hb916b936),
	.w2(32'h3b17905e),
	.w3(32'h3bc20377),
	.w4(32'hba8f0c7c),
	.w5(32'hbb9353e3),
	.w6(32'h3bc4dc41),
	.w7(32'hb9e16f95),
	.w8(32'h3b1812bf),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa496d3),
	.w1(32'hbad179bc),
	.w2(32'h3bbce2da),
	.w3(32'h3aa4cf2b),
	.w4(32'hb98a0029),
	.w5(32'h3b86dca4),
	.w6(32'hb9f2f51e),
	.w7(32'hba5d763a),
	.w8(32'h3b56402c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee66c),
	.w1(32'h3aa51388),
	.w2(32'hba726b60),
	.w3(32'h3a6c391d),
	.w4(32'h3bed816d),
	.w5(32'hbb128749),
	.w6(32'h3978cdaf),
	.w7(32'hb865419d),
	.w8(32'hb95bbf20),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237eb6),
	.w1(32'hbbd39b06),
	.w2(32'hb998abb4),
	.w3(32'hbb317f13),
	.w4(32'h3ab138c3),
	.w5(32'h3c40ea4c),
	.w6(32'hbbaf52e4),
	.w7(32'hb938a170),
	.w8(32'h3c0dc393),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32d737),
	.w1(32'h3b42a33e),
	.w2(32'h3b1d0348),
	.w3(32'h3bf4688e),
	.w4(32'h3b59cb0e),
	.w5(32'h3cc44ac2),
	.w6(32'h3b6e6588),
	.w7(32'h3aa3eab2),
	.w8(32'h3c253e1b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3979a3),
	.w1(32'h3aff5a68),
	.w2(32'h3ae4583d),
	.w3(32'h3c6a55cd),
	.w4(32'h3aa7673c),
	.w5(32'hbacd4b97),
	.w6(32'h3b9b7fcc),
	.w7(32'h3ab6aca0),
	.w8(32'h3a0f1869),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e7068),
	.w1(32'h3ba2f027),
	.w2(32'h3bef2765),
	.w3(32'h3ababc4c),
	.w4(32'h3b5be484),
	.w5(32'h39bce5b0),
	.w6(32'h3ac292e1),
	.w7(32'h3bdeca08),
	.w8(32'h3b9cbbbc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90bded),
	.w1(32'h3a0d2113),
	.w2(32'hbaccec4e),
	.w3(32'hbad2e183),
	.w4(32'hbb6cb2c2),
	.w5(32'hbba8e0e3),
	.w6(32'h3935516a),
	.w7(32'hbb9597d2),
	.w8(32'hb9a86025),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a388ab),
	.w1(32'h3b33d30d),
	.w2(32'hbad7cd6b),
	.w3(32'h3aea9ccb),
	.w4(32'h3b7b48c8),
	.w5(32'hbad33c2b),
	.w6(32'h3b998aa3),
	.w7(32'h3bb3b277),
	.w8(32'h3bd31814),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f5038),
	.w1(32'hba93ab51),
	.w2(32'hba44fb60),
	.w3(32'h3a38910e),
	.w4(32'h3915d533),
	.w5(32'h3b382132),
	.w6(32'h3b940d21),
	.w7(32'hba0b5edb),
	.w8(32'hba14fd4d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eff1d),
	.w1(32'h3a9b1a8b),
	.w2(32'h3a7d5b6d),
	.w3(32'h3ade8159),
	.w4(32'hbb3e4666),
	.w5(32'hbb11a933),
	.w6(32'h3b70c021),
	.w7(32'h3926725e),
	.w8(32'h3b9bbeef),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fe7d4),
	.w1(32'h3baaf553),
	.w2(32'h3c6f4020),
	.w3(32'h3adb8cce),
	.w4(32'h3b718939),
	.w5(32'h3d388ab6),
	.w6(32'h3aed6c99),
	.w7(32'hbb31d230),
	.w8(32'h3b8d9dad),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb5384),
	.w1(32'hbb72301d),
	.w2(32'hbb1e5e1e),
	.w3(32'h3cb141ab),
	.w4(32'hbb479fde),
	.w5(32'hb8c6a359),
	.w6(32'h3c01aeba),
	.w7(32'hbc346f9a),
	.w8(32'hbc2ccb8e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a166bfd),
	.w1(32'hbbbeb276),
	.w2(32'h3b1c0237),
	.w3(32'h3af7f867),
	.w4(32'hbbb6aa0e),
	.w5(32'h3ab819a2),
	.w6(32'h3a8cc506),
	.w7(32'hbbb96624),
	.w8(32'h3b45e1a9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfea8b),
	.w1(32'h3b1ddcaa),
	.w2(32'hbbf52251),
	.w3(32'h3b68d7d2),
	.w4(32'hba6f040b),
	.w5(32'hbc1aeb32),
	.w6(32'hb95b3a15),
	.w7(32'hbb7f9842),
	.w8(32'hbbf34288),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f300),
	.w1(32'h3c649d82),
	.w2(32'h3c86a646),
	.w3(32'hbc018b2e),
	.w4(32'h3caab3d6),
	.w5(32'h3cbb724e),
	.w6(32'hbbb0afd6),
	.w7(32'h3c7991d8),
	.w8(32'h3c5e3f70),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c416483),
	.w1(32'hbb0474b5),
	.w2(32'hbb157c70),
	.w3(32'h3c89287d),
	.w4(32'hbb0b18ff),
	.w5(32'h3adda20f),
	.w6(32'h3bc947e1),
	.w7(32'h3bba7828),
	.w8(32'h3bbca406),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010c1a),
	.w1(32'h3c08e5cd),
	.w2(32'h3b351eb9),
	.w3(32'hbabef8dd),
	.w4(32'h3a2755f4),
	.w5(32'hbbbff296),
	.w6(32'hbb968c7a),
	.w7(32'hbb9a84b2),
	.w8(32'hbbb689b1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7901da),
	.w1(32'h3b746327),
	.w2(32'hb934903b),
	.w3(32'hbad24a02),
	.w4(32'hbbcdabac),
	.w5(32'hbc04d905),
	.w6(32'hbb0da76d),
	.w7(32'h3c464568),
	.w8(32'h3b88ef98),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b416cf5),
	.w1(32'hbba29b9c),
	.w2(32'hba0c2396),
	.w3(32'hbbb278ae),
	.w4(32'hbbb19454),
	.w5(32'hbc0a3322),
	.w6(32'h3c456cc9),
	.w7(32'h3a5a302c),
	.w8(32'h39263775),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf3f0),
	.w1(32'h3b08def9),
	.w2(32'h3b8739e3),
	.w3(32'hb84aa009),
	.w4(32'h3b90b545),
	.w5(32'h3be133d3),
	.w6(32'h3b13292e),
	.w7(32'hbaafb0c9),
	.w8(32'h3b145687),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5db869),
	.w1(32'hbccc0222),
	.w2(32'hbce6b098),
	.w3(32'hbb24c42a),
	.w4(32'hbd022f18),
	.w5(32'hbd35dd54),
	.w6(32'hba9e56a9),
	.w7(32'hbc518274),
	.w8(32'hbd117bd2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba59fe5),
	.w1(32'hbbd5b527),
	.w2(32'hba00d240),
	.w3(32'hbcdb9903),
	.w4(32'hbc0424e0),
	.w5(32'h3bd6a159),
	.w6(32'hbceaba52),
	.w7(32'hbc4f75eb),
	.w8(32'hbb0ee2b9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba551f9a),
	.w1(32'hbb7d4b21),
	.w2(32'h3a0fd60a),
	.w3(32'hba4daa6d),
	.w4(32'hbbadc462),
	.w5(32'h39ba0499),
	.w6(32'hba3c72f0),
	.w7(32'hbb9be177),
	.w8(32'hbb7d5cce),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09d946),
	.w1(32'hbbf58987),
	.w2(32'h3b312b2c),
	.w3(32'h3b18b20e),
	.w4(32'h3ba42053),
	.w5(32'h3cc14a4b),
	.w6(32'hbac369b0),
	.w7(32'hbbff18c2),
	.w8(32'h3c030aad),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84d3fe),
	.w1(32'h3b5e0543),
	.w2(32'h3acb3d15),
	.w3(32'hba1f5772),
	.w4(32'hbaadc1de),
	.w5(32'hbb02611e),
	.w6(32'hbc288a4a),
	.w7(32'hb9b3ebe2),
	.w8(32'h3a3c43f1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2db560),
	.w1(32'h3b5c6fa7),
	.w2(32'hbaf6c0b0),
	.w3(32'hbb2603b0),
	.w4(32'hbb9a1422),
	.w5(32'hbc101b5b),
	.w6(32'h3b79d2ef),
	.w7(32'hbbad3eac),
	.w8(32'hbc00a886),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3624dd),
	.w1(32'h3a02334e),
	.w2(32'h3aa62f2f),
	.w3(32'hbc0b5f0c),
	.w4(32'hbad76662),
	.w5(32'hbab07343),
	.w6(32'hbb17d3f0),
	.w7(32'hbb1d3b48),
	.w8(32'hba8b0172),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac30f7f),
	.w1(32'h3c158857),
	.w2(32'h3c9e4e1b),
	.w3(32'h39a6c5a9),
	.w4(32'h3b640f55),
	.w5(32'h3c29d2b6),
	.w6(32'hbbadf0f9),
	.w7(32'h3c1206c4),
	.w8(32'h3c6a4ca3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82b75d),
	.w1(32'h38447824),
	.w2(32'hbbacc2ca),
	.w3(32'h3c7b30a5),
	.w4(32'hbb86dc65),
	.w5(32'hbc4c7d30),
	.w6(32'h3c7e229a),
	.w7(32'hbb7a95b5),
	.w8(32'hbae0d305),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc255b5e),
	.w1(32'h3c808770),
	.w2(32'h3cb0aa5c),
	.w3(32'hbbb27a0a),
	.w4(32'h3cb3a454),
	.w5(32'h3cdebde1),
	.w6(32'hbb088b03),
	.w7(32'h3c2d7693),
	.w8(32'h3c9db9bf),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3068fa),
	.w1(32'h3c675e30),
	.w2(32'h3c2dbe37),
	.w3(32'h3caeea3a),
	.w4(32'h3cb180cc),
	.w5(32'h3c7a4702),
	.w6(32'h3c715337),
	.w7(32'h3c974000),
	.w8(32'h3c1e3ee8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fac8e),
	.w1(32'hbad3dc8c),
	.w2(32'h3a18ea01),
	.w3(32'h3c202014),
	.w4(32'h38ab27fd),
	.w5(32'h3b142bf5),
	.w6(32'h3b9c370c),
	.w7(32'hbb001121),
	.w8(32'h397c708d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5a8f8),
	.w1(32'hbb4c3029),
	.w2(32'hba807c9d),
	.w3(32'h38c06e61),
	.w4(32'hbb8d9c9a),
	.w5(32'hbc1f8fbb),
	.w6(32'h3aa49fa4),
	.w7(32'h3abab08d),
	.w8(32'hbb62a5ce),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad80d30),
	.w1(32'h3c673c93),
	.w2(32'h3b53d07d),
	.w3(32'hbb53542c),
	.w4(32'h3a36cdb4),
	.w5(32'hbbe99aa0),
	.w6(32'hba3631c7),
	.w7(32'h3c0fca0a),
	.w8(32'h3b9681bc),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dc9cd),
	.w1(32'h3c1c9b00),
	.w2(32'h3c015ca8),
	.w3(32'h3b846218),
	.w4(32'h3c167bfc),
	.w5(32'h3b3fb689),
	.w6(32'h3b4a8134),
	.w7(32'hbb08cd9e),
	.w8(32'h3b051c70),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad23ed),
	.w1(32'hbc0ad575),
	.w2(32'h3b19ef0d),
	.w3(32'hbac24030),
	.w4(32'hbbb718c1),
	.w5(32'h3c185ba6),
	.w6(32'hbaa03cfb),
	.w7(32'hbbc3335e),
	.w8(32'h3b9ce3c9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17d993),
	.w1(32'hbbd78452),
	.w2(32'h3a1881f2),
	.w3(32'h3bb47075),
	.w4(32'hbb831e35),
	.w5(32'h3b8fdad8),
	.w6(32'h3b5d2454),
	.w7(32'hbbec43d4),
	.w8(32'h3a301636),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14021d),
	.w1(32'h3b117d49),
	.w2(32'h3b36dc66),
	.w3(32'hbb7a315a),
	.w4(32'hba98d32a),
	.w5(32'h39d00087),
	.w6(32'hba4766f4),
	.w7(32'hbc15cd6b),
	.w8(32'hbc00cc71),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1689c9),
	.w1(32'hbc81ef29),
	.w2(32'hbcf93646),
	.w3(32'h3b22b735),
	.w4(32'hbcea6cae),
	.w5(32'hbd46d8a4),
	.w6(32'hbb6e449f),
	.w7(32'hbd024d01),
	.w8(32'hbd29047e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfd8f3a),
	.w1(32'hba0cc192),
	.w2(32'h3bf4a050),
	.w3(32'hbceeeb5a),
	.w4(32'h3c449537),
	.w5(32'h3c57fd4b),
	.w6(32'hbcc843af),
	.w7(32'h3ca6003a),
	.w8(32'h3cbd4fcd),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23380c),
	.w1(32'h3aca40cd),
	.w2(32'h3b34e7b6),
	.w3(32'h3c78f69d),
	.w4(32'h3b836d05),
	.w5(32'h3b51b99e),
	.w6(32'h3ca372ac),
	.w7(32'h3ab36a40),
	.w8(32'h3b30781c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9149f0),
	.w1(32'h3a1a4c7b),
	.w2(32'hba915126),
	.w3(32'h3c072d8c),
	.w4(32'h3beac2b7),
	.w5(32'h3b840302),
	.w6(32'h3c23cc0d),
	.w7(32'h3b6f1c1c),
	.w8(32'h3bef893f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1af18),
	.w1(32'hbb19b0f1),
	.w2(32'h389ecc49),
	.w3(32'h3b824483),
	.w4(32'hbbb115ed),
	.w5(32'hbba8f27b),
	.w6(32'h3b871326),
	.w7(32'h3b5ad88c),
	.w8(32'hba52b66a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75049f),
	.w1(32'h3c39cc3e),
	.w2(32'h3c4a2579),
	.w3(32'hba14fcc7),
	.w4(32'h3c7313d2),
	.w5(32'h3c956e39),
	.w6(32'hbb1625d6),
	.w7(32'h3c2d7866),
	.w8(32'h3c1c118b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27dd83),
	.w1(32'h3c66453b),
	.w2(32'h3c3e0fa5),
	.w3(32'h3c8e2b0c),
	.w4(32'h3beccf39),
	.w5(32'h3b4c6600),
	.w6(32'h3c09eb62),
	.w7(32'h3c3608ae),
	.w8(32'h3c36c7ca),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e7f23),
	.w1(32'hba4306ed),
	.w2(32'h3a4a7c7a),
	.w3(32'h3bb03980),
	.w4(32'hbacc59aa),
	.w5(32'hbc0faebd),
	.w6(32'h3c14b825),
	.w7(32'hbc264d60),
	.w8(32'hbc201365),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fad67),
	.w1(32'hbad68f76),
	.w2(32'h3b101ccf),
	.w3(32'hbc6109f9),
	.w4(32'h3a914034),
	.w5(32'hbb58df8e),
	.w6(32'hbbb466e8),
	.w7(32'hbb92d397),
	.w8(32'hbb078a37),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99764c3),
	.w1(32'hbc012739),
	.w2(32'hbc59a759),
	.w3(32'h3b398305),
	.w4(32'hbcf4fce3),
	.w5(32'hbd0e3a1b),
	.w6(32'hb8804e4c),
	.w7(32'hbce6c26a),
	.w8(32'hbce36f84),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca06111),
	.w1(32'hbb4af72a),
	.w2(32'hba14649c),
	.w3(32'hbcf6ecdf),
	.w4(32'hbb4c37d5),
	.w5(32'hbbca620c),
	.w6(32'hbccf5724),
	.w7(32'h38e71a6a),
	.w8(32'h3b5bbd68),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b961ed),
	.w1(32'hbc4922eb),
	.w2(32'hbc2acbbc),
	.w3(32'hbb422f4b),
	.w4(32'hbc3d0efe),
	.w5(32'hbc1de36a),
	.w6(32'h3bfb5ddd),
	.w7(32'hbbea6054),
	.w8(32'hbc25731c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15fb75),
	.w1(32'h3b5d7bc9),
	.w2(32'hb9ad9149),
	.w3(32'hbbeeb754),
	.w4(32'h3b32e981),
	.w5(32'hbba131a5),
	.w6(32'hbc169d62),
	.w7(32'h3c08c3f8),
	.w8(32'h3ad27e2d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97b797),
	.w1(32'hba1321fa),
	.w2(32'h399a823d),
	.w3(32'h39c48fbe),
	.w4(32'hbac97150),
	.w5(32'hbb8c2d59),
	.w6(32'h3a2f485e),
	.w7(32'hbb5a9efb),
	.w8(32'h39295a16),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad49abc),
	.w1(32'hbc963bcb),
	.w2(32'hbcb963b9),
	.w3(32'hbb0767e0),
	.w4(32'hbcdfb6ff),
	.w5(32'hbd11963d),
	.w6(32'h3a00376f),
	.w7(32'hbc4cf584),
	.w8(32'hbcd1a800),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3be5bc),
	.w1(32'hbbbaeb80),
	.w2(32'h3a19de19),
	.w3(32'hbc9d510d),
	.w4(32'h3ae2db12),
	.w5(32'hbbce2ae1),
	.w6(32'hbcda2f0f),
	.w7(32'h3b4e16da),
	.w8(32'h3b35c6d7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1599bf),
	.w1(32'h397e6703),
	.w2(32'h3bf313a4),
	.w3(32'h3bed0631),
	.w4(32'h3a60528d),
	.w5(32'h3bbb2594),
	.w6(32'h3c0b73b2),
	.w7(32'hbbad7701),
	.w8(32'h3b756744),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2572),
	.w1(32'hbb720c9c),
	.w2(32'hba5ac744),
	.w3(32'h3b93c1a1),
	.w4(32'h3a99dd8a),
	.w5(32'h3b731aef),
	.w6(32'h3b669780),
	.w7(32'hb911be08),
	.w8(32'h3b62edee),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d196),
	.w1(32'hb98d473c),
	.w2(32'h3bce2b36),
	.w3(32'h3b102dfb),
	.w4(32'hbb3d879c),
	.w5(32'h3b4c4a8b),
	.w6(32'hb83556c6),
	.w7(32'hbaf884ec),
	.w8(32'h3c01881a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65a0c8),
	.w1(32'hbb9a038b),
	.w2(32'h397636a4),
	.w3(32'hbb4491b0),
	.w4(32'hbbefe879),
	.w5(32'h3c319a1f),
	.w6(32'hbb9731c7),
	.w7(32'hbc07a7df),
	.w8(32'h3c157490),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29bc90),
	.w1(32'hbc1c64d2),
	.w2(32'hbb2228e8),
	.w3(32'h3c06c0ee),
	.w4(32'hbc297c12),
	.w5(32'hbb9bdc9e),
	.w6(32'h3b77a7f5),
	.w7(32'hbbcf391f),
	.w8(32'hb9b78b49),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe93e80),
	.w1(32'hbb309458),
	.w2(32'hbbb36fe4),
	.w3(32'hbbbe6c40),
	.w4(32'h3b1e5adb),
	.w5(32'h3b417062),
	.w6(32'hb95cc290),
	.w7(32'h3b230bc5),
	.w8(32'h3ba2c47b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e6f3),
	.w1(32'hba8aa72b),
	.w2(32'hbb7f233c),
	.w3(32'h3bc31ded),
	.w4(32'h3bd0fa10),
	.w5(32'h3c1415d8),
	.w6(32'h3b2e9688),
	.w7(32'h3b71bf18),
	.w8(32'h3b2579dd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d4423),
	.w1(32'h3af99278),
	.w2(32'hba6b8b64),
	.w3(32'h3b2c0b34),
	.w4(32'hbc1788c7),
	.w5(32'hbc72a04d),
	.w6(32'h3b98ff71),
	.w7(32'hbb338264),
	.w8(32'hbc1af7b6),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4c1db),
	.w1(32'hbaad5022),
	.w2(32'hbbf949ba),
	.w3(32'hbc5c9560),
	.w4(32'h3b2663e2),
	.w5(32'hbc3a25da),
	.w6(32'hbc07ed2e),
	.w7(32'h3a8ca982),
	.w8(32'hbbef2436),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb13d47),
	.w1(32'hbba15424),
	.w2(32'h392a721f),
	.w3(32'hbbba1dd6),
	.w4(32'hbab95801),
	.w5(32'h3bacd61e),
	.w6(32'hba37fac5),
	.w7(32'hbb9621f4),
	.w8(32'h3a367ae3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba58ad1),
	.w1(32'hb984974e),
	.w2(32'h3b7ad7a9),
	.w3(32'h39a9ca01),
	.w4(32'hbb527778),
	.w5(32'hbbe9ad7e),
	.w6(32'hbc1aaa40),
	.w7(32'hbb8026ae),
	.w8(32'hbb33c2d0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e9d91),
	.w1(32'h3a81a229),
	.w2(32'hba24a087),
	.w3(32'hbb19629b),
	.w4(32'h3c2f3500),
	.w5(32'h3c956413),
	.w6(32'h3af10ace),
	.w7(32'h3c1e6c5e),
	.w8(32'h3c2cbda6),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6bbf6),
	.w1(32'h3b36c2ce),
	.w2(32'h3bade9a6),
	.w3(32'h3c3d4325),
	.w4(32'h3c2f5a07),
	.w5(32'h3c67e553),
	.w6(32'h3b1b6164),
	.w7(32'h3b3fddf1),
	.w8(32'h3c65b5e9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0fa62),
	.w1(32'h3c389f07),
	.w2(32'h3c25deb4),
	.w3(32'h3ba766cd),
	.w4(32'h3ccfa2ad),
	.w5(32'h3ce53c3d),
	.w6(32'h3b37a0c2),
	.w7(32'h3c3e0170),
	.w8(32'h3c8571d0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a831b),
	.w1(32'h3bd2db5d),
	.w2(32'hbbeeb259),
	.w3(32'h3cf1f361),
	.w4(32'hbb8fc9f4),
	.w5(32'hbc8de956),
	.w6(32'h3c84a2f9),
	.w7(32'h3aeba772),
	.w8(32'hbb1b453b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5202e8),
	.w1(32'h39f3cfe8),
	.w2(32'hbb4ff3b7),
	.w3(32'hbc19d7c0),
	.w4(32'hbb9f4be9),
	.w5(32'hbbc8b5b1),
	.w6(32'hbb3bf3d2),
	.w7(32'hbba991c1),
	.w8(32'hbb2afb41),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06333a),
	.w1(32'h3bd826c0),
	.w2(32'hba96e403),
	.w3(32'h3bf2a307),
	.w4(32'hb9bf3808),
	.w5(32'hbbae06f9),
	.w6(32'h3c1df270),
	.w7(32'h3b145c91),
	.w8(32'hbb24e2a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule