module layer_10_featuremap_15(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc747fa),
	.w1(32'h3bf0d53a),
	.w2(32'h3b622aea),
	.w3(32'hbcb44aee),
	.w4(32'hbbfc5f7c),
	.w5(32'h3a734297),
	.w6(32'hbc8e5d49),
	.w7(32'hbba084d2),
	.w8(32'hbaafc544),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb36bcf),
	.w1(32'hbc1fdb92),
	.w2(32'h3c0f54bd),
	.w3(32'hba545110),
	.w4(32'hbc2d6e37),
	.w5(32'h3bdaebdb),
	.w6(32'hbb922c73),
	.w7(32'h3ba88ec9),
	.w8(32'h3bcfa5bf),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f2a2d),
	.w1(32'h3c317b96),
	.w2(32'hbc5fea39),
	.w3(32'h3b0a0322),
	.w4(32'hbb85dc87),
	.w5(32'hbc73422e),
	.w6(32'hba641a22),
	.w7(32'hbbf2b46f),
	.w8(32'hbc2856b9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e25fc),
	.w1(32'hbc6c8939),
	.w2(32'h3b26c9e0),
	.w3(32'hbd07a3fa),
	.w4(32'hbc8948dc),
	.w5(32'hba9d7c36),
	.w6(32'hbc45423b),
	.w7(32'hbc5036d2),
	.w8(32'h39ec67fe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba28da3),
	.w1(32'hbba1fa57),
	.w2(32'h3988dfda),
	.w3(32'hbc09a9cf),
	.w4(32'hbc5df2f9),
	.w5(32'h3bb38d1a),
	.w6(32'h3c002fc3),
	.w7(32'h3b880928),
	.w8(32'h3a787d0f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169785),
	.w1(32'h3c06c0b0),
	.w2(32'h39e80788),
	.w3(32'h3c7b8ded),
	.w4(32'h3be6cad0),
	.w5(32'hbb3c5a7f),
	.w6(32'h3c1d4cdf),
	.w7(32'h3b84d94f),
	.w8(32'hbba59e67),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76247),
	.w1(32'hba207643),
	.w2(32'h3bbcf971),
	.w3(32'hbc097ccc),
	.w4(32'hbb07df08),
	.w5(32'h3b76bca0),
	.w6(32'hbc346820),
	.w7(32'hbbd37656),
	.w8(32'h3b94ba4d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c089c1d),
	.w1(32'hba83739b),
	.w2(32'h3aea3c53),
	.w3(32'h39b9b6d5),
	.w4(32'hbb539168),
	.w5(32'hbb87ae7a),
	.w6(32'h3b10d9a2),
	.w7(32'hbb9a0d0d),
	.w8(32'hbc6a7319),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71862b),
	.w1(32'h3bba4f16),
	.w2(32'h3b7ea4c3),
	.w3(32'hbc50039a),
	.w4(32'hbc0b03e3),
	.w5(32'hbaf9bfa3),
	.w6(32'hbc940519),
	.w7(32'hbc24d1e5),
	.w8(32'hbbd6c028),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea9f3a),
	.w1(32'h3c317bb7),
	.w2(32'h3bf339b8),
	.w3(32'h39f54eb6),
	.w4(32'h391b13d4),
	.w5(32'h3c2709fc),
	.w6(32'hbbd655c6),
	.w7(32'h3b7cde5b),
	.w8(32'h3c3cb6c7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebb4c4),
	.w1(32'hbba15f25),
	.w2(32'hbc14171d),
	.w3(32'hbaf3ee73),
	.w4(32'hbb8449c6),
	.w5(32'hbc7783ba),
	.w6(32'h3b77a568),
	.w7(32'hb8b5c8ec),
	.w8(32'hbbb850e9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87a886),
	.w1(32'hbc5626ba),
	.w2(32'h3b83efd7),
	.w3(32'hbcea593b),
	.w4(32'hbccaa2ad),
	.w5(32'h3bdddcd5),
	.w6(32'hbc962b6b),
	.w7(32'hbca47727),
	.w8(32'h3bbd065d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818837),
	.w1(32'h3b9a70df),
	.w2(32'h3cc82b4c),
	.w3(32'h3abc053c),
	.w4(32'h3ad94e1a),
	.w5(32'h3caf68d6),
	.w6(32'h3b1af93c),
	.w7(32'h3b85ce5e),
	.w8(32'h3c4fce9e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf89c4),
	.w1(32'h3c749211),
	.w2(32'h3c16e573),
	.w3(32'h3cffcd49),
	.w4(32'h3c70dd00),
	.w5(32'h3c02ba76),
	.w6(32'h3cd8352e),
	.w7(32'h3c69c0cb),
	.w8(32'h3c60032c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33072c),
	.w1(32'h3ba8b72e),
	.w2(32'h38845aee),
	.w3(32'h3c7ff821),
	.w4(32'h3c1b29ba),
	.w5(32'h3b8a31b4),
	.w6(32'h3c6bb176),
	.w7(32'hba08db13),
	.w8(32'h3afb29b3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b049718),
	.w1(32'h37c6003e),
	.w2(32'h3c2181ff),
	.w3(32'h3c7feaa0),
	.w4(32'h3b3e6b7c),
	.w5(32'h3c38f949),
	.w6(32'h3c465e2b),
	.w7(32'h3bd72923),
	.w8(32'h3c57f9ce),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d05711),
	.w1(32'hbb0e5b87),
	.w2(32'hb91cd97a),
	.w3(32'hbaaec408),
	.w4(32'hbb475925),
	.w5(32'hbaba7a0d),
	.w6(32'h3b3ee952),
	.w7(32'hb93a4376),
	.w8(32'hb8085e76),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b738aba),
	.w1(32'h3c49dab6),
	.w2(32'h3c56c92e),
	.w3(32'hb9d2f681),
	.w4(32'h3b98a397),
	.w5(32'h3c5ce44a),
	.w6(32'h3b5be5e1),
	.w7(32'h3bf0ba02),
	.w8(32'h3c34f9c8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cedb8),
	.w1(32'h3bf86a00),
	.w2(32'hbc117ec8),
	.w3(32'h3c621e2d),
	.w4(32'h3aa8effa),
	.w5(32'h3a40d02f),
	.w6(32'h39c7a550),
	.w7(32'hba818049),
	.w8(32'h3c1aaaf7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7f394),
	.w1(32'hbc57e299),
	.w2(32'h3a2c022a),
	.w3(32'hbcabb0c2),
	.w4(32'hbc985d7e),
	.w5(32'h39ffd916),
	.w6(32'hbbdf26f8),
	.w7(32'hbc9b7f3b),
	.w8(32'hb977dc67),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf109a7),
	.w1(32'hba61f3ef),
	.w2(32'hbb132e95),
	.w3(32'h3a969113),
	.w4(32'h3aa8c6f8),
	.w5(32'hbba6cd01),
	.w6(32'h3aac77a5),
	.w7(32'hba5470c0),
	.w8(32'hb8dcd1d8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc863061),
	.w1(32'hbc3fac59),
	.w2(32'hbc186673),
	.w3(32'hbcc7eaee),
	.w4(32'hbcaadbdb),
	.w5(32'hbbdb7fec),
	.w6(32'hbc2cfedd),
	.w7(32'hbbcfb905),
	.w8(32'h3b85a104),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2654ae),
	.w1(32'hbc53f017),
	.w2(32'h3c5115f1),
	.w3(32'hbc04cd1e),
	.w4(32'hbc718c58),
	.w5(32'h3c1da0c9),
	.w6(32'hba4788c1),
	.w7(32'hbc004f68),
	.w8(32'h3c4d2823),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad00e09),
	.w1(32'hbb625e84),
	.w2(32'h3c66239d),
	.w3(32'hbb27d408),
	.w4(32'hbb5d44ab),
	.w5(32'h3c8b5537),
	.w6(32'h3b445f9b),
	.w7(32'h3a8b18a8),
	.w8(32'h3bf1eb7e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb874bd),
	.w1(32'h392316e7),
	.w2(32'hbc4d98f0),
	.w3(32'h3cdbb03b),
	.w4(32'h3c12c264),
	.w5(32'hbb996099),
	.w6(32'h3cbeecc7),
	.w7(32'h3c2f543d),
	.w8(32'hbc10d822),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8c0c),
	.w1(32'hbc0b54e5),
	.w2(32'h3c07ba72),
	.w3(32'hbc1da5d2),
	.w4(32'hbc736a04),
	.w5(32'h3a2a78b9),
	.w6(32'hbc35e43c),
	.w7(32'hbc326025),
	.w8(32'h3ae3a246),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f87b),
	.w1(32'hbac9d188),
	.w2(32'h37079b61),
	.w3(32'hb74e554d),
	.w4(32'hbc85673a),
	.w5(32'h3a4bdb3d),
	.w6(32'h3ba4728b),
	.w7(32'h3b9b2e0e),
	.w8(32'h39c9219a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894b06a),
	.w1(32'hbbfbbf19),
	.w2(32'h3b905b37),
	.w3(32'h3c083734),
	.w4(32'hbab76347),
	.w5(32'h3b72477d),
	.w6(32'h3bf6685c),
	.w7(32'hbaf4375b),
	.w8(32'h3bbdc447),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c243193),
	.w1(32'h3b8bbb6a),
	.w2(32'hbc1842cd),
	.w3(32'h3b85fe71),
	.w4(32'h3b93efd8),
	.w5(32'h3bed63a8),
	.w6(32'hbbeb235f),
	.w7(32'h3b494ce4),
	.w8(32'h3afc14c7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec1d61),
	.w1(32'hbce18850),
	.w2(32'hbb78d6fe),
	.w3(32'hbcd14cf1),
	.w4(32'hbce4e1ec),
	.w5(32'hbb1a3b9e),
	.w6(32'hbba2a1d5),
	.w7(32'hbcd03569),
	.w8(32'hba597381),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aba612),
	.w1(32'hbb32ecb8),
	.w2(32'hbbcd4bc9),
	.w3(32'h3b4e9bfa),
	.w4(32'hba8201da),
	.w5(32'hbb41e268),
	.w6(32'h3af0041c),
	.w7(32'hba89f6aa),
	.w8(32'h3b1a70ed),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558c24),
	.w1(32'h3baf0f37),
	.w2(32'h3aeaf46e),
	.w3(32'h3bdde82b),
	.w4(32'h39d6c953),
	.w5(32'h3c8c95b7),
	.w6(32'h3ab1b07c),
	.w7(32'h3b03bf4c),
	.w8(32'h3c2f1a55),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2efbc9),
	.w1(32'h3ba2b166),
	.w2(32'hbac55424),
	.w3(32'h3c011736),
	.w4(32'hbc0b252b),
	.w5(32'hba4c6337),
	.w6(32'hbb40522c),
	.w7(32'hbc836b3c),
	.w8(32'hbb6306fa),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0d18),
	.w1(32'hbaf32d08),
	.w2(32'h3be07f30),
	.w3(32'hba9b6a3d),
	.w4(32'h3a6acf6e),
	.w5(32'hbc4a41ff),
	.w6(32'h3b1b6fe1),
	.w7(32'h3b1b0748),
	.w8(32'hbc6c3ef1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a76c9),
	.w1(32'hbc9af48c),
	.w2(32'hba6f1c13),
	.w3(32'hbd2fff4c),
	.w4(32'hbcf7a9f8),
	.w5(32'hbaf9d37d),
	.w6(32'hbca76846),
	.w7(32'hbc7d9eb8),
	.w8(32'hbbd220e4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a4fdc),
	.w1(32'h3b7f98dd),
	.w2(32'hbbb05055),
	.w3(32'hbbdb4386),
	.w4(32'hbbe26555),
	.w5(32'hbcbd5bb7),
	.w6(32'hbc1abf28),
	.w7(32'hbbee4d3e),
	.w8(32'hbca79205),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd5ae7),
	.w1(32'hbd1f183a),
	.w2(32'hbb366401),
	.w3(32'hbd203342),
	.w4(32'hbce5da6e),
	.w5(32'h3b6a58dd),
	.w6(32'hbccc8c1c),
	.w7(32'hbcab43a6),
	.w8(32'hb8e8d5ef),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfcd42),
	.w1(32'hbb08dd73),
	.w2(32'hbbbd742e),
	.w3(32'h3c0160d3),
	.w4(32'hb8c8ab78),
	.w5(32'hbb9d0622),
	.w6(32'h3c525a28),
	.w7(32'h3b255808),
	.w8(32'h3b68fea4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81fb046),
	.w1(32'hbc4a9d80),
	.w2(32'hbbbd21df),
	.w3(32'hbc1cebec),
	.w4(32'hbc5dda49),
	.w5(32'hbb16252d),
	.w6(32'h3c2028b3),
	.w7(32'h3c056701),
	.w8(32'hbc473202),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01943e),
	.w1(32'h3bdf96a7),
	.w2(32'hbc016e42),
	.w3(32'h3b9b8379),
	.w4(32'h3b8494db),
	.w5(32'hbc463eee),
	.w6(32'hbc915fa7),
	.w7(32'hbae9f9b0),
	.w8(32'hbbf7f043),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03e5af),
	.w1(32'hba6392b4),
	.w2(32'hb973e527),
	.w3(32'hbc15bb05),
	.w4(32'hbba10923),
	.w5(32'h3b881f41),
	.w6(32'hbbd5dd9d),
	.w7(32'hbb19355b),
	.w8(32'h3c303643),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480421),
	.w1(32'h3bff2ce1),
	.w2(32'h3bd5602a),
	.w3(32'h3b9f93c5),
	.w4(32'h3bbef607),
	.w5(32'h3cbe7fa7),
	.w6(32'h3a780f52),
	.w7(32'h3bc384f3),
	.w8(32'h3c16d21d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a970),
	.w1(32'hbbbebd87),
	.w2(32'h3a85e8d3),
	.w3(32'h3ca391ba),
	.w4(32'hbbcfbea0),
	.w5(32'hb94e6f20),
	.w6(32'h3ba09686),
	.w7(32'hbac110e5),
	.w8(32'hbb988e7f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ad40),
	.w1(32'h3b7cc158),
	.w2(32'h38c2cd62),
	.w3(32'h3a3ac405),
	.w4(32'hbb40f611),
	.w5(32'h3bed0118),
	.w6(32'hbbdb5778),
	.w7(32'hbc10503d),
	.w8(32'h3b807d30),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb169590),
	.w1(32'h3bafd2b8),
	.w2(32'hbb65a007),
	.w3(32'h3c29d946),
	.w4(32'h3c3dfd17),
	.w5(32'h3cd79e5b),
	.w6(32'h3c0e4559),
	.w7(32'h3bc5e4a2),
	.w8(32'h3cd45d69),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c05a8),
	.w1(32'h3c883508),
	.w2(32'h3c881be1),
	.w3(32'h3cc9b6f7),
	.w4(32'h3c22f9af),
	.w5(32'h3c458533),
	.w6(32'h3cb7f5a7),
	.w7(32'hbbce5e9f),
	.w8(32'h3bffc339),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d24760e),
	.w1(32'h3c9148f2),
	.w2(32'h3cc23dbe),
	.w3(32'h3cd9552b),
	.w4(32'hb93a3dbc),
	.w5(32'h3cc87c31),
	.w6(32'hbc0c0e4f),
	.w7(32'hbcc12d58),
	.w8(32'h3c1d3d17),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99d30f),
	.w1(32'h3bac6c09),
	.w2(32'h3c47e53d),
	.w3(32'hbb9600b5),
	.w4(32'hbc3ffe83),
	.w5(32'h3c1bf211),
	.w6(32'hbc007294),
	.w7(32'hbc976216),
	.w8(32'h3bd6ed34),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9b925),
	.w1(32'h3b45067a),
	.w2(32'hbaf771ce),
	.w3(32'hba6a9723),
	.w4(32'hbb66f862),
	.w5(32'hbbe027bd),
	.w6(32'hbb50ac30),
	.w7(32'hbaf5f907),
	.w8(32'hbc27209e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9066f),
	.w1(32'h3c0083ee),
	.w2(32'hbaa3279f),
	.w3(32'h3bb26057),
	.w4(32'h3c25233b),
	.w5(32'hbb7cf3f6),
	.w6(32'h3aac3d51),
	.w7(32'hbadf059e),
	.w8(32'hba7f8e8b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1acf8e),
	.w1(32'hbbcb5bda),
	.w2(32'hbd07b865),
	.w3(32'hbb74f93a),
	.w4(32'h3b9c29e6),
	.w5(32'hbcbb5821),
	.w6(32'h3c808160),
	.w7(32'h3c499df9),
	.w8(32'hbb9117ea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cfe7b),
	.w1(32'h3c2511e9),
	.w2(32'h3c4c4f28),
	.w3(32'hbad939ae),
	.w4(32'h3c53f04d),
	.w5(32'h3b4d8e4a),
	.w6(32'h3a5500a8),
	.w7(32'h3ba9c1ec),
	.w8(32'h3c89659c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72656c),
	.w1(32'hbb6e850d),
	.w2(32'h3aeff5c2),
	.w3(32'h3bdecc32),
	.w4(32'h3c0468df),
	.w5(32'h3ba03428),
	.w6(32'h3cb96cbb),
	.w7(32'h3c91a893),
	.w8(32'h3952676c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40bfb8),
	.w1(32'h3a6af0c9),
	.w2(32'h3a0c9cd1),
	.w3(32'hba3819f1),
	.w4(32'h3a59e3eb),
	.w5(32'h3c85e165),
	.w6(32'hbbd7dee0),
	.w7(32'hbac6e2e8),
	.w8(32'hba56ab57),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec3772),
	.w1(32'hbc13e84d),
	.w2(32'hbb58f17d),
	.w3(32'hbcdfa396),
	.w4(32'hbc515248),
	.w5(32'hbbe3b56a),
	.w6(32'h3bb5127e),
	.w7(32'hb95660b4),
	.w8(32'hbaa7b461),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca6782),
	.w1(32'hbb223f65),
	.w2(32'h3c276b0c),
	.w3(32'hbc77c674),
	.w4(32'hbc3521d7),
	.w5(32'h3c6d6ad1),
	.w6(32'hbc4100c2),
	.w7(32'hbbf244c5),
	.w8(32'hbbb30ecd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb32e75),
	.w1(32'h3a33b2e9),
	.w2(32'hbbcc9e35),
	.w3(32'hbb6bf9bd),
	.w4(32'hbc3892b6),
	.w5(32'hbb92c161),
	.w6(32'hbc895ba9),
	.w7(32'hbc496c3a),
	.w8(32'hba0fbf68),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7f755),
	.w1(32'hba7f7d0f),
	.w2(32'hbafd34ff),
	.w3(32'h3b9fab56),
	.w4(32'h3b5fd327),
	.w5(32'hba478c86),
	.w6(32'h3b9d896a),
	.w7(32'h3b720523),
	.w8(32'h3bf23180),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031377),
	.w1(32'h3c16bfba),
	.w2(32'hbb8b1455),
	.w3(32'hba5e0cf7),
	.w4(32'h3c26c984),
	.w5(32'hba4c2553),
	.w6(32'h3c12f6f8),
	.w7(32'h3ca788cd),
	.w8(32'hbbc54f34),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a0c1),
	.w1(32'hbb2c2cb0),
	.w2(32'hbc12758b),
	.w3(32'h3aea86ea),
	.w4(32'hbb635c86),
	.w5(32'hbbb9e30c),
	.w6(32'hbb7676e4),
	.w7(32'hbb8cdb94),
	.w8(32'h3bf38548),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06fd0a),
	.w1(32'h3aedb4ab),
	.w2(32'h3ce51b3c),
	.w3(32'h3ba857f5),
	.w4(32'h3c3f523d),
	.w5(32'h3d184ef4),
	.w6(32'h3c4a7a79),
	.w7(32'h3c2a42c4),
	.w8(32'h3bfc4001),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00a057),
	.w1(32'h39e11ec7),
	.w2(32'h3ce65586),
	.w3(32'h3cc9c8dc),
	.w4(32'hbc85780d),
	.w5(32'h3c7526c0),
	.w6(32'hbc86374f),
	.w7(32'hbcec8562),
	.w8(32'hb9f34d8d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f3c69),
	.w1(32'hbb3419ba),
	.w2(32'hbc923d2e),
	.w3(32'h3a876500),
	.w4(32'hbcb61f2f),
	.w5(32'hbc5c2bc0),
	.w6(32'hbcc1b56a),
	.w7(32'hbd006b86),
	.w8(32'hbc2902af),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d7a91),
	.w1(32'hbc0caf6b),
	.w2(32'h3bc87fe3),
	.w3(32'hbc464862),
	.w4(32'hbb92a94b),
	.w5(32'hbb53b7c2),
	.w6(32'hbbf12313),
	.w7(32'hbb72dec4),
	.w8(32'h3bf360fc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc029cd),
	.w1(32'h3c4e8875),
	.w2(32'hbb905b0b),
	.w3(32'hbbd54059),
	.w4(32'h3c10f2c4),
	.w5(32'h3a92b6fe),
	.w6(32'hbb069ce2),
	.w7(32'h3bb6cf24),
	.w8(32'h3bd187ca),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85435a),
	.w1(32'h3b5f6feb),
	.w2(32'h3b9350be),
	.w3(32'h3bc4d4b4),
	.w4(32'h3bfd5904),
	.w5(32'h3b694ee9),
	.w6(32'h3c2ab0a1),
	.w7(32'h3c20f0be),
	.w8(32'hbb1ea768),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028ca0),
	.w1(32'h39366c11),
	.w2(32'h3a710fff),
	.w3(32'h3c15cdd9),
	.w4(32'h3bbb086f),
	.w5(32'hbb86cc6e),
	.w6(32'hbb651233),
	.w7(32'hbbc75da5),
	.w8(32'hbb2578ce),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca58ff),
	.w1(32'h3ca588ff),
	.w2(32'h3c1eefdb),
	.w3(32'hbbca64bd),
	.w4(32'h3c0cb1fe),
	.w5(32'h3c7a259d),
	.w6(32'hbaa392fc),
	.w7(32'h3c69396b),
	.w8(32'h3cb6570e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c453),
	.w1(32'h3ba413ac),
	.w2(32'hba87fc74),
	.w3(32'h3c9ec020),
	.w4(32'h3cc33531),
	.w5(32'h3aade53b),
	.w6(32'h3d01bc07),
	.w7(32'h3cdf6fb8),
	.w8(32'h3a9d6382),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8572cd),
	.w1(32'hbc431926),
	.w2(32'h3be3342f),
	.w3(32'h3a96121b),
	.w4(32'hbc0ac43c),
	.w5(32'hbb9219d5),
	.w6(32'h3b9ea91f),
	.w7(32'hbb3aa88d),
	.w8(32'hbbfd9a83),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52ea54),
	.w1(32'h3b2ec304),
	.w2(32'hbbc95287),
	.w3(32'hbbe8d95a),
	.w4(32'hbc0ccb89),
	.w5(32'hbb7c9894),
	.w6(32'hbc6b50da),
	.w7(32'hbbb58a09),
	.w8(32'hbba14251),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38c4bd),
	.w1(32'hbaf9bc8a),
	.w2(32'h3c9c2bd0),
	.w3(32'hbabae6cd),
	.w4(32'hbbe0ab8d),
	.w5(32'h3be7ace6),
	.w6(32'hbc0812c9),
	.w7(32'hbaced4a3),
	.w8(32'hbb0517a1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3b50c),
	.w1(32'h3cef0808),
	.w2(32'hbb9a7979),
	.w3(32'h3c8d0423),
	.w4(32'h3c104dfb),
	.w5(32'h3c752586),
	.w6(32'hbca3e031),
	.w7(32'hbc79a502),
	.w8(32'h3cbfd39b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40c0e7),
	.w1(32'hbd13937e),
	.w2(32'hb637063e),
	.w3(32'h3be61b84),
	.w4(32'hbca12fa2),
	.w5(32'h3b8a0742),
	.w6(32'h3cd253cb),
	.w7(32'h3bdd5c9a),
	.w8(32'h3b943785),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3f21),
	.w1(32'h3ac87e4f),
	.w2(32'hbc007ea7),
	.w3(32'h3ba74b6f),
	.w4(32'hbb699a1f),
	.w5(32'hbc00560f),
	.w6(32'h3b8b01ae),
	.w7(32'h3b109ab1),
	.w8(32'hba131c7c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d77b8),
	.w1(32'hbb9f62a9),
	.w2(32'h3c9f1eae),
	.w3(32'hbbb60e92),
	.w4(32'hbbf17d55),
	.w5(32'h3c94e68f),
	.w6(32'hbb30c846),
	.w7(32'hbbf5bd34),
	.w8(32'h3c837ee2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c858344),
	.w1(32'h3c53ca43),
	.w2(32'h3bd11ff8),
	.w3(32'h3c8461b3),
	.w4(32'h3c8b60ca),
	.w5(32'h3bd56c1a),
	.w6(32'h3c4aae5e),
	.w7(32'h3c2aab68),
	.w8(32'h3b4929d0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf982ff),
	.w1(32'hbaa12d4a),
	.w2(32'h3c6626bd),
	.w3(32'h3b8e5db4),
	.w4(32'h3ab276da),
	.w5(32'h3c941339),
	.w6(32'h3b7398ea),
	.w7(32'hbb664d8a),
	.w8(32'h3b46e787),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc4351),
	.w1(32'h3bec53a6),
	.w2(32'h3b86c61f),
	.w3(32'h3c972cc7),
	.w4(32'hbbe3eeed),
	.w5(32'h3b357010),
	.w6(32'hbbb6f40d),
	.w7(32'hbc592a1f),
	.w8(32'h3b07da5c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f271fc),
	.w1(32'hba304d23),
	.w2(32'h3c10eb81),
	.w3(32'h3b0c9005),
	.w4(32'h3bb9cefe),
	.w5(32'h37ba95b5),
	.w6(32'h3ab369b0),
	.w7(32'hba799d3f),
	.w8(32'h3c28d3b1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a848609),
	.w1(32'h3bb4ccf5),
	.w2(32'hba426323),
	.w3(32'hbb9b2abf),
	.w4(32'hbb2a9546),
	.w5(32'h3b22a8e7),
	.w6(32'h3c044297),
	.w7(32'h3bd757db),
	.w8(32'hba0ccfc1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac367),
	.w1(32'hbaa14c29),
	.w2(32'h3b9be755),
	.w3(32'h3c1e0c9b),
	.w4(32'h3b5b532a),
	.w5(32'hbc77249f),
	.w6(32'h3b3fea86),
	.w7(32'hbaf31acd),
	.w8(32'hbb17f53e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f233c),
	.w1(32'h3bfa4a1e),
	.w2(32'h3cc40a2a),
	.w3(32'hbcdc8ae0),
	.w4(32'hb957e685),
	.w5(32'h3c78f254),
	.w6(32'hbc925b30),
	.w7(32'h3bc13855),
	.w8(32'hbb68eaab),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda37ca),
	.w1(32'h3c4367d3),
	.w2(32'h3cc55a2a),
	.w3(32'h3cb8c905),
	.w4(32'hbb9221d3),
	.w5(32'h3c869399),
	.w6(32'hbc11f97c),
	.w7(32'hbcf5e0ee),
	.w8(32'h3ab3af0d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce31536),
	.w1(32'h3c20a1cd),
	.w2(32'hbbaa72b3),
	.w3(32'h3cbcf82c),
	.w4(32'h3b78f804),
	.w5(32'hbd058a1d),
	.w6(32'hbc922933),
	.w7(32'hbcc8b433),
	.w8(32'hbc285908),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb831da8),
	.w1(32'h3b476b03),
	.w2(32'hba9a20df),
	.w3(32'hbc84b030),
	.w4(32'h3c0cf607),
	.w5(32'h3b0b5bd6),
	.w6(32'h3b7ffe93),
	.w7(32'h3c6f792e),
	.w8(32'h3b7fd974),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278886),
	.w1(32'h3b5f6639),
	.w2(32'hbb8ceccd),
	.w3(32'h3a3bcdf0),
	.w4(32'h3a286279),
	.w5(32'hb9cc6e9e),
	.w6(32'h3ac9ea76),
	.w7(32'h3aefbef2),
	.w8(32'h3ba201d5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81b7a6),
	.w1(32'hba542b55),
	.w2(32'hbaf70701),
	.w3(32'h3b35ff0a),
	.w4(32'hb9f2f253),
	.w5(32'hbc4ff24a),
	.w6(32'h3b8c4483),
	.w7(32'hba6556b8),
	.w8(32'hba61855e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fd96),
	.w1(32'hbbca7279),
	.w2(32'h3b3c6eec),
	.w3(32'hbbcef0e1),
	.w4(32'h3b474d4c),
	.w5(32'hbb91cc1a),
	.w6(32'h3c8a3543),
	.w7(32'h3c15520e),
	.w8(32'hbb274514),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a0058),
	.w1(32'h3b0ab589),
	.w2(32'hb90838cf),
	.w3(32'hbc837e90),
	.w4(32'hbc431977),
	.w5(32'h3ad4a3f2),
	.w6(32'hbc2131cf),
	.w7(32'hbc826cfa),
	.w8(32'h3b05de76),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b423106),
	.w1(32'h3c2cb472),
	.w2(32'hbb5cf06c),
	.w3(32'h3b73e2ee),
	.w4(32'h3a6eb67f),
	.w5(32'hb9da038d),
	.w6(32'h3bb97894),
	.w7(32'hbb93bf5d),
	.w8(32'h3ace0b11),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74996b),
	.w1(32'h3941bc6a),
	.w2(32'hb9c23b4b),
	.w3(32'h3ba59e6e),
	.w4(32'h3bfb4c0b),
	.w5(32'h3be812e5),
	.w6(32'h3b437729),
	.w7(32'h3c3a96a7),
	.w8(32'h3c023435),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae186e9),
	.w1(32'hbbc0b367),
	.w2(32'hbbe460ab),
	.w3(32'h3b24ba22),
	.w4(32'hb80a7514),
	.w5(32'hbb76ebe3),
	.w6(32'h3c01dfbd),
	.w7(32'h3b3a0bfb),
	.w8(32'hba8c96ec),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9beec1),
	.w1(32'h3ba146fd),
	.w2(32'h3c7a8252),
	.w3(32'h3ae5e0f2),
	.w4(32'h3a99b37f),
	.w5(32'h3c9b1d28),
	.w6(32'hb9ed2e4f),
	.w7(32'h3ad140af),
	.w8(32'h3ce93b6a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fabb),
	.w1(32'h3c1f36c2),
	.w2(32'hbc46e19d),
	.w3(32'h3caf43bd),
	.w4(32'h3cacbe4d),
	.w5(32'hbca77fab),
	.w6(32'h3cf534c5),
	.w7(32'h3cd97424),
	.w8(32'hbc16c529),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5dd23c),
	.w1(32'hbb2a6231),
	.w2(32'hbcdc4332),
	.w3(32'hbbb680aa),
	.w4(32'h3c19920f),
	.w5(32'hbd0c47e0),
	.w6(32'h3bb4d085),
	.w7(32'h3c54f369),
	.w8(32'hbc6ea624),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbecb7e),
	.w1(32'hbc31d6b8),
	.w2(32'h3d0354ee),
	.w3(32'hbcde5ff5),
	.w4(32'hbc5b2f69),
	.w5(32'h3cb378e9),
	.w6(32'hbc862861),
	.w7(32'hbbb92ff3),
	.w8(32'hbb6a526c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfdcbae),
	.w1(32'hbb65af9c),
	.w2(32'h3b7897ac),
	.w3(32'h3c85930a),
	.w4(32'hbc93f155),
	.w5(32'hbc55c454),
	.w6(32'hbc435e80),
	.w7(32'hbd0bab15),
	.w8(32'hbbaae61a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89c9f7),
	.w1(32'hbc9235a2),
	.w2(32'h3afbfb02),
	.w3(32'hbce3e616),
	.w4(32'hbb8ec650),
	.w5(32'h3be8d398),
	.w6(32'hbccc7b83),
	.w7(32'hbc8679a8),
	.w8(32'h3c59bf37),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085658),
	.w1(32'hbb930b02),
	.w2(32'hbbe2bef8),
	.w3(32'hbbae0bcd),
	.w4(32'hb943a960),
	.w5(32'hba5dd88d),
	.w6(32'h3bbe3dce),
	.w7(32'h3bafc66b),
	.w8(32'h3bb4c44b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0c82f),
	.w1(32'h3bc74f63),
	.w2(32'hbbf37686),
	.w3(32'h3b3e3f75),
	.w4(32'hbc38addc),
	.w5(32'hbc172d56),
	.w6(32'h3bbdcc4d),
	.w7(32'hba964ec8),
	.w8(32'hbbfd7641),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51dcde),
	.w1(32'h3c7c9ce3),
	.w2(32'h3c157db0),
	.w3(32'h3b31d677),
	.w4(32'h3c1388d7),
	.w5(32'h3c23e778),
	.w6(32'h3a88642d),
	.w7(32'h3c25aaa3),
	.w8(32'h3bb3ccea),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dd9e8),
	.w1(32'hbadedb5c),
	.w2(32'h3b22d44a),
	.w3(32'hbaa874b5),
	.w4(32'hbb8d99d1),
	.w5(32'h3b95c5db),
	.w6(32'hbc63523f),
	.w7(32'hbc01c235),
	.w8(32'h3a0e7fa7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cdfd6),
	.w1(32'h3bbd04ad),
	.w2(32'h3bf0fdca),
	.w3(32'hbafce25f),
	.w4(32'h3b3c7b0a),
	.w5(32'hbc2efdff),
	.w6(32'hbbbb4162),
	.w7(32'hbb2eec19),
	.w8(32'hbbacd22a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82810e),
	.w1(32'h3c477534),
	.w2(32'hbc3fb227),
	.w3(32'h3b8740db),
	.w4(32'h3c2819c5),
	.w5(32'hbc2ec90a),
	.w6(32'hbac4a59c),
	.w7(32'h3a595e47),
	.w8(32'hbaec03b6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2a7a),
	.w1(32'hbb9dc038),
	.w2(32'h3b80d795),
	.w3(32'hbbf7e0ff),
	.w4(32'h3b17acdf),
	.w5(32'hbb14235f),
	.w6(32'hbc15313a),
	.w7(32'h3b81d835),
	.w8(32'hbb8efa8e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29f2e5),
	.w1(32'h3c0880c9),
	.w2(32'h3bf598eb),
	.w3(32'hba7dd4b4),
	.w4(32'h3b1aee21),
	.w5(32'h3c3498cc),
	.w6(32'hbbb1ca8c),
	.w7(32'h3b389bc5),
	.w8(32'h3a843b5c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc3089),
	.w1(32'hbaa29b68),
	.w2(32'h3ce15c80),
	.w3(32'h3c499673),
	.w4(32'hbb613d89),
	.w5(32'h3c9168bb),
	.w6(32'hba574423),
	.w7(32'hbb37ea63),
	.w8(32'hbbc7af9c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce58367),
	.w1(32'hbb1e0206),
	.w2(32'h3b9a8331),
	.w3(32'h3c2aa842),
	.w4(32'hbc3aeb40),
	.w5(32'h3c7e2a2c),
	.w6(32'hbcd051d8),
	.w7(32'hbcc8af0e),
	.w8(32'h3b21e771),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b894d25),
	.w1(32'hbc046290),
	.w2(32'h3caea163),
	.w3(32'h3c1cce24),
	.w4(32'hbbf76d2b),
	.w5(32'h3ce6e536),
	.w6(32'hbb8d516e),
	.w7(32'hbbf532c2),
	.w8(32'h3bec8c30),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabc8aa),
	.w1(32'h3b253f50),
	.w2(32'hbbac8ccf),
	.w3(32'h3cb78550),
	.w4(32'hbbc310f0),
	.w5(32'hbc643c92),
	.w6(32'h3b52f902),
	.w7(32'hbbb8c50c),
	.w8(32'hbaf1264f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c646dd2),
	.w1(32'h3c837173),
	.w2(32'h3bc8f957),
	.w3(32'hbbf89f01),
	.w4(32'hba00ee8a),
	.w5(32'hbbfc1598),
	.w6(32'hba1f9db4),
	.w7(32'hba9d0ba3),
	.w8(32'hbbaed8cf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc325f2),
	.w1(32'h3a44167a),
	.w2(32'h3bbf657d),
	.w3(32'hbccc6bbb),
	.w4(32'hbc3cc4ac),
	.w5(32'h3d102995),
	.w6(32'hbaba0704),
	.w7(32'hba40d2ae),
	.w8(32'h3c444964),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b9d82),
	.w1(32'hbc43a084),
	.w2(32'hbb831b77),
	.w3(32'h3ce72226),
	.w4(32'hbcb08a28),
	.w5(32'hbc0174b4),
	.w6(32'h3bdd90ee),
	.w7(32'hbc88193d),
	.w8(32'hbbc208f7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab51e4),
	.w1(32'hbb6a123a),
	.w2(32'h3a5afccc),
	.w3(32'hbc1248b1),
	.w4(32'hbbf99dc8),
	.w5(32'hbb64ff97),
	.w6(32'hbc4c382b),
	.w7(32'hbbeeec72),
	.w8(32'hbb38f5e4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a636641),
	.w1(32'h3b5b161c),
	.w2(32'h3ac387bc),
	.w3(32'h3b2a2262),
	.w4(32'h3b990cf2),
	.w5(32'h39ef749e),
	.w6(32'h3b2ef81b),
	.w7(32'h3c231323),
	.w8(32'hba825537),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed5a0f),
	.w1(32'hbafc3f51),
	.w2(32'hba06e344),
	.w3(32'hbba3a2f7),
	.w4(32'hbc192659),
	.w5(32'h3baca5ef),
	.w6(32'hbb1d13f0),
	.w7(32'hbbb18daa),
	.w8(32'h3b9536ed),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14b7ae),
	.w1(32'hbb049cb5),
	.w2(32'hbc9f3eef),
	.w3(32'h3aaf6190),
	.w4(32'hbacc3e34),
	.w5(32'hbca266f4),
	.w6(32'hba2d60fa),
	.w7(32'h3b6d1b84),
	.w8(32'hbac29215),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88a2c5),
	.w1(32'hbbac59d4),
	.w2(32'h3b9b8d55),
	.w3(32'hbcaeec56),
	.w4(32'hbc277f2c),
	.w5(32'h3bf640a0),
	.w6(32'hbc230dc0),
	.w7(32'hbbd81674),
	.w8(32'h3bdd61c3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1216d6),
	.w1(32'h3c3caed8),
	.w2(32'h3bc5d9ba),
	.w3(32'hba51be7a),
	.w4(32'h3bf22569),
	.w5(32'h3c27ad32),
	.w6(32'hba83e76a),
	.w7(32'h3bc12400),
	.w8(32'hba9c38c4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c411d46),
	.w1(32'hbb04248b),
	.w2(32'hbade4d2b),
	.w3(32'h3b823e48),
	.w4(32'hbc640a19),
	.w5(32'hbb014c61),
	.w6(32'hbbb8612c),
	.w7(32'hbcb3ec20),
	.w8(32'hbacc697e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6660ad),
	.w1(32'hbb5c5775),
	.w2(32'h3a80098c),
	.w3(32'hb8e65a9e),
	.w4(32'hbb656964),
	.w5(32'hba29dada),
	.w6(32'hbb396f46),
	.w7(32'hbb9112cd),
	.w8(32'h39dd85c5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab24998),
	.w1(32'h3aa35f93),
	.w2(32'h3b175a58),
	.w3(32'h3ae13eb6),
	.w4(32'hbb0c85a5),
	.w5(32'h3ad3e35b),
	.w6(32'h3bdd30e0),
	.w7(32'hba154a26),
	.w8(32'h3b736aa8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6909ea),
	.w1(32'h3c06a7ba),
	.w2(32'h3c1ac4e7),
	.w3(32'hbabdeadc),
	.w4(32'h38bc7d5e),
	.w5(32'h3b575666),
	.w6(32'h3af03cf0),
	.w7(32'hbc2a8113),
	.w8(32'hb9ab817f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd71e8e),
	.w1(32'hbb71c7ef),
	.w2(32'hbba04376),
	.w3(32'hbad6cc7c),
	.w4(32'hbc260265),
	.w5(32'hbcda06a8),
	.w6(32'hbbafe4ce),
	.w7(32'hbbd7e8c5),
	.w8(32'hbc28effd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c5617),
	.w1(32'h3afb09be),
	.w2(32'hbc562aea),
	.w3(32'hbc9e4b77),
	.w4(32'h3ba812ae),
	.w5(32'hbc3b90cd),
	.w6(32'hbc3d812b),
	.w7(32'hbb0c6c66),
	.w8(32'hbbf2b011),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010ece),
	.w1(32'h3c8ae827),
	.w2(32'hba28fcce),
	.w3(32'hbc07c2d5),
	.w4(32'h3c31aa75),
	.w5(32'hbc3b3f99),
	.w6(32'hba7e6859),
	.w7(32'h3c4a754a),
	.w8(32'hbbcd7ef2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cbe1a),
	.w1(32'h3cf2c77f),
	.w2(32'h3cc8a887),
	.w3(32'h3be920f6),
	.w4(32'h3c88d04f),
	.w5(32'h3cb89f04),
	.w6(32'hb8f1fb8e),
	.w7(32'h3c518116),
	.w8(32'h3b39b93c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c209066),
	.w1(32'h3c5890cb),
	.w2(32'h3c8e3f1b),
	.w3(32'h3ba8441d),
	.w4(32'hba9e1ddb),
	.w5(32'h3b15df82),
	.w6(32'hbc5d765a),
	.w7(32'hbc47af02),
	.w8(32'hbc03520d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb19f30),
	.w1(32'h3aa76404),
	.w2(32'h3c1b151c),
	.w3(32'h3a9a9ee7),
	.w4(32'hbb91612f),
	.w5(32'h3c49b8f6),
	.w6(32'hbbd2acf1),
	.w7(32'hbc2259b5),
	.w8(32'hba0284b1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd77b18),
	.w1(32'hbbbccd8e),
	.w2(32'h3c478bf4),
	.w3(32'h3b01b0c4),
	.w4(32'hbca13219),
	.w5(32'h3cc206de),
	.w6(32'hbc5b2485),
	.w7(32'hbc79d8c2),
	.w8(32'h3bc385b0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27419a),
	.w1(32'hba278789),
	.w2(32'hbc35193c),
	.w3(32'h3ca51432),
	.w4(32'hbbf38869),
	.w5(32'hbbc2e5cf),
	.w6(32'h3bbc6fc7),
	.w7(32'hbbb38d60),
	.w8(32'h3b81c790),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37d91a),
	.w1(32'hba9350ec),
	.w2(32'h3a56312b),
	.w3(32'h3b19d4ba),
	.w4(32'h3caacf2c),
	.w5(32'hbae2af84),
	.w6(32'h3c4e1e3b),
	.w7(32'h3c67703f),
	.w8(32'hbc41378c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c255198),
	.w1(32'h3c3cd003),
	.w2(32'h3aa53204),
	.w3(32'h3b95e190),
	.w4(32'h3bfbdf79),
	.w5(32'h39c0e6b0),
	.w6(32'h3bd75cfc),
	.w7(32'h3c1e0e35),
	.w8(32'h3a0e3276),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09c7f7),
	.w1(32'h3badb67f),
	.w2(32'h3ad15d7d),
	.w3(32'h3bf555e2),
	.w4(32'h3b832401),
	.w5(32'h3b71d830),
	.w6(32'hbb9deb2b),
	.w7(32'hbbe3cace),
	.w8(32'h3bde8ee1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ea835),
	.w1(32'hbc1984df),
	.w2(32'h3b20ebc6),
	.w3(32'hbb99c392),
	.w4(32'hb9c88cf7),
	.w5(32'h3b10763c),
	.w6(32'h3b669a42),
	.w7(32'h3c06041b),
	.w8(32'h38bcd84e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0c07e),
	.w1(32'h3b234001),
	.w2(32'hbc20505c),
	.w3(32'h3be7ae27),
	.w4(32'hbb855542),
	.w5(32'hbc2756ba),
	.w6(32'hbbda7a9f),
	.w7(32'hbc4bb980),
	.w8(32'hbb6a15f7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc278ec),
	.w1(32'hbbdfd7c9),
	.w2(32'h3bfe9fbc),
	.w3(32'hbc83d2f4),
	.w4(32'h3b33b0f2),
	.w5(32'h3be94a4a),
	.w6(32'hbc02e1a6),
	.w7(32'h3b94b773),
	.w8(32'h3be4c7ff),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49681c),
	.w1(32'h3b20164c),
	.w2(32'h3b16be8c),
	.w3(32'h3b9da763),
	.w4(32'h3b959f9f),
	.w5(32'h3c5c3c83),
	.w6(32'h3bc480aa),
	.w7(32'h3bccdd2e),
	.w8(32'h3bea6fca),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badf1ec),
	.w1(32'h3bd63122),
	.w2(32'h3b438627),
	.w3(32'h3c90086b),
	.w4(32'hbbc99a26),
	.w5(32'h3b04efad),
	.w6(32'h3c0b5d2f),
	.w7(32'hbb7f46a4),
	.w8(32'h3b82533f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01e349),
	.w1(32'h3b86891e),
	.w2(32'h3ba828f0),
	.w3(32'hba957323),
	.w4(32'hba91b251),
	.w5(32'h3be5282d),
	.w6(32'h3b366135),
	.w7(32'hb8cbabc9),
	.w8(32'h3c170d4f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cecd6),
	.w1(32'h3a4dba8c),
	.w2(32'hbc1d09a4),
	.w3(32'h3caa10aa),
	.w4(32'hbb1906e9),
	.w5(32'hbbad4ae1),
	.w6(32'h3c9cef66),
	.w7(32'h3bc2bc6b),
	.w8(32'h3b13b6d1),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02aa43),
	.w1(32'h3a8c4a6a),
	.w2(32'hbb1c5b26),
	.w3(32'hbb8e94f2),
	.w4(32'h3c014953),
	.w5(32'h3b92e302),
	.w6(32'h3c4cd909),
	.w7(32'h3b784101),
	.w8(32'h3aa02e25),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8260ae8),
	.w1(32'h3b2e7eec),
	.w2(32'h3acd46e4),
	.w3(32'h3c039f5f),
	.w4(32'h3b2b19a6),
	.w5(32'h3b3ea4d8),
	.w6(32'h3b92dfcd),
	.w7(32'h3b21ba94),
	.w8(32'h3b36c03a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51d721),
	.w1(32'h3b12f013),
	.w2(32'hbbeb9dce),
	.w3(32'h3b9bdbb7),
	.w4(32'h3b9165fe),
	.w5(32'hbc16c310),
	.w6(32'h3b5f17e3),
	.w7(32'h3b870e77),
	.w8(32'hbbadeb47),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07e98a),
	.w1(32'hbbac49ca),
	.w2(32'h3af13863),
	.w3(32'hbc49067c),
	.w4(32'hbc235db0),
	.w5(32'h3b8faf9a),
	.w6(32'hbbaf7d79),
	.w7(32'hbb2d1191),
	.w8(32'hbb2a4a5e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd72aa8),
	.w1(32'hbba044fd),
	.w2(32'h3c81819c),
	.w3(32'h3b89de47),
	.w4(32'hbc14beb5),
	.w5(32'h3c37fb5d),
	.w6(32'hbbfe39dc),
	.w7(32'hbc18c809),
	.w8(32'h39af7caf),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c671410),
	.w1(32'hbc031b3a),
	.w2(32'h39f6cd49),
	.w3(32'h3b4e62c9),
	.w4(32'hbcac1159),
	.w5(32'h3a233a00),
	.w6(32'hbc0904a3),
	.w7(32'hbcbeb01d),
	.w8(32'h3baa58d4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba806883),
	.w1(32'h3b8811f3),
	.w2(32'h3cecbecd),
	.w3(32'hbb2d3bef),
	.w4(32'h3bc479de),
	.w5(32'h3d0fb1bf),
	.w6(32'h3bd7e052),
	.w7(32'h39da45d6),
	.w8(32'h3a5db675),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d029e99),
	.w1(32'h3ba476bc),
	.w2(32'h3b5cc92d),
	.w3(32'h3cd1be53),
	.w4(32'hbc9fe933),
	.w5(32'h3c26d4bd),
	.w6(32'hbcc9db9b),
	.w7(32'hbd027ded),
	.w8(32'h3aa3f854),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55a34a),
	.w1(32'hbc143702),
	.w2(32'hbb68a772),
	.w3(32'hbb41c13d),
	.w4(32'hbc0b8da8),
	.w5(32'hba72a718),
	.w6(32'hbb838c40),
	.w7(32'hbc1126da),
	.w8(32'h38b8d716),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a370),
	.w1(32'hbbb5ec71),
	.w2(32'h3bcc628e),
	.w3(32'hbac9a54f),
	.w4(32'hbb97c399),
	.w5(32'h3c4a7873),
	.w6(32'hbb1adcb2),
	.w7(32'hbb52721e),
	.w8(32'h3c5262c6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be39c38),
	.w1(32'h3b44a13e),
	.w2(32'h3c9098e3),
	.w3(32'h3c8a2dc1),
	.w4(32'h3c76b29a),
	.w5(32'h3c288d85),
	.w6(32'h3cc0329c),
	.w7(32'h3c5bb3e3),
	.w8(32'h3bdaec38),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca92cae),
	.w1(32'hbc33ad38),
	.w2(32'h3c776a05),
	.w3(32'hbba9435c),
	.w4(32'hbcaaaa3a),
	.w5(32'h3c165929),
	.w6(32'h3c6c71fe),
	.w7(32'hbb9cf935),
	.w8(32'h3c33d7e5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89926b),
	.w1(32'h3baf78cc),
	.w2(32'hbad5159f),
	.w3(32'h3c326c74),
	.w4(32'h3c70c72b),
	.w5(32'hbb77905c),
	.w6(32'h3c4c4624),
	.w7(32'h3be4d1ca),
	.w8(32'hbaf31e55),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe77b7),
	.w1(32'h3a825157),
	.w2(32'hbb0c4405),
	.w3(32'hbb387bcd),
	.w4(32'hbb1a4a54),
	.w5(32'hbc59259b),
	.w6(32'h396615b2),
	.w7(32'h3a440f14),
	.w8(32'h3a0622de),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ef509),
	.w1(32'h3c3e7fbb),
	.w2(32'h3bb30c97),
	.w3(32'hbbd40c5c),
	.w4(32'h3be9982c),
	.w5(32'hbb65f91c),
	.w6(32'hb8a20185),
	.w7(32'h3c0d2f82),
	.w8(32'hbc5d17f1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab166bc),
	.w1(32'h3b071d40),
	.w2(32'h3aa02cae),
	.w3(32'h39920f1f),
	.w4(32'hbafbd127),
	.w5(32'hbaa25ad9),
	.w6(32'h393b50a9),
	.w7(32'hbbdc1d05),
	.w8(32'h39a6a1a0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a853e53),
	.w1(32'hbb3ec973),
	.w2(32'h390f542c),
	.w3(32'hbb562189),
	.w4(32'hbbc971aa),
	.w5(32'hbbbc260c),
	.w6(32'h394f2d54),
	.w7(32'hbb640603),
	.w8(32'hbc3b5fb1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e63d3),
	.w1(32'h3c014c23),
	.w2(32'h3a12fdc7),
	.w3(32'hbc814f70),
	.w4(32'h3b9d16ed),
	.w5(32'hbc34e791),
	.w6(32'hbc1d7696),
	.w7(32'h3a906b15),
	.w8(32'hbc072a51),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cedea),
	.w1(32'h3cab8803),
	.w2(32'h3bade003),
	.w3(32'h3c8eb558),
	.w4(32'h3cc32f7d),
	.w5(32'hbbbe86e2),
	.w6(32'hbb70d21a),
	.w7(32'h3b052025),
	.w8(32'hbb194f5a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b56b),
	.w1(32'h3bced0f4),
	.w2(32'h3c049baa),
	.w3(32'h3a2cbc44),
	.w4(32'h3b78134b),
	.w5(32'hbb719f8f),
	.w6(32'hb82edc76),
	.w7(32'hb9fd8e90),
	.w8(32'hbc161b90),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27dad0),
	.w1(32'hb951d753),
	.w2(32'h3b27c576),
	.w3(32'hbb87d8ec),
	.w4(32'hb9a3e9e3),
	.w5(32'hbab86ce1),
	.w6(32'hbbb1ffc2),
	.w7(32'hbc236ff1),
	.w8(32'hbba64eae),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d66ae),
	.w1(32'h3c50dbff),
	.w2(32'h3c99e5d6),
	.w3(32'h3c174124),
	.w4(32'h3c3db89d),
	.w5(32'h3ca04ae0),
	.w6(32'h3928f83b),
	.w7(32'h3b675978),
	.w8(32'h3b85a636),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9a4d),
	.w1(32'hba3a0b04),
	.w2(32'h3b964cba),
	.w3(32'h3c73d27d),
	.w4(32'hba84efd6),
	.w5(32'hbb8efb03),
	.w6(32'hbc65eb1c),
	.w7(32'hbca005b2),
	.w8(32'hbae7b821),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6472e),
	.w1(32'h3bb8db76),
	.w2(32'h3be4cfd0),
	.w3(32'hbad014d4),
	.w4(32'hba403eb7),
	.w5(32'hbc4f53db),
	.w6(32'hbb65cb56),
	.w7(32'hbbad07dc),
	.w8(32'hbb5cf0cb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d3648),
	.w1(32'h3c40baf9),
	.w2(32'h3c16b701),
	.w3(32'hbb88a4cc),
	.w4(32'hba7a660b),
	.w5(32'h3c05c5f0),
	.w6(32'hbb69265c),
	.w7(32'hbbbcd364),
	.w8(32'hbb01a12e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba484b6),
	.w1(32'hbba3c108),
	.w2(32'h3a7fc532),
	.w3(32'h3aebca8f),
	.w4(32'hbc3d4388),
	.w5(32'hbbc8897d),
	.w6(32'h3b80025e),
	.w7(32'hbb4f0469),
	.w8(32'hbaafa82c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e89f),
	.w1(32'h3a9b0709),
	.w2(32'hbba7efb1),
	.w3(32'h3b134165),
	.w4(32'hb868c1e0),
	.w5(32'hbc45f0f1),
	.w6(32'h3b079241),
	.w7(32'h3c3b2833),
	.w8(32'hbc5c4ce7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa58d),
	.w1(32'hbb9e967a),
	.w2(32'h3a96ac56),
	.w3(32'hbc40db8d),
	.w4(32'hbb0f12e1),
	.w5(32'hbb0ce895),
	.w6(32'hbc15e920),
	.w7(32'h3a650772),
	.w8(32'hbc1df410),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c728e18),
	.w1(32'h3c75f8a8),
	.w2(32'h3af0dea0),
	.w3(32'h3ac97c89),
	.w4(32'h3c203154),
	.w5(32'h3a4a783b),
	.w6(32'hbbd8f033),
	.w7(32'h3a5923d6),
	.w8(32'hbb4f2520),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170e5a),
	.w1(32'h3c1fa593),
	.w2(32'h3b908273),
	.w3(32'h3c05541d),
	.w4(32'h3c174c76),
	.w5(32'hbb154762),
	.w6(32'hbb55e44d),
	.w7(32'hb9a16165),
	.w8(32'hbc7111f0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba370e08),
	.w1(32'hbbb84639),
	.w2(32'h3b87125d),
	.w3(32'hbb8f0a00),
	.w4(32'hbb9ba0ac),
	.w5(32'hbb27616a),
	.w6(32'hbb3917fb),
	.w7(32'hba87b7c8),
	.w8(32'h3b3f3466),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d96f4),
	.w1(32'h3be1ae3a),
	.w2(32'h3b98a600),
	.w3(32'hbbc55174),
	.w4(32'h3a9f875d),
	.w5(32'hbba79359),
	.w6(32'h3b93c703),
	.w7(32'h38bbbada),
	.w8(32'h3ab96f07),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8080c6),
	.w1(32'h3b8ed719),
	.w2(32'h3c20d408),
	.w3(32'hbbd5859c),
	.w4(32'h3b27e561),
	.w5(32'h3b54eb53),
	.w6(32'hbbac2435),
	.w7(32'h3b390033),
	.w8(32'h3ae1dbef),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb8351),
	.w1(32'h3c8172c1),
	.w2(32'hbb393d15),
	.w3(32'h3c431560),
	.w4(32'h3c5710d8),
	.w5(32'hbb2fe02e),
	.w6(32'hbb1532fb),
	.w7(32'h3beea7db),
	.w8(32'hbbf87308),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7731ac),
	.w1(32'h3bd4abc4),
	.w2(32'hbcf433db),
	.w3(32'hbb1cd5fc),
	.w4(32'h3b1de7d0),
	.w5(32'hbd2ff828),
	.w6(32'hbc291088),
	.w7(32'hbbc27032),
	.w8(32'hbcb6b18f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd42450b),
	.w1(32'hbce43e7d),
	.w2(32'h3ab74d9c),
	.w3(32'hbd8ef2db),
	.w4(32'hbd25ee87),
	.w5(32'h3bfe0b68),
	.w6(32'hbd3c7498),
	.w7(32'hbce476c7),
	.w8(32'hb7bb5ceb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbbe74),
	.w1(32'h3c54a436),
	.w2(32'h3ba9ea17),
	.w3(32'h3c546376),
	.w4(32'h3c4bc393),
	.w5(32'h3c851f08),
	.w6(32'hb9aa1bf3),
	.w7(32'hbbb61aac),
	.w8(32'h3bbf7254),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc24e4),
	.w1(32'h3c20c0e7),
	.w2(32'hbbd440f6),
	.w3(32'h3becb7d0),
	.w4(32'hbb0e2c03),
	.w5(32'hbbd656be),
	.w6(32'h3ab83ebe),
	.w7(32'hbb8f85fc),
	.w8(32'hbb56a138),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8a1a7),
	.w1(32'h3c2fa073),
	.w2(32'hbc0d8ee2),
	.w3(32'h3b81d76c),
	.w4(32'h3c17a216),
	.w5(32'hbbd6c189),
	.w6(32'hbc0af529),
	.w7(32'h3b9543b3),
	.w8(32'h3b274da3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba28b4c),
	.w1(32'h39937988),
	.w2(32'hbcb325c0),
	.w3(32'hbc72a6ec),
	.w4(32'hbc3ddc98),
	.w5(32'hbd07106c),
	.w6(32'hbc484b53),
	.w7(32'hbb8e778e),
	.w8(32'hbd01604b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd306697),
	.w1(32'hbcf46f44),
	.w2(32'hbbd80cc1),
	.w3(32'hbd8309b0),
	.w4(32'hbd3fbed6),
	.w5(32'hbb0531b4),
	.w6(32'hbd39baf5),
	.w7(32'hbcd2eb1b),
	.w8(32'hbbd27517),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5acfe),
	.w1(32'hbb727f3f),
	.w2(32'hbc860144),
	.w3(32'hbc0e1f1e),
	.w4(32'hbaadf68d),
	.w5(32'hbcd6add5),
	.w6(32'hbb6a402f),
	.w7(32'h3bf3daad),
	.w8(32'hbccb93cc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27a5c5),
	.w1(32'h3c0b5415),
	.w2(32'h3b85b93c),
	.w3(32'hbcf09b13),
	.w4(32'h3af28bf4),
	.w5(32'hbb20e91d),
	.w6(32'hbd015337),
	.w7(32'hbc6c9798),
	.w8(32'h3bbf4de6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebd29),
	.w1(32'hbc12ada3),
	.w2(32'hbba5b5a7),
	.w3(32'hbc64a404),
	.w4(32'hbc054a91),
	.w5(32'hbb84531a),
	.w6(32'hbc1759ed),
	.w7(32'hbc872982),
	.w8(32'h3c08abd4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0efc36),
	.w1(32'h3bb52661),
	.w2(32'h3b4300ce),
	.w3(32'hbaf14bde),
	.w4(32'h3b402954),
	.w5(32'hba78c9eb),
	.w6(32'h3c10a4b3),
	.w7(32'h3c24101d),
	.w8(32'h3ad5babc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabdea3),
	.w1(32'h3b87193d),
	.w2(32'h3b87afb2),
	.w3(32'hba74dc39),
	.w4(32'h3bbe85d1),
	.w5(32'h3b7a3331),
	.w6(32'h3b369d4f),
	.w7(32'h3b4a2957),
	.w8(32'h3c5e4a5b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8fc53),
	.w1(32'hbc8e2fa7),
	.w2(32'hbb46e374),
	.w3(32'hbcedb21e),
	.w4(32'hbd10a87d),
	.w5(32'hbbec0111),
	.w6(32'hbb7609b4),
	.w7(32'hbc7bdc8f),
	.w8(32'h3b71dea2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bb6ae),
	.w1(32'hbadc9970),
	.w2(32'hbb6db611),
	.w3(32'h3a1c58b3),
	.w4(32'hbb6eca2a),
	.w5(32'hbac5af2a),
	.w6(32'h3826c126),
	.w7(32'hb9107e0b),
	.w8(32'h3ba00852),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc076134),
	.w1(32'hbb61bc80),
	.w2(32'hbc19ab41),
	.w3(32'hbb854719),
	.w4(32'h3ad204b2),
	.w5(32'hbb6232b0),
	.w6(32'hbb8d6419),
	.w7(32'hbb62adc4),
	.w8(32'h3c071dcc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebdc9d),
	.w1(32'h3b0b644a),
	.w2(32'h3b3c3760),
	.w3(32'h3a98eb40),
	.w4(32'h3ba60d2f),
	.w5(32'hba71fe87),
	.w6(32'h3c3279d8),
	.w7(32'h3bfe0268),
	.w8(32'hbbcbc509),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f4eb),
	.w1(32'h3b48107a),
	.w2(32'hbb347a9e),
	.w3(32'h3aec48fd),
	.w4(32'h3b957303),
	.w5(32'hbbe04b47),
	.w6(32'hbb8179ca),
	.w7(32'h3c4af730),
	.w8(32'h3b5c91c2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2264d1),
	.w1(32'hbba5f9db),
	.w2(32'hba3a4b9a),
	.w3(32'hbc1e5e66),
	.w4(32'hbbfe467f),
	.w5(32'h3b8a0b7b),
	.w6(32'hbb943894),
	.w7(32'hbb742bdb),
	.w8(32'hba99c689),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33643a),
	.w1(32'hbc0902c7),
	.w2(32'hbb441daa),
	.w3(32'h3bb1f881),
	.w4(32'hbac71fee),
	.w5(32'hbbb350f8),
	.w6(32'h39e5962a),
	.w7(32'hbba13c12),
	.w8(32'hbb86f835),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1da683),
	.w1(32'h3a695f89),
	.w2(32'hbba0ac8b),
	.w3(32'hbaee084d),
	.w4(32'hba715e9b),
	.w5(32'hbc10fed0),
	.w6(32'hbb472e08),
	.w7(32'hbbaf3e8f),
	.w8(32'hbc5f4f6d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3463),
	.w1(32'h3b3266c1),
	.w2(32'hbbf57c51),
	.w3(32'hbc07de14),
	.w4(32'hbb2d4810),
	.w5(32'hbb1d8ea2),
	.w6(32'hbc401a7b),
	.w7(32'hbab8bb26),
	.w8(32'h3bb4ffdb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aa15a),
	.w1(32'hbc645d07),
	.w2(32'h3c965759),
	.w3(32'hbb6b176b),
	.w4(32'hbc368722),
	.w5(32'h3ca8a903),
	.w6(32'h3b987c21),
	.w7(32'hbb6aa421),
	.w8(32'h3b0090bc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01b795),
	.w1(32'hb9a21b05),
	.w2(32'hbc0271a3),
	.w3(32'h3be2a416),
	.w4(32'hb9d5c142),
	.w5(32'hbc214ad0),
	.w6(32'hbb08dc85),
	.w7(32'h3c16ef78),
	.w8(32'hbb2771a0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf4b98),
	.w1(32'h3b4ad94b),
	.w2(32'hbb062c37),
	.w3(32'hbc6c4736),
	.w4(32'hbc0ebaaf),
	.w5(32'hbb41ea2c),
	.w6(32'hbc20c051),
	.w7(32'hbb9285f5),
	.w8(32'hbb3083a0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5750),
	.w1(32'h3c02ca79),
	.w2(32'h3bc0d70e),
	.w3(32'h3c5a6271),
	.w4(32'h3c4bd8c2),
	.w5(32'h3b5f18b9),
	.w6(32'h3c02911c),
	.w7(32'h3b298498),
	.w8(32'hbc14fe21),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c333cd9),
	.w1(32'h3bfe52d8),
	.w2(32'h3b6bf514),
	.w3(32'h3b32e808),
	.w4(32'h3c09a15d),
	.w5(32'h3ac84c43),
	.w6(32'hbb904092),
	.w7(32'hbb5fa01e),
	.w8(32'hbb963ef0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a90d5),
	.w1(32'h3b220b1b),
	.w2(32'hbb0a939d),
	.w3(32'hbbdd022a),
	.w4(32'hbb8c5a76),
	.w5(32'hbd06a14d),
	.w6(32'hbc0c9337),
	.w7(32'hbbcc18fe),
	.w8(32'hbd228441),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd9fd0),
	.w1(32'h3c9a8543),
	.w2(32'h3b0c6c64),
	.w3(32'hbc8c4eba),
	.w4(32'h3ba6d858),
	.w5(32'hba83e856),
	.w6(32'hbd2096d2),
	.w7(32'hbcb5e818),
	.w8(32'hbc5c08eb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18243d),
	.w1(32'h3c8e901a),
	.w2(32'hbc2c9fed),
	.w3(32'h3b479dee),
	.w4(32'h3bd44a46),
	.w5(32'h3abfbc6b),
	.w6(32'hbb1787ed),
	.w7(32'h3c168ce5),
	.w8(32'h3ba43081),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16be66),
	.w1(32'h3c65e1f9),
	.w2(32'hbcd93a79),
	.w3(32'h3c1c91fc),
	.w4(32'h3c761075),
	.w5(32'hbd00e015),
	.w6(32'h3aef006a),
	.w7(32'h3c6ab3e0),
	.w8(32'hbc85cd99),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd09f3ad),
	.w1(32'hbc1dbd4f),
	.w2(32'hbb99d402),
	.w3(32'hbd4a488b),
	.w4(32'hbd084d47),
	.w5(32'hbc0b17e5),
	.w6(32'hbd017b7a),
	.w7(32'hbcd0e1a3),
	.w8(32'hba3b6788),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88f1f5),
	.w1(32'h3a77fc00),
	.w2(32'h3b2403d6),
	.w3(32'h3b0ba265),
	.w4(32'hbbd26167),
	.w5(32'hba15daa7),
	.w6(32'h3be8911c),
	.w7(32'hb98bd58d),
	.w8(32'hbb787a2e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982c53f),
	.w1(32'h3b3792da),
	.w2(32'h3beb7f6f),
	.w3(32'h3a289702),
	.w4(32'hbb1cfff0),
	.w5(32'h3b5e673d),
	.w6(32'hbb6c66e5),
	.w7(32'hbbb63f30),
	.w8(32'h3baf58a2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a31bc),
	.w1(32'hba0ae599),
	.w2(32'h3b894703),
	.w3(32'h3a55874e),
	.w4(32'hba3f2979),
	.w5(32'h3b96543e),
	.w6(32'h3b9580c9),
	.w7(32'h3af7b854),
	.w8(32'h3b484e32),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca61a82),
	.w1(32'h3b3ebd5b),
	.w2(32'hbc33742c),
	.w3(32'h3c196e8a),
	.w4(32'hb9745d03),
	.w5(32'hbc93c8e3),
	.w6(32'h3b9a0e30),
	.w7(32'hbba001b3),
	.w8(32'hbb89d5b5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7443d),
	.w1(32'h3b32fd03),
	.w2(32'h3ade1a69),
	.w3(32'hbc9a5ac5),
	.w4(32'hbbbe87b7),
	.w5(32'h3ac9903d),
	.w6(32'hbc0fe4df),
	.w7(32'h3b1a118b),
	.w8(32'h39e96c4f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa25b3),
	.w1(32'h3c308ae1),
	.w2(32'h3bdee4d1),
	.w3(32'h3b3137a6),
	.w4(32'h3ad674eb),
	.w5(32'h3c77f4fc),
	.w6(32'hbb92760c),
	.w7(32'h3bf1aa7c),
	.w8(32'h3c412fe0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe3061),
	.w1(32'h3c6d186d),
	.w2(32'hbc060019),
	.w3(32'h3c989d63),
	.w4(32'h3cc284cd),
	.w5(32'hbc1970c2),
	.w6(32'h3bf411a8),
	.w7(32'h3c8462bc),
	.w8(32'hbb1f2f41),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f9fc8),
	.w1(32'hbbc51be7),
	.w2(32'h3b6dade7),
	.w3(32'hbc54fcd8),
	.w4(32'hbb6d0f5e),
	.w5(32'h3b5d2f66),
	.w6(32'hbc3dde23),
	.w7(32'hbba79349),
	.w8(32'h383042be),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39a1d7),
	.w1(32'h3b2d8df5),
	.w2(32'h3adef258),
	.w3(32'hbad2e4a0),
	.w4(32'h3b4c09de),
	.w5(32'h3ba0d2a4),
	.w6(32'hbaded9d1),
	.w7(32'hbb49397b),
	.w8(32'hbad4d478),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e5e35),
	.w1(32'h3c1f8374),
	.w2(32'h3c05d10a),
	.w3(32'h3be1afb8),
	.w4(32'h3bf9586b),
	.w5(32'h3c047b67),
	.w6(32'hbade7686),
	.w7(32'hbbbe5660),
	.w8(32'h3b9671d9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97ef31),
	.w1(32'h3bd54d47),
	.w2(32'h3b7a943c),
	.w3(32'hbb58d98c),
	.w4(32'hbaa9e96e),
	.w5(32'hba470374),
	.w6(32'h3a84942c),
	.w7(32'hbbc07797),
	.w8(32'hbae980c7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb91f),
	.w1(32'h3c1c4f6e),
	.w2(32'h3c8bc0ec),
	.w3(32'hbc724036),
	.w4(32'hbb995654),
	.w5(32'h3cca2d15),
	.w6(32'hbcbac46e),
	.w7(32'hbc82c346),
	.w8(32'h3d16f64c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa0c7e),
	.w1(32'hbcc309e2),
	.w2(32'h3a1232c1),
	.w3(32'hbbdfdc04),
	.w4(32'hbc50e962),
	.w5(32'hbb7a28f8),
	.w6(32'h3c9168cd),
	.w7(32'h3c0da01b),
	.w8(32'hbbce26e5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e875c),
	.w1(32'h3b8caf6b),
	.w2(32'h39b3eaa7),
	.w3(32'h3b1071d1),
	.w4(32'hbabb433d),
	.w5(32'hba88cd1e),
	.w6(32'hbb74b12b),
	.w7(32'hbb54e335),
	.w8(32'hbae3aa3e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00da42),
	.w1(32'hbb86de34),
	.w2(32'h3adf2edd),
	.w3(32'hb9edad04),
	.w4(32'hbc16abd2),
	.w5(32'hbc038e7a),
	.w6(32'h3b269045),
	.w7(32'hbb8de3dd),
	.w8(32'h3a17a137),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a0cf),
	.w1(32'h3bb794bd),
	.w2(32'h3c154413),
	.w3(32'h3a1024a5),
	.w4(32'h3985128b),
	.w5(32'h3c4ecd50),
	.w6(32'hbbc434e5),
	.w7(32'h3ac1e210),
	.w8(32'h3c4bde23),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee033),
	.w1(32'h3bde53d5),
	.w2(32'hbcf349c2),
	.w3(32'h3cc7f34f),
	.w4(32'h3c86b7ea),
	.w5(32'hbd2d9fbb),
	.w6(32'h3c346633),
	.w7(32'h3ac402c2),
	.w8(32'hbd1bfd92),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd286950),
	.w1(32'hbc9817c8),
	.w2(32'h3a3cfd1e),
	.w3(32'hbd8c8eb5),
	.w4(32'hbd2afed6),
	.w5(32'h3a0c7933),
	.w6(32'hbd60fe16),
	.w7(32'hbd316fa9),
	.w8(32'h3b961977),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba8b46),
	.w1(32'h3c272bfa),
	.w2(32'hbb9391ec),
	.w3(32'h3b79dc9a),
	.w4(32'h3c86e235),
	.w5(32'hbc1c2d35),
	.w6(32'hb9afb10a),
	.w7(32'h3b543120),
	.w8(32'hbb724823),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cd74a),
	.w1(32'h3bf44137),
	.w2(32'h3997b4ef),
	.w3(32'hbc199761),
	.w4(32'h3c0d8716),
	.w5(32'h3bb34297),
	.w6(32'hbb1691f6),
	.w7(32'h3bac1de7),
	.w8(32'hbb5d18c0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aeb66),
	.w1(32'hbbde7659),
	.w2(32'h3a737fa6),
	.w3(32'hbbec56cc),
	.w4(32'hbc959037),
	.w5(32'hbbd9cf74),
	.w6(32'hbc2b27db),
	.w7(32'hbc81e6db),
	.w8(32'hbb1c1fb8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93e0be),
	.w1(32'h3c2e9751),
	.w2(32'h3907a3d6),
	.w3(32'hbab61189),
	.w4(32'h3adfdff6),
	.w5(32'hbb3ae070),
	.w6(32'hbb6f6412),
	.w7(32'h3a9ed3af),
	.w8(32'hbb96ba0a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44732a),
	.w1(32'h3bcae413),
	.w2(32'hbbdbc61a),
	.w3(32'h3c496ba8),
	.w4(32'h3c6ff795),
	.w5(32'hbbea4b6c),
	.w6(32'h3be32d91),
	.w7(32'h3bde2fb2),
	.w8(32'h3a269e16),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f96c9),
	.w1(32'h3c29145f),
	.w2(32'hbabac49d),
	.w3(32'h3a94ae83),
	.w4(32'h3c3aba97),
	.w5(32'h3b37a21f),
	.w6(32'hba6e3808),
	.w7(32'h3ba92e2b),
	.w8(32'h3b270b5a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399438d2),
	.w1(32'h3bac353a),
	.w2(32'h3ba40b90),
	.w3(32'h3b1716d0),
	.w4(32'h3b0d5c48),
	.w5(32'h3b1a82f8),
	.w6(32'hbb08d705),
	.w7(32'h3b09d6fa),
	.w8(32'hbbb95e13),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aedf2),
	.w1(32'h3bcb4853),
	.w2(32'hbb809554),
	.w3(32'hba61ecb0),
	.w4(32'hbbb9d0af),
	.w5(32'hbc443a4b),
	.w6(32'hbc1af368),
	.w7(32'hbac2c9ce),
	.w8(32'hbb2f36ed),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ed316),
	.w1(32'h3b8bd780),
	.w2(32'hbbc4f778),
	.w3(32'hbbebc4ab),
	.w4(32'hbad555c8),
	.w5(32'hbc80c51d),
	.w6(32'hbb9eb5df),
	.w7(32'h3acb095e),
	.w8(32'hbc51dca2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa66265),
	.w1(32'h3c3282b9),
	.w2(32'hbb8a8aa8),
	.w3(32'hbbf3c849),
	.w4(32'h3bba0b49),
	.w5(32'hbc2f17d8),
	.w6(32'hbc23057c),
	.w7(32'hbae8c969),
	.w8(32'hbbf8a987),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d226fb),
	.w1(32'h3bb0b7cf),
	.w2(32'h3b7278f6),
	.w3(32'hbc3c807a),
	.w4(32'hbb62f8a3),
	.w5(32'h3aa6c7a8),
	.w6(32'hbb5d98fe),
	.w7(32'h3b62d972),
	.w8(32'hbc148d7a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e558),
	.w1(32'h3b7461bc),
	.w2(32'hbb690576),
	.w3(32'h3c285ba2),
	.w4(32'h3bcf0cf3),
	.w5(32'hbc1f91c8),
	.w6(32'h3b4a9e1b),
	.w7(32'hba91f56a),
	.w8(32'hbbf81ea8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32889a),
	.w1(32'hbba1d647),
	.w2(32'h3a8cf104),
	.w3(32'hbc90a739),
	.w4(32'hbbd2b8a4),
	.w5(32'h3a963840),
	.w6(32'hbc997b32),
	.w7(32'hbb84e84c),
	.w8(32'h3a6a6841),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5064b2),
	.w1(32'h3c7409f9),
	.w2(32'h3b82c719),
	.w3(32'h3b81985a),
	.w4(32'h3c4fb74d),
	.w5(32'h3c1f114d),
	.w6(32'h3a79069a),
	.w7(32'h3b967e76),
	.w8(32'h3a926935),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07fa2d),
	.w1(32'h3b9a6fad),
	.w2(32'h3c2e7af3),
	.w3(32'h3bc7e4aa),
	.w4(32'h3b98c5d5),
	.w5(32'h39794fc4),
	.w6(32'h39f8b14d),
	.w7(32'hbabd631c),
	.w8(32'h3b4a1765),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cfc93),
	.w1(32'h3c3ffcf9),
	.w2(32'h3b816ea4),
	.w3(32'h3abc7883),
	.w4(32'hbbe01bbe),
	.w5(32'hbb2fae80),
	.w6(32'hbbbe87fb),
	.w7(32'hbc250451),
	.w8(32'hbc1bd783),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110c65),
	.w1(32'hbae25ba5),
	.w2(32'h3bf5ada4),
	.w3(32'hbb808a0f),
	.w4(32'h3bfddd2b),
	.w5(32'hbbc6999a),
	.w6(32'hbbdba52f),
	.w7(32'h3b00744d),
	.w8(32'hbbd3ec34),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0ab9),
	.w1(32'hbb1742b2),
	.w2(32'hbb3f2940),
	.w3(32'hbc37963d),
	.w4(32'h3b946a5e),
	.w5(32'hbab1dd88),
	.w6(32'hbb00acd7),
	.w7(32'h3c4a7df2),
	.w8(32'hbc196903),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c78ee),
	.w1(32'hbbd8349a),
	.w2(32'hbb4971d8),
	.w3(32'hbc078cd1),
	.w4(32'hbbc539a7),
	.w5(32'hbc6e6031),
	.w6(32'hbbe01061),
	.w7(32'hbc09f309),
	.w8(32'hbba0815c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37a1de),
	.w1(32'hbb6bf304),
	.w2(32'hbba4180a),
	.w3(32'hbd16f247),
	.w4(32'hbcfbec44),
	.w5(32'hbbbc38fe),
	.w6(32'hbcbf7965),
	.w7(32'hbc710ddf),
	.w8(32'h3ad3e2d4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc213779),
	.w1(32'hbb788831),
	.w2(32'hbb7986e1),
	.w3(32'hbb762080),
	.w4(32'h3b542f0c),
	.w5(32'h3b04d08d),
	.w6(32'h3bf423e6),
	.w7(32'h3c0023b0),
	.w8(32'h3b8efc43),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf1868),
	.w1(32'h3c9f1abb),
	.w2(32'h3a94a11a),
	.w3(32'h3c836097),
	.w4(32'h3cacdef0),
	.w5(32'h3b9ae87e),
	.w6(32'h3c7e25c7),
	.w7(32'h3c2c638e),
	.w8(32'h3ae3a8e8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62e372),
	.w1(32'h3b8d3457),
	.w2(32'hbc3085a0),
	.w3(32'hba936579),
	.w4(32'h3c4e75bf),
	.w5(32'hbc56fb6c),
	.w6(32'hbbd9d769),
	.w7(32'h3c10ca0f),
	.w8(32'hbbd173c4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36818a),
	.w1(32'h3ac8eab5),
	.w2(32'h3af81782),
	.w3(32'hbc077cd3),
	.w4(32'hbad27d62),
	.w5(32'h3abf0824),
	.w6(32'hbc22f4cd),
	.w7(32'hbac85429),
	.w8(32'h3aab849c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8859fed),
	.w1(32'hbb11a407),
	.w2(32'h3bd58ec3),
	.w3(32'hbae92927),
	.w4(32'hbb8832d1),
	.w5(32'h38830e4d),
	.w6(32'h3b54ccc8),
	.w7(32'h392ef23f),
	.w8(32'hbb49d3a3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ff7ff),
	.w1(32'h3bfae30a),
	.w2(32'hbc421f16),
	.w3(32'hb94ae470),
	.w4(32'h3ab00e10),
	.w5(32'hbcd84020),
	.w6(32'hbb2bea8e),
	.w7(32'hbb192433),
	.w8(32'hbc61913d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b084),
	.w1(32'hb9747d49),
	.w2(32'hbb8d7a75),
	.w3(32'hbcf52280),
	.w4(32'hbcb2673f),
	.w5(32'hbbf760e1),
	.w6(32'hbc85850f),
	.w7(32'hbbef56c6),
	.w8(32'h3ae83a6b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb760207),
	.w1(32'hba5b2278),
	.w2(32'hbc1f2559),
	.w3(32'hbbb5309f),
	.w4(32'hb970b909),
	.w5(32'hbc0d89ba),
	.w6(32'h3b28d8eb),
	.w7(32'h3b1e36e7),
	.w8(32'hbc0bf69f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae80f77),
	.w1(32'hba91f76e),
	.w2(32'h3c2f67a7),
	.w3(32'hbbcf4175),
	.w4(32'h3a60312f),
	.w5(32'h3c3618a1),
	.w6(32'h3a6bc8f3),
	.w7(32'hba9360c4),
	.w8(32'h3c4ead9b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bdfe9),
	.w1(32'h3c43a047),
	.w2(32'h3c6ae6c9),
	.w3(32'h3c447b27),
	.w4(32'hbbb706a1),
	.w5(32'h3b8d3aa4),
	.w6(32'h3c232a73),
	.w7(32'hbbac5759),
	.w8(32'hbb574ab1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe4df5),
	.w1(32'h3c84114b),
	.w2(32'h3c9138d6),
	.w3(32'h3c357b22),
	.w4(32'h3c4835c1),
	.w5(32'hbac01457),
	.w6(32'h3bd9d882),
	.w7(32'h3b8522e1),
	.w8(32'h3a338f71),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule