module layer_10_featuremap_63(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa095),
	.w1(32'h3b418a73),
	.w2(32'h3aeeb823),
	.w3(32'hbc0d53c0),
	.w4(32'h3af24dc1),
	.w5(32'h3b3c7d9b),
	.w6(32'hbc5686b7),
	.w7(32'hbc23bcb4),
	.w8(32'hba91c6a5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993341),
	.w1(32'hbb3fb085),
	.w2(32'h3b91f89a),
	.w3(32'hbc0f1017),
	.w4(32'h3a9fef44),
	.w5(32'h3b8a744b),
	.w6(32'h3b974aae),
	.w7(32'h3b2e1944),
	.w8(32'hbbd34dd5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2138a9),
	.w1(32'h3b726288),
	.w2(32'h3c5cbb8b),
	.w3(32'hbc5cb1e1),
	.w4(32'h3bd1e759),
	.w5(32'h3c857bf3),
	.w6(32'hbc6f20c7),
	.w7(32'h3b593bb0),
	.w8(32'h3ae0bf2a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba32af4),
	.w1(32'h3a9b4f7d),
	.w2(32'hbb168c59),
	.w3(32'h3bc67bd6),
	.w4(32'hbbe9e623),
	.w5(32'hbc8a7e3c),
	.w6(32'hbbb8ee55),
	.w7(32'hbc8578f2),
	.w8(32'hbcb67f5f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed73ed),
	.w1(32'h3c4b81e1),
	.w2(32'hbcd5a8ca),
	.w3(32'hbc4fac9d),
	.w4(32'h3bcc1210),
	.w5(32'h3a90621e),
	.w6(32'hbca30de6),
	.w7(32'hbbda6855),
	.w8(32'h3d2ef643),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf8e7fc),
	.w1(32'h3af1b86a),
	.w2(32'hbbeb292c),
	.w3(32'hbbc7fa35),
	.w4(32'hbb69167b),
	.w5(32'hbc40064c),
	.w6(32'h3d1052a4),
	.w7(32'h3a44d45d),
	.w8(32'hbc0261bc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ea98d),
	.w1(32'hb98c4b72),
	.w2(32'hbacc9287),
	.w3(32'h3aa24fe3),
	.w4(32'h3a072985),
	.w5(32'hbb8537db),
	.w6(32'h3bbeccd8),
	.w7(32'h3ba3b145),
	.w8(32'hbbfebde3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bfd1e),
	.w1(32'h3bdc23e1),
	.w2(32'hbbebc7cb),
	.w3(32'h3bd33eb6),
	.w4(32'h391c0e23),
	.w5(32'hbbe09e60),
	.w6(32'hbbe3d841),
	.w7(32'hbb35266d),
	.w8(32'hbb4cda81),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2142ce),
	.w1(32'h39a2f333),
	.w2(32'h3bbab60e),
	.w3(32'hbc7d472c),
	.w4(32'hbb8d058c),
	.w5(32'h3b30ebc6),
	.w6(32'hbb89fc94),
	.w7(32'hbbd89983),
	.w8(32'hbbacf520),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c07d6),
	.w1(32'h3bfd5225),
	.w2(32'hbab1f69b),
	.w3(32'h3be7bff3),
	.w4(32'h3b62ad0c),
	.w5(32'hb91604a1),
	.w6(32'hbb94ebfb),
	.w7(32'hbc262b94),
	.w8(32'h3b3ea247),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160125),
	.w1(32'h3b5db1d6),
	.w2(32'h3c11d026),
	.w3(32'h3aa5792d),
	.w4(32'h3b06cc23),
	.w5(32'h3c400eba),
	.w6(32'hb9027d66),
	.w7(32'hb8c46efa),
	.w8(32'h3bb8c935),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba6ab3),
	.w1(32'h3bdfb37e),
	.w2(32'hb9cc4ce7),
	.w3(32'h3c72c6ba),
	.w4(32'h3bebdb0c),
	.w5(32'hbb9ae576),
	.w6(32'hbb3dc2d4),
	.w7(32'hbb5ec185),
	.w8(32'hbbe013b4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b646e7b),
	.w1(32'h3af97205),
	.w2(32'h3a393ea5),
	.w3(32'h39d1e731),
	.w4(32'h3a8b8c11),
	.w5(32'h39972559),
	.w6(32'h381bb386),
	.w7(32'h3b6f3f06),
	.w8(32'hbbda641c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf55769),
	.w1(32'h3baaf35d),
	.w2(32'hbca20163),
	.w3(32'h3b7fb7a5),
	.w4(32'h3bd9f847),
	.w5(32'hbc91ba41),
	.w6(32'hbbe47ce1),
	.w7(32'h3b92f61a),
	.w8(32'h3bf0c0ff),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8c7d),
	.w1(32'h3a716934),
	.w2(32'hb99c1731),
	.w3(32'hbcf0f818),
	.w4(32'h3b19d6ed),
	.w5(32'hbbd40618),
	.w6(32'h3ae6f07c),
	.w7(32'h3b20a168),
	.w8(32'hbb581377),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b67c4),
	.w1(32'h3bb73c66),
	.w2(32'hbb8fb0cc),
	.w3(32'hbb8ab9be),
	.w4(32'hb9a2cd22),
	.w5(32'hbb477059),
	.w6(32'hbb28a893),
	.w7(32'hbb7b0c3d),
	.w8(32'h39de91ac),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafee98e),
	.w1(32'h3b08c815),
	.w2(32'hbb409bb3),
	.w3(32'hb9e9ce26),
	.w4(32'h3aac5494),
	.w5(32'hbb9e79ec),
	.w6(32'h3ada5e9a),
	.w7(32'h3a9809d5),
	.w8(32'hba91109d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9044e),
	.w1(32'hbbcbf1cb),
	.w2(32'h3ad08310),
	.w3(32'hbb987154),
	.w4(32'hbb782851),
	.w5(32'h3b231f51),
	.w6(32'h3bba452c),
	.w7(32'h3b948c73),
	.w8(32'hb899c353),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3600c9),
	.w1(32'h3c0cc5fc),
	.w2(32'h3bdf7293),
	.w3(32'h3b27f7e7),
	.w4(32'h3c0e934c),
	.w5(32'hbb2a0fcd),
	.w6(32'hbb2519d2),
	.w7(32'h3ae1d34a),
	.w8(32'hba1e6d08),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf632c9),
	.w1(32'hbc41f9d4),
	.w2(32'hbb4663b1),
	.w3(32'hbbc13508),
	.w4(32'hbc5b6631),
	.w5(32'hbb0b0041),
	.w6(32'hbbd7cae2),
	.w7(32'hbc19eee6),
	.w8(32'h3a0f5a3b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5617ac),
	.w1(32'h3b745114),
	.w2(32'h3c2a1234),
	.w3(32'h39340ca9),
	.w4(32'hba5d9268),
	.w5(32'h3880af21),
	.w6(32'hbb51fdb0),
	.w7(32'hbb5aae7f),
	.w8(32'hbbbcb71b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93ab5c),
	.w1(32'h3c23d233),
	.w2(32'h3b5dbb58),
	.w3(32'h3b816692),
	.w4(32'h3bfb8a52),
	.w5(32'h3b0a6942),
	.w6(32'hbc076b8e),
	.w7(32'hbc2f19f9),
	.w8(32'hbb985ab7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58ef86),
	.w1(32'h3bd75495),
	.w2(32'hbc0d72a5),
	.w3(32'hbbdd208a),
	.w4(32'h3b17e4ce),
	.w5(32'hbc35c58c),
	.w6(32'hbc0fdf51),
	.w7(32'hbc137755),
	.w8(32'hbc08b48c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe82df5),
	.w1(32'hbbb9eedb),
	.w2(32'hbb25c7ac),
	.w3(32'hbbb57ed0),
	.w4(32'hbb955a31),
	.w5(32'hba7285e1),
	.w6(32'hbb4e46d9),
	.w7(32'hbb46ed96),
	.w8(32'hbb5f035f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c058d7c),
	.w1(32'h3bd48137),
	.w2(32'h3b3232cb),
	.w3(32'h3a1d8eb7),
	.w4(32'h3aa98b5d),
	.w5(32'h3b81e7be),
	.w6(32'hbbd0aecd),
	.w7(32'hb9ccb7fc),
	.w8(32'h3c0fc395),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc193616),
	.w1(32'hbc6a1063),
	.w2(32'h3beebe9d),
	.w3(32'hbc13953a),
	.w4(32'hbc2fba1e),
	.w5(32'hbc79172c),
	.w6(32'h3c17d6ec),
	.w7(32'h3c21d3c1),
	.w8(32'hbcb16315),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb915e9),
	.w1(32'h3c930e1c),
	.w2(32'h3ae920b0),
	.w3(32'h3b8d922b),
	.w4(32'h3c61f013),
	.w5(32'h3b4f5200),
	.w6(32'hbca4d552),
	.w7(32'hbb717b2c),
	.w8(32'h3a811abe),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba434912),
	.w1(32'h3a95c8fe),
	.w2(32'h3b00c287),
	.w3(32'hba124cc5),
	.w4(32'h3b81c889),
	.w5(32'hbb0277eb),
	.w6(32'hba5909ed),
	.w7(32'h3b01c9c7),
	.w8(32'hbb135b92),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ba9eb),
	.w1(32'hbc7ac014),
	.w2(32'h3ba857f3),
	.w3(32'hbc98754e),
	.w4(32'hbcb3b441),
	.w5(32'h3d1f57a7),
	.w6(32'hbce3de45),
	.w7(32'hbcb091e8),
	.w8(32'h3c8767f4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0201e),
	.w1(32'hbcbdb0a3),
	.w2(32'h3bea65f9),
	.w3(32'h3c82eece),
	.w4(32'hbb918c3b),
	.w5(32'h3bff2927),
	.w6(32'h3c1ccf38),
	.w7(32'h3c1f23ca),
	.w8(32'h3b83e43d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c107989),
	.w1(32'h3a30bb7e),
	.w2(32'hbb93c476),
	.w3(32'h3c2bdc42),
	.w4(32'h3bbf91b7),
	.w5(32'hbba01b3c),
	.w6(32'h3be438c7),
	.w7(32'h3b0fb7a5),
	.w8(32'hbb4faf61),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61071f),
	.w1(32'h3bc5f1fa),
	.w2(32'hba8a144a),
	.w3(32'hbb55a078),
	.w4(32'h3c69509c),
	.w5(32'h3a936a18),
	.w6(32'hbaf78c55),
	.w7(32'h3cad0393),
	.w8(32'hbb76f81e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac817d2),
	.w1(32'h3b915d6b),
	.w2(32'hbb17feb6),
	.w3(32'h3c42bafd),
	.w4(32'h3c82aa81),
	.w5(32'hbb66416b),
	.w6(32'h3aafdd30),
	.w7(32'h3c8aec92),
	.w8(32'hbadf52e3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5093),
	.w1(32'hbb09a0ea),
	.w2(32'hba9448b0),
	.w3(32'hbb2ae2ed),
	.w4(32'hbb8c4a67),
	.w5(32'hbc17361a),
	.w6(32'hbbbc91c3),
	.w7(32'hbbc33a5a),
	.w8(32'hbb2319e3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a979b97),
	.w1(32'hbbc16d98),
	.w2(32'hbbaa9d05),
	.w3(32'hbcccfe05),
	.w4(32'hbb94fb14),
	.w5(32'hbb96734a),
	.w6(32'hbb5e6dc5),
	.w7(32'h3c1b39be),
	.w8(32'hbb4b7e01),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb17a2),
	.w1(32'hbb0ff667),
	.w2(32'hbc2cedfa),
	.w3(32'hbc1a8345),
	.w4(32'hbbfd9ce7),
	.w5(32'h3b7db7ab),
	.w6(32'hbc2ca8b2),
	.w7(32'hbc0bc456),
	.w8(32'h3c511df5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa39ca),
	.w1(32'h3b01fbfc),
	.w2(32'hbb384c77),
	.w3(32'h3c827ce0),
	.w4(32'h3c81cb52),
	.w5(32'h3b1fb9e5),
	.w6(32'h3ba84bee),
	.w7(32'h3cb1b3bc),
	.w8(32'hbbbace44),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ab76),
	.w1(32'hbb95321a),
	.w2(32'h3b805604),
	.w3(32'h3b322e05),
	.w4(32'hbb966425),
	.w5(32'h3beceb41),
	.w6(32'hbc063e2a),
	.w7(32'hbbd0da11),
	.w8(32'hbbc5b5ad),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b2205),
	.w1(32'hbb2de481),
	.w2(32'hbc101afc),
	.w3(32'hbb2f6c26),
	.w4(32'hbb6efe3e),
	.w5(32'hbb487a65),
	.w6(32'hbb5333f7),
	.w7(32'h3b4ac96a),
	.w8(32'hb9e8e2ee),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb996d33),
	.w1(32'hbc4238d4),
	.w2(32'hbbc79aa6),
	.w3(32'hbbd33e22),
	.w4(32'hbc15ad90),
	.w5(32'hbc27b79c),
	.w6(32'hbc0f6c14),
	.w7(32'hbbd4c46b),
	.w8(32'hbc4e5fed),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08afd1),
	.w1(32'hbada6086),
	.w2(32'h3c4271c8),
	.w3(32'hbc35fc9e),
	.w4(32'hbbf23903),
	.w5(32'h3c228bba),
	.w6(32'hbc379261),
	.w7(32'hbc0779c0),
	.w8(32'h3adede38),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda2e1a),
	.w1(32'h3b8f20c6),
	.w2(32'hb8be4ac3),
	.w3(32'h3b90b120),
	.w4(32'h3c1e8439),
	.w5(32'h3b94b4f2),
	.w6(32'h3a9f65bb),
	.w7(32'hbac0dea5),
	.w8(32'hbb375f9d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b184850),
	.w1(32'h3b65082d),
	.w2(32'hbb6e1dc8),
	.w3(32'hbaf001a7),
	.w4(32'h3ca383a8),
	.w5(32'h3a8e7bf9),
	.w6(32'h3b97b99d),
	.w7(32'h3cbdc185),
	.w8(32'h3a7f7e43),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074264),
	.w1(32'h3a97a8c3),
	.w2(32'h3c71dc60),
	.w3(32'h3b0fa6c3),
	.w4(32'h3bcc4545),
	.w5(32'h3cde0e7b),
	.w6(32'h3bb93590),
	.w7(32'h3c1a0036),
	.w8(32'h3cae6462),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc245f44),
	.w1(32'hbca510a5),
	.w2(32'hbae904a8),
	.w3(32'hbaa17c15),
	.w4(32'hbc896304),
	.w5(32'h3b6a6d02),
	.w6(32'hbaffab5e),
	.w7(32'hbcb925b0),
	.w8(32'h3bbe560c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2afc1),
	.w1(32'h3af11ef0),
	.w2(32'h3c124c1e),
	.w3(32'h3cae16e7),
	.w4(32'hbb5e8f0e),
	.w5(32'h3c2105b0),
	.w6(32'h3bf302d2),
	.w7(32'hbc3c5538),
	.w8(32'h3bb085e8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a3a5b),
	.w1(32'h393d6e8d),
	.w2(32'hba9a7c5c),
	.w3(32'h3c179d20),
	.w4(32'h3b7886c6),
	.w5(32'hbbc36e8d),
	.w6(32'h3c3decfe),
	.w7(32'h3c89c1ed),
	.w8(32'hbb8de7e2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3be64),
	.w1(32'hbc597060),
	.w2(32'h3b1f94da),
	.w3(32'h39ece428),
	.w4(32'hbc582b67),
	.w5(32'h3b9b82c1),
	.w6(32'h3c475eb5),
	.w7(32'h3b13d688),
	.w8(32'h3b43dba3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b943162),
	.w1(32'h3af6a28f),
	.w2(32'hbb9eda7e),
	.w3(32'h3bb9d052),
	.w4(32'h3bc485d8),
	.w5(32'hbc1105a9),
	.w6(32'h3bb40c53),
	.w7(32'h3bae7615),
	.w8(32'hbc398c92),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e088e),
	.w1(32'h3c01a688),
	.w2(32'hbc6bcc00),
	.w3(32'hbc5ae72d),
	.w4(32'h3bb4f169),
	.w5(32'hbcc8da8a),
	.w6(32'hbc6af8f3),
	.w7(32'h3b30e60d),
	.w8(32'hbaf6ae18),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7ae34),
	.w1(32'hba376e28),
	.w2(32'hbc465cbb),
	.w3(32'hbd428c71),
	.w4(32'hbc07b35e),
	.w5(32'hbbaaa803),
	.w6(32'hbc6adbba),
	.w7(32'h3aebeee6),
	.w8(32'h3ba18590),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb362ed4),
	.w1(32'h3c42e528),
	.w2(32'hbc9ff266),
	.w3(32'h3c309361),
	.w4(32'h3c49c04d),
	.w5(32'hbcd66388),
	.w6(32'h3cc13557),
	.w7(32'h3cafada0),
	.w8(32'hbbdeb3d4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce06f72),
	.w1(32'hba9b6c43),
	.w2(32'hbbf05206),
	.w3(32'hbd347208),
	.w4(32'hbc64009e),
	.w5(32'hbc24817e),
	.w6(32'hbcb591c3),
	.w7(32'hbb0425ca),
	.w8(32'hbbe3c600),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ec54f),
	.w1(32'h3c45528d),
	.w2(32'hbc46d9fb),
	.w3(32'h3bec445e),
	.w4(32'h3c517123),
	.w5(32'h3c044b12),
	.w6(32'h3c0b543c),
	.w7(32'h3c86a697),
	.w8(32'h3ac26c70),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e2646),
	.w1(32'hb991a02f),
	.w2(32'hbb4673ec),
	.w3(32'hbc5df41d),
	.w4(32'hbc4ba093),
	.w5(32'hb9c534fe),
	.w6(32'hba23752b),
	.w7(32'h3b17b30c),
	.w8(32'hba51f995),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93a37),
	.w1(32'hbc17091a),
	.w2(32'h3b8673d2),
	.w3(32'h3c310a1c),
	.w4(32'h3c0c4ace),
	.w5(32'h3b1c87a6),
	.w6(32'hbb430cbc),
	.w7(32'h3c3243fc),
	.w8(32'h3b604371),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75510b),
	.w1(32'hbb8c70ac),
	.w2(32'hbc392eca),
	.w3(32'h3a1d4c1a),
	.w4(32'hbba913fc),
	.w5(32'hbc1651f1),
	.w6(32'h3a85c329),
	.w7(32'h3a50ce75),
	.w8(32'hbbf99d04),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b496b4c),
	.w1(32'hba4b6773),
	.w2(32'hbb8f1d0c),
	.w3(32'h3bb12d4b),
	.w4(32'h3c68aafc),
	.w5(32'hbb87f520),
	.w6(32'h3c232c4b),
	.w7(32'h3c3354d7),
	.w8(32'hbc9c1165),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e24ad),
	.w1(32'hbc82b770),
	.w2(32'hbc167c3a),
	.w3(32'hbb70fff5),
	.w4(32'hbc770ff1),
	.w5(32'hbbb42bdb),
	.w6(32'hbc9cb278),
	.w7(32'hbcecff9a),
	.w8(32'h3b8529c3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a015),
	.w1(32'hbbb4b802),
	.w2(32'hbba7671d),
	.w3(32'h3a3daa39),
	.w4(32'h3c1ec9df),
	.w5(32'h3b2906a0),
	.w6(32'h3c360bc6),
	.w7(32'h3c11dddf),
	.w8(32'h3af22e4b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3aa340),
	.w1(32'h3b6e5505),
	.w2(32'h3c18ea8f),
	.w3(32'h3bc5727f),
	.w4(32'h3ae999e1),
	.w5(32'hb897d40e),
	.w6(32'h3b3ba0b7),
	.w7(32'h3b4a6bb4),
	.w8(32'hbc021a34),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe899d),
	.w1(32'hbb82addd),
	.w2(32'hbbe9d080),
	.w3(32'h3bad664f),
	.w4(32'hbb57e683),
	.w5(32'hbb8a8c14),
	.w6(32'hbb648417),
	.w7(32'hba7c6253),
	.w8(32'hbbf80bb5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20648),
	.w1(32'hbb86f057),
	.w2(32'h3a207b7a),
	.w3(32'hbc5ac307),
	.w4(32'hbc5d7ae3),
	.w5(32'h3a03a6e0),
	.w6(32'hbc618156),
	.w7(32'hbc57efde),
	.w8(32'hba2d7292),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becaeb6),
	.w1(32'h3c14ddcf),
	.w2(32'hbbe95e39),
	.w3(32'h3c77a7ca),
	.w4(32'h3ca2a5de),
	.w5(32'hbcae9d47),
	.w6(32'h3c76a68f),
	.w7(32'h3ca8dfe6),
	.w8(32'hbc3f3f9d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf69f68),
	.w1(32'hbb1d8511),
	.w2(32'h3b19b12e),
	.w3(32'hbcd1e7fb),
	.w4(32'hbc4e7067),
	.w5(32'h3c0666fd),
	.w6(32'hbcd24fc3),
	.w7(32'hbc205d52),
	.w8(32'h3c2b3282),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3794bc83),
	.w1(32'hbadf2605),
	.w2(32'hbc1cdfef),
	.w3(32'h3b89a1a6),
	.w4(32'h3b3d7b38),
	.w5(32'hbbbdcce1),
	.w6(32'h3b7cbe84),
	.w7(32'hb74d367c),
	.w8(32'hbbbe6b6f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5583ec),
	.w1(32'hbaf5c6d6),
	.w2(32'hbc68ff3a),
	.w3(32'h3b80bc3c),
	.w4(32'h3b96cb91),
	.w5(32'hbc653a74),
	.w6(32'h3b573997),
	.w7(32'h3bdd0d01),
	.w8(32'h3c119d08),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc841d89),
	.w1(32'h3aa1b27a),
	.w2(32'hbc9409da),
	.w3(32'hbcae105d),
	.w4(32'h3b262acc),
	.w5(32'hbcbd9ad0),
	.w6(32'h3b43cfd2),
	.w7(32'h3b9f01d9),
	.w8(32'hbc947ac0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6850a),
	.w1(32'hbca960cb),
	.w2(32'h3c098aa0),
	.w3(32'hbd3991f9),
	.w4(32'hbd116c2d),
	.w5(32'h3c510761),
	.w6(32'hbd1a673e),
	.w7(32'hbca22d1c),
	.w8(32'h3bbf8464),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c873888),
	.w1(32'h3c46eb46),
	.w2(32'h39a3041b),
	.w3(32'h3cc2d264),
	.w4(32'h3ca73805),
	.w5(32'h3c659d07),
	.w6(32'h3c8b197b),
	.w7(32'h3c665b1d),
	.w8(32'h3c08eb3e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07c575),
	.w1(32'hbbe0a6f0),
	.w2(32'h3aa504a5),
	.w3(32'hba3cf9ed),
	.w4(32'hbb71d7ec),
	.w5(32'hbaa43d50),
	.w6(32'h3b5b1c96),
	.w7(32'hbb93b38f),
	.w8(32'h3a0cbee8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1885f),
	.w1(32'hbb63aaad),
	.w2(32'h3b2054a2),
	.w3(32'hbb8fb0dd),
	.w4(32'hbc0246b6),
	.w5(32'hbb037518),
	.w6(32'hbbf70efb),
	.w7(32'hbc3188a6),
	.w8(32'h39ea273d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08fe44),
	.w1(32'h3b938d42),
	.w2(32'h3b922f4e),
	.w3(32'h3c0aa8bc),
	.w4(32'h3ba818a4),
	.w5(32'hbb60e3b4),
	.w6(32'h3c98bad3),
	.w7(32'h3be6541a),
	.w8(32'hbb834235),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0bec3),
	.w1(32'h3bdd05e8),
	.w2(32'h3b9f9238),
	.w3(32'hbbd4fd8b),
	.w4(32'h3c3cd2d2),
	.w5(32'h3c0eeabe),
	.w6(32'hbbd777f7),
	.w7(32'h3bd1ecf0),
	.w8(32'h3b2563a8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08b7bd),
	.w1(32'hbb1b90a1),
	.w2(32'hbc98b469),
	.w3(32'h3b210ca4),
	.w4(32'hba3ee841),
	.w5(32'hbcc3f935),
	.w6(32'hbac28bc8),
	.w7(32'hbb4ba391),
	.w8(32'hbc710a15),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca19b1),
	.w1(32'hbc828e09),
	.w2(32'hbcc6df43),
	.w3(32'hbd114529),
	.w4(32'hbca0ad30),
	.w5(32'hbd19039b),
	.w6(32'hbcbb39b0),
	.w7(32'hbca597b7),
	.w8(32'hbccdef9f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05c3ed),
	.w1(32'hbc92c1d8),
	.w2(32'hbce7ee83),
	.w3(32'hbd6505b1),
	.w4(32'hbce3cb9f),
	.w5(32'hbcdd61fb),
	.w6(32'hbd0711b0),
	.w7(32'hbc1280ad),
	.w8(32'hbc02efcb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5bf4b),
	.w1(32'hbbec3223),
	.w2(32'h3a7905fa),
	.w3(32'hbd43d6d7),
	.w4(32'hbc43a3d5),
	.w5(32'h3c166c75),
	.w6(32'hbc00eebc),
	.w7(32'h3b8c747b),
	.w8(32'h3b5863fe),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b43b),
	.w1(32'hbc13add1),
	.w2(32'hba43a66b),
	.w3(32'hbbd20106),
	.w4(32'hbb98f632),
	.w5(32'hb9e4d105),
	.w6(32'h3b024f25),
	.w7(32'hbae56ab8),
	.w8(32'hbac6a4c8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13021e),
	.w1(32'h3b18522e),
	.w2(32'hbb9682d2),
	.w3(32'hbb61d67e),
	.w4(32'h3b270a92),
	.w5(32'hbbea6d5d),
	.w6(32'h3aaaeb62),
	.w7(32'h3b135f69),
	.w8(32'hb9eabcab),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01b98),
	.w1(32'hbbe4575d),
	.w2(32'h39b26d91),
	.w3(32'hbbbd6f24),
	.w4(32'h3b29b0a0),
	.w5(32'hb9ae36bc),
	.w6(32'h3b4cb74d),
	.w7(32'h3c1ab1f3),
	.w8(32'h39462493),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ddb1),
	.w1(32'h3b450272),
	.w2(32'hbb8bc488),
	.w3(32'h3bba96e3),
	.w4(32'h3b8ae378),
	.w5(32'hbbe44335),
	.w6(32'h3b3d9239),
	.w7(32'h3b688dd9),
	.w8(32'hbb81945c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce68790),
	.w1(32'h3c8b2b39),
	.w2(32'h3c04dc23),
	.w3(32'h3cc3fc3e),
	.w4(32'h3c82c954),
	.w5(32'h3aa73e99),
	.w6(32'h3b98990c),
	.w7(32'h3c8826fc),
	.w8(32'hbb8107a5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a95ac),
	.w1(32'hbc179c60),
	.w2(32'hba228c1f),
	.w3(32'hbbe32338),
	.w4(32'hbb12e003),
	.w5(32'h3be9c38a),
	.w6(32'h3a30ab14),
	.w7(32'h3be85dfe),
	.w8(32'hb9382428),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b389a8a),
	.w1(32'hbbe5cfcb),
	.w2(32'hbbe8335e),
	.w3(32'h3c491c46),
	.w4(32'hbb25b0c2),
	.w5(32'hbc8f2eb9),
	.w6(32'h3b05827c),
	.w7(32'hbb094358),
	.w8(32'h3c0df491),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa67370),
	.w1(32'hbb6443b5),
	.w2(32'h3a858f31),
	.w3(32'hb8b6a815),
	.w4(32'h3c24cc27),
	.w5(32'h3a06dff3),
	.w6(32'h3cc9012b),
	.w7(32'h3c9dfefb),
	.w8(32'h3b289507),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a933c67),
	.w1(32'hbb95c15d),
	.w2(32'hbb63b8f9),
	.w3(32'hbba8630e),
	.w4(32'hbb784eba),
	.w5(32'hbbe077bf),
	.w6(32'hba7e886b),
	.w7(32'hbb8b18b2),
	.w8(32'hbbfe70fb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5255c),
	.w1(32'hbb1dea35),
	.w2(32'hbc6f858e),
	.w3(32'hbba1e75c),
	.w4(32'hbb355cc5),
	.w5(32'hbccb197a),
	.w6(32'hbb56e124),
	.w7(32'hba446f46),
	.w8(32'hba109ffd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a282e),
	.w1(32'h3b31395a),
	.w2(32'h3bb3004a),
	.w3(32'hbd081a81),
	.w4(32'h3b05f785),
	.w5(32'h3a87384c),
	.w6(32'hbc2e549e),
	.w7(32'h3b96bfbb),
	.w8(32'h3bb27d7e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f1b3b),
	.w1(32'h3a9220cd),
	.w2(32'hbc55065d),
	.w3(32'hbba03ae6),
	.w4(32'h3b74b497),
	.w5(32'hb9e22904),
	.w6(32'h3b5a206e),
	.w7(32'h3c14f382),
	.w8(32'h3bac2043),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2ac1),
	.w1(32'hbc1c0faa),
	.w2(32'hbc487c97),
	.w3(32'h3b84a0b0),
	.w4(32'hba17f6d7),
	.w5(32'hbb45ade2),
	.w6(32'hba9b3503),
	.w7(32'hbbc5310a),
	.w8(32'hbc468b22),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00687b),
	.w1(32'hbc3db533),
	.w2(32'hbbcfd669),
	.w3(32'hbbc8725f),
	.w4(32'hbc90e394),
	.w5(32'hbbcfba6e),
	.w6(32'hbcbf7960),
	.w7(32'hbcc6a52e),
	.w8(32'hbc7fa3c2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84b505),
	.w1(32'hbbbd74ff),
	.w2(32'hbb18c120),
	.w3(32'hbbb299eb),
	.w4(32'hbb3db1d1),
	.w5(32'hb9aa1f5a),
	.w6(32'hbc16bba8),
	.w7(32'hbb9d1758),
	.w8(32'hbb40633a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39610d33),
	.w1(32'hbb02c0e2),
	.w2(32'hbc49585f),
	.w3(32'hb8e8ed02),
	.w4(32'hbaafc50d),
	.w5(32'hbcfcdb2f),
	.w6(32'hbb851df7),
	.w7(32'hbbaa2446),
	.w8(32'hbcdd1dbf),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced450f),
	.w1(32'hbc62937b),
	.w2(32'hbad307a0),
	.w3(32'hbd4668ec),
	.w4(32'hbd154670),
	.w5(32'hbc6259d2),
	.w6(32'hbd26b7c4),
	.w7(32'hbcf9cecc),
	.w8(32'hbc82122d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0cbc7),
	.w1(32'h3b741f4d),
	.w2(32'hbb667016),
	.w3(32'hbb325ec2),
	.w4(32'hbc3a4e7b),
	.w5(32'hbb8925d6),
	.w6(32'hbc5abffb),
	.w7(32'hbc51a76b),
	.w8(32'h3b8e85dc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd249df),
	.w1(32'h3a2e4310),
	.w2(32'h3b1bddb9),
	.w3(32'hbbe400a4),
	.w4(32'hb7f944f9),
	.w5(32'h3b8426b5),
	.w6(32'h3a892698),
	.w7(32'hbbfc2c34),
	.w8(32'h39cafe7c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290f6b),
	.w1(32'h3b197b8b),
	.w2(32'hbc77ebeb),
	.w3(32'hbc4401b7),
	.w4(32'hbc23c469),
	.w5(32'hbc219b56),
	.w6(32'hbb603a6f),
	.w7(32'h3b1f18c0),
	.w8(32'h3c92b10b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ffe3),
	.w1(32'h3cc9899c),
	.w2(32'hbc25e5a4),
	.w3(32'hbbad918e),
	.w4(32'h3cced117),
	.w5(32'hbbecf83b),
	.w6(32'h3c8c13bc),
	.w7(32'h3d2078b1),
	.w8(32'hbc1553f6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b77ef),
	.w1(32'h3b4b29aa),
	.w2(32'hbc091fd2),
	.w3(32'h3b6f9c14),
	.w4(32'hba63d076),
	.w5(32'hbb6d458d),
	.w6(32'hb947e32b),
	.w7(32'hbb85447d),
	.w8(32'hbc2b1ecc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dbb1e),
	.w1(32'h3af852f9),
	.w2(32'hbc7adf92),
	.w3(32'hbc80402b),
	.w4(32'h3b034816),
	.w5(32'hbc94f714),
	.w6(32'hbc41bce0),
	.w7(32'h3bf02d15),
	.w8(32'hbc7685da),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32176b),
	.w1(32'h3bd38616),
	.w2(32'hbaf417da),
	.w3(32'hbc6ab9bd),
	.w4(32'h3bd84c68),
	.w5(32'h3b40bfad),
	.w6(32'hbaf00b4a),
	.w7(32'h3c82747b),
	.w8(32'h3b5dd145),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125d1d),
	.w1(32'h37d2a4bc),
	.w2(32'hbc35ea5d),
	.w3(32'h3c40f3ca),
	.w4(32'h3c140760),
	.w5(32'hbb8da343),
	.w6(32'h3bd3ab40),
	.w7(32'h3c53b6d9),
	.w8(32'h3b9fa27e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7a69),
	.w1(32'h3bb16c6a),
	.w2(32'hbba6bb91),
	.w3(32'h3c16db28),
	.w4(32'h3c84a66f),
	.w5(32'hbb0e1810),
	.w6(32'h3c97968f),
	.w7(32'h3caa5152),
	.w8(32'hbae19f46),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc396e87),
	.w1(32'hb9e6cc7f),
	.w2(32'hbc34beff),
	.w3(32'hbb42d629),
	.w4(32'h3b8d7633),
	.w5(32'hbc380925),
	.w6(32'h3c7247b2),
	.w7(32'h3c96a6ca),
	.w8(32'h3aceeeaa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44667d),
	.w1(32'h3a946831),
	.w2(32'hbbab88a6),
	.w3(32'hbaaac027),
	.w4(32'h3c20a6c3),
	.w5(32'hbb1c0803),
	.w6(32'h3c18e360),
	.w7(32'h3c72884e),
	.w8(32'h3bd4e654),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ba249),
	.w1(32'hbbf07114),
	.w2(32'h3b30fcf1),
	.w3(32'h3a4167fe),
	.w4(32'h3b1307ff),
	.w5(32'h3b85a570),
	.w6(32'h3afbfc98),
	.w7(32'h3adb8e36),
	.w8(32'hbb4f6356),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd74608),
	.w1(32'h3bfbd821),
	.w2(32'h3be9212d),
	.w3(32'h3bcd38c7),
	.w4(32'h3c693843),
	.w5(32'h3b7a4b86),
	.w6(32'h3b7d1388),
	.w7(32'h3a319dd7),
	.w8(32'h3b42e91b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b91c),
	.w1(32'h3a2dc334),
	.w2(32'hbb9c9ed9),
	.w3(32'hbb217b30),
	.w4(32'hbbc7282f),
	.w5(32'hbb1ec37c),
	.w6(32'h3a89b6dc),
	.w7(32'h3bae7b79),
	.w8(32'hbb876898),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bf3cb),
	.w1(32'h3a92f61c),
	.w2(32'h3b051cd9),
	.w3(32'h3b8a3a35),
	.w4(32'h3c9c0eb6),
	.w5(32'hbbd1cbb6),
	.w6(32'h3bc7bc4a),
	.w7(32'h3cba643d),
	.w8(32'h3b7a27e1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0883a1),
	.w1(32'hbb726c2e),
	.w2(32'hbb4ca741),
	.w3(32'hbc916475),
	.w4(32'hbc1e1099),
	.w5(32'hbc0d5258),
	.w6(32'hbc6f77a7),
	.w7(32'hbae90f4a),
	.w8(32'hbb13aa5f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952abdc),
	.w1(32'h3bad65fb),
	.w2(32'h3bab8634),
	.w3(32'h3b25c14c),
	.w4(32'h3c49271f),
	.w5(32'hbb8b6452),
	.w6(32'h3bcfb4c2),
	.w7(32'h3bbfd369),
	.w8(32'hbbea5f54),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b3605),
	.w1(32'h3aaad2b7),
	.w2(32'h3bb932f3),
	.w3(32'hbbbb4854),
	.w4(32'hbba6c5c7),
	.w5(32'h3b8e651d),
	.w6(32'hbc361b6f),
	.w7(32'h3a270c61),
	.w8(32'hbb5ab84d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6703a3),
	.w1(32'h3b29430e),
	.w2(32'h39525c63),
	.w3(32'h3be46829),
	.w4(32'h3c960b7d),
	.w5(32'hbb44871d),
	.w6(32'h3c10cb5b),
	.w7(32'h3cbf911b),
	.w8(32'h3b50da45),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7fca),
	.w1(32'hbc106325),
	.w2(32'h3a83dadb),
	.w3(32'hbc4e6720),
	.w4(32'hbbb90e26),
	.w5(32'h3b2a0561),
	.w6(32'hbc87703d),
	.w7(32'hbbc95ed4),
	.w8(32'hbba8a38e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21c2ad),
	.w1(32'h3bf2a7a8),
	.w2(32'hbaced2d8),
	.w3(32'h3a7fe170),
	.w4(32'hbbb71dd1),
	.w5(32'hbbfde2d8),
	.w6(32'hbbf5d7d2),
	.w7(32'hbc4bf33e),
	.w8(32'hbc214bd6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c209979),
	.w1(32'h3bae97f7),
	.w2(32'h3bc4874b),
	.w3(32'h39d895b6),
	.w4(32'h3ae75c51),
	.w5(32'hbbb477b0),
	.w6(32'hbc14df4b),
	.w7(32'hbbd0946b),
	.w8(32'hbc065cb2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0d7eb),
	.w1(32'h3bbfef3d),
	.w2(32'hbc7ae558),
	.w3(32'hbbd88933),
	.w4(32'hbb748f55),
	.w5(32'hbc5a0e23),
	.w6(32'hbb96a5a6),
	.w7(32'hbb4e2f97),
	.w8(32'hb84e39b3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31c9ba),
	.w1(32'h3bab4466),
	.w2(32'hbb9b77b7),
	.w3(32'hbc1f69fb),
	.w4(32'h3c923016),
	.w5(32'hbc200d16),
	.w6(32'h3c1ecedd),
	.w7(32'h3cb64b84),
	.w8(32'hbb21a83f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc338f9),
	.w1(32'h3b60ae5a),
	.w2(32'hbb3bd35c),
	.w3(32'hba6c1250),
	.w4(32'h3b8730e7),
	.w5(32'hbc38368d),
	.w6(32'hbb8e30a4),
	.w7(32'h3c1949c3),
	.w8(32'hbc265316),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ae7de),
	.w1(32'hbbbb1557),
	.w2(32'h3adcba70),
	.w3(32'hbc869baf),
	.w4(32'hbc8443d7),
	.w5(32'h3b55b3ec),
	.w6(32'hbcbe5410),
	.w7(32'hbcdda119),
	.w8(32'h3b7a4dac),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10ff3c),
	.w1(32'h3b27c1fd),
	.w2(32'h3b7fa6fe),
	.w3(32'h3b902690),
	.w4(32'h3b33ba5c),
	.w5(32'h3b68efb3),
	.w6(32'h3b3c4ffc),
	.w7(32'h3a100dda),
	.w8(32'h3bbcc02e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e6c57),
	.w1(32'hba9292cc),
	.w2(32'hbb9b8b81),
	.w3(32'hbb45db66),
	.w4(32'hbb3acb05),
	.w5(32'h3b112688),
	.w6(32'hbad17065),
	.w7(32'hbb3e5a50),
	.w8(32'h3c1b21d5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374dc8),
	.w1(32'hbba76678),
	.w2(32'h3c13411e),
	.w3(32'hba1dac3e),
	.w4(32'hbb45a73c),
	.w5(32'h3bf4b6af),
	.w6(32'h3c08d5e7),
	.w7(32'h3bf2d56f),
	.w8(32'h3ad011c3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb8527),
	.w1(32'h3a3a84a0),
	.w2(32'hbca651e4),
	.w3(32'h3bd49dea),
	.w4(32'h3980ecab),
	.w5(32'hbc0e5d71),
	.w6(32'h3a7641a3),
	.w7(32'hba6ee264),
	.w8(32'h3c1bba0c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc183acf),
	.w1(32'h3c0cf705),
	.w2(32'hbc616836),
	.w3(32'hbc7f62ff),
	.w4(32'h3c4aa0c2),
	.w5(32'hbbbe1590),
	.w6(32'h3c39c313),
	.w7(32'h3cea9a5b),
	.w8(32'h3b59c191),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ee8c8),
	.w1(32'hbb7b08a9),
	.w2(32'hbc103f80),
	.w3(32'hbc45e09b),
	.w4(32'hbabe0303),
	.w5(32'hbc34e57c),
	.w6(32'h3c3cb952),
	.w7(32'h3c2b2a3b),
	.w8(32'h3a54f504),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce39f9),
	.w1(32'h3a9cf403),
	.w2(32'h3bdd5140),
	.w3(32'hbbdc5dae),
	.w4(32'h3b3a23a4),
	.w5(32'hbbcec50c),
	.w6(32'h3bd3ff37),
	.w7(32'h3c1389f3),
	.w8(32'hbc1f7380),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f301),
	.w1(32'hba2fd5b9),
	.w2(32'h3c34743c),
	.w3(32'h3ba5422e),
	.w4(32'h3ba2d56e),
	.w5(32'hbc7d6abc),
	.w6(32'hbbca6113),
	.w7(32'hb98ce325),
	.w8(32'hbce1e0ff),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d016c2f),
	.w1(32'h3ca3ecff),
	.w2(32'h3caca39d),
	.w3(32'h3bdfd1f8),
	.w4(32'h3cc29cf2),
	.w5(32'h3c3fe22a),
	.w6(32'hbb8f656f),
	.w7(32'h3bbaf92d),
	.w8(32'h3b17d042),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5e0ea),
	.w1(32'h3a9d2b0d),
	.w2(32'hbb49a2b9),
	.w3(32'h3cd8a2e8),
	.w4(32'h3bf2f24a),
	.w5(32'h3b84032b),
	.w6(32'h3bd7fe71),
	.w7(32'hbb7c4989),
	.w8(32'hbbd60d5d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6ba4e),
	.w1(32'h3b28c31e),
	.w2(32'hbc4ff2eb),
	.w3(32'hbc140295),
	.w4(32'h3b693b88),
	.w5(32'hbae48045),
	.w6(32'hbc731254),
	.w7(32'h3b35192e),
	.w8(32'h3bbfeae0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc360537),
	.w1(32'h3c1a4e61),
	.w2(32'h3c2b570e),
	.w3(32'hbb7a6cc2),
	.w4(32'h3caec890),
	.w5(32'h3c527a6d),
	.w6(32'h3c61180c),
	.w7(32'h3c51478d),
	.w8(32'h3c8539e3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c817963),
	.w1(32'h3ac11e0e),
	.w2(32'hbb1b2135),
	.w3(32'h3c6f546a),
	.w4(32'hbafe97a3),
	.w5(32'h3a4ba99c),
	.w6(32'h3c421afc),
	.w7(32'hb9ad7443),
	.w8(32'hb9b3d105),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e63e2),
	.w1(32'hbaaa9674),
	.w2(32'hbc0f09a2),
	.w3(32'hbb497260),
	.w4(32'hb98a188d),
	.w5(32'hbb332ba9),
	.w6(32'hbb43b81e),
	.w7(32'hbb1355db),
	.w8(32'hbadb57bf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee6e25),
	.w1(32'hbb3f544e),
	.w2(32'h3b4c8643),
	.w3(32'h3a8555ed),
	.w4(32'h3b18fac9),
	.w5(32'h3c2b4282),
	.w6(32'h3b95fb66),
	.w7(32'h3ba96526),
	.w8(32'h3c0d4c28),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d93fe),
	.w1(32'hbb3526d0),
	.w2(32'hbc2f5366),
	.w3(32'h3c001f42),
	.w4(32'h3b31b0c2),
	.w5(32'hbc319393),
	.w6(32'h3b795a62),
	.w7(32'hbba6dd5a),
	.w8(32'hbc3e5e80),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ce6ad),
	.w1(32'hbc087cf4),
	.w2(32'hbc11d732),
	.w3(32'hbcb8ae6d),
	.w4(32'hbcaf155d),
	.w5(32'hbbff6e7f),
	.w6(32'hbcfde236),
	.w7(32'hbcd54db3),
	.w8(32'hbb831547),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec19f),
	.w1(32'hbb86c5f4),
	.w2(32'hb993a40a),
	.w3(32'hbbbc9f4a),
	.w4(32'hbbb58f0d),
	.w5(32'hbae22842),
	.w6(32'hbba9ad39),
	.w7(32'hbb4b5475),
	.w8(32'hbc6b5f3f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce4941),
	.w1(32'h39925358),
	.w2(32'h3c4f70a0),
	.w3(32'h3b1f8f75),
	.w4(32'h3c5bb3ae),
	.w5(32'h3c7c8aa4),
	.w6(32'hbbccdbca),
	.w7(32'h3bc37b43),
	.w8(32'h3c0a3ab7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c824586),
	.w1(32'h3c5d55f9),
	.w2(32'h3b90e95e),
	.w3(32'h3c871d84),
	.w4(32'h3c2a480c),
	.w5(32'h3b3dc968),
	.w6(32'h3bfbf728),
	.w7(32'h3b8c5caa),
	.w8(32'hbb3cfbac),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba301eb9),
	.w1(32'hba9ee9e7),
	.w2(32'hbae73335),
	.w3(32'hbc671ad9),
	.w4(32'hbbd7b6ab),
	.w5(32'h3c2f0203),
	.w6(32'hbc469b64),
	.w7(32'hbaeab439),
	.w8(32'hb9a7ffc7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251e5d),
	.w1(32'h3ba4f2fd),
	.w2(32'h3bb5988d),
	.w3(32'h3bcbb35e),
	.w4(32'h3c5fcb8e),
	.w5(32'h3bc1b85c),
	.w6(32'h3c83cfcf),
	.w7(32'h3c59fb51),
	.w8(32'h3a7d0145),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b344b39),
	.w1(32'h3b6feb9c),
	.w2(32'h3afbbbd0),
	.w3(32'h3b56fa2a),
	.w4(32'hba1eab39),
	.w5(32'h3b4de020),
	.w6(32'hba869522),
	.w7(32'hbbf138c6),
	.w8(32'h3b43ab78),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2cf07),
	.w1(32'h3a0dada8),
	.w2(32'h3b18ca44),
	.w3(32'h3b922ce5),
	.w4(32'h3a84bd9f),
	.w5(32'h3bbae0da),
	.w6(32'h3b76493c),
	.w7(32'h39d338b5),
	.w8(32'h3ad32111),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8d8e4),
	.w1(32'h3b0a17a3),
	.w2(32'h3b0beb6a),
	.w3(32'h3c8a6024),
	.w4(32'h3c254772),
	.w5(32'h3b6aedb0),
	.w6(32'h3c2c18cc),
	.w7(32'h3ba23966),
	.w8(32'hbad73727),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814c0e),
	.w1(32'hbadd25ab),
	.w2(32'h3bcc966e),
	.w3(32'h3b8adab5),
	.w4(32'hba909e60),
	.w5(32'hbae2420f),
	.w6(32'hbc069796),
	.w7(32'hbc0da15b),
	.w8(32'hbbd02158),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390d60),
	.w1(32'hbc09fc6d),
	.w2(32'hb9bb80cc),
	.w3(32'h3c2b2bd8),
	.w4(32'h3c4f0dff),
	.w5(32'h3b34945b),
	.w6(32'h3b9abc09),
	.w7(32'h3c7bf515),
	.w8(32'h3c02da12),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8b183),
	.w1(32'h3b99c26f),
	.w2(32'hbbb0bf35),
	.w3(32'h3befc038),
	.w4(32'h3c275e03),
	.w5(32'h3b66738f),
	.w6(32'h3c3eebb1),
	.w7(32'h3c3ffe1c),
	.w8(32'hbb2f4630),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb5c61),
	.w1(32'hba92f74a),
	.w2(32'hbbc5ce92),
	.w3(32'hbc02d92b),
	.w4(32'hbb231b3d),
	.w5(32'hbb9baaeb),
	.w6(32'hbc1bcc3d),
	.w7(32'hbbda3074),
	.w8(32'hba61bc5f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa894),
	.w1(32'hbbe8305f),
	.w2(32'h3b77caec),
	.w3(32'h3bf7e257),
	.w4(32'h3c1f2244),
	.w5(32'h3ba864dd),
	.w6(32'h3c045d6b),
	.w7(32'h3bbb7e47),
	.w8(32'hba27b1f9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe94c),
	.w1(32'hb91d2b48),
	.w2(32'hbb2ebcc5),
	.w3(32'h3b4a0ebf),
	.w4(32'hbafb68f6),
	.w5(32'hbb48b199),
	.w6(32'hbaae4880),
	.w7(32'hbbc9b30e),
	.w8(32'hbb63c967),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb412),
	.w1(32'h3a8d265a),
	.w2(32'h3c83db88),
	.w3(32'hbc150ce6),
	.w4(32'hbad6b45c),
	.w5(32'h3bd860b2),
	.w6(32'hbc087abd),
	.w7(32'hb9e01d02),
	.w8(32'hbbb00cb3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd11c6e),
	.w1(32'h3c426a27),
	.w2(32'hbc42cbb5),
	.w3(32'h3c51ee3e),
	.w4(32'h3bfd2347),
	.w5(32'hbcef2d5e),
	.w6(32'hbaf0735f),
	.w7(32'h3c96f256),
	.w8(32'hbc4e12ff),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf3e8e3),
	.w1(32'hbc986d02),
	.w2(32'h3a535ef3),
	.w3(32'hbd47233a),
	.w4(32'hbd00bff5),
	.w5(32'h394527a4),
	.w6(32'hbce103b8),
	.w7(32'hbb8b58d6),
	.w8(32'hb9e1fee8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31a887),
	.w1(32'hbabd7cce),
	.w2(32'hbae608b3),
	.w3(32'hba54b233),
	.w4(32'hbb1d9175),
	.w5(32'h3aff173e),
	.w6(32'hb856533d),
	.w7(32'hbb1bf62f),
	.w8(32'h3bf6ec6b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c54e3),
	.w1(32'hbbefe435),
	.w2(32'h3b9bbf8b),
	.w3(32'hbac1c225),
	.w4(32'hbabb838c),
	.w5(32'hbbb3e756),
	.w6(32'hb9b301f0),
	.w7(32'h3c2fe41d),
	.w8(32'h3aa65769),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902fc3e),
	.w1(32'hbbbc80f9),
	.w2(32'hb8fe53e1),
	.w3(32'hbcb4cfa9),
	.w4(32'hbc4a6662),
	.w5(32'hba292148),
	.w6(32'hbb3ad838),
	.w7(32'h3b772d9c),
	.w8(32'hbaf4a236),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9642),
	.w1(32'h3b3048cc),
	.w2(32'hbc2c69ca),
	.w3(32'h3af2e44a),
	.w4(32'hb9c81050),
	.w5(32'hbc30acfd),
	.w6(32'hb9d7d5fc),
	.w7(32'hbac20b0a),
	.w8(32'hbc00983e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc221e3d),
	.w1(32'hbbebd065),
	.w2(32'hbb47faa6),
	.w3(32'hbc2f05cf),
	.w4(32'hbc6d5aad),
	.w5(32'hbc2bb901),
	.w6(32'hbba05de6),
	.w7(32'hbc068fbb),
	.w8(32'hbc7e0fa6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05b794),
	.w1(32'h3a57845f),
	.w2(32'hb9e808b7),
	.w3(32'hbc3e8b20),
	.w4(32'h3b340b4a),
	.w5(32'h3b0c67ab),
	.w6(32'hba0ccdd4),
	.w7(32'hbbe794d9),
	.w8(32'h3a5aaca9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc10ae),
	.w1(32'h3b0c4313),
	.w2(32'hbc1c57c3),
	.w3(32'h3b18b312),
	.w4(32'h3b77a7e4),
	.w5(32'hb9ec790d),
	.w6(32'h3b168cf4),
	.w7(32'h3b317868),
	.w8(32'h3b51adc1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b9758),
	.w1(32'h3b8e1f4e),
	.w2(32'h3adaa603),
	.w3(32'h3b64065a),
	.w4(32'h3c640cad),
	.w5(32'hbb1cb865),
	.w6(32'h3c11b4a3),
	.w7(32'h3bab1c01),
	.w8(32'hbb9524fc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804a5a),
	.w1(32'h3b9318bf),
	.w2(32'hba41ecfe),
	.w3(32'hbaca269d),
	.w4(32'hbae843be),
	.w5(32'hbcc6ac9a),
	.w6(32'hbb9dd383),
	.w7(32'hbbb2cab4),
	.w8(32'hbb992c67),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4e109),
	.w1(32'h3b6113d0),
	.w2(32'hba9a2957),
	.w3(32'hbd27a29b),
	.w4(32'hbc97110c),
	.w5(32'hbba808bd),
	.w6(32'hbc8e74c7),
	.w7(32'hbc07a3a2),
	.w8(32'hbba17aed),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52f884),
	.w1(32'h3b8f98c3),
	.w2(32'hbad065ad),
	.w3(32'hba976160),
	.w4(32'hbb186ce7),
	.w5(32'h3b8c4607),
	.w6(32'hbae8ba2e),
	.w7(32'hbb9a0575),
	.w8(32'hbac35cd4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fac15),
	.w1(32'h3c57ba74),
	.w2(32'h3aad8b97),
	.w3(32'h3cb72a51),
	.w4(32'h3cbca936),
	.w5(32'hb9b27d02),
	.w6(32'h3a7695f6),
	.w7(32'h3a1ed776),
	.w8(32'h3b07ea6b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6de47),
	.w1(32'h3ab293ad),
	.w2(32'hbba22684),
	.w3(32'hbafee2d1),
	.w4(32'hbc0af09c),
	.w5(32'hbba36fb9),
	.w6(32'h3bcdc122),
	.w7(32'h3b3c31f8),
	.w8(32'hbc0c65a6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920821a),
	.w1(32'h3b2a6aa7),
	.w2(32'h3a9434fb),
	.w3(32'hbaad5921),
	.w4(32'hbadb982f),
	.w5(32'hbaac7cf9),
	.w6(32'hbc224efb),
	.w7(32'hbbbbbeb2),
	.w8(32'hbc9d1aa7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c957a0c),
	.w1(32'h3c2c2de5),
	.w2(32'hbc965c18),
	.w3(32'h3b8b54b2),
	.w4(32'h3a5fd6d1),
	.w5(32'hbc88c256),
	.w6(32'hbc8345db),
	.w7(32'hbc9ae752),
	.w8(32'hbb8c350c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe5718),
	.w1(32'hbc16c3fa),
	.w2(32'h3a57ad15),
	.w3(32'hbb7b25a6),
	.w4(32'h39d4486c),
	.w5(32'hbb6504bb),
	.w6(32'hbac0ccc5),
	.w7(32'h3bdefede),
	.w8(32'h3a071ef2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72592e),
	.w1(32'h3b092679),
	.w2(32'h3cb19f01),
	.w3(32'hba9d38a8),
	.w4(32'hbaef023e),
	.w5(32'h3b61c40d),
	.w6(32'hbac11d99),
	.w7(32'hbb79c021),
	.w8(32'hbc92e6ad),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc45b30),
	.w1(32'hbb869331),
	.w2(32'hbc2740a9),
	.w3(32'h3b4a7ad7),
	.w4(32'h3bc9153d),
	.w5(32'h3b5ad6e7),
	.w6(32'hbc0c5af2),
	.w7(32'h3c867c39),
	.w8(32'h3c2d6a39),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47be13),
	.w1(32'hbc8a9a10),
	.w2(32'h3c79f7a6),
	.w3(32'hbb3f583b),
	.w4(32'hbadfd7be),
	.w5(32'h3bef7424),
	.w6(32'h3c76ff0e),
	.w7(32'h3c996e5c),
	.w8(32'h3c0c63f2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dd0a7),
	.w1(32'h3b9c0263),
	.w2(32'hbbf7181b),
	.w3(32'hba6a1e04),
	.w4(32'hbc08e9ae),
	.w5(32'h3bce4641),
	.w6(32'hbc00bd5f),
	.w7(32'h3ab2d7da),
	.w8(32'h3c814449),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c336c9f),
	.w1(32'h3b932891),
	.w2(32'h3a86c14a),
	.w3(32'h3be78fea),
	.w4(32'h3b9d6b56),
	.w5(32'hb9917829),
	.w6(32'h3b3b3658),
	.w7(32'hb9f12908),
	.w8(32'h3b553b72),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b965d51),
	.w1(32'h3ac1f17f),
	.w2(32'hbb36f8e9),
	.w3(32'h3a2fd9db),
	.w4(32'h381c9dab),
	.w5(32'h3b0b6ee1),
	.w6(32'h3abbc1c7),
	.w7(32'h3af7a5c1),
	.w8(32'h3bba3f8b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9c4f4),
	.w1(32'h3b99f227),
	.w2(32'hbb2529f7),
	.w3(32'h3c64d51b),
	.w4(32'h3bc33bb2),
	.w5(32'h3b9cf04f),
	.w6(32'h3c20da16),
	.w7(32'h3c249ca9),
	.w8(32'h3bd3d2aa),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea8a75),
	.w1(32'hbb85bbdb),
	.w2(32'hbb70fe8a),
	.w3(32'h3c5089c0),
	.w4(32'h3c83fe6e),
	.w5(32'hbae92692),
	.w6(32'h3c7ec336),
	.w7(32'h3c66d22e),
	.w8(32'hbb9f7e1a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc303f40),
	.w1(32'hbc6efd61),
	.w2(32'hbbefbf5c),
	.w3(32'h3c0338b8),
	.w4(32'h39ba8ac2),
	.w5(32'hbad274ab),
	.w6(32'h3a3f22eb),
	.w7(32'h3c288ddf),
	.w8(32'h3bdf52c8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdb487),
	.w1(32'hbc4b576d),
	.w2(32'hbbc20601),
	.w3(32'h3c73328e),
	.w4(32'h3c193914),
	.w5(32'hbb4f1d81),
	.w6(32'h3c16ecd8),
	.w7(32'h3c75069f),
	.w8(32'h3acd0551),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc321865),
	.w1(32'hbbd4cde4),
	.w2(32'hbb4953e5),
	.w3(32'hbb6eed7d),
	.w4(32'hbbdf68c8),
	.w5(32'h3bbbb46d),
	.w6(32'h3b0b6900),
	.w7(32'hba6e2eef),
	.w8(32'h3ba2d5ab),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca62f78),
	.w1(32'hbbcdf5d9),
	.w2(32'h3bb14d88),
	.w3(32'hbc51e59c),
	.w4(32'h3c2a17f7),
	.w5(32'hbb039fe7),
	.w6(32'h3bce4c8f),
	.w7(32'h3a319953),
	.w8(32'hbc606602),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b700b98),
	.w1(32'h3b970c64),
	.w2(32'h3b448bfe),
	.w3(32'hbcbf2434),
	.w4(32'hbc304abd),
	.w5(32'h3b970a6c),
	.w6(32'hbc8b6e75),
	.w7(32'hbca39713),
	.w8(32'h3b7757bc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fe0c3),
	.w1(32'hbbb47be8),
	.w2(32'hbb90f631),
	.w3(32'h3c1aadd2),
	.w4(32'hbc0e0f9c),
	.w5(32'hbba4c418),
	.w6(32'h3b1c2cae),
	.w7(32'h3c1a88c6),
	.w8(32'h3b52beff),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86aae3),
	.w1(32'hbbd604b1),
	.w2(32'hbb2da581),
	.w3(32'hb95b81ab),
	.w4(32'hbb34e0bb),
	.w5(32'hbb7b4830),
	.w6(32'h3a94e239),
	.w7(32'hb966f454),
	.w8(32'hbc16f8c5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc548d0),
	.w1(32'h3b7b114f),
	.w2(32'hbaf695fe),
	.w3(32'hbb9a79c5),
	.w4(32'h39d0a6f7),
	.w5(32'hbbe5c56f),
	.w6(32'hba47a94a),
	.w7(32'h3b0d493b),
	.w8(32'h3b0b94eb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf88edf),
	.w1(32'hba52fbed),
	.w2(32'hbc752469),
	.w3(32'h3b907bdb),
	.w4(32'h3b66099c),
	.w5(32'h3b7681a3),
	.w6(32'h3c9ca891),
	.w7(32'h3c977f08),
	.w8(32'h3c233d7f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1267b1),
	.w1(32'hbb8735ef),
	.w2(32'hbac32d0e),
	.w3(32'hba1ac582),
	.w4(32'hbb1fdfbe),
	.w5(32'h3b00c074),
	.w6(32'h3b833f51),
	.w7(32'h3c054c3a),
	.w8(32'h3a8e6937),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3529d),
	.w1(32'hbae6e831),
	.w2(32'hbc5b5232),
	.w3(32'hbb67815d),
	.w4(32'hbaedd21e),
	.w5(32'hbc18ba3d),
	.w6(32'h3bb52506),
	.w7(32'h38a6327a),
	.w8(32'h3c285e1a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc396cb2),
	.w1(32'hbbe1fa5a),
	.w2(32'h3b005407),
	.w3(32'h3c223053),
	.w4(32'h3bfb0e50),
	.w5(32'hbc345a57),
	.w6(32'h3cd4f4ce),
	.w7(32'h3cd799a5),
	.w8(32'hbbb8ced2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0abdf7),
	.w1(32'hb9f436be),
	.w2(32'h37fc2378),
	.w3(32'hbbcece70),
	.w4(32'hbc201eb0),
	.w5(32'hbb8a52ca),
	.w6(32'hbb4e3336),
	.w7(32'hbc38f3f0),
	.w8(32'hbb7319a8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4cf3),
	.w1(32'hbb5f06c9),
	.w2(32'hbb664665),
	.w3(32'hbc37a7dd),
	.w4(32'hbc3ff581),
	.w5(32'hbb3acd77),
	.w6(32'h3ae49ebc),
	.w7(32'hbc258fdd),
	.w8(32'h3aa8f63a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e1514),
	.w1(32'hbb1ee84b),
	.w2(32'h3af93582),
	.w3(32'hbaa02745),
	.w4(32'hbb28d4e8),
	.w5(32'hbb08fd0c),
	.w6(32'h3aa05737),
	.w7(32'hbaf7f828),
	.w8(32'h3b0910cf),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d1860),
	.w1(32'h3ab66948),
	.w2(32'h3ba006bd),
	.w3(32'h399a44b2),
	.w4(32'hba9131ea),
	.w5(32'hbc13da0e),
	.w6(32'h3bbc882c),
	.w7(32'h3b6e051b),
	.w8(32'hbc9d0e90),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d054761),
	.w1(32'h3ce5c784),
	.w2(32'hbc14a7c1),
	.w3(32'h3c8c12a0),
	.w4(32'h3c696822),
	.w5(32'h3bf8fcf2),
	.w6(32'hbc920d99),
	.w7(32'hbbe9c01b),
	.w8(32'h3c87ebf8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8df8bf),
	.w1(32'hbc877edd),
	.w2(32'hbb53d469),
	.w3(32'h39ea0ac5),
	.w4(32'hbba57f25),
	.w5(32'hbaafc74a),
	.w6(32'h3c472c3b),
	.w7(32'h3bb3872c),
	.w8(32'hb8f0b6fd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d039a),
	.w1(32'hbb75b2d0),
	.w2(32'h3bcffcfa),
	.w3(32'hba915960),
	.w4(32'hbaa9e368),
	.w5(32'h3b722610),
	.w6(32'h3a4958c4),
	.w7(32'h3b3b88cc),
	.w8(32'hbb735fdf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfcd0e),
	.w1(32'h3b8c1216),
	.w2(32'h3a8cd9c8),
	.w3(32'h3bd7cfce),
	.w4(32'h3b8463f7),
	.w5(32'h3ba8ef85),
	.w6(32'hbafbfb85),
	.w7(32'h3c15ba3b),
	.w8(32'h3b70e9e3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95aa5b),
	.w1(32'h39b24f4c),
	.w2(32'h3cd52725),
	.w3(32'h3b376746),
	.w4(32'h3b9e0120),
	.w5(32'h3b056b4c),
	.w6(32'h3a8f0c40),
	.w7(32'h3afcf607),
	.w8(32'hbc85f2a2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07d00e),
	.w1(32'h3cb7e71b),
	.w2(32'hbc226934),
	.w3(32'hbb7c0b8c),
	.w4(32'hbc1f52a4),
	.w5(32'h3b9f3d87),
	.w6(32'hbcf63d51),
	.w7(32'hbd18317c),
	.w8(32'h3c899e10),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1643bd),
	.w1(32'hbcd5b16c),
	.w2(32'hbb1444d9),
	.w3(32'h3c02cfb7),
	.w4(32'h3c4ed44d),
	.w5(32'hbb8e2882),
	.w6(32'h3d063266),
	.w7(32'h3ce54bbf),
	.w8(32'hba233e8b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68b9fa),
	.w1(32'h38e63832),
	.w2(32'h3b192dda),
	.w3(32'hb983eb69),
	.w4(32'hbb3b1b51),
	.w5(32'hb8e8be3f),
	.w6(32'h3b35a3a6),
	.w7(32'hbade12c3),
	.w8(32'hbb3ea2aa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f180cb),
	.w1(32'hba93c14e),
	.w2(32'hbbfde042),
	.w3(32'hbaaabdb5),
	.w4(32'hbbcd3ed3),
	.w5(32'h3a30c41a),
	.w6(32'hbc518dad),
	.w7(32'hbc3fd6f7),
	.w8(32'h3c8526db),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabc8e5),
	.w1(32'hbce6cb24),
	.w2(32'hbc1659b8),
	.w3(32'hb9b8139e),
	.w4(32'hbc4ba516),
	.w5(32'h3b816f3d),
	.w6(32'h3c1debf0),
	.w7(32'h3b53e5be),
	.w8(32'h3c47bb1d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca62933),
	.w1(32'hbcc47d96),
	.w2(32'hba861d8f),
	.w3(32'hbafaae60),
	.w4(32'hbca3559c),
	.w5(32'hbb082c78),
	.w6(32'h3b575813),
	.w7(32'hbc6cd5d3),
	.w8(32'h3bc8992a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaf624),
	.w1(32'hbbd4fe78),
	.w2(32'hba6f42ac),
	.w3(32'hbbc0baa1),
	.w4(32'hbbc615fd),
	.w5(32'hbae2483c),
	.w6(32'hba287978),
	.w7(32'hba9c6c22),
	.w8(32'hbb0b8f28),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3b448),
	.w1(32'hba98dcb0),
	.w2(32'hbb19cdaa),
	.w3(32'hbb13c0f5),
	.w4(32'hbb36c128),
	.w5(32'hb909965f),
	.w6(32'hbb3b17c1),
	.w7(32'h39a33d80),
	.w8(32'h3ba36139),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0363bd),
	.w1(32'h3c1084e1),
	.w2(32'hbaa06119),
	.w3(32'h3bfa5dbc),
	.w4(32'h3bfb085c),
	.w5(32'hbaa8bb58),
	.w6(32'h3bfc9aac),
	.w7(32'h3c1ce89c),
	.w8(32'hbb332bf3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f68f5),
	.w1(32'h3adaeb99),
	.w2(32'hbbd8eea7),
	.w3(32'h3ab1606b),
	.w4(32'hbb99c854),
	.w5(32'hbbcc92d6),
	.w6(32'hbb104fe0),
	.w7(32'hbbc683ca),
	.w8(32'h3c92f923),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb87b3f),
	.w1(32'h3d015873),
	.w2(32'hba7aa58b),
	.w3(32'h3b70f133),
	.w4(32'h3ac03e4b),
	.w5(32'hb859488c),
	.w6(32'hbc3984d6),
	.w7(32'hbbeca30a),
	.w8(32'h3bf47bb8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d681f),
	.w1(32'hbbd8bdf8),
	.w2(32'h3c1dd904),
	.w3(32'hbb9cc1ec),
	.w4(32'hbbdcffe7),
	.w5(32'h3c2982ed),
	.w6(32'hb941eb39),
	.w7(32'h3b8e0f88),
	.w8(32'h3c479dd9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85e7c1),
	.w1(32'h3b89027d),
	.w2(32'hbb02d70a),
	.w3(32'h3c32239e),
	.w4(32'hbb63c278),
	.w5(32'hbbcaed14),
	.w6(32'h3ae9d755),
	.w7(32'hbc0e42ff),
	.w8(32'hbc98ad90),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85656d),
	.w1(32'h3b756812),
	.w2(32'hbba4e848),
	.w3(32'h3be3b061),
	.w4(32'h3bc5dd01),
	.w5(32'hbb6692c8),
	.w6(32'hbc2dbe1a),
	.w7(32'hba3a4f46),
	.w8(32'h3bb8a5ed),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08fd84),
	.w1(32'hbb435837),
	.w2(32'hbb20987f),
	.w3(32'hbaa072ab),
	.w4(32'hbae253a7),
	.w5(32'hbbf38819),
	.w6(32'h397ebb0c),
	.w7(32'hbb27fa20),
	.w8(32'hbbd37b0d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb324de),
	.w1(32'hbb25fd2a),
	.w2(32'hbbc1cd6a),
	.w3(32'hbb7a76cf),
	.w4(32'hbb998aeb),
	.w5(32'h3b2e60c5),
	.w6(32'hbbdbc786),
	.w7(32'hbb7dd70b),
	.w8(32'h3bcc719a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aa2af),
	.w1(32'hbc123cb4),
	.w2(32'h3bfef652),
	.w3(32'h3c7f43ff),
	.w4(32'h3c55116c),
	.w5(32'hbb5e9d12),
	.w6(32'h3cb9561d),
	.w7(32'h3bdc5228),
	.w8(32'hbc570f4a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b806),
	.w1(32'h3c41a6b7),
	.w2(32'hbb0489d5),
	.w3(32'h3aa490d7),
	.w4(32'hbb8f9153),
	.w5(32'hbb2179ea),
	.w6(32'hbc432030),
	.w7(32'hbc25eb45),
	.w8(32'h3be5fdbe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4b3b8),
	.w1(32'h3afc273b),
	.w2(32'h3aca3948),
	.w3(32'hbac2a5a2),
	.w4(32'hbb1f0bfd),
	.w5(32'h3b3a2a8f),
	.w6(32'h3c807112),
	.w7(32'h3c6d3ffa),
	.w8(32'h3c8d6a3d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e33a9b),
	.w1(32'h3ba04762),
	.w2(32'hbb3f0a91),
	.w3(32'h3b3be9a4),
	.w4(32'h3bc6f388),
	.w5(32'hbb72f27f),
	.w6(32'h3ce171a4),
	.w7(32'h3cd35f5a),
	.w8(32'hbc099875),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf5371),
	.w1(32'hbc2c8804),
	.w2(32'h3a4b69c7),
	.w3(32'hbc08b81d),
	.w4(32'hbc15d045),
	.w5(32'hbb5c3095),
	.w6(32'hbc656eda),
	.w7(32'hbc4afea9),
	.w8(32'hbb896a41),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a299906),
	.w1(32'h3a832524),
	.w2(32'hba510a83),
	.w3(32'hbacdc57d),
	.w4(32'hbb1e2a7d),
	.w5(32'h3ba9cad4),
	.w6(32'hbb52d5fa),
	.w7(32'hbb01e9e3),
	.w8(32'h3bde8aca),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7edb91),
	.w1(32'hbc930841),
	.w2(32'h3c468b47),
	.w3(32'h3acd4f86),
	.w4(32'hbb1209a7),
	.w5(32'h3c6b4dac),
	.w6(32'h3c64116e),
	.w7(32'h3bd6c0ec),
	.w8(32'h3bb9975d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d88d1),
	.w1(32'h3b94dcd3),
	.w2(32'hb94f1a82),
	.w3(32'h3caf98d7),
	.w4(32'h3b9874b9),
	.w5(32'h3b3fa2e4),
	.w6(32'h3c562e81),
	.w7(32'h3b542d0c),
	.w8(32'hbb888aa3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cd14f),
	.w1(32'h3aadbfe8),
	.w2(32'hbbe421fb),
	.w3(32'hbbaea812),
	.w4(32'hbb07c733),
	.w5(32'hbba0bab5),
	.w6(32'hbc281bf7),
	.w7(32'hba9de083),
	.w8(32'h3b5edacb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91beea),
	.w1(32'hbc3049f2),
	.w2(32'hbc2f1be8),
	.w3(32'h3bc80346),
	.w4(32'h3a89741c),
	.w5(32'h3c086791),
	.w6(32'h3cf86deb),
	.w7(32'h3cc5c8c3),
	.w8(32'h3c27a1b6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7986dd),
	.w1(32'hbcbdf564),
	.w2(32'h3b46d0a5),
	.w3(32'hbb9059ac),
	.w4(32'hbb9f5093),
	.w5(32'hbafe9db5),
	.w6(32'h3c8f9a2b),
	.w7(32'h3c520cc2),
	.w8(32'hbb672276),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb709de39),
	.w1(32'hbb883d52),
	.w2(32'hbc266112),
	.w3(32'hba37be86),
	.w4(32'hbb9d35f0),
	.w5(32'hbc26b583),
	.w6(32'h3b215ff8),
	.w7(32'h3b306a6d),
	.w8(32'hbc3d5073),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fffeb),
	.w1(32'h3bd20994),
	.w2(32'h3b77e9a6),
	.w3(32'hbb862fe5),
	.w4(32'h3b6fa458),
	.w5(32'hbab6650e),
	.w6(32'hbc507bfc),
	.w7(32'hbc0cb549),
	.w8(32'hbc1f1035),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f4b2f),
	.w1(32'h39d2008c),
	.w2(32'h3c189ab6),
	.w3(32'hbbd72a26),
	.w4(32'hbac71815),
	.w5(32'h3b2e5b0a),
	.w6(32'hbb468404),
	.w7(32'hbc1fd718),
	.w8(32'hbb554fd0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf33e06),
	.w1(32'h3ba75d71),
	.w2(32'h3bce5980),
	.w3(32'h3c0fd592),
	.w4(32'h3bfa44f3),
	.w5(32'h3b16fc99),
	.w6(32'hbab4b329),
	.w7(32'h3b57f247),
	.w8(32'h3af3be4a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8f1e7),
	.w1(32'h3b8ff939),
	.w2(32'h3bfd3e76),
	.w3(32'h3bece57a),
	.w4(32'h3b5791bd),
	.w5(32'hbbad7925),
	.w6(32'hbb021a41),
	.w7(32'h3b5e7ba5),
	.w8(32'hbc0fb0d2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96150f),
	.w1(32'h3c7e4388),
	.w2(32'hbb6fd08b),
	.w3(32'h3b7a9758),
	.w4(32'h3ade8b88),
	.w5(32'h3b817736),
	.w6(32'hbc85aedf),
	.w7(32'hbb6fd035),
	.w8(32'h3bbd030d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90b9e),
	.w1(32'hbb955b43),
	.w2(32'h3b0201d0),
	.w3(32'h3be12f6b),
	.w4(32'h3bb6ef3f),
	.w5(32'h3a39bee1),
	.w6(32'h39e41831),
	.w7(32'h3b675062),
	.w8(32'h3bb8ab8d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886c69),
	.w1(32'hbb886e92),
	.w2(32'h3b2b6922),
	.w3(32'h3b86ad56),
	.w4(32'hb872cc04),
	.w5(32'hb9e8a432),
	.w6(32'h3ace33b3),
	.w7(32'h3bb0b5ef),
	.w8(32'h3b8757ae),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50865c),
	.w1(32'hbc168911),
	.w2(32'h3c7dbf5d),
	.w3(32'hbb1b5421),
	.w4(32'hbbd4356a),
	.w5(32'h3c96ebf2),
	.w6(32'h3c0abd6a),
	.w7(32'h3aacebcf),
	.w8(32'hbb1f8e37),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41ec8b),
	.w1(32'h3aa41550),
	.w2(32'hbbf42138),
	.w3(32'h3b89386b),
	.w4(32'hbb48e01b),
	.w5(32'h38a147cd),
	.w6(32'h3aee650d),
	.w7(32'h3acf7d07),
	.w8(32'hbb3d65e0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8a33d),
	.w1(32'hbb1a551a),
	.w2(32'hbce82c9a),
	.w3(32'h3ba7bf50),
	.w4(32'h3c0a3e5a),
	.w5(32'hbc7537e5),
	.w6(32'hb941d7d4),
	.w7(32'hbbfaadeb),
	.w8(32'hbb727b34),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8cca3),
	.w1(32'hbc37d102),
	.w2(32'hbc5e34ed),
	.w3(32'h3a772c2c),
	.w4(32'h3a53e12a),
	.w5(32'hbc5bd292),
	.w6(32'h3ca50ca5),
	.w7(32'h3ccf9994),
	.w8(32'hbb54225f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20664e),
	.w1(32'h3be33117),
	.w2(32'hbc356481),
	.w3(32'h3a752959),
	.w4(32'h3b445104),
	.w5(32'hbc1fd45e),
	.w6(32'h3ac22b94),
	.w7(32'hba90bc8c),
	.w8(32'h3aa27f3d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf99d5c),
	.w1(32'h3bd9c16e),
	.w2(32'hbc8e6327),
	.w3(32'h3c81cc63),
	.w4(32'h3c92354b),
	.w5(32'hbc96e751),
	.w6(32'h3b895e96),
	.w7(32'h3b1eb664),
	.w8(32'h3ab105bb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc867eca),
	.w1(32'hbc10c0d7),
	.w2(32'hba1d2a9c),
	.w3(32'hbbdab365),
	.w4(32'h3b0a2ba9),
	.w5(32'hbb803c9d),
	.w6(32'h3c1970a3),
	.w7(32'h3c524ef8),
	.w8(32'hbc3fdc6e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25e8f),
	.w1(32'hbbf9bccf),
	.w2(32'h389d5c24),
	.w3(32'hbc937207),
	.w4(32'hbc471083),
	.w5(32'h3b3f09cf),
	.w6(32'hbc083e69),
	.w7(32'hbb9b3939),
	.w8(32'hba5ee941),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2b6ea),
	.w1(32'h3a559d73),
	.w2(32'h3acbc906),
	.w3(32'hb9b6f263),
	.w4(32'hbaca3ea5),
	.w5(32'hbaf740a1),
	.w6(32'hbb5d41f2),
	.w7(32'hbb7695dd),
	.w8(32'h3b3f8c80),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376334),
	.w1(32'h3bc45768),
	.w2(32'hbb47cfd4),
	.w3(32'hbbf687ba),
	.w4(32'hbb9c8159),
	.w5(32'hbb00af78),
	.w6(32'hbb138b45),
	.w7(32'hbb6d3052),
	.w8(32'h3a5323cd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafb22a),
	.w1(32'hbb330297),
	.w2(32'hbc68bc8d),
	.w3(32'hbad3b39a),
	.w4(32'hbb214797),
	.w5(32'hbc0ebb31),
	.w6(32'h3bc6ebb7),
	.w7(32'h3b72117f),
	.w8(32'h3a38a34e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc994238),
	.w1(32'hbc947119),
	.w2(32'hbae13cb7),
	.w3(32'hbbe8caf4),
	.w4(32'hbc4b6001),
	.w5(32'hbbbcedde),
	.w6(32'hbb9b9585),
	.w7(32'hbbf3cc3d),
	.w8(32'hbc04a795),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17cde3),
	.w1(32'hb9a7d8e4),
	.w2(32'hbc39088e),
	.w3(32'hbb9c664b),
	.w4(32'h3b305493),
	.w5(32'hbc105f83),
	.w6(32'hbbf7f165),
	.w7(32'hbc11b287),
	.w8(32'hbb3b23e6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52bec2),
	.w1(32'hbb87350a),
	.w2(32'h3a01152e),
	.w3(32'hbc2de104),
	.w4(32'h3b6510fe),
	.w5(32'h3a658f78),
	.w6(32'h3c60d264),
	.w7(32'h3cb7de06),
	.w8(32'hbb255be1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c0f53),
	.w1(32'hbadccccc),
	.w2(32'h3baaa1b1),
	.w3(32'hba393c94),
	.w4(32'hb8dcb30d),
	.w5(32'h3a3057a9),
	.w6(32'hbb9704df),
	.w7(32'hbb3e87cd),
	.w8(32'hbb49b808),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3ce7f),
	.w1(32'h3bbb06ea),
	.w2(32'hbc1f7687),
	.w3(32'h3b8f74ed),
	.w4(32'h3a79d583),
	.w5(32'h38975913),
	.w6(32'hbbccc453),
	.w7(32'hbc032967),
	.w8(32'h3cbbdfb8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2f2f7),
	.w1(32'h3b882215),
	.w2(32'h3b14cadc),
	.w3(32'hbb54bcd0),
	.w4(32'hbb9d4c01),
	.w5(32'h3a419a90),
	.w6(32'h3a2e3d21),
	.w7(32'hbadc3987),
	.w8(32'h3b541370),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3071b4),
	.w1(32'hbc075a6f),
	.w2(32'hbc7d8c6d),
	.w3(32'hba8ac050),
	.w4(32'hbb88867c),
	.w5(32'hb9c45664),
	.w6(32'h3951394f),
	.w7(32'h3b8cbafc),
	.w8(32'h3be9dcfa),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d3b23),
	.w1(32'hbbb04131),
	.w2(32'h3c049528),
	.w3(32'h3bcf53f0),
	.w4(32'h3ba7f4d4),
	.w5(32'hbbb52804),
	.w6(32'h3be50867),
	.w7(32'h3bd8ef77),
	.w8(32'hbcbe575f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4d58f),
	.w1(32'h3cb38f5d),
	.w2(32'h3c5e36c5),
	.w3(32'hbbc9f57e),
	.w4(32'h3b679bb6),
	.w5(32'hbb6b6dc9),
	.w6(32'hbd22d13f),
	.w7(32'hbcb32f3b),
	.w8(32'hbcd38412),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf9c4ed),
	.w1(32'h3d131f09),
	.w2(32'h3b1a9d86),
	.w3(32'h3b737a7c),
	.w4(32'h3ad804a9),
	.w5(32'h3a961262),
	.w6(32'hbd48e072),
	.w7(32'hbcf8c743),
	.w8(32'h3b8bbfc3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule