module layer_10_featuremap_221(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbefb9618),
	.w1(32'hbece2bc4),
	.w2(32'hbf534d0a),
	.w3(32'hbf065677),
	.w4(32'hbf3b3e04),
	.w5(32'hbed31428),
	.w6(32'hbd0cbaff),
	.w7(32'h3ef8c9e7),
	.w8(32'hbed369e5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea43ead),
	.w1(32'hbe3366d6),
	.w2(32'hbebce1d6),
	.w3(32'hbead9fcb),
	.w4(32'hbec0073d),
	.w5(32'hbf03ce92),
	.w6(32'hbf5a9a38),
	.w7(32'hbece707b),
	.w8(32'hbe9d4048),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbedf9aa1),
	.w1(32'hbe4ae067),
	.w2(32'hbe724acc),
	.w3(32'hbe69c7e9),
	.w4(32'h3dcc221d),
	.w5(32'hbec90cc6),
	.w6(32'hbe310b22),
	.w7(32'hbe87156d),
	.w8(32'h3dd430ae),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf50daaa),
	.w1(32'h3d844f4f),
	.w2(32'hbefaccf8),
	.w3(32'hbe7a42ab),
	.w4(32'hbdec6560),
	.w5(32'hbea837cf),
	.w6(32'hbea55ae9),
	.w7(32'hbeac53ec),
	.w8(32'h3e7aeaac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf08f819),
	.w1(32'hbda79205),
	.w2(32'hbf3fef23),
	.w3(32'hbed8e64d),
	.w4(32'hbec584af),
	.w5(32'hbed3a14a),
	.w6(32'hbf0b906c),
	.w7(32'hbea8d01f),
	.w8(32'hbeb97766),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbee9f225),
	.w1(32'hbf43121c),
	.w2(32'hbe57d019),
	.w3(32'hbf205379),
	.w4(32'hbeae2364),
	.w5(32'hbed02a10),
	.w6(32'hbe7fb777),
	.w7(32'hbedd07ff),
	.w8(32'h3d5a7451),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec18e53),
	.w1(32'hbe99ec30),
	.w2(32'hbe166ad3),
	.w3(32'hbd55bb6c),
	.w4(32'hbe533a1d),
	.w5(32'h3f256c4e),
	.w6(32'hbdf786f1),
	.w7(32'hbea237f2),
	.w8(32'hbe52e000),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eaa6460),
	.w1(32'hbf2be71e),
	.w2(32'hbf212e1d),
	.w3(32'hbf183391),
	.w4(32'hbee89013),
	.w5(32'hbe8af37d),
	.w6(32'hbec1e402),
	.w7(32'hbedf7cbe),
	.w8(32'hbeecaac6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e906478),
	.w1(32'hbdca39e5),
	.w2(32'hbf355468),
	.w3(32'hbc2bb1a5),
	.w4(32'hbf3d49e2),
	.w5(32'hbf06a693),
	.w6(32'hbeae3a24),
	.w7(32'hbee8e401),
	.w8(32'hbe12c95b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf520b1c),
	.w1(32'hbdab418f),
	.w2(32'hbe8d9f3d),
	.w3(32'hbf7c451f),
	.w4(32'hbe864f00),
	.w5(32'hbe6d2283),
	.w6(32'hbec1d541),
	.w7(32'hbede9fc5),
	.w8(32'h3ef1d67b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbef52938),
	.w1(32'h3c9e7566),
	.w2(32'hbf39a3c3),
	.w3(32'hbdf6e1e4),
	.w4(32'h3d0a1fd8),
	.w5(32'hbf5cdc7e),
	.w6(32'hbd1c6653),
	.w7(32'hbe5eb51b),
	.w8(32'hbf16860e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe47f37b),
	.w1(32'h3c8c8409),
	.w2(32'hbf2637a1),
	.w3(32'hbefa2d77),
	.w4(32'hbf0ec502),
	.w5(32'hbec65a7f),
	.w6(32'hbee85da2),
	.w7(32'hbe9b5b57),
	.w8(32'hbf5094e9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea007b9),
	.w1(32'hbf0ca98f),
	.w2(32'h3f7ec318),
	.w3(32'hbedbf37a),
	.w4(32'h3f3eb244),
	.w5(32'h3f8877ca),
	.w6(32'h3e43af44),
	.w7(32'h3f61529e),
	.w8(32'h3f4a2468),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f417656),
	.w1(32'h3f70015f),
	.w2(32'h3f775970),
	.w3(32'h3f8eec08),
	.w4(32'h3f295113),
	.w5(32'h3f2f83af),
	.w6(32'h3f3c058d),
	.w7(32'h3f87477a),
	.w8(32'h3f71010c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2497ab),
	.w1(32'h3f60e28e),
	.w2(32'h3f896cef),
	.w3(32'h3f6f7489),
	.w4(32'h3f257fd9),
	.w5(32'h3f5fc495),
	.w6(32'h3f830b05),
	.w7(32'h3f77a2df),
	.w8(32'h3f8b61c7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3e22be),
	.w1(32'h3f396110),
	.w2(32'h3f452a30),
	.w3(32'h3f56ca1e),
	.w4(32'h3f8fb31b),
	.w5(32'h3f724bf8),
	.w6(32'h3f279be7),
	.w7(32'h3f25fd8a),
	.w8(32'h3f2c3274),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f86ff73),
	.w1(32'h3f2fde3d),
	.w2(32'h3f131633),
	.w3(32'h3f30d519),
	.w4(32'h3f296ff2),
	.w5(32'h3f2c5748),
	.w6(32'h3fa60e0a),
	.w7(32'h3f574be2),
	.w8(32'h3f1f9e96),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f7882e7),
	.w1(32'h3f23d8d1),
	.w2(32'h3ef0d0c6),
	.w3(32'h3f41ce99),
	.w4(32'h3f36d839),
	.w5(32'h3f461a3c),
	.w6(32'h3f8dd53a),
	.w7(32'h3f1cd465),
	.w8(32'h3f67889e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f347ca5),
	.w1(32'h3f64f82e),
	.w2(32'h3f4d44e4),
	.w3(32'h3f063711),
	.w4(32'h3f82c773),
	.w5(32'h3f7116a3),
	.w6(32'h3f6916cc),
	.w7(32'h3f25c230),
	.w8(32'h3f89e0c2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3a04a5),
	.w1(32'h3f9ba71d),
	.w2(32'h3f4c0074),
	.w3(32'h3f87bdc8),
	.w4(32'h3f355938),
	.w5(32'h3f816b83),
	.w6(32'h3f87b281),
	.w7(32'h3f90ef08),
	.w8(32'h3f3d8727),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f344148),
	.w1(32'h3f2df474),
	.w2(32'h3f7839d4),
	.w3(32'h3f8266a4),
	.w4(32'h3f43193d),
	.w5(32'h3f52c812),
	.w6(32'h3f5c7f8f),
	.w7(32'h3f856483),
	.w8(32'h3f42b544),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f08a1a3),
	.w1(32'h3f92c4fc),
	.w2(32'h3f8d826c),
	.w3(32'h3f231bd1),
	.w4(32'h3f43cb2a),
	.w5(32'h3f44c229),
	.w6(32'h3f0ea099),
	.w7(32'h3f86c698),
	.w8(32'h3f5e0971),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f37afbd),
	.w1(32'h3f8b550b),
	.w2(32'h3f86c7ef),
	.w3(32'h3f4f31b6),
	.w4(32'h3f1b51b6),
	.w5(32'h3f43d811),
	.w6(32'h3f10e639),
	.w7(32'h3f2778ae),
	.w8(32'h3f808eac),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6a2c05),
	.w1(32'h3fa20553),
	.w2(32'h3f38aee5),
	.w3(32'h3f2ceba3),
	.w4(32'h3f674615),
	.w5(32'h3f4b2bcd),
	.w6(32'h3fb5a729),
	.w7(32'h3f135287),
	.w8(32'h3f3ce317),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3b5165),
	.w1(32'h3f2c08c6),
	.w2(32'h3f549f63),
	.w3(32'h3f19b402),
	.w4(32'h3f181905),
	.w5(32'h3f2a0af4),
	.w6(32'h3f596196),
	.w7(32'h3f2fdb1c),
	.w8(32'h3f68b968),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fbb8281),
	.w1(32'h3f8c8207),
	.w2(32'h3f86f07d),
	.w3(32'h3f4f4c0e),
	.w4(32'h3f4bc641),
	.w5(32'h3f3d65f9),
	.w6(32'h3f31da21),
	.w7(32'h3f1a9119),
	.w8(32'h3f7e9387),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f8e4575),
	.w1(32'h3f859d55),
	.w2(32'h3bb3435d),
	.w3(32'h3f9150b5),
	.w4(32'h3f415f80),
	.w5(32'hbe9c0571),
	.w6(32'h3f315412),
	.w7(32'h3fa4fb1b),
	.w8(32'hbdb63433),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe255c90),
	.w1(32'h3bce3e13),
	.w2(32'h3d197c6f),
	.w3(32'h3dcb5a75),
	.w4(32'hbc2fb8ed),
	.w5(32'hbe957282),
	.w6(32'hbeca33a7),
	.w7(32'hbe032962),
	.w8(32'hbd141e2b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d713d40),
	.w1(32'hbeeeb6cd),
	.w2(32'hbe4c9ed0),
	.w3(32'hbe521457),
	.w4(32'hbe2c1bdc),
	.w5(32'hbe69d4d3),
	.w6(32'h3d523e8e),
	.w7(32'hbebd5f9e),
	.w8(32'h3e853e40),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe4a26ce),
	.w1(32'hbcd85481),
	.w2(32'hbe5e4a6f),
	.w3(32'hbe825d53),
	.w4(32'hbc27e85b),
	.w5(32'h3dd4e288),
	.w6(32'h3b8bf71a),
	.w7(32'h3cb61993),
	.w8(32'hbdd37fa3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e6c354c),
	.w1(32'h3d6aa0d6),
	.w2(32'h3d9c64fa),
	.w3(32'hbaef3d05),
	.w4(32'h3ed7e925),
	.w5(32'h3dd60508),
	.w6(32'h3e1cc492),
	.w7(32'h3caa55da),
	.w8(32'h3db4a645),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd247dae),
	.w1(32'hbce9fd88),
	.w2(32'h3e0be5de),
	.w3(32'h3e96e7c0),
	.w4(32'h3df286d4),
	.w5(32'h3dbaea86),
	.w6(32'hbe5a8920),
	.w7(32'h3e13f318),
	.w8(32'h3d2b4973),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdab90da),
	.w1(32'hbe80ed1d),
	.w2(32'hbec680ef),
	.w3(32'hbe53da2c),
	.w4(32'hbe8150a6),
	.w5(32'h3e0acfa1),
	.w6(32'h3cd0d17f),
	.w7(32'h3e5f7a10),
	.w8(32'hbe5e5f5a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de1a81e),
	.w1(32'h3d2cc336),
	.w2(32'h3d8602b6),
	.w3(32'hbd8aacbb),
	.w4(32'hbe50ff40),
	.w5(32'hbeb426a1),
	.w6(32'hbb12e4c3),
	.w7(32'hbe236819),
	.w8(32'hbe251018),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5b40bf),
	.w1(32'hbe2afa9e),
	.w2(32'hbe4ac1ad),
	.w3(32'h3d8fe6ef),
	.w4(32'hbe736147),
	.w5(32'h3e2fbcb2),
	.w6(32'hbda242b6),
	.w7(32'h3e811642),
	.w8(32'hbd932d86),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd35d0fe),
	.w1(32'h3e3c2300),
	.w2(32'hbd42234a),
	.w3(32'hbe101275),
	.w4(32'h3d96567d),
	.w5(32'hbd9cb244),
	.w6(32'hbdafd1c9),
	.w7(32'hbe95e599),
	.w8(32'h3d3aa8c1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe29bb31),
	.w1(32'h3e9c3b69),
	.w2(32'h3d279ff7),
	.w3(32'h3df1dcfd),
	.w4(32'h3e55f5f3),
	.w5(32'h3e15a5e1),
	.w6(32'hbebf0a52),
	.w7(32'h3d57d27e),
	.w8(32'hbdd5b8b3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdfd82d5),
	.w1(32'h3d7968ae),
	.w2(32'hbe4ff0f6),
	.w3(32'hbd53be15),
	.w4(32'h3d9294ec),
	.w5(32'hbdf2e485),
	.w6(32'hbe6bb17c),
	.w7(32'h3dadc657),
	.w8(32'h3de67515),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf9134b),
	.w1(32'hbc8afb04),
	.w2(32'h3dd32ef5),
	.w3(32'h3d3d4f5c),
	.w4(32'hbdcc04ef),
	.w5(32'h3cb503ac),
	.w6(32'h3de85387),
	.w7(32'hbe23415d),
	.w8(32'hbe79f377),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d095a5e),
	.w1(32'hbe7e08e1),
	.w2(32'hbc988ce3),
	.w3(32'hbb0e2930),
	.w4(32'h3e286d04),
	.w5(32'h3d991e59),
	.w6(32'hbdab3b09),
	.w7(32'h3d506291),
	.w8(32'hbb4b9f99),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1025d),
	.w1(32'h3ee6a824),
	.w2(32'hbe44aa4b),
	.w3(32'h3e1f4f99),
	.w4(32'h3de7d759),
	.w5(32'h3e3a20e5),
	.w6(32'h3e42fa17),
	.w7(32'hbbd42770),
	.w8(32'h3ccee4ce),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbce31),
	.w1(32'h3caa97d7),
	.w2(32'h3c9bffea),
	.w3(32'h3cdc69a9),
	.w4(32'h3daf1c64),
	.w5(32'h3cce5a6a),
	.w6(32'h3d05db82),
	.w7(32'h3c9fa258),
	.w8(32'h3c56f447),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0330eb),
	.w1(32'h3d07692d),
	.w2(32'h3cddfe5a),
	.w3(32'h3d1fb941),
	.w4(32'h3d0a1641),
	.w5(32'h3cc06ec9),
	.w6(32'h3c5dee37),
	.w7(32'h3c8b17a7),
	.w8(32'h3ce9efe3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caefc0c),
	.w1(32'h3cf29be5),
	.w2(32'h3c7f0c28),
	.w3(32'h3cafc886),
	.w4(32'h3c70c65f),
	.w5(32'h3c7f8c51),
	.w6(32'h3dd55504),
	.w7(32'h3cc379fe),
	.w8(32'h3d178e8a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f810),
	.w1(32'h3c376b0a),
	.w2(32'h3ce10797),
	.w3(32'h3c2c5da1),
	.w4(32'h3cc4907c),
	.w5(32'h3cafcb51),
	.w6(32'h3cc761d1),
	.w7(32'h3c1ce04a),
	.w8(32'h3c8af201),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd13c80),
	.w1(32'h3c2512b1),
	.w2(32'h3cff3a3e),
	.w3(32'h3cbf064c),
	.w4(32'h3c7e858a),
	.w5(32'h3c1f2aec),
	.w6(32'h3c555548),
	.w7(32'h3d326daf),
	.w8(32'h3c703c32),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1f262),
	.w1(32'h3cdadf5e),
	.w2(32'h3cacefa3),
	.w3(32'h3c59c569),
	.w4(32'h3c426fe0),
	.w5(32'h3ca65855),
	.w6(32'h3cc9c74e),
	.w7(32'h3cbdd850),
	.w8(32'h3cec3677),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4408ec),
	.w1(32'h3d155f77),
	.w2(32'h3c8fdaa9),
	.w3(32'h3c38cb61),
	.w4(32'h3c7d5a27),
	.w5(32'h3cc5d1be),
	.w6(32'h3d451fe5),
	.w7(32'h3cc72d3a),
	.w8(32'h3cec32a8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d155a71),
	.w1(32'h3c3e9d90),
	.w2(32'h3cb5c941),
	.w3(32'h3ca99aef),
	.w4(32'h3c88122a),
	.w5(32'h3c8d350c),
	.w6(32'h3ca2e8d4),
	.w7(32'h3d1c8eb5),
	.w8(32'h3ce5dd38),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ce2b2),
	.w1(32'h3cb377da),
	.w2(32'h3cd599b7),
	.w3(32'h3d580a7b),
	.w4(32'h3d0b8dfe),
	.w5(32'h3cb2bb5f),
	.w6(32'h3cae6022),
	.w7(32'h3ca9ebfd),
	.w8(32'h3ca5ba3c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfee85a),
	.w1(32'h3cd8cdd3),
	.w2(32'h3cf6f7ac),
	.w3(32'h3cbecc2b),
	.w4(32'h3c74e4ff),
	.w5(32'h3d0d57d9),
	.w6(32'h3cc92b58),
	.w7(32'h3c3d1306),
	.w8(32'h3c3329b6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7dee59),
	.w1(32'h3cda3bf6),
	.w2(32'h3d1f801e),
	.w3(32'h3cfd6a1f),
	.w4(32'h3cf121be),
	.w5(32'h3d238679),
	.w6(32'h3ca3a1e6),
	.w7(32'h3c60faa8),
	.w8(32'h3cbe1035),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d8814),
	.w1(32'h3cb695ec),
	.w2(32'h3caa8c9d),
	.w3(32'h3c318b5f),
	.w4(32'h3c870a79),
	.w5(32'h3c8b7166),
	.w6(32'h3c60a53a),
	.w7(32'h3d58b524),
	.w8(32'h3c5e9ff9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd1f49),
	.w1(32'h3ca47f6b),
	.w2(32'h3c46504e),
	.w3(32'h3cf33014),
	.w4(32'h3d19c3fa),
	.w5(32'h3cc4a35b),
	.w6(32'h3cceccc5),
	.w7(32'h3c8d2025),
	.w8(32'h3ccf7cc6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc35ff0),
	.w1(32'h3cea775d),
	.w2(32'h3c1d53ae),
	.w3(32'h3cd9074a),
	.w4(32'h3ccc5ef2),
	.w5(32'h3cee2673),
	.w6(32'h3c2433c2),
	.w7(32'h3c8ad430),
	.w8(32'h3d18d741),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d04f137),
	.w1(32'h3b772a2f),
	.w2(32'h3b0c834b),
	.w3(32'h3bcb77f7),
	.w4(32'h3b0673db),
	.w5(32'h3ad205a5),
	.w6(32'h3be9134e),
	.w7(32'h3acd30a9),
	.w8(32'hbc198c5e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18dcc6),
	.w1(32'h3b601fb9),
	.w2(32'h3c7662fc),
	.w3(32'hbb9af74d),
	.w4(32'hbc40cfea),
	.w5(32'h3c26d242),
	.w6(32'h3bcb533e),
	.w7(32'h3c8ccc03),
	.w8(32'hbc3cfe7b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e80a),
	.w1(32'h3b6519e2),
	.w2(32'h3cb321ba),
	.w3(32'h3ab2ab3d),
	.w4(32'h3af59bd2),
	.w5(32'hbbfcd328),
	.w6(32'hbcacdb8e),
	.w7(32'hbb6cf943),
	.w8(32'hbb5866eb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd8ff5),
	.w1(32'h3bb8b021),
	.w2(32'hbaec53e8),
	.w3(32'h3a588200),
	.w4(32'hb94555d7),
	.w5(32'h3c117251),
	.w6(32'h39b92387),
	.w7(32'hbbaee830),
	.w8(32'h3b899202),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6eee9),
	.w1(32'h3b0d2887),
	.w2(32'hbc05982e),
	.w3(32'h3a81f180),
	.w4(32'hbb3bd21b),
	.w5(32'h3b78d5e0),
	.w6(32'hbc1fb587),
	.w7(32'hbc02aa37),
	.w8(32'h3d011699),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfda2f),
	.w1(32'h3afe88fe),
	.w2(32'h3ad12b82),
	.w3(32'h3c8673f1),
	.w4(32'h3afd0c3d),
	.w5(32'hbbfb2a55),
	.w6(32'h3ac92dcc),
	.w7(32'h3b3fcbe4),
	.w8(32'h3b50bd55),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba453b45),
	.w1(32'h3bdbc0d9),
	.w2(32'h3bea8bd1),
	.w3(32'hbbd2732d),
	.w4(32'hbbbff3a7),
	.w5(32'h3b6a8a49),
	.w6(32'hbc3d305e),
	.w7(32'hbbc28651),
	.w8(32'h3b5eb891),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9b4a),
	.w1(32'h3ba61b19),
	.w2(32'h3c2169a0),
	.w3(32'hb9d013a1),
	.w4(32'hbbf6fca9),
	.w5(32'hbc3d3dc3),
	.w6(32'hbbc9b59f),
	.w7(32'hbb651c88),
	.w8(32'hbab82073),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5b12c),
	.w1(32'h3b3869ba),
	.w2(32'h3ad8d785),
	.w3(32'h3c2e1be3),
	.w4(32'hbca93dd1),
	.w5(32'h3c0d4dcc),
	.w6(32'h3d1f4f81),
	.w7(32'hbc036d16),
	.w8(32'hbb586cb0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24ad34),
	.w1(32'hbbacfe59),
	.w2(32'hbb8b5bcb),
	.w3(32'hbc19a134),
	.w4(32'hbc0c7cad),
	.w5(32'hbc0623b0),
	.w6(32'h3cd5dc58),
	.w7(32'hba872838),
	.w8(32'hbb0f8556),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6d343),
	.w1(32'h3d266f0c),
	.w2(32'h3bbfbbf0),
	.w3(32'h3bac8274),
	.w4(32'h3c427e11),
	.w5(32'h3b4d791b),
	.w6(32'hbb0e3f14),
	.w7(32'hbbbb0fc0),
	.w8(32'h3b0ea132),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d7745),
	.w1(32'hba92153c),
	.w2(32'h3b55f079),
	.w3(32'h391ddf47),
	.w4(32'h3b5c3e3d),
	.w5(32'h3d224775),
	.w6(32'hba61e3eb),
	.w7(32'h3b0474ff),
	.w8(32'hbb2953b8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f2dbe),
	.w1(32'hbb24aae6),
	.w2(32'h3b49f178),
	.w3(32'hbbf3bd09),
	.w4(32'hbc047a68),
	.w5(32'h3c6d5b34),
	.w6(32'h3bd6a4a8),
	.w7(32'hbb811fa8),
	.w8(32'hbc06e7de),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eabf4),
	.w1(32'h3bee7bcd),
	.w2(32'hb99576fe),
	.w3(32'h3ba69037),
	.w4(32'h38013393),
	.w5(32'hbb6028dc),
	.w6(32'h3aab3176),
	.w7(32'h393c2ab4),
	.w8(32'h3b81a912),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd064),
	.w1(32'hbb0255e6),
	.w2(32'hbc461822),
	.w3(32'h3be3f65f),
	.w4(32'hbb3bf61d),
	.w5(32'hbb7e6ccc),
	.w6(32'h3b51f1ff),
	.w7(32'hbbd8f9d7),
	.w8(32'hbb791bba),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba90f),
	.w1(32'h3bc2b94e),
	.w2(32'hbaff3423),
	.w3(32'hba9e69c4),
	.w4(32'h3c13697d),
	.w5(32'h3b7ce398),
	.w6(32'hba9301b9),
	.w7(32'hbbb45fa1),
	.w8(32'hbc58e417),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b95a),
	.w1(32'h3ad0a4fb),
	.w2(32'h3c270850),
	.w3(32'h3c4502b6),
	.w4(32'h3c20f191),
	.w5(32'hba237ff7),
	.w6(32'hbc3ca9be),
	.w7(32'h3bef4eba),
	.w8(32'h3bc6e66a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb54a13),
	.w1(32'hba790d4a),
	.w2(32'h3a3d0428),
	.w3(32'hba154654),
	.w4(32'hbc94b157),
	.w5(32'h3b0030fd),
	.w6(32'h3b14f319),
	.w7(32'hbbe401b7),
	.w8(32'h3c205f44),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9cdcf),
	.w1(32'h37a504df),
	.w2(32'hbb4fe04e),
	.w3(32'hbbcfdca0),
	.w4(32'h3c011ea8),
	.w5(32'h3bd44943),
	.w6(32'h3c289677),
	.w7(32'h3be5f936),
	.w8(32'hbb90a254),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56425d),
	.w1(32'h3ad74388),
	.w2(32'h3ae4e920),
	.w3(32'hbbfdd13e),
	.w4(32'hb880659a),
	.w5(32'hbbdaf87f),
	.w6(32'h3b6aef78),
	.w7(32'hbc196c2e),
	.w8(32'h3c8e7f6f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de4b66),
	.w1(32'h3b53e96a),
	.w2(32'hbb97bc46),
	.w3(32'hbbbf95d1),
	.w4(32'h3c3d2ae4),
	.w5(32'hbc36b231),
	.w6(32'h3bcfb999),
	.w7(32'hba8c6c6d),
	.w8(32'hbb552dc5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c3981),
	.w1(32'h3c08240c),
	.w2(32'h3a9a0020),
	.w3(32'h3c651324),
	.w4(32'hbb90c458),
	.w5(32'hbb25c7fd),
	.w6(32'h3b85a179),
	.w7(32'h3c9ee50a),
	.w8(32'h3ab1ab57),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc5c7c),
	.w1(32'h3a2099ff),
	.w2(32'h3b7a015e),
	.w3(32'hbbeaafb6),
	.w4(32'hba0ee3e7),
	.w5(32'hba50a4b7),
	.w6(32'h3b870f7e),
	.w7(32'h3c2257a4),
	.w8(32'hbad29038),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a54448),
	.w1(32'h3bc02fcf),
	.w2(32'hbbcf5f53),
	.w3(32'hbbf25a7f),
	.w4(32'hb96824a4),
	.w5(32'h3c03130c),
	.w6(32'hbaa7d58e),
	.w7(32'hbbec7110),
	.w8(32'h3cb093d6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e3568),
	.w1(32'hbbbdee36),
	.w2(32'hba86a627),
	.w3(32'h3bca09b6),
	.w4(32'hbb4debdf),
	.w5(32'h3bdcf6e1),
	.w6(32'hba83c83c),
	.w7(32'h3b7992c5),
	.w8(32'hbbcb1e37),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc702038),
	.w1(32'hbbe4d648),
	.w2(32'hbb1f62d9),
	.w3(32'hbb6ce176),
	.w4(32'hbc0a26f9),
	.w5(32'h3c02c862),
	.w6(32'hbcbdfe1e),
	.w7(32'h390b006c),
	.w8(32'h3bc31601),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce27dd),
	.w1(32'h3bc67d39),
	.w2(32'hb9b906a6),
	.w3(32'hbb35a8f6),
	.w4(32'h3b2ed2e9),
	.w5(32'hbb8b292a),
	.w6(32'hbc035212),
	.w7(32'h3c931d32),
	.w8(32'h3c3f971f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc391015),
	.w1(32'hbc9133d6),
	.w2(32'h3c381cb2),
	.w3(32'hba9f6276),
	.w4(32'h3c01d7fb),
	.w5(32'hbbbfedb3),
	.w6(32'hbd1b5c85),
	.w7(32'h3cac1ad2),
	.w8(32'hbce4b250),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87857d),
	.w1(32'hbb31df78),
	.w2(32'h3b3479f6),
	.w3(32'h3cae88d0),
	.w4(32'hbae717c4),
	.w5(32'hbb412002),
	.w6(32'hbc1de933),
	.w7(32'hbc2b153c),
	.w8(32'hb8dd03af),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03ddf),
	.w1(32'hbc879e61),
	.w2(32'hbc2c5b49),
	.w3(32'hbbe4eb9d),
	.w4(32'hbbb1ccbe),
	.w5(32'hbb082206),
	.w6(32'h3b9e8290),
	.w7(32'hbc0aed03),
	.w8(32'hbc9d7135),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b687cce),
	.w1(32'hbc4d7aff),
	.w2(32'h3c407f3d),
	.w3(32'hb9d8af7f),
	.w4(32'hbbe89f2c),
	.w5(32'hbbee1b65),
	.w6(32'h3b672f0c),
	.w7(32'h3af06dae),
	.w8(32'hbb0d8569),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c995b81),
	.w1(32'hb99b1bc3),
	.w2(32'h3b831328),
	.w3(32'hbc07166b),
	.w4(32'hbb8251b2),
	.w5(32'hbbf0c8ce),
	.w6(32'h3b395ae6),
	.w7(32'h3c216892),
	.w8(32'hbc600941),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb738d2f),
	.w1(32'h3b7f58c3),
	.w2(32'h39e32451),
	.w3(32'hbba4b488),
	.w4(32'hbb00f1ec),
	.w5(32'h3c54994f),
	.w6(32'h3ba244cb),
	.w7(32'hbc253d5b),
	.w8(32'hbbbf8a9b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b091fa4),
	.w1(32'h3cd816fc),
	.w2(32'hbb8f5855),
	.w3(32'h39ed09fe),
	.w4(32'h3a463cd6),
	.w5(32'h3b922230),
	.w6(32'hb9783713),
	.w7(32'h3cb23dc7),
	.w8(32'h3b904a6f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc092c2c),
	.w1(32'h39be67d2),
	.w2(32'hb999873a),
	.w3(32'h3c4fad0e),
	.w4(32'h3c268eef),
	.w5(32'hbbb0ce74),
	.w6(32'hbae696ee),
	.w7(32'hbbdca705),
	.w8(32'hbc5ffc8a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92be93),
	.w1(32'hbc017900),
	.w2(32'h3c037cb5),
	.w3(32'hb98c2494),
	.w4(32'hbbbac2cf),
	.w5(32'h39069095),
	.w6(32'hbb83d182),
	.w7(32'hbbd0494d),
	.w8(32'hbac87e6d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe604eb),
	.w1(32'hbaaf6e0f),
	.w2(32'h3b180b38),
	.w3(32'hbca075d0),
	.w4(32'hbc9f455a),
	.w5(32'h3ad25d39),
	.w6(32'h3c5bb192),
	.w7(32'h3cd44aeb),
	.w8(32'hbb23f977),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109d28),
	.w1(32'h3b6012cb),
	.w2(32'h3c9e3f24),
	.w3(32'h39a18f7f),
	.w4(32'h3b5ba0cb),
	.w5(32'hbc004e7c),
	.w6(32'hbc54dc2f),
	.w7(32'hbc3c0c60),
	.w8(32'hbcbcf281),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a123f7d),
	.w1(32'h3c1ed4e3),
	.w2(32'hbaa4e0ee),
	.w3(32'hbbe07758),
	.w4(32'h3bed3717),
	.w5(32'hbbf9433f),
	.w6(32'hbc3edc3c),
	.w7(32'hbbc664b3),
	.w8(32'h3bd9aae3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59032b),
	.w1(32'h3b3001a4),
	.w2(32'h3819d160),
	.w3(32'h3be00ad2),
	.w4(32'h391d896c),
	.w5(32'hbbe1f06d),
	.w6(32'hba938c3b),
	.w7(32'h3beab075),
	.w8(32'h3b832d7a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5a4ae3),
	.w1(32'hbc45a290),
	.w2(32'h3b213cc7),
	.w3(32'hbc768b73),
	.w4(32'h3b26d7d7),
	.w5(32'h3aa56f26),
	.w6(32'h3d0d03fd),
	.w7(32'hbbf17d8c),
	.w8(32'hb978aebb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b914b),
	.w1(32'hbab030a9),
	.w2(32'h3911a9a6),
	.w3(32'hbc27799c),
	.w4(32'hbc5f522c),
	.w5(32'h3b50cc72),
	.w6(32'hbc10a57d),
	.w7(32'hbc8e7098),
	.w8(32'h35343f29),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61abf),
	.w1(32'hbca96d92),
	.w2(32'h3c1372f4),
	.w3(32'h3ae76f36),
	.w4(32'hbc02882d),
	.w5(32'h3b83becd),
	.w6(32'hbd375432),
	.w7(32'hbb99422c),
	.w8(32'hbc1608a9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7db8ee),
	.w1(32'hbba1aa55),
	.w2(32'hbbd69bc4),
	.w3(32'hbaa28dc3),
	.w4(32'hbb7ca17e),
	.w5(32'hbbca0747),
	.w6(32'hbb6d2c12),
	.w7(32'h3c748b23),
	.w8(32'hb945ff59),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fb5c9),
	.w1(32'h38ff0862),
	.w2(32'h3ad19826),
	.w3(32'h3c7fa745),
	.w4(32'hbb8dc447),
	.w5(32'h3c432ad6),
	.w6(32'h3bf6e790),
	.w7(32'h3cba7d14),
	.w8(32'h3a71f6fd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd643),
	.w1(32'h3bdb2f85),
	.w2(32'h3bfc7a13),
	.w3(32'hbc29ed2e),
	.w4(32'hbc8135d8),
	.w5(32'hbb68044b),
	.w6(32'hba99399a),
	.w7(32'h39921afa),
	.w8(32'hbbf5dd76),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f402b),
	.w1(32'h3b8ecdfa),
	.w2(32'h3b071c20),
	.w3(32'h3bfe905e),
	.w4(32'hbc2afa50),
	.w5(32'hba03773e),
	.w6(32'hbb46bd10),
	.w7(32'hbadb9d21),
	.w8(32'h3b6cb9bc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15fab9),
	.w1(32'hb9d45565),
	.w2(32'h3bfa7219),
	.w3(32'h3ad18bd5),
	.w4(32'h3ad54aee),
	.w5(32'h3a084915),
	.w6(32'hbc078e89),
	.w7(32'hbcc18686),
	.w8(32'h3a7bc312),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7529df),
	.w1(32'h3bc3ae8b),
	.w2(32'hbbeba2a3),
	.w3(32'h38c10fc2),
	.w4(32'h3cb0d02b),
	.w5(32'hbbb9aaf1),
	.w6(32'h3b855a18),
	.w7(32'hbc1b4390),
	.w8(32'h3c4778d6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2672c),
	.w1(32'h3bddc5d8),
	.w2(32'hbc169159),
	.w3(32'hbac565c5),
	.w4(32'h391c37dd),
	.w5(32'h3af08f09),
	.w6(32'h3c48d78e),
	.w7(32'h3b1ebc47),
	.w8(32'h3b4c3895),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293405),
	.w1(32'hbc922de8),
	.w2(32'h3b5ed339),
	.w3(32'hbc106b10),
	.w4(32'hbbf8ab32),
	.w5(32'hbb3b9691),
	.w6(32'hbbb145b1),
	.w7(32'hbc0da0e5),
	.w8(32'hbb92236d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98e04d),
	.w1(32'h3c0aecc6),
	.w2(32'h3b496638),
	.w3(32'h3bd1a76f),
	.w4(32'h39c66640),
	.w5(32'h3bf04e78),
	.w6(32'h3b4fce4d),
	.w7(32'h3be638bc),
	.w8(32'hb96a25a0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10a3f7),
	.w1(32'hbb258ad4),
	.w2(32'h39e160d1),
	.w3(32'hbbd9467b),
	.w4(32'hba8219dd),
	.w5(32'hbb6c4c3c),
	.w6(32'h3c49ab8a),
	.w7(32'h3b6bd833),
	.w8(32'hbc8a9628),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac25ba3),
	.w1(32'h3c65f091),
	.w2(32'hbc84c278),
	.w3(32'hbb9d82f3),
	.w4(32'hbb2992e4),
	.w5(32'hba94bf01),
	.w6(32'h3b0dc675),
	.w7(32'h3c0cb5ff),
	.w8(32'h3c57f147),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40559f),
	.w1(32'h3b96e350),
	.w2(32'hbc772a18),
	.w3(32'hbc131fa8),
	.w4(32'h3c31c0d5),
	.w5(32'h3bb14202),
	.w6(32'h3a1e7cfd),
	.w7(32'h3b52ac58),
	.w8(32'hbc345509),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9065df),
	.w1(32'hbc0ba7dd),
	.w2(32'hbcd7b5c2),
	.w3(32'hbb2ef6ac),
	.w4(32'hbb3651af),
	.w5(32'hbc87c3ac),
	.w6(32'h3ca6ca2a),
	.w7(32'h39bdf462),
	.w8(32'h3bba8399),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ae1d8),
	.w1(32'hbc96058b),
	.w2(32'hbbe27bcc),
	.w3(32'hba753fbe),
	.w4(32'h3b18f250),
	.w5(32'hbb7f3460),
	.w6(32'hb92baf26),
	.w7(32'h3b3f03cb),
	.w8(32'hbbba7b5c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c976fdc),
	.w1(32'hbc5a4ba6),
	.w2(32'hbc8feea7),
	.w3(32'hbb91860e),
	.w4(32'hb99f0518),
	.w5(32'hbb17d2f0),
	.w6(32'hbb97a5db),
	.w7(32'h3b3ab61b),
	.w8(32'hbb13b4ef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90d2d7),
	.w1(32'h3b6f35bf),
	.w2(32'hbc13f3d3),
	.w3(32'h3b3caa39),
	.w4(32'hbbc34710),
	.w5(32'h3b318afc),
	.w6(32'hbc451fa1),
	.w7(32'hbc2e824a),
	.w8(32'hbabe4b0a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aeeba),
	.w1(32'hbb2196bd),
	.w2(32'h3c5526d8),
	.w3(32'h3c4420b1),
	.w4(32'hbc1e9a1f),
	.w5(32'h3b88c616),
	.w6(32'h3af54147),
	.w7(32'h3cb9f507),
	.w8(32'hbb3e5517),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2d841),
	.w1(32'hbac5b5bc),
	.w2(32'h3c1552eb),
	.w3(32'hbc5dc461),
	.w4(32'hbbdc6707),
	.w5(32'hbb48b22c),
	.w6(32'h3b79fa7c),
	.w7(32'h3ab97d95),
	.w8(32'h3bae5300),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dc85e),
	.w1(32'h3c8904a1),
	.w2(32'h3c3f1bef),
	.w3(32'h3c58c5d2),
	.w4(32'hbc7cb012),
	.w5(32'h3a6da27c),
	.w6(32'hbaca8395),
	.w7(32'h3c448e22),
	.w8(32'h3bb53f49),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0fdc),
	.w1(32'h3ba4ffff),
	.w2(32'hbcbbd2b5),
	.w3(32'h3a2a90e3),
	.w4(32'h3bc333c7),
	.w5(32'hbcb578cb),
	.w6(32'hbc0e8ee1),
	.w7(32'h3ba0bb46),
	.w8(32'h3b209e96),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba12a0c),
	.w1(32'h3ae62743),
	.w2(32'hbb92f4df),
	.w3(32'hba3aa78c),
	.w4(32'h3b7e1282),
	.w5(32'h3be4f9a7),
	.w6(32'h3b98b884),
	.w7(32'hbb0787b1),
	.w8(32'h3b9fb0a8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3ab7a),
	.w1(32'hbadd8372),
	.w2(32'h3b453a77),
	.w3(32'hbc5f28bf),
	.w4(32'h3c9556f8),
	.w5(32'hba802ca0),
	.w6(32'h3a786518),
	.w7(32'hbcca699f),
	.w8(32'h3c70e91e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8decde),
	.w1(32'h3be6acf0),
	.w2(32'hbc38fb2b),
	.w3(32'h3cd7b89b),
	.w4(32'hbbcbd372),
	.w5(32'h3c81162b),
	.w6(32'hbbe85007),
	.w7(32'hbbba4339),
	.w8(32'hbbcdb49e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7b14c),
	.w1(32'hbbebf566),
	.w2(32'hbb62d7c5),
	.w3(32'h3a1f615c),
	.w4(32'hbba5fa1e),
	.w5(32'hbb1d9a05),
	.w6(32'hbc16791a),
	.w7(32'h3c24b8ba),
	.w8(32'h3ca9c7ef),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46b242),
	.w1(32'hb8bd7a8c),
	.w2(32'hbb130174),
	.w3(32'hbc0aab5b),
	.w4(32'h3b04f25f),
	.w5(32'h39b7e10a),
	.w6(32'h3c7af125),
	.w7(32'hbc258ed8),
	.w8(32'hbb8f06df),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7089b8),
	.w1(32'hbc2e67e3),
	.w2(32'h3cdf1f4a),
	.w3(32'hb9951811),
	.w4(32'hbc0bb4b9),
	.w5(32'hbbfdcb76),
	.w6(32'hbb8c0ff3),
	.w7(32'hbbccca7f),
	.w8(32'h3d232048),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7955),
	.w1(32'h3b3c0d20),
	.w2(32'h3c0f1690),
	.w3(32'hbb49dd49),
	.w4(32'h3cc61f4f),
	.w5(32'hbb04e87b),
	.w6(32'hbc35bdb6),
	.w7(32'hb944fba9),
	.w8(32'h3c55a35b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12297f),
	.w1(32'h332aeb8c),
	.w2(32'hbc556fcc),
	.w3(32'hbb0a9f0f),
	.w4(32'h3bdaa90d),
	.w5(32'hbc3325ce),
	.w6(32'h3bc04cc9),
	.w7(32'hbaf431be),
	.w8(32'hbbeec090),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39514448),
	.w1(32'hb8840bb3),
	.w2(32'h3a99cc3c),
	.w3(32'hbba022ad),
	.w4(32'hbc005a91),
	.w5(32'hba9f07e7),
	.w6(32'hba59dbe7),
	.w7(32'h3bf6ec4c),
	.w8(32'hbbece68e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ee18f),
	.w1(32'hbc00f659),
	.w2(32'h3bacda9f),
	.w3(32'hbb88ca67),
	.w4(32'hbc14bf4d),
	.w5(32'hbc964c92),
	.w6(32'h39798498),
	.w7(32'hbb813f64),
	.w8(32'hbb2b29be),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc809d),
	.w1(32'hbc8148d5),
	.w2(32'h3ba6c488),
	.w3(32'h3b24df0a),
	.w4(32'hba28279a),
	.w5(32'hbaaae914),
	.w6(32'h3b2fd07c),
	.w7(32'hbb10344f),
	.w8(32'h3bc5de14),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c51e4),
	.w1(32'hbbadd284),
	.w2(32'hbbf1125f),
	.w3(32'h3a9ff59a),
	.w4(32'h3c442d78),
	.w5(32'h3c185e33),
	.w6(32'h3bf35655),
	.w7(32'hbb557366),
	.w8(32'h3aa4c06a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2e385),
	.w1(32'hbb3f7fa0),
	.w2(32'h3ba4c0d0),
	.w3(32'hbbc78a00),
	.w4(32'hb9e0a386),
	.w5(32'hbc5561cd),
	.w6(32'h38df5197),
	.w7(32'hbb52e9d2),
	.w8(32'hbb0c30e2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2adee),
	.w1(32'h3acd05f7),
	.w2(32'h3b827610),
	.w3(32'hbc65be8d),
	.w4(32'h38e7fd78),
	.w5(32'h3b82c004),
	.w6(32'h3b5329b8),
	.w7(32'h398b2b08),
	.w8(32'hbc12ddac),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f51af),
	.w1(32'hbc18b98b),
	.w2(32'h3c0ade4b),
	.w3(32'h3bec72d4),
	.w4(32'h3bcdefd5),
	.w5(32'hbbb4319e),
	.w6(32'h3b813f81),
	.w7(32'hbb819ff7),
	.w8(32'hbb1c9225),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42dbc9),
	.w1(32'h3b53fcf1),
	.w2(32'hbbde5969),
	.w3(32'h3bf69f23),
	.w4(32'hbbfb222d),
	.w5(32'hbc209ec6),
	.w6(32'h3b06e6ed),
	.w7(32'hbb3e937e),
	.w8(32'hbc3d69d6),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40d3a2),
	.w1(32'hbacc3730),
	.w2(32'hbb7710b8),
	.w3(32'h3bce18ff),
	.w4(32'hb8ba1420),
	.w5(32'hbc699601),
	.w6(32'h3c257fc8),
	.w7(32'hbcf79a04),
	.w8(32'h3ba18a9c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d2439),
	.w1(32'hb915c101),
	.w2(32'hbb1246d3),
	.w3(32'h3ba957df),
	.w4(32'h3c833828),
	.w5(32'hbc2c7eb9),
	.w6(32'h3b0aaee9),
	.w7(32'hbaf965a9),
	.w8(32'h3afcbb2d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e77dd4),
	.w1(32'hbc498412),
	.w2(32'hbc429ffd),
	.w3(32'hba710e50),
	.w4(32'h3c2840fd),
	.w5(32'hbc7c2d09),
	.w6(32'hbae39a89),
	.w7(32'h3b86c6ca),
	.w8(32'h3bbc2f37),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddcda5),
	.w1(32'hbbf88459),
	.w2(32'h3bbf612e),
	.w3(32'h3cb06a74),
	.w4(32'hbc6be494),
	.w5(32'h3b95c727),
	.w6(32'h3b93bead),
	.w7(32'hbbe979be),
	.w8(32'h3c2aea8e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e73c4),
	.w1(32'h3ba3b0a4),
	.w2(32'hbbd89b12),
	.w3(32'hbb739eb0),
	.w4(32'hbb7b20af),
	.w5(32'hbb22fdf0),
	.w6(32'hbbc872a4),
	.w7(32'h3c47f910),
	.w8(32'hbbfad74c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb697b12),
	.w1(32'h3c48b73e),
	.w2(32'h3bb6051e),
	.w3(32'hbc9eabb0),
	.w4(32'h3d4d4876),
	.w5(32'h3baca439),
	.w6(32'h3d101b2f),
	.w7(32'h3c1e2063),
	.w8(32'h3a83c004),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3185de),
	.w1(32'h3b5393ff),
	.w2(32'h3b93a8d9),
	.w3(32'hbc8d21f7),
	.w4(32'hba7058b7),
	.w5(32'hbba7f5a4),
	.w6(32'h3bae926a),
	.w7(32'hbb9b84be),
	.w8(32'h3a26c4d4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09e32f),
	.w1(32'h3b7f3739),
	.w2(32'h3b991ea6),
	.w3(32'h3a1648a5),
	.w4(32'hbc9a1cac),
	.w5(32'h39e52dbd),
	.w6(32'hbae758f2),
	.w7(32'hbc88f5bc),
	.w8(32'h3b1dd2ef),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64947),
	.w1(32'h3ba159d2),
	.w2(32'h3c1e6101),
	.w3(32'hbaae2be9),
	.w4(32'h3c4ddb94),
	.w5(32'h3b9120d6),
	.w6(32'h3c144303),
	.w7(32'hbc030bb7),
	.w8(32'hbb8043a7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49c947),
	.w1(32'hbbc3d35d),
	.w2(32'h3b88f582),
	.w3(32'h3b4eb8ff),
	.w4(32'h3c47f0f7),
	.w5(32'hbca77913),
	.w6(32'hbd489422),
	.w7(32'hbbba9a13),
	.w8(32'hbc590758),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bd59f),
	.w1(32'hbaa6aa75),
	.w2(32'hbb3bf9cb),
	.w3(32'hbbc1f400),
	.w4(32'h3c19f011),
	.w5(32'hbbb7a455),
	.w6(32'h3c292675),
	.w7(32'h3be908ac),
	.w8(32'h3c470ac4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a702),
	.w1(32'h3ce1a83b),
	.w2(32'hbc676972),
	.w3(32'hbb590493),
	.w4(32'hbbaf325d),
	.w5(32'hbc0cb19d),
	.w6(32'hbbbff033),
	.w7(32'hbc3fed77),
	.w8(32'h3a2bb724),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c191da3),
	.w1(32'hbb6de56f),
	.w2(32'hbaf0f7f7),
	.w3(32'hbbd2d99b),
	.w4(32'h3b549ac6),
	.w5(32'h3b4e6be7),
	.w6(32'h3c0f9c47),
	.w7(32'h3bbb808b),
	.w8(32'hbb3c49fe),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b4265),
	.w1(32'h3b807f6c),
	.w2(32'hbb10223e),
	.w3(32'hbbdd0ac0),
	.w4(32'h3b57bfbb),
	.w5(32'h3b8ed5e6),
	.w6(32'h3a22e605),
	.w7(32'h3c143b8a),
	.w8(32'hbaf60e0a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfca9b4),
	.w1(32'hb854b7a3),
	.w2(32'h3c8f9070),
	.w3(32'hbbb692f9),
	.w4(32'h3b139003),
	.w5(32'h3c5fe66d),
	.w6(32'h3a4e0cf3),
	.w7(32'hbbb693e2),
	.w8(32'hbbc5676d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800296),
	.w1(32'hbb2a73fe),
	.w2(32'hbb8a153c),
	.w3(32'h3c339349),
	.w4(32'hbb932a5c),
	.w5(32'hbbbaa985),
	.w6(32'h3b2986ba),
	.w7(32'h3b35fd5e),
	.w8(32'h3ad078e5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccc77d),
	.w1(32'h3b81af75),
	.w2(32'hbbaa5460),
	.w3(32'hbcaae605),
	.w4(32'h3b044620),
	.w5(32'hbb8ecf16),
	.w6(32'hbc069ce3),
	.w7(32'hbaa000ca),
	.w8(32'hbc126ed3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c6b11),
	.w1(32'hbbeac7b1),
	.w2(32'h3c314ae7),
	.w3(32'hbaeac02e),
	.w4(32'hbc3b9847),
	.w5(32'h3b025425),
	.w6(32'hbd43ca6b),
	.w7(32'hba03cc8d),
	.w8(32'hbb0726ea),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c98ea),
	.w1(32'hb989097e),
	.w2(32'h3c29c2f1),
	.w3(32'hbb4c9e8e),
	.w4(32'h3bc4d2c4),
	.w5(32'hbb8c1176),
	.w6(32'hbc004ca1),
	.w7(32'hbbfdbb63),
	.w8(32'h3b574df1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51ee47),
	.w1(32'h3c4ba9d7),
	.w2(32'hbc8b5fd7),
	.w3(32'hbc087a41),
	.w4(32'h3aa96abf),
	.w5(32'h38b60003),
	.w6(32'hba89db05),
	.w7(32'h373ccf71),
	.w8(32'hbca71012),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ade2b1),
	.w1(32'hb961f7f4),
	.w2(32'h3ac25d95),
	.w3(32'hba51e20d),
	.w4(32'h3c455d72),
	.w5(32'h3bb71252),
	.w6(32'hbc6a4473),
	.w7(32'h3c27254d),
	.w8(32'h3b0ef666),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4545b),
	.w1(32'h3c81369d),
	.w2(32'h3ce825c6),
	.w3(32'h3b5866db),
	.w4(32'hbb36163a),
	.w5(32'h3b12070c),
	.w6(32'h3d043d1e),
	.w7(32'hbc6ec725),
	.w8(32'h3babcebb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b58d5),
	.w1(32'hbac279f7),
	.w2(32'h3c3737c1),
	.w3(32'h3b679f67),
	.w4(32'hbc96875e),
	.w5(32'hbb6cff0f),
	.w6(32'h3d187dd4),
	.w7(32'h3a3527cb),
	.w8(32'h3c4f40e0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86bd3f),
	.w1(32'hbadbb798),
	.w2(32'hbb9ccff4),
	.w3(32'hb8d7bd9c),
	.w4(32'hbbb1addc),
	.w5(32'hbb37acbf),
	.w6(32'h3abc21c5),
	.w7(32'h3acda6ba),
	.w8(32'h3c2fb88a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc22c4),
	.w1(32'h3a70a7dd),
	.w2(32'h3919abf9),
	.w3(32'h389d9eea),
	.w4(32'h3ba98f7c),
	.w5(32'h3b8fe1c5),
	.w6(32'hb985ec45),
	.w7(32'h3c08c6ff),
	.w8(32'h3aed9047),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53da3e),
	.w1(32'hbb9659cc),
	.w2(32'hbbaef5cd),
	.w3(32'hbb527a4f),
	.w4(32'h3c2df264),
	.w5(32'hbcb208d2),
	.w6(32'hb897e508),
	.w7(32'h3b0a41f5),
	.w8(32'hbc2d2372),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5b2b1),
	.w1(32'h3ab9f902),
	.w2(32'hb91c101a),
	.w3(32'h3bd6e0e6),
	.w4(32'hbae54783),
	.w5(32'hba037cb4),
	.w6(32'hbc5c5dc9),
	.w7(32'hbc7121d5),
	.w8(32'h3badab37),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05a136),
	.w1(32'hbb949722),
	.w2(32'hbaa385d5),
	.w3(32'h3bf393b1),
	.w4(32'h3be28f10),
	.w5(32'h3b30529c),
	.w6(32'h3cc337c4),
	.w7(32'h3a5fd38d),
	.w8(32'hbc3d393e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8687d9),
	.w1(32'hbc02a41b),
	.w2(32'h3aa7cbd1),
	.w3(32'h3c184e83),
	.w4(32'hbc0dcf60),
	.w5(32'h3a10114d),
	.w6(32'h3c89dc33),
	.w7(32'hbadb9051),
	.w8(32'h3bd23d96),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27034f),
	.w1(32'h3b2a45aa),
	.w2(32'hbbd0acfa),
	.w3(32'h3c66eb04),
	.w4(32'hbc21c0e3),
	.w5(32'hb8aa18a3),
	.w6(32'h3c3026fb),
	.w7(32'h3a6793c2),
	.w8(32'hbb1b8118),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb055c43),
	.w1(32'hbc1ab032),
	.w2(32'hbb971c5d),
	.w3(32'h3b340697),
	.w4(32'hb98c92d8),
	.w5(32'hbb778c81),
	.w6(32'hbb66adc5),
	.w7(32'h396428ec),
	.w8(32'hb993d4c7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6da57),
	.w1(32'hbb955231),
	.w2(32'h3c29bf1f),
	.w3(32'h3ce089d0),
	.w4(32'hbb667f44),
	.w5(32'h3a89a2c1),
	.w6(32'hbbb5c8e9),
	.w7(32'h3c51c4c5),
	.w8(32'hbc60081d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55c0ff),
	.w1(32'hbc985228),
	.w2(32'h3d2e153c),
	.w3(32'hbba546e7),
	.w4(32'hbab0c9d2),
	.w5(32'h3c1b0d27),
	.w6(32'h3b1f6480),
	.w7(32'hbc04e784),
	.w8(32'hbc3810f2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf0ccf),
	.w1(32'hbc0f805b),
	.w2(32'hbcf65131),
	.w3(32'hbcd5c946),
	.w4(32'h3b32f483),
	.w5(32'hba66efdd),
	.w6(32'hbbf88981),
	.w7(32'hbc4c74fd),
	.w8(32'h3bffe9f6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3bc2b),
	.w1(32'hbbe23bb6),
	.w2(32'hbbdfbc3f),
	.w3(32'hbbb02fab),
	.w4(32'h3b0acedc),
	.w5(32'h3c03d1d9),
	.w6(32'hbbd21fe1),
	.w7(32'hb9355286),
	.w8(32'hbbaed53c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe956c),
	.w1(32'h3b20590f),
	.w2(32'hbbdf9b81),
	.w3(32'hbb5bc052),
	.w4(32'hb9440fd5),
	.w5(32'h3bad98a3),
	.w6(32'hbb2b6d0a),
	.w7(32'h3c1449db),
	.w8(32'h3c598c35),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce4c32),
	.w1(32'h3ba65f48),
	.w2(32'hbbed77b6),
	.w3(32'h3a51b7a5),
	.w4(32'h3b3549c1),
	.w5(32'hbabfdb1e),
	.w6(32'h3a4e81b6),
	.w7(32'hbab58c66),
	.w8(32'h3cfdc03f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35da95),
	.w1(32'hbb7e67a8),
	.w2(32'hbce44795),
	.w3(32'hbbbc9608),
	.w4(32'h3c40409d),
	.w5(32'hbb143636),
	.w6(32'h3a40d093),
	.w7(32'h3b42c7d8),
	.w8(32'h3ab8d2a6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65bb0),
	.w1(32'hbc30bb86),
	.w2(32'h3b997ca5),
	.w3(32'h3b844150),
	.w4(32'hbb491d7a),
	.w5(32'hbb0e5f1b),
	.w6(32'hbbb35fae),
	.w7(32'hbbc945bb),
	.w8(32'hbc077626),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315511),
	.w1(32'hbc0e4866),
	.w2(32'h3a455ee0),
	.w3(32'h3c0bcf23),
	.w4(32'h3b819fb2),
	.w5(32'hbbbd0ee2),
	.w6(32'hbb57ec15),
	.w7(32'h39291b1c),
	.w8(32'hbb88071b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ef0c),
	.w1(32'hbb27dd2f),
	.w2(32'h3ba60b18),
	.w3(32'hbc04a0c1),
	.w4(32'hbbe49113),
	.w5(32'h3a01673a),
	.w6(32'h3a8a1300),
	.w7(32'hba61471a),
	.w8(32'hbba8da26),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d39f3),
	.w1(32'hb9b375f7),
	.w2(32'h3ba98828),
	.w3(32'hbba0b3f7),
	.w4(32'h3a67933f),
	.w5(32'h396388a9),
	.w6(32'hbb1a1db7),
	.w7(32'h3c16dfd7),
	.w8(32'hba7bd10d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c651719),
	.w1(32'hbaca6dfd),
	.w2(32'h3b3e171e),
	.w3(32'hba6dc254),
	.w4(32'h3b272012),
	.w5(32'hbb8eace3),
	.w6(32'hbb678907),
	.w7(32'hbb2508cf),
	.w8(32'hb96e3c6d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b170b77),
	.w1(32'h3adcd3d6),
	.w2(32'h3b2e6105),
	.w3(32'hb98673df),
	.w4(32'hbbe21dbf),
	.w5(32'h3bac5eef),
	.w6(32'h3a495f42),
	.w7(32'hbb35df91),
	.w8(32'hbc7b802b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06e8b9),
	.w1(32'hbb447430),
	.w2(32'hbba2c5d6),
	.w3(32'hbb8b4125),
	.w4(32'hba244e00),
	.w5(32'h3ba58763),
	.w6(32'h3b6a6d88),
	.w7(32'hbbf2e383),
	.w8(32'hb9bff69a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c11eb),
	.w1(32'h3b6c07e9),
	.w2(32'h3bb72e38),
	.w3(32'h3b064f13),
	.w4(32'h3b29b65a),
	.w5(32'h3bf4efba),
	.w6(32'h3c0f1b7c),
	.w7(32'h3a12b2dd),
	.w8(32'h3c8bcfbd),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f17251),
	.w1(32'h3bd4b6f3),
	.w2(32'hbc0a7be8),
	.w3(32'hbb4bedb5),
	.w4(32'hbb90afc4),
	.w5(32'h3ae2b93d),
	.w6(32'h3bcdf2b3),
	.w7(32'h3bcd509c),
	.w8(32'h3b7b1cea),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31d2a8),
	.w1(32'h3adb9820),
	.w2(32'h39d83763),
	.w3(32'h3a4249be),
	.w4(32'h3cf86124),
	.w5(32'h3b4b4b1c),
	.w6(32'hbba864df),
	.w7(32'hbba7386d),
	.w8(32'h3a7fcb60),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8324bc),
	.w1(32'h3c4d7f2b),
	.w2(32'hbc2c7cc9),
	.w3(32'hba5da682),
	.w4(32'hba968866),
	.w5(32'h3b09e5a6),
	.w6(32'hb6320f3f),
	.w7(32'hbad1d6a8),
	.w8(32'h3b67721e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37cc7b),
	.w1(32'h3a48033f),
	.w2(32'h3c82eaea),
	.w3(32'h3b41a2d6),
	.w4(32'h397c9e6d),
	.w5(32'hbb9ac1f8),
	.w6(32'hb98ca861),
	.w7(32'hbc3f56fa),
	.w8(32'h3c81e00a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84862b),
	.w1(32'h3b378567),
	.w2(32'hbc662369),
	.w3(32'hbc276e8d),
	.w4(32'h3a9dccfe),
	.w5(32'hbb186aab),
	.w6(32'hbb772a30),
	.w7(32'hbb908f75),
	.w8(32'hbafbf5b8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafbc60),
	.w1(32'h37d69ca4),
	.w2(32'hbb8d6dab),
	.w3(32'h3b7c67a1),
	.w4(32'h397789d8),
	.w5(32'hbc4b228f),
	.w6(32'h390a3c81),
	.w7(32'hbb486253),
	.w8(32'hba96836b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36b4d4),
	.w1(32'hbb1e0c37),
	.w2(32'hb9be9e0a),
	.w3(32'h3b7e10f7),
	.w4(32'hba28ff63),
	.w5(32'h3b1c473b),
	.w6(32'hbbac4771),
	.w7(32'h3d263418),
	.w8(32'hbb912057),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9dcfb),
	.w1(32'hbb14aa42),
	.w2(32'hbb265d6b),
	.w3(32'hb9526f22),
	.w4(32'h3b7eca83),
	.w5(32'hba7e3f5b),
	.w6(32'h3b6edafa),
	.w7(32'hbb8a01ad),
	.w8(32'hbb771652),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca06246),
	.w1(32'hbbeec904),
	.w2(32'h3c1fe57f),
	.w3(32'h3bce767c),
	.w4(32'h39e9ac20),
	.w5(32'h3aa18d86),
	.w6(32'h3cb0c888),
	.w7(32'h3a745cec),
	.w8(32'hbbfda177),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc231df9),
	.w1(32'hbc011c37),
	.w2(32'hbbe22391),
	.w3(32'h3b85b1b6),
	.w4(32'hbcce1b89),
	.w5(32'hb8a171fb),
	.w6(32'hbaafe56e),
	.w7(32'h3b1c98ff),
	.w8(32'h3983c119),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1027),
	.w1(32'h390cabd2),
	.w2(32'h3bcec682),
	.w3(32'hbc7ef215),
	.w4(32'h3afff1a8),
	.w5(32'hbb1f69bc),
	.w6(32'hbaa5881b),
	.w7(32'h3bc7429b),
	.w8(32'hbc864a75),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5ac33),
	.w1(32'hbcc724d6),
	.w2(32'h3b699ca9),
	.w3(32'hbb3817a9),
	.w4(32'hbb7a9d48),
	.w5(32'hb9b4f4c2),
	.w6(32'hbbcece70),
	.w7(32'h3b9e65c3),
	.w8(32'hbc1d9b8a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5ce3),
	.w1(32'hb9fa4cbb),
	.w2(32'h3aec03e0),
	.w3(32'h3a7a4d1d),
	.w4(32'hbb3a82b3),
	.w5(32'h3b8f363a),
	.w6(32'h38be4b73),
	.w7(32'hbb0f68aa),
	.w8(32'h3b052710),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f98a8),
	.w1(32'h3d0b62af),
	.w2(32'hbbedf782),
	.w3(32'hbb33b4b4),
	.w4(32'hb966f02f),
	.w5(32'hba4c8ec5),
	.w6(32'hbba41b74),
	.w7(32'h3c6d9f2d),
	.w8(32'hba1a7f8d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a092),
	.w1(32'hbbf23cc2),
	.w2(32'h39245d7a),
	.w3(32'h3b3e6bbc),
	.w4(32'hbb55e9fb),
	.w5(32'hbb873428),
	.w6(32'hbc985f7d),
	.w7(32'h3a0ed460),
	.w8(32'hbb56caaa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe32def),
	.w1(32'h3c31d205),
	.w2(32'h3b5482cd),
	.w3(32'h3cf79a78),
	.w4(32'h37e1b731),
	.w5(32'hbba6e8bd),
	.w6(32'h3c1cb4e0),
	.w7(32'h3c990475),
	.w8(32'h3940ae39),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf84897),
	.w1(32'h3bcb3dde),
	.w2(32'hbb854959),
	.w3(32'hbb514409),
	.w4(32'hba8b81d7),
	.w5(32'hbb26f009),
	.w6(32'h385b9e95),
	.w7(32'h3b533d7d),
	.w8(32'h3b3fe71e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11e6fc),
	.w1(32'h3b8cb19d),
	.w2(32'hbb981316),
	.w3(32'h3b04c196),
	.w4(32'hb78fed5a),
	.w5(32'hbcdb4e3d),
	.w6(32'h3afdfa34),
	.w7(32'h3b8616b2),
	.w8(32'h3af4296c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e8d63),
	.w1(32'hbbb7e543),
	.w2(32'h3cdd689d),
	.w3(32'h3bbc3fc6),
	.w4(32'hbbb296f6),
	.w5(32'hbc0fe068),
	.w6(32'hbc078441),
	.w7(32'hbb5d9d0a),
	.w8(32'hba353839),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb1104),
	.w1(32'hbb507f0f),
	.w2(32'h3bdaf3eb),
	.w3(32'hbc32ce55),
	.w4(32'h3c07b33e),
	.w5(32'h3c3a7e11),
	.w6(32'hbb5c9df6),
	.w7(32'h3c1078b8),
	.w8(32'hbcabfecb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b84f9),
	.w1(32'h3c82560e),
	.w2(32'h3be87593),
	.w3(32'hbb9b1e8a),
	.w4(32'h3bd13f7b),
	.w5(32'hbbbfc57b),
	.w6(32'hba74d109),
	.w7(32'hbd003855),
	.w8(32'h3abbe52f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c431c),
	.w1(32'h3b72c746),
	.w2(32'h3c3caec8),
	.w3(32'h3c53c004),
	.w4(32'h3b62dfd5),
	.w5(32'hbca5c446),
	.w6(32'hbaded7da),
	.w7(32'h3b538f13),
	.w8(32'h3c09c804),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c0915),
	.w1(32'h3cc763d4),
	.w2(32'h3c622ff8),
	.w3(32'h3cffb8e8),
	.w4(32'hbb22ac54),
	.w5(32'hbb95a378),
	.w6(32'hbc21c119),
	.w7(32'hbc6aa48d),
	.w8(32'h3ad9a2fa),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6308fd),
	.w1(32'hbc59ab4f),
	.w2(32'hbbff645b),
	.w3(32'h3c78a15b),
	.w4(32'h3c49e4d7),
	.w5(32'hbc03e362),
	.w6(32'h3be2d4c5),
	.w7(32'h3817b63d),
	.w8(32'hbb4f6ff2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb3256),
	.w1(32'hbc947024),
	.w2(32'hbca59af1),
	.w3(32'h3bb8ceda),
	.w4(32'hbb17f9b5),
	.w5(32'hb8402689),
	.w6(32'h3b804d5f),
	.w7(32'hbb6a1b7e),
	.w8(32'hbda301c3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf23a76),
	.w1(32'h3bfce006),
	.w2(32'h3c927e37),
	.w3(32'hbbbf2d38),
	.w4(32'h3d9ae761),
	.w5(32'h3c889b81),
	.w6(32'h3b102a06),
	.w7(32'hbb031c4b),
	.w8(32'hbc2ae5a7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b4a6b),
	.w1(32'hbd0395fa),
	.w2(32'h3c39227a),
	.w3(32'h3b5a9d1a),
	.w4(32'h3c1d1e42),
	.w5(32'h3c0d32f7),
	.w6(32'hba915ed9),
	.w7(32'hbb46386b),
	.w8(32'h3b9e7222),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22e18b),
	.w1(32'h3bf3f5cf),
	.w2(32'hbb9e5094),
	.w3(32'hbb2369ca),
	.w4(32'hba3c3764),
	.w5(32'h3bad070b),
	.w6(32'h3cb3a250),
	.w7(32'h3d0b68f1),
	.w8(32'hbc2aac73),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54e29f),
	.w1(32'hbb2df28e),
	.w2(32'hbbec1faf),
	.w3(32'h3c30e632),
	.w4(32'hba1b61f5),
	.w5(32'h3d628f25),
	.w6(32'hbc21dfd2),
	.w7(32'h3bd2fba6),
	.w8(32'hbbdad5db),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74b63c),
	.w1(32'hbc4de4cf),
	.w2(32'hbad98bf8),
	.w3(32'hbbef1b2f),
	.w4(32'hbaab052d),
	.w5(32'h3c17e728),
	.w6(32'hbc1b76dc),
	.w7(32'h3c72e64c),
	.w8(32'hbbe7ef0e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced7b03),
	.w1(32'hbc173af1),
	.w2(32'hb5eeeb2f),
	.w3(32'hba9a6172),
	.w4(32'h3c8d0798),
	.w5(32'hbbf5e554),
	.w6(32'hbbc98254),
	.w7(32'h3b9c0cb6),
	.w8(32'hbab1f876),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6109db),
	.w1(32'hbb951d4d),
	.w2(32'h3b137f45),
	.w3(32'h3cc92c4c),
	.w4(32'h3bec505f),
	.w5(32'hbc22ec01),
	.w6(32'hbb993337),
	.w7(32'hbb78d26f),
	.w8(32'hbab404e2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f1090),
	.w1(32'h3b36af38),
	.w2(32'hbb64fd8d),
	.w3(32'hbbdb10d5),
	.w4(32'h3bb1c2bd),
	.w5(32'h3c14af05),
	.w6(32'h399a6d54),
	.w7(32'h3bc12dd0),
	.w8(32'hbbd6b11c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc725bd),
	.w1(32'hbd0c9605),
	.w2(32'hbc8b53e2),
	.w3(32'hba9cae85),
	.w4(32'h3b9b4f42),
	.w5(32'hbc52ad1b),
	.w6(32'h3b1e23a2),
	.w7(32'h3bacd2e2),
	.w8(32'hbc274e1f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd725da),
	.w1(32'hbaa5537e),
	.w2(32'h3b13a16e),
	.w3(32'hbbe3aeb9),
	.w4(32'hbbea8d6c),
	.w5(32'hbc2f566f),
	.w6(32'hbc2e237e),
	.w7(32'hbc20887a),
	.w8(32'h3bd593a8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6b3ff),
	.w1(32'h3bc50085),
	.w2(32'h3b41658b),
	.w3(32'hbc4083dd),
	.w4(32'hbc4aa1f9),
	.w5(32'hbc0248ba),
	.w6(32'hbbfebde3),
	.w7(32'h38b1dc69),
	.w8(32'h3bc22b2c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9a31d),
	.w1(32'hbc2c81f7),
	.w2(32'h3bcce61c),
	.w3(32'hbd2e5a10),
	.w4(32'hba0559ef),
	.w5(32'hbc2ba64c),
	.w6(32'h3afb4341),
	.w7(32'hbcde5a16),
	.w8(32'hbb000d22),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb734030),
	.w1(32'hbb4d8467),
	.w2(32'hbc50f477),
	.w3(32'hbc13348e),
	.w4(32'hbc04df37),
	.w5(32'h3be7a9ec),
	.w6(32'hbc87c86c),
	.w7(32'h3b444c79),
	.w8(32'hbb65e630),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41e8eb),
	.w1(32'hbc43f3e3),
	.w2(32'hbc90218a),
	.w3(32'hbab4e7ca),
	.w4(32'h3b412634),
	.w5(32'hba84fad3),
	.w6(32'h3b5f512e),
	.w7(32'h3acd602d),
	.w8(32'h3a931af4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1792f0),
	.w1(32'h3bf84ab2),
	.w2(32'h39f3cfe8),
	.w3(32'hbbf82cd0),
	.w4(32'hba96a941),
	.w5(32'h3be640ce),
	.w6(32'h3cadf11e),
	.w7(32'hbc3657ae),
	.w8(32'h3ced6524),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fff5e),
	.w1(32'h3bf7b237),
	.w2(32'h395d880b),
	.w3(32'hbc13c978),
	.w4(32'h3bd6c4d7),
	.w5(32'h3bdacc62),
	.w6(32'h3be7a64a),
	.w7(32'h3b947b0e),
	.w8(32'hbc43d8a5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7aec62),
	.w1(32'h3b0da74b),
	.w2(32'hbc861971),
	.w3(32'hbcac622d),
	.w4(32'h374c9644),
	.w5(32'hbb5b50eb),
	.w6(32'hb946dbb1),
	.w7(32'hbb69af87),
	.w8(32'h3b9652b5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e037f),
	.w1(32'hbbebd0bd),
	.w2(32'hba9b808f),
	.w3(32'hbb006498),
	.w4(32'hbd2b7750),
	.w5(32'h3b05dc84),
	.w6(32'hbbb6061d),
	.w7(32'hbc0c5368),
	.w8(32'hbbfe5fbe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba309bc3),
	.w1(32'h3c81d066),
	.w2(32'h3c2fa150),
	.w3(32'hbbddce8b),
	.w4(32'hba9bbd8f),
	.w5(32'hbbf63ad1),
	.w6(32'hbc813c60),
	.w7(32'hbc849fff),
	.w8(32'hbc1cecdf),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ef00),
	.w1(32'hba35a838),
	.w2(32'hbb99a535),
	.w3(32'h3c53a039),
	.w4(32'hbd7e614a),
	.w5(32'h3cb4ac66),
	.w6(32'h3c8538a9),
	.w7(32'h3c1a9401),
	.w8(32'h3c29d318),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb1db9),
	.w1(32'hbc99c78d),
	.w2(32'hba26815f),
	.w3(32'hbda33cc0),
	.w4(32'h3b1470dd),
	.w5(32'hbc00464c),
	.w6(32'h3a342709),
	.w7(32'h3c125314),
	.w8(32'h3a9fd23c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb456ea9),
	.w1(32'h3c3ad355),
	.w2(32'h3c64a420),
	.w3(32'h3c39ebfd),
	.w4(32'h3af0cf49),
	.w5(32'h3c1dcff0),
	.w6(32'h3a2e0436),
	.w7(32'hbbda74a5),
	.w8(32'hbc2f4bf7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870e80),
	.w1(32'hbc138979),
	.w2(32'h3b5bd3e5),
	.w3(32'h3bb331da),
	.w4(32'hbbfcdd61),
	.w5(32'hbbf53d62),
	.w6(32'h3c01d821),
	.w7(32'h3c43a2af),
	.w8(32'h3b9d9ec6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba2be9),
	.w1(32'h3c594961),
	.w2(32'h3c58f052),
	.w3(32'h3b8cf346),
	.w4(32'h3b76ed50),
	.w5(32'hbcab1a0a),
	.w6(32'hbc847a4a),
	.w7(32'h3c347cc7),
	.w8(32'hbc0463a7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03492e),
	.w1(32'h3cfc1af6),
	.w2(32'h3c129043),
	.w3(32'hb9db867e),
	.w4(32'h3ab23a82),
	.w5(32'hbb741ce4),
	.w6(32'h3be6db01),
	.w7(32'hbc7f56a8),
	.w8(32'h3c0bc125),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1d265),
	.w1(32'hba4150c0),
	.w2(32'h3cb204ca),
	.w3(32'h3c86db37),
	.w4(32'h3b1ca03e),
	.w5(32'hbbfd0696),
	.w6(32'h3b6e64af),
	.w7(32'hbc6c47ef),
	.w8(32'h3c362d91),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15f29d),
	.w1(32'hbc0e0e1c),
	.w2(32'hbbd42e0a),
	.w3(32'hbbfd7a15),
	.w4(32'h3c94d7a1),
	.w5(32'h3cbfec11),
	.w6(32'hbb6754d3),
	.w7(32'hbb25b033),
	.w8(32'hbb960799),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5627b),
	.w1(32'h3b0e47ef),
	.w2(32'h3d11ac92),
	.w3(32'h3cd0e1b2),
	.w4(32'h39cb0aee),
	.w5(32'hbc190a6a),
	.w6(32'h3c997f08),
	.w7(32'hba7f1944),
	.w8(32'h39cc7429),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6a334),
	.w1(32'h3bd2545b),
	.w2(32'h39b84783),
	.w3(32'h3c203e93),
	.w4(32'h3c9dc545),
	.w5(32'hbbc57554),
	.w6(32'h3caced87),
	.w7(32'hb5b5650c),
	.w8(32'hbc7a05ac),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf68213),
	.w1(32'h3b1591aa),
	.w2(32'h3bfb6202),
	.w3(32'hbb22fd03),
	.w4(32'h3b34297b),
	.w5(32'hbc9965fd),
	.w6(32'h3cbc79ce),
	.w7(32'hb9f88cb8),
	.w8(32'h3b76c17b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44a41a),
	.w1(32'h3bd3e745),
	.w2(32'h3b75aac4),
	.w3(32'hbbce816a),
	.w4(32'hbcac383e),
	.w5(32'h388d2181),
	.w6(32'hbbdbd819),
	.w7(32'hbbbaba2e),
	.w8(32'hbc0a2850),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc761126),
	.w1(32'h3c60bc4a),
	.w2(32'h3a1f8f01),
	.w3(32'hba2211e7),
	.w4(32'h3b0dd08e),
	.w5(32'h3b8757c0),
	.w6(32'hbc311682),
	.w7(32'h3be815fa),
	.w8(32'hb899dc22),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c3d3a),
	.w1(32'h3c013704),
	.w2(32'h3c97e251),
	.w3(32'hb92f5ff5),
	.w4(32'hbbb289ff),
	.w5(32'hbbca2773),
	.w6(32'hbca867f3),
	.w7(32'hbc2a5b2d),
	.w8(32'hbba979bf),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d555),
	.w1(32'hba199325),
	.w2(32'hbc331cd5),
	.w3(32'h3c1fba27),
	.w4(32'hbc2aa2d0),
	.w5(32'h3c30c3d8),
	.w6(32'h3bfc072f),
	.w7(32'hba8b1a52),
	.w8(32'h3b0e9318),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc106ee4),
	.w1(32'h3b3b8361),
	.w2(32'h3c14a1ad),
	.w3(32'h3928dd65),
	.w4(32'hbca7f632),
	.w5(32'h3c99772c),
	.w6(32'h3ba8dc7b),
	.w7(32'hbb1d1e14),
	.w8(32'h3af62197),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad55519),
	.w1(32'hbc6cd593),
	.w2(32'hbbd3b417),
	.w3(32'hbabf4ac1),
	.w4(32'h3b97adb1),
	.w5(32'h3a5d6bf0),
	.w6(32'h3c5de0b4),
	.w7(32'hb93a05fa),
	.w8(32'h3c3d30a3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b8999),
	.w1(32'h3b0484f1),
	.w2(32'hbb59ce3b),
	.w3(32'hb7999efe),
	.w4(32'hbc0f5f39),
	.w5(32'h3a152921),
	.w6(32'hbc78a706),
	.w7(32'h3c76cbe5),
	.w8(32'h3ce9135d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a3d56),
	.w1(32'h3bd75790),
	.w2(32'h3b47f67d),
	.w3(32'h3c2344c6),
	.w4(32'h3b1dbada),
	.w5(32'hbbd4ac02),
	.w6(32'h3c10eb4c),
	.w7(32'hbc4e1c4b),
	.w8(32'h3c6b11f1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d0c1),
	.w1(32'hbbb142a7),
	.w2(32'h3c89556f),
	.w3(32'h3cb44b1c),
	.w4(32'h3b456801),
	.w5(32'h3c1631ff),
	.w6(32'hba6e15e4),
	.w7(32'h3b1eb400),
	.w8(32'hbbf78b06),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b46975),
	.w1(32'hbc39d585),
	.w2(32'h3bebf3b7),
	.w3(32'h3b3d499a),
	.w4(32'hbc1420ff),
	.w5(32'hbc39b571),
	.w6(32'h3ace0aac),
	.w7(32'h3b3f9c6d),
	.w8(32'hbb1e6a02),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69750f),
	.w1(32'h3a5ea1fb),
	.w2(32'h3d07632a),
	.w3(32'h3b34c16e),
	.w4(32'h3b909e25),
	.w5(32'h3b8c7cd8),
	.w6(32'h3bb80018),
	.w7(32'h3c0da550),
	.w8(32'h3aeb8e67),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc248f90),
	.w1(32'h3c1a0ae9),
	.w2(32'hb9b685c4),
	.w3(32'hbc47fd64),
	.w4(32'h3d00f6c7),
	.w5(32'h3b756c45),
	.w6(32'hba908b86),
	.w7(32'hbac045c8),
	.w8(32'hbb960df9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc6be3),
	.w1(32'h3d2d90dc),
	.w2(32'hbc8743b3),
	.w3(32'h3b3941f3),
	.w4(32'hbaba5043),
	.w5(32'hbbe71cda),
	.w6(32'h3abd4c56),
	.w7(32'hba88614d),
	.w8(32'h3c0d44a9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3b15),
	.w1(32'hbc8606c8),
	.w2(32'hb8a5ec6b),
	.w3(32'hbc55a637),
	.w4(32'hbba10884),
	.w5(32'h3aebe246),
	.w6(32'h3b4e2d04),
	.w7(32'hbb14002a),
	.w8(32'hbbdb1ae1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f5d40),
	.w1(32'h3c0ec0aa),
	.w2(32'h3bf5aafb),
	.w3(32'h398e5b75),
	.w4(32'hbbc40f25),
	.w5(32'h3b3fab40),
	.w6(32'h3ca2313d),
	.w7(32'h3cd6be8b),
	.w8(32'hb951e77c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a32ee),
	.w1(32'h3b381d91),
	.w2(32'hbbf44e0e),
	.w3(32'hbaae43bd),
	.w4(32'h3ad54160),
	.w5(32'h3ae9cb7b),
	.w6(32'hbbd110ef),
	.w7(32'hbb83e6e4),
	.w8(32'h3c39d625),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d5680),
	.w1(32'h3c9d6ba4),
	.w2(32'hbb436318),
	.w3(32'h3c9e8746),
	.w4(32'h3b09e7b2),
	.w5(32'h3b2077af),
	.w6(32'hbbc83fe4),
	.w7(32'h3c03991b),
	.w8(32'h3bf68c46),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdec71d),
	.w1(32'hbbde3794),
	.w2(32'hbbf38710),
	.w3(32'h3bf21b0b),
	.w4(32'hbbfe07da),
	.w5(32'h3b78a187),
	.w6(32'h3c02a2f5),
	.w7(32'hbc18e5ef),
	.w8(32'h3c0c55e4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f96db),
	.w1(32'hbb857de3),
	.w2(32'hbbc8de6a),
	.w3(32'h3c8ffd42),
	.w4(32'h3be692bb),
	.w5(32'h3c4f8d98),
	.w6(32'hbbe81780),
	.w7(32'h3c9a7b61),
	.w8(32'hbb9f78f9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc452b61),
	.w1(32'h3a9ecb25),
	.w2(32'hbb49f595),
	.w3(32'hbb8c4afa),
	.w4(32'h3bcff160),
	.w5(32'hbb56009f),
	.w6(32'h3c5a44b9),
	.w7(32'hbc421688),
	.w8(32'hbc1536e1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c265d3e),
	.w1(32'hbb56fed8),
	.w2(32'h3ac20cc9),
	.w3(32'hbb21356c),
	.w4(32'h3a935048),
	.w5(32'hbb90f9b1),
	.w6(32'hbc0f25e3),
	.w7(32'hbc1b0395),
	.w8(32'h3a805b74),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule