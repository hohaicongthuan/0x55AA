module layer_10_featuremap_128(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3178c),
	.w1(32'h39bf19d9),
	.w2(32'hb99b8ef2),
	.w3(32'h38377a58),
	.w4(32'h3a22658d),
	.w5(32'hb806654c),
	.w6(32'hba30a3f8),
	.w7(32'hb9aa7caa),
	.w8(32'hb91c5696),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5057fe),
	.w1(32'hba8e7887),
	.w2(32'hbb09dc7b),
	.w3(32'hbb25b224),
	.w4(32'hb92598f6),
	.w5(32'hbad23d3d),
	.w6(32'hbb09f90d),
	.w7(32'hba676c08),
	.w8(32'hbb1a90ac),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982d1e9),
	.w1(32'hb9a493ea),
	.w2(32'hb9b1effc),
	.w3(32'hb8bac9dd),
	.w4(32'hba20a379),
	.w5(32'hba5d1538),
	.w6(32'hb9a808a4),
	.w7(32'hb98a9e24),
	.w8(32'h39ab5cf7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a8936),
	.w1(32'h3b6e232a),
	.w2(32'h3b718967),
	.w3(32'hba21b1ab),
	.w4(32'h3a0780fc),
	.w5(32'hba74a753),
	.w6(32'h39e2b7ac),
	.w7(32'h39fad428),
	.w8(32'h3a14849f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c11b),
	.w1(32'h39ca14fc),
	.w2(32'h3810ed00),
	.w3(32'hb9a31921),
	.w4(32'h3a6281bc),
	.w5(32'h39edcfc9),
	.w6(32'hba26cfa9),
	.w7(32'hb95a932c),
	.w8(32'hb9e8ff24),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9778f33),
	.w1(32'h3a0b5bfb),
	.w2(32'h3aa3ae36),
	.w3(32'hba064016),
	.w4(32'h39a042c4),
	.w5(32'h3a2abe40),
	.w6(32'h3904db9a),
	.w7(32'h3a127e52),
	.w8(32'h3a5ccb52),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393db9ec),
	.w1(32'hbb453df5),
	.w2(32'hbb681c8c),
	.w3(32'hba24aa01),
	.w4(32'hbb965842),
	.w5(32'hbbb3da10),
	.w6(32'h3a874526),
	.w7(32'hbb0d51a9),
	.w8(32'hbb5a25bd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30bc41),
	.w1(32'hbbd12096),
	.w2(32'hbb55aed7),
	.w3(32'hbc2a44c0),
	.w4(32'hbbe2a94d),
	.w5(32'hbb127412),
	.w6(32'hbbd6d06c),
	.w7(32'hbae5c312),
	.w8(32'hba8e44f3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1082a),
	.w1(32'h3a4ee8e1),
	.w2(32'h3a161797),
	.w3(32'hb8cc4131),
	.w4(32'h39dacc0d),
	.w5(32'h3929856f),
	.w6(32'h37d337c5),
	.w7(32'h398ce507),
	.w8(32'h39989cd2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb597e56),
	.w1(32'hba86d53b),
	.w2(32'hbbdd3d89),
	.w3(32'hbb3627cf),
	.w4(32'hb9fe5085),
	.w5(32'hbb93c192),
	.w6(32'hbb3931b3),
	.w7(32'hbae8c989),
	.w8(32'hbba4403e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998bf6a),
	.w1(32'h3987c59d),
	.w2(32'h3a3fbfca),
	.w3(32'h378d2e43),
	.w4(32'h39128132),
	.w5(32'h392ab6bb),
	.w6(32'h3a0b2d12),
	.w7(32'h3aef2dfc),
	.w8(32'h3adc75f7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5350e),
	.w1(32'h393e273e),
	.w2(32'h3a27eff2),
	.w3(32'hba3aeb4f),
	.w4(32'hba99b5b8),
	.w5(32'hbb4716b5),
	.w6(32'h3a5d1679),
	.w7(32'h3ab913c2),
	.w8(32'hba9b1a8e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8bd6),
	.w1(32'hbaa472a4),
	.w2(32'hbb8e34d4),
	.w3(32'hbb3825e3),
	.w4(32'h38b62ffa),
	.w5(32'hbb13d404),
	.w6(32'hbadfeb65),
	.w7(32'hb92335d2),
	.w8(32'hbb24474f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882a50),
	.w1(32'hbb8dfbbf),
	.w2(32'hbba73327),
	.w3(32'hba2018ab),
	.w4(32'hbb71166a),
	.w5(32'hbb84422c),
	.w6(32'hba9c3707),
	.w7(32'hbae20cc6),
	.w8(32'hbb2156c0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f48ca),
	.w1(32'h3a530682),
	.w2(32'hba17e819),
	.w3(32'hbb17b65f),
	.w4(32'h3ac13095),
	.w5(32'hba283fe4),
	.w6(32'hbab9bc7b),
	.w7(32'h3a80f2e7),
	.w8(32'hbac1281e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad9812),
	.w1(32'hbb45c2e5),
	.w2(32'hbbc3fc3c),
	.w3(32'hbba8779b),
	.w4(32'hba8bd2ff),
	.w5(32'hbb234f5f),
	.w6(32'hbbb9c535),
	.w7(32'hbb21c4dc),
	.w8(32'hbb800a92),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d16d3),
	.w1(32'h39f2e801),
	.w2(32'h3a4a3c81),
	.w3(32'h399c44f2),
	.w4(32'h3a5f4c7e),
	.w5(32'h3a62c755),
	.w6(32'h39a20e37),
	.w7(32'h3a9e3955),
	.w8(32'h3a362ed8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0433e),
	.w1(32'hbb4034cd),
	.w2(32'hbbae9d8e),
	.w3(32'hbb85106c),
	.w4(32'hbb33beaa),
	.w5(32'hbb8724c1),
	.w6(32'hbb83f035),
	.w7(32'h398a61c4),
	.w8(32'hbb27ac52),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b97b6),
	.w1(32'hba4af612),
	.w2(32'hbb298eee),
	.w3(32'hbab1909b),
	.w4(32'hba81898a),
	.w5(32'hbb1db48e),
	.w6(32'hba9c47a5),
	.w7(32'h39abcd70),
	.w8(32'hbac70721),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980ef9c),
	.w1(32'h3a374146),
	.w2(32'h3a06aeb7),
	.w3(32'h37d025d6),
	.w4(32'h399f5830),
	.w5(32'h3822c765),
	.w6(32'h3a10f37e),
	.w7(32'h3a2d260f),
	.w8(32'h3a00702f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f45d00),
	.w1(32'hb960c44e),
	.w2(32'hba18dd1d),
	.w3(32'h390f5075),
	.w4(32'hb915f3b6),
	.w5(32'hb7edcc29),
	.w6(32'hb9868a1b),
	.w7(32'hb9bddb0d),
	.w8(32'hb887cc2b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a810d1b),
	.w1(32'h3b4e5e26),
	.w2(32'h3b4b8911),
	.w3(32'h3a8d4286),
	.w4(32'h3a8d0a1e),
	.w5(32'h38c918b8),
	.w6(32'h3b4bbf48),
	.w7(32'h3b84c58f),
	.w8(32'h3b6413cc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3ed15),
	.w1(32'hbb415cfd),
	.w2(32'hbb8d8faf),
	.w3(32'hbbe70da7),
	.w4(32'hba9897c3),
	.w5(32'hbb8b9af6),
	.w6(32'hbc1c9e98),
	.w7(32'hbb6b6d75),
	.w8(32'hbc0896eb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa29cb1),
	.w1(32'h3794ca6d),
	.w2(32'hbbb1580f),
	.w3(32'hb9bab563),
	.w4(32'h3aaecf9c),
	.w5(32'hbb797294),
	.w6(32'hbb1f1434),
	.w7(32'hb8fd947b),
	.w8(32'hbb770dc2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabec573),
	.w1(32'h3b0941a9),
	.w2(32'hbaf6100d),
	.w3(32'hbb6e7983),
	.w4(32'h3b2ae1c1),
	.w5(32'hbaac6be6),
	.w6(32'hbbcbb014),
	.w7(32'hba9c31d5),
	.w8(32'hbb7738e4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9e647),
	.w1(32'h3a71d356),
	.w2(32'h3aac7a77),
	.w3(32'h39c226f7),
	.w4(32'h3a101ac9),
	.w5(32'h39aa7cbd),
	.w6(32'h3a79a269),
	.w7(32'h3acef1d5),
	.w8(32'h3accbef5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9888cd),
	.w1(32'h3a1385c1),
	.w2(32'h3a0c514e),
	.w3(32'h3ab66141),
	.w4(32'h3995cc26),
	.w5(32'h398bb10e),
	.w6(32'h3a0a6b6b),
	.w7(32'h3a094c08),
	.w8(32'h3a16e35d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ef30),
	.w1(32'hb98b9c3c),
	.w2(32'hbb5125ba),
	.w3(32'h3abc43f2),
	.w4(32'hb9917e58),
	.w5(32'hbb088a32),
	.w6(32'h3ad51bb3),
	.w7(32'h3a65ec63),
	.w8(32'h3a4e41bf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f09c13),
	.w1(32'h3ad0a873),
	.w2(32'hb9a07e1a),
	.w3(32'hba1aec9c),
	.w4(32'h3af747a3),
	.w5(32'hb8532ec1),
	.w6(32'hb87ddaff),
	.w7(32'hb860c48e),
	.w8(32'h391754ee),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517b40),
	.w1(32'h3b5ae8b5),
	.w2(32'hba9eafaa),
	.w3(32'hba6e8eec),
	.w4(32'h3adec12c),
	.w5(32'hbb09823c),
	.w6(32'hba4c9c31),
	.w7(32'hba21acb3),
	.w8(32'hbb5acb46),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fa3c3),
	.w1(32'h390b0105),
	.w2(32'hb853eb73),
	.w3(32'h3a8ec8df),
	.w4(32'h398b8ada),
	.w5(32'h39818f5b),
	.w6(32'hb68e73fe),
	.w7(32'hb7e6a649),
	.w8(32'h3604ee20),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f03552),
	.w1(32'h39a0df94),
	.w2(32'h39c9ca13),
	.w3(32'h39ac209e),
	.w4(32'h3935851a),
	.w5(32'h37214eef),
	.w6(32'h396bdf68),
	.w7(32'h39905a3a),
	.w8(32'h39d0f9ae),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50925a),
	.w1(32'h3aa28738),
	.w2(32'hbada8751),
	.w3(32'hb7eb18d6),
	.w4(32'h3a68ab5c),
	.w5(32'hbb00225a),
	.w6(32'h3abcc6c8),
	.w7(32'h3aca0133),
	.w8(32'hba4d0f76),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcebbb),
	.w1(32'hba021c3e),
	.w2(32'hba8a69df),
	.w3(32'hbad5794f),
	.w4(32'hbabdac88),
	.w5(32'hbafc77f5),
	.w6(32'hb9a83a1d),
	.w7(32'h3a2021d7),
	.w8(32'hba0fa130),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89145c),
	.w1(32'h397d94a6),
	.w2(32'h3a2433fc),
	.w3(32'h38c3c7ee),
	.w4(32'hb9b283b7),
	.w5(32'hb9b6b71f),
	.w6(32'h3980043b),
	.w7(32'h39d5db8e),
	.w8(32'h3a276748),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d17212),
	.w1(32'hbaa79d1f),
	.w2(32'hba80e810),
	.w3(32'hb9bb334b),
	.w4(32'hbaa8f970),
	.w5(32'hbac97635),
	.w6(32'h39d97ec8),
	.w7(32'h3a06c4b8),
	.w8(32'h3a7e07d5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc254ec4),
	.w1(32'hbb645c72),
	.w2(32'hbafad965),
	.w3(32'hbb9e0b38),
	.w4(32'hba01e3a0),
	.w5(32'h3ab84fb3),
	.w6(32'hba9a86ee),
	.w7(32'h3b4d81d0),
	.w8(32'h3a5f9c16),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e867),
	.w1(32'h3b68d1b6),
	.w2(32'hbaaa078e),
	.w3(32'hbaf06e06),
	.w4(32'h3bb080e8),
	.w5(32'h39aea9e9),
	.w6(32'hbbacc9b4),
	.w7(32'h39eb25c6),
	.w8(32'hbb65d1dd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e3b3),
	.w1(32'h3b9305ee),
	.w2(32'hbb2e4f00),
	.w3(32'hb9b43fd6),
	.w4(32'h3af5721c),
	.w5(32'hbb8e9723),
	.w6(32'hbb254f35),
	.w7(32'hbab8d60b),
	.w8(32'hbbbc29cb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4602e8),
	.w1(32'h3984108c),
	.w2(32'h39985bd9),
	.w3(32'hba520022),
	.w4(32'h3a2bad1e),
	.w5(32'h39f835e1),
	.w6(32'hbab5eb04),
	.w7(32'h392ce468),
	.w8(32'h3802befe),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392aba5a),
	.w1(32'h3a4dd1e2),
	.w2(32'h3a2497fa),
	.w3(32'hb914cde2),
	.w4(32'h3a9da92f),
	.w5(32'h3a9d96db),
	.w6(32'h3a0b3b69),
	.w7(32'h3a1fe450),
	.w8(32'h39d6733d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd6f7c),
	.w1(32'h395bb025),
	.w2(32'h3a0899a2),
	.w3(32'h3a912223),
	.w4(32'hba02d9d7),
	.w5(32'hba2cdfb4),
	.w6(32'h39e59801),
	.w7(32'h3a1aa346),
	.w8(32'h3a1c8dd8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a9f4),
	.w1(32'h39b59840),
	.w2(32'hb9846afe),
	.w3(32'hba07aad1),
	.w4(32'h3a21b13c),
	.w5(32'hba257ee6),
	.w6(32'h3a1b664f),
	.w7(32'h3a896496),
	.w8(32'hb797d8db),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83bc9),
	.w1(32'hba9445a0),
	.w2(32'hbbf9e38d),
	.w3(32'hbb959a65),
	.w4(32'hb9354ba6),
	.w5(32'hbba2434f),
	.w6(32'hbb999ceb),
	.w7(32'hba58a3b8),
	.w8(32'hbb92ceb8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f20de),
	.w1(32'hba941b43),
	.w2(32'hbbbdece3),
	.w3(32'hb95197a7),
	.w4(32'hba37357d),
	.w5(32'hbba9f533),
	.w6(32'hbb8244d8),
	.w7(32'hbaf2ad9a),
	.w8(32'hbbb2c8aa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba490d5),
	.w1(32'hba7732be),
	.w2(32'hbb8b2a3b),
	.w3(32'hbba79b0e),
	.w4(32'h38f92091),
	.w5(32'hbb5da46a),
	.w6(32'hbb7d9651),
	.w7(32'hb9b98822),
	.w8(32'hbb34b70f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36a947),
	.w1(32'h3a9cff2b),
	.w2(32'hbafbbf9b),
	.w3(32'hbb72fffb),
	.w4(32'h3b6754df),
	.w5(32'hb9cb3f25),
	.w6(32'hbb2e1a10),
	.w7(32'h398e95c1),
	.w8(32'hbb3736bb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb64c3),
	.w1(32'hbb7ac338),
	.w2(32'hbbb558ad),
	.w3(32'hbb6597ba),
	.w4(32'hbb67b7be),
	.w5(32'hbb91dca7),
	.w6(32'hbb9ccf69),
	.w7(32'hba213d18),
	.w8(32'hbb785658),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f3e6cf),
	.w1(32'h39d453f0),
	.w2(32'h39980a0b),
	.w3(32'h3908dd11),
	.w4(32'h3876f144),
	.w5(32'hb96d74a8),
	.w6(32'h39bf0d89),
	.w7(32'h39e6fa01),
	.w8(32'h3a1caa8c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84301ab),
	.w1(32'hba077236),
	.w2(32'hb9b8281a),
	.w3(32'hb93c3132),
	.w4(32'hba1bd4c8),
	.w5(32'hba058a4b),
	.w6(32'hba187a5f),
	.w7(32'hba2ddcea),
	.w8(32'hba2ac1ec),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba010183),
	.w1(32'hbac167d6),
	.w2(32'hbac66d73),
	.w3(32'hba12b596),
	.w4(32'hbad4e772),
	.w5(32'hbade09d5),
	.w6(32'hbac01010),
	.w7(32'hbac54c58),
	.w8(32'hba89d376),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ac4b),
	.w1(32'hb9ee3df4),
	.w2(32'hbb2306b6),
	.w3(32'hbb52ec34),
	.w4(32'hbb1d1b85),
	.w5(32'hbb8d6b42),
	.w6(32'hb9620a5d),
	.w7(32'hba2ff607),
	.w8(32'hbb099564),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b37ec),
	.w1(32'h39e81a3b),
	.w2(32'h3a10ac71),
	.w3(32'hbaeb6925),
	.w4(32'h386144ba),
	.w5(32'hb95dc02b),
	.w6(32'hb97f30a5),
	.w7(32'h3a1fc4b2),
	.w8(32'h395ef084),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55114),
	.w1(32'hbb01b49f),
	.w2(32'hbba2c31f),
	.w3(32'hbb96de8c),
	.w4(32'hbb0e2f5a),
	.w5(32'hbb2d2f6b),
	.w6(32'hbb60891b),
	.w7(32'h39fdb064),
	.w8(32'hbb7319e2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba872633),
	.w1(32'h3816b993),
	.w2(32'hba849133),
	.w3(32'hbab752f6),
	.w4(32'hb95677f3),
	.w5(32'hbac2a684),
	.w6(32'hba032421),
	.w7(32'h3a8b48ed),
	.w8(32'hb98acd45),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d7230),
	.w1(32'h3a176bf5),
	.w2(32'h34be871b),
	.w3(32'h397d9e87),
	.w4(32'h3a6cb00b),
	.w5(32'h38ed067c),
	.w6(32'h387c27c4),
	.w7(32'h39277e62),
	.w8(32'h35e95ff7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b0c69),
	.w1(32'hbac79410),
	.w2(32'hbab7307b),
	.w3(32'h3945c11a),
	.w4(32'hbad3657a),
	.w5(32'hbad9d95f),
	.w6(32'hbac9e46d),
	.w7(32'hbacb5914),
	.w8(32'hba91408b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f797ba),
	.w1(32'h397da977),
	.w2(32'hba34a388),
	.w3(32'hba8e16ee),
	.w4(32'hb9cca0e0),
	.w5(32'hbaa2a7d7),
	.w6(32'h3a4ce7ac),
	.w7(32'hb78cbad5),
	.w8(32'h398e9177),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a371bc1),
	.w1(32'h3a4a1038),
	.w2(32'h39d0e4d9),
	.w3(32'hba646a95),
	.w4(32'h39d381c8),
	.w5(32'hb815b0b6),
	.w6(32'hb916a60c),
	.w7(32'h38f0dcfe),
	.w8(32'hb88484a3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df1440),
	.w1(32'hb872d8e4),
	.w2(32'hb81b2549),
	.w3(32'hb9a18340),
	.w4(32'hb9db2e9b),
	.w5(32'hba16ef47),
	.w6(32'hba138e15),
	.w7(32'hba074b18),
	.w8(32'hb95bfcf9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb312f7d),
	.w1(32'hbadfdf5b),
	.w2(32'hbb1d4916),
	.w3(32'hbaf7ac85),
	.w4(32'hba5e0e9f),
	.w5(32'hbb2088ca),
	.w6(32'hbb005789),
	.w7(32'h3a021d23),
	.w8(32'hba1414d7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e8323),
	.w1(32'hb9cfa2b0),
	.w2(32'hbb2d3028),
	.w3(32'hbb80ce06),
	.w4(32'hb99d1b45),
	.w5(32'hbaf027ca),
	.w6(32'hbb12f075),
	.w7(32'h39c58603),
	.w8(32'hba25494c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe7259),
	.w1(32'h3aabfa61),
	.w2(32'h39fa1e0b),
	.w3(32'hb82c85a7),
	.w4(32'hb8ba4b26),
	.w5(32'hba6698e4),
	.w6(32'h3a8e675b),
	.w7(32'h3ac5c26d),
	.w8(32'h3a8f4b54),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38edb490),
	.w1(32'h399833d8),
	.w2(32'h38e99b81),
	.w3(32'hba7da38f),
	.w4(32'hb4de8f23),
	.w5(32'hb874392c),
	.w6(32'h396be0b1),
	.w7(32'hb9c433ec),
	.w8(32'h3929700e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ff596),
	.w1(32'hb96b7c46),
	.w2(32'hb74ebe0e),
	.w3(32'h3a135500),
	.w4(32'hb9caa451),
	.w5(32'hba6050a7),
	.w6(32'hb92008db),
	.w7(32'h3928ea84),
	.w8(32'h3a3f84df),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a063ada),
	.w1(32'hb9d21c67),
	.w2(32'hba2f67e9),
	.w3(32'hba09bfab),
	.w4(32'hba72a87a),
	.w5(32'hba9c4238),
	.w6(32'h3a38f1ab),
	.w7(32'h38eb8a95),
	.w8(32'h3a231f07),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba190c2),
	.w1(32'hba73835c),
	.w2(32'hbb9365c0),
	.w3(32'hbba78083),
	.w4(32'h39f7c6c8),
	.w5(32'h3a259f9f),
	.w6(32'hbb1ce625),
	.w7(32'h3a9f539e),
	.w8(32'hbaa65827),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa60957),
	.w1(32'h3857ed2e),
	.w2(32'hbb45b04f),
	.w3(32'hba842c93),
	.w4(32'h3a9b5cdc),
	.w5(32'hbb84ba39),
	.w6(32'hbbb07569),
	.w7(32'hba976e4d),
	.w8(32'hbbad4fc3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaff19f),
	.w1(32'h39f47f80),
	.w2(32'hbb6d5d19),
	.w3(32'hbb5ab921),
	.w4(32'h3a8d94b0),
	.w5(32'hbb5150e9),
	.w6(32'hbb8f9484),
	.w7(32'h3a88a293),
	.w8(32'hbb5b7435),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c266d),
	.w1(32'h3aaf4069),
	.w2(32'hbbcd7784),
	.w3(32'hbb17f853),
	.w4(32'h3ab850eb),
	.w5(32'hbb80a790),
	.w6(32'hbbf4c2cb),
	.w7(32'hbb1b6091),
	.w8(32'hbbfd8916),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c9522),
	.w1(32'hb99b2bd8),
	.w2(32'hb8225a5e),
	.w3(32'hbae22c3a),
	.w4(32'hba10036d),
	.w5(32'hba31da2c),
	.w6(32'h380bab35),
	.w7(32'h38f85f16),
	.w8(32'h383d3997),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f538f0),
	.w1(32'hb88f0de5),
	.w2(32'h394a23de),
	.w3(32'hb8e02c95),
	.w4(32'hb91b4d59),
	.w5(32'hb6dd006a),
	.w6(32'hb882102e),
	.w7(32'h3921588d),
	.w8(32'h39d68430),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a040466),
	.w1(32'hb90ca090),
	.w2(32'hb6aa6d65),
	.w3(32'h393ee166),
	.w4(32'hb982af13),
	.w5(32'hb97dfceb),
	.w6(32'hb9c3d0b9),
	.w7(32'hb9a8e9c6),
	.w8(32'h38d8e6a3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad451b),
	.w1(32'h3a778388),
	.w2(32'h39de8a58),
	.w3(32'hba008e56),
	.w4(32'h3a559ef1),
	.w5(32'h38fd0770),
	.w6(32'hb9ae2522),
	.w7(32'h3a696a05),
	.w8(32'h3a0aedba),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d14d0),
	.w1(32'hb889306c),
	.w2(32'hb90ddccf),
	.w3(32'h399e19ff),
	.w4(32'hba18d61b),
	.w5(32'hba3ae3f6),
	.w6(32'h38841a52),
	.w7(32'hb88c8798),
	.w8(32'h38a3fe70),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb752c8c),
	.w1(32'hbaacf3fd),
	.w2(32'h391aa687),
	.w3(32'hbb27dd9f),
	.w4(32'hbb6b58e0),
	.w5(32'hbb110aed),
	.w6(32'h3a2dba3b),
	.w7(32'h3b029753),
	.w8(32'h3a847bb2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee5712),
	.w1(32'hbb7309e1),
	.w2(32'hbb86aef4),
	.w3(32'hbb3f70f2),
	.w4(32'hbb698abd),
	.w5(32'hbb55a3b8),
	.w6(32'hbb9e2615),
	.w7(32'hb8edb371),
	.w8(32'hbb152308),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabafc46),
	.w1(32'hba2ddec2),
	.w2(32'hbb3a0853),
	.w3(32'hbb309571),
	.w4(32'hba0d823f),
	.w5(32'hbae02189),
	.w6(32'hbb2dc884),
	.w7(32'hba249261),
	.w8(32'hbb2d0603),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aac25),
	.w1(32'hb962f04f),
	.w2(32'hbaea7013),
	.w3(32'hbb17a1a3),
	.w4(32'hba4243cb),
	.w5(32'hbb109081),
	.w6(32'hba9a7065),
	.w7(32'h3aa4930f),
	.w8(32'hb9b79beb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22eefb),
	.w1(32'hbaa86463),
	.w2(32'hbb0b9811),
	.w3(32'hba8bcb26),
	.w4(32'hbad11ce9),
	.w5(32'hbaa3a915),
	.w6(32'hba7bccde),
	.w7(32'hba9bd61d),
	.w8(32'hbaa70d9d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75bb0f),
	.w1(32'h3a27237e),
	.w2(32'hbb071b0c),
	.w3(32'hba47e8df),
	.w4(32'h3aa77112),
	.w5(32'hb9d3183c),
	.w6(32'hb9b86e49),
	.w7(32'h3a68bebf),
	.w8(32'hbae125e2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb3277),
	.w1(32'hbaa0f844),
	.w2(32'hbac9c2e8),
	.w3(32'hb9d883ce),
	.w4(32'hbabf11e2),
	.w5(32'hbaf68aac),
	.w6(32'hba82ea84),
	.w7(32'hb9649519),
	.w8(32'hbaa47620),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857af41),
	.w1(32'h3a697453),
	.w2(32'h3a113826),
	.w3(32'hb93796ef),
	.w4(32'h3a33203c),
	.w5(32'h39e8ab35),
	.w6(32'h3a2a9cfd),
	.w7(32'h3a19b0ca),
	.w8(32'h39ea1a51),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aee29c),
	.w1(32'hb9648431),
	.w2(32'hb7aae7b6),
	.w3(32'h3a1503e6),
	.w4(32'hb981b092),
	.w5(32'hb801a594),
	.w6(32'hb890e373),
	.w7(32'h38b5bfc5),
	.w8(32'h38a5ac6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9292ef9),
	.w1(32'hb9f61164),
	.w2(32'h3a462262),
	.w3(32'hb95183dc),
	.w4(32'hba0cd707),
	.w5(32'h39c1349d),
	.w6(32'hb9eedbce),
	.w7(32'h3a63ac4f),
	.w8(32'hb9365345),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a863920),
	.w1(32'h3886ba65),
	.w2(32'h39561265),
	.w3(32'h3963602d),
	.w4(32'hb912f13a),
	.w5(32'hb8de4508),
	.w6(32'hb8f185e0),
	.w7(32'hb918634c),
	.w8(32'hb8bd8788),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158b06),
	.w1(32'hbabb666c),
	.w2(32'hbb4c868a),
	.w3(32'hbb00dc09),
	.w4(32'hb9d2a171),
	.w5(32'hbac7f634),
	.w6(32'hbb678724),
	.w7(32'h35014dd9),
	.w8(32'hbb2bb793),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f316af),
	.w1(32'h3a68fd68),
	.w2(32'h39ba6ec2),
	.w3(32'hba3817e7),
	.w4(32'h3a7b5003),
	.w5(32'h3a319db7),
	.w6(32'hba2c224a),
	.w7(32'h39608f71),
	.w8(32'h37a5f179),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61bcba),
	.w1(32'hba055f95),
	.w2(32'hba81b5e4),
	.w3(32'hba5e9161),
	.w4(32'h3a139148),
	.w5(32'hb9d50094),
	.w6(32'hbad0a745),
	.w7(32'h39557f82),
	.w8(32'hba6430d3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1ebb6),
	.w1(32'hbad8501d),
	.w2(32'hbb600fc2),
	.w3(32'hbb370612),
	.w4(32'hbaae0eea),
	.w5(32'hbb1cd312),
	.w6(32'hbba468cd),
	.w7(32'hba2acb7c),
	.w8(32'hbb342af2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b143e58),
	.w1(32'h3b52aced),
	.w2(32'hb924bb0c),
	.w3(32'h39a369ea),
	.w4(32'h3ab7ba3a),
	.w5(32'hbaa63b5a),
	.w6(32'hb91acfb7),
	.w7(32'h39a1d536),
	.w8(32'hbae3c530),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe310a2),
	.w1(32'hbb971727),
	.w2(32'hbb837671),
	.w3(32'hbb86a0e5),
	.w4(32'hbac00bca),
	.w5(32'hba72094a),
	.w6(32'hbb782084),
	.w7(32'hbb1209e2),
	.w8(32'hbb2cef17),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab153bf),
	.w1(32'h3ae88c03),
	.w2(32'h38fa10a3),
	.w3(32'hb908be4a),
	.w4(32'h39ae73a7),
	.w5(32'hba9c9d64),
	.w6(32'hb9cdd4d5),
	.w7(32'h3a7f6135),
	.w8(32'hb957db0a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3451f),
	.w1(32'hbb75801a),
	.w2(32'hbbe0e774),
	.w3(32'hbb89f8ae),
	.w4(32'hb7e5ac6d),
	.w5(32'hbac9e746),
	.w6(32'hbbbdc34e),
	.w7(32'hbaa56409),
	.w8(32'hbb558125),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea8ad6),
	.w1(32'hba4c69f7),
	.w2(32'hbb28a2e1),
	.w3(32'hbaa2ce76),
	.w4(32'h3a2481a8),
	.w5(32'hba8ec7b9),
	.w6(32'hbac7ef84),
	.w7(32'hb9499a11),
	.w8(32'hbb065694),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c9bba),
	.w1(32'hba5799d5),
	.w2(32'hbad63b32),
	.w3(32'hbaf42819),
	.w4(32'h3a33e88c),
	.w5(32'hb97cc56b),
	.w6(32'hbb333aeb),
	.w7(32'hba434149),
	.w8(32'hbadd1593),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1944b6),
	.w1(32'hb9a7a2a9),
	.w2(32'h3a422f18),
	.w3(32'h3a6501f7),
	.w4(32'hba52ae7a),
	.w5(32'h388b04eb),
	.w6(32'hba0f0523),
	.w7(32'h3a014159),
	.w8(32'h3a15de1e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dd312),
	.w1(32'hba35b8be),
	.w2(32'hbbd81a91),
	.w3(32'hbb0fbdad),
	.w4(32'hb9b16907),
	.w5(32'hbba71047),
	.w6(32'hbb1a5841),
	.w7(32'hbabe607d),
	.w8(32'hbb75bd45),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb027df4),
	.w1(32'hb7cbcbf2),
	.w2(32'hbb0adc79),
	.w3(32'hbaf8bb52),
	.w4(32'hb9f8f8d2),
	.w5(32'hbaec67ba),
	.w6(32'hba7c8ca4),
	.w7(32'h38512e33),
	.w8(32'hbb01615d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d13f8),
	.w1(32'hbbb2a211),
	.w2(32'hba602079),
	.w3(32'hbbcfc8ff),
	.w4(32'hbaf1d8c4),
	.w5(32'h3a8d14d6),
	.w6(32'hbbdad3e1),
	.w7(32'h3aea8a80),
	.w8(32'h3b100d26),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fdd8d),
	.w1(32'h3b40c899),
	.w2(32'hb8404736),
	.w3(32'hbb327253),
	.w4(32'h3bd5b4dc),
	.w5(32'h3b4d4d25),
	.w6(32'hbb297aab),
	.w7(32'h3ba9e657),
	.w8(32'h3b1408f2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5bcc9),
	.w1(32'h3a5d0b60),
	.w2(32'hbb381058),
	.w3(32'hbae975ba),
	.w4(32'h3a76db1c),
	.w5(32'hbb04a5f4),
	.w6(32'hbad4fef9),
	.w7(32'h3878bc29),
	.w8(32'hbb5b9215),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3aedf),
	.w1(32'hbb4eed2c),
	.w2(32'hbb19b8bd),
	.w3(32'hbb3e8064),
	.w4(32'hbacfedd0),
	.w5(32'hba4b763f),
	.w6(32'hba12f657),
	.w7(32'h3aa87cf5),
	.w8(32'h388bf6af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f43e4b),
	.w1(32'hb937848e),
	.w2(32'h3922acd6),
	.w3(32'hb9126027),
	.w4(32'hb89a69a4),
	.w5(32'h3931e8ca),
	.w6(32'hb9d5b92f),
	.w7(32'h379905d3),
	.w8(32'h3a04d5c8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e877e),
	.w1(32'hbbe489c3),
	.w2(32'hbbde0094),
	.w3(32'hbbc4cc90),
	.w4(32'hbb7863e9),
	.w5(32'hbb73f94b),
	.w6(32'hbbb66739),
	.w7(32'h3a644ed1),
	.w8(32'hbab02d1c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba551707),
	.w1(32'hba947f92),
	.w2(32'hbb71a715),
	.w3(32'hbafa6a1f),
	.w4(32'hbb0f0d50),
	.w5(32'hbb96921f),
	.w6(32'h39bec601),
	.w7(32'hba8187de),
	.w8(32'hbb5e34e4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05ca43),
	.w1(32'hb90268b3),
	.w2(32'hb99a7609),
	.w3(32'h395ccf54),
	.w4(32'hb9edf126),
	.w5(32'hba01d6de),
	.w6(32'hb7abc96e),
	.w7(32'hb9172055),
	.w8(32'h393f4c18),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf2111),
	.w1(32'hba8e44ff),
	.w2(32'hbb0490b1),
	.w3(32'hbaed6f59),
	.w4(32'hba0426dc),
	.w5(32'hba34b8ba),
	.w6(32'hbae9c4cd),
	.w7(32'hba718ca9),
	.w8(32'hbad1716a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac628aa),
	.w1(32'hbac495e2),
	.w2(32'hbba1ce1a),
	.w3(32'hba26b397),
	.w4(32'hba9cb0ff),
	.w5(32'hbb77a52d),
	.w6(32'hbb10828f),
	.w7(32'hbb07c58a),
	.w8(32'hbb810092),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b88179),
	.w1(32'hbaa77c43),
	.w2(32'hbb855190),
	.w3(32'hba8c7615),
	.w4(32'hbae9ce10),
	.w5(32'hbb95f9c7),
	.w6(32'hbb5ca669),
	.w7(32'hbb295f9b),
	.w8(32'hbb7525cf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dfe9b),
	.w1(32'h39db7e9b),
	.w2(32'hbb3f6e77),
	.w3(32'hbb3f6031),
	.w4(32'h3928cd26),
	.w5(32'hbb5fee17),
	.w6(32'hbaba96c5),
	.w7(32'hba94faa7),
	.w8(32'hbb6d2605),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba076fd4),
	.w1(32'h371a6d79),
	.w2(32'hbb00ab32),
	.w3(32'hba101231),
	.w4(32'hba909aee),
	.w5(32'hbb41116f),
	.w6(32'hba660cdf),
	.w7(32'hb933cda3),
	.w8(32'hbb3e2385),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac33e09),
	.w1(32'h3a5d2c3b),
	.w2(32'h3a1cc1dc),
	.w3(32'hbb527188),
	.w4(32'h3a426eff),
	.w5(32'hb97b1b20),
	.w6(32'hbb42275b),
	.w7(32'h39a06e0d),
	.w8(32'h3a41108e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0240),
	.w1(32'hbb93cefa),
	.w2(32'hbbadd616),
	.w3(32'hbb856795),
	.w4(32'hbb0eb814),
	.w5(32'hbadf142c),
	.w6(32'hbb85880c),
	.w7(32'hbac8e722),
	.w8(32'hbb0f6a8c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fcea9),
	.w1(32'hb83ba5ca),
	.w2(32'hbb0ff09b),
	.w3(32'hbaa8e96d),
	.w4(32'hba183808),
	.w5(32'hbb42d461),
	.w6(32'hbad8eef1),
	.w7(32'hba2d943a),
	.w8(32'hbb0d4277),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ad73),
	.w1(32'hb88bb28f),
	.w2(32'hb99b88de),
	.w3(32'hbac422a3),
	.w4(32'hba07738f),
	.w5(32'hba23bcd2),
	.w6(32'hba0045ad),
	.w7(32'hba04eb87),
	.w8(32'h38f78d52),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f7dce),
	.w1(32'hba00b234),
	.w2(32'hb949b7e2),
	.w3(32'hba1045b8),
	.w4(32'hba1e034f),
	.w5(32'hb9ea9fd8),
	.w6(32'hba37387b),
	.w7(32'hb9a5b468),
	.w8(32'hb89d0124),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a091dae),
	.w1(32'h399db3ae),
	.w2(32'h39a5493e),
	.w3(32'hb882a0b7),
	.w4(32'hb95dc34c),
	.w5(32'hb98a78a4),
	.w6(32'h37ee449a),
	.w7(32'h39971147),
	.w8(32'h39cd13a5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21fd42),
	.w1(32'h3a0e7248),
	.w2(32'h3a83dcf4),
	.w3(32'hb81bccbb),
	.w4(32'hb9d639d1),
	.w5(32'hba0a1112),
	.w6(32'h39de1c34),
	.w7(32'h39bb49b6),
	.w8(32'h3aa103bf),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b97560),
	.w1(32'h39e17507),
	.w2(32'hbb318bb5),
	.w3(32'hba779d87),
	.w4(32'h3a1eeedf),
	.w5(32'hbb24e158),
	.w6(32'hba346f43),
	.w7(32'h39e057dc),
	.w8(32'hbaaa990f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf3f9e),
	.w1(32'h3a31e947),
	.w2(32'h3a2c72ea),
	.w3(32'hba5a4fb5),
	.w4(32'h39d0c3af),
	.w5(32'h39ce8d90),
	.w6(32'h3a33ba47),
	.w7(32'h3a6f2891),
	.w8(32'h3a92656e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a3272),
	.w1(32'hb913b43e),
	.w2(32'hba5deab0),
	.w3(32'hba8bef16),
	.w4(32'hba7e56ee),
	.w5(32'hba4f597e),
	.w6(32'hb99c2c53),
	.w7(32'h38c3eaf6),
	.w8(32'hb99bda0a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bd273),
	.w1(32'hba1bdb9a),
	.w2(32'hbb26e8de),
	.w3(32'hbb1db86c),
	.w4(32'hb9930519),
	.w5(32'hbb213a25),
	.w6(32'hbb87e8d1),
	.w7(32'hbb1806a6),
	.w8(32'hbb9f8136),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eefb06),
	.w1(32'hb9c222f9),
	.w2(32'h3a50c570),
	.w3(32'hb6e09c36),
	.w4(32'h39c689fa),
	.w5(32'h3abf4f9d),
	.w6(32'h395ee311),
	.w7(32'h3952c71a),
	.w8(32'h39f2499b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3996d),
	.w1(32'h3a07e535),
	.w2(32'h3aca32ed),
	.w3(32'h3aad9b94),
	.w4(32'h3a33802f),
	.w5(32'h3a7ff6e4),
	.w6(32'h39a5e442),
	.w7(32'h3a54f1a4),
	.w8(32'h3a33a593),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb74d8),
	.w1(32'h39a2cc74),
	.w2(32'h39ac4612),
	.w3(32'h3a79adef),
	.w4(32'h39e9dfd8),
	.w5(32'h3a01feb4),
	.w6(32'h36289e1f),
	.w7(32'h391d0bf6),
	.w8(32'h38add267),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d810ed),
	.w1(32'hb951dc93),
	.w2(32'hb6fe4cb2),
	.w3(32'h38ce680d),
	.w4(32'hb9d084f1),
	.w5(32'hb914354d),
	.w6(32'hba858163),
	.w7(32'hb683e3cb),
	.w8(32'hba12d2d8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1d5de),
	.w1(32'hbb54aaaa),
	.w2(32'hbb1fdf40),
	.w3(32'hbad7fa44),
	.w4(32'hbb6ccbeb),
	.w5(32'hbb87e26f),
	.w6(32'hb9d22af5),
	.w7(32'h39158fb4),
	.w8(32'hbaa37574),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28098e),
	.w1(32'hbb75f245),
	.w2(32'hbb89e156),
	.w3(32'hbb162791),
	.w4(32'hbb208aad),
	.w5(32'hbb6bf4f3),
	.w6(32'hbb10258c),
	.w7(32'hb96063c7),
	.w8(32'hbb249c8a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa21ad),
	.w1(32'hb9946b1f),
	.w2(32'hb9720b12),
	.w3(32'h388e0a72),
	.w4(32'h39129c31),
	.w5(32'hb8421987),
	.w6(32'hb8ffab97),
	.w7(32'h3868b892),
	.w8(32'hba1c868e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1949c4),
	.w1(32'hba8a55ff),
	.w2(32'hb900fc4d),
	.w3(32'hbb0393ba),
	.w4(32'hb830e017),
	.w5(32'hb9fc3274),
	.w6(32'hbaaf1f25),
	.w7(32'h37e41a5d),
	.w8(32'hb96e66bb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c844a2),
	.w1(32'h3a451a3f),
	.w2(32'hb96864c6),
	.w3(32'hb947cba3),
	.w4(32'hb9a35e82),
	.w5(32'h3a171e45),
	.w6(32'hbaaa7016),
	.w7(32'hb8deacbc),
	.w8(32'hba0f1adf),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd5518),
	.w1(32'hba2a3b24),
	.w2(32'hbb1a604c),
	.w3(32'hb963586c),
	.w4(32'h39a3d418),
	.w5(32'hb9d78885),
	.w6(32'hbb0a076d),
	.w7(32'hb9a96659),
	.w8(32'hb92bdc35),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb269d97),
	.w1(32'hb9f8bf6d),
	.w2(32'hbb37ddce),
	.w3(32'hbadaa733),
	.w4(32'h3b02dd6d),
	.w5(32'h3a1d0e3b),
	.w6(32'hba16c2a1),
	.w7(32'h39436a71),
	.w8(32'hbae42dbd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45ba6b),
	.w1(32'hbaa63ebc),
	.w2(32'hbba89a54),
	.w3(32'hbb28af90),
	.w4(32'hbb12295f),
	.w5(32'hbb8ade97),
	.w6(32'hbaae86bf),
	.w7(32'hba8450b7),
	.w8(32'hbb91f68b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a4429),
	.w1(32'h3a190404),
	.w2(32'hba88a349),
	.w3(32'hbad1b371),
	.w4(32'h39cbab97),
	.w5(32'hba6b6491),
	.w6(32'hbae9bbe8),
	.w7(32'hb9aa8e65),
	.w8(32'hbb0834ca),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e540e),
	.w1(32'hba0f99c7),
	.w2(32'hbb193e1a),
	.w3(32'hbaa792c7),
	.w4(32'h3a946940),
	.w5(32'h39a308e4),
	.w6(32'hbad09624),
	.w7(32'hb88680ed),
	.w8(32'hbb02e649),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e41cd),
	.w1(32'hbaf075a6),
	.w2(32'hbb3a665a),
	.w3(32'hbb453ae1),
	.w4(32'hbabc79c7),
	.w5(32'hbb23aa65),
	.w6(32'hbac8404f),
	.w7(32'h39334f45),
	.w8(32'hbb1f32ee),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19f850),
	.w1(32'h3ab0816e),
	.w2(32'h3a96d821),
	.w3(32'hbae98010),
	.w4(32'h3b61a0e7),
	.w5(32'h3b40b9e2),
	.w6(32'hbaa66b6d),
	.w7(32'h3ab55200),
	.w8(32'h3a50d5eb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d40ec),
	.w1(32'hba95df71),
	.w2(32'hbb8f13cd),
	.w3(32'h3a18d7b6),
	.w4(32'hba1b9af1),
	.w5(32'hbb0a6c65),
	.w6(32'hbaf52927),
	.w7(32'hbadb5876),
	.w8(32'hbb550a79),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3da279),
	.w1(32'hb912ab6f),
	.w2(32'hba39ed29),
	.w3(32'h37a40d65),
	.w4(32'hb7952431),
	.w5(32'hba1036af),
	.w6(32'hba5c79a8),
	.w7(32'hb9cee7bd),
	.w8(32'hba8f4941),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab85ed2),
	.w1(32'h3a42feb7),
	.w2(32'hba647ac5),
	.w3(32'hbb1bf423),
	.w4(32'hbb26c6ad),
	.w5(32'hbb8ef88d),
	.w6(32'hbb76482e),
	.w7(32'hbb81ee9a),
	.w8(32'hbbb9581f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491bd0),
	.w1(32'hba2b9dda),
	.w2(32'hbaaae73e),
	.w3(32'hbb30d387),
	.w4(32'h391cc2db),
	.w5(32'h391a6a1b),
	.w6(32'hbb760361),
	.w7(32'hba9de78a),
	.w8(32'hbaace75e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8c7ad),
	.w1(32'h38ba5035),
	.w2(32'h3742e274),
	.w3(32'hb95f622f),
	.w4(32'h38434756),
	.w5(32'h3925a94d),
	.w6(32'hb80e60c0),
	.w7(32'h36867bcd),
	.w8(32'h39538e6b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398abaf5),
	.w1(32'h39f16d40),
	.w2(32'h39c693e0),
	.w3(32'h39b70939),
	.w4(32'h3a6a9e77),
	.w5(32'hb9cd4165),
	.w6(32'h3a0869e3),
	.w7(32'h39877c81),
	.w8(32'h3a5c3f6c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c37ce),
	.w1(32'hba5fafb3),
	.w2(32'hba683b34),
	.w3(32'hb9f8a35d),
	.w4(32'h38499ae4),
	.w5(32'hb9421fde),
	.w6(32'hbabb3d70),
	.w7(32'hba0dcac4),
	.w8(32'hbacd51c0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d46e),
	.w1(32'hba24a221),
	.w2(32'hbb240be2),
	.w3(32'hbb485c9e),
	.w4(32'h3a94c70e),
	.w5(32'hba490433),
	.w6(32'hba9e7533),
	.w7(32'hb8e80d36),
	.w8(32'hbb021722),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2bd67),
	.w1(32'h3a8db97b),
	.w2(32'hbb02159f),
	.w3(32'hbb091f03),
	.w4(32'h3a940305),
	.w5(32'hb964019c),
	.w6(32'hbb03c14f),
	.w7(32'hb9893a65),
	.w8(32'hbaf013f7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc1b00),
	.w1(32'hba02fb8d),
	.w2(32'hb99c8fd5),
	.w3(32'h39dc3592),
	.w4(32'hba4ee0da),
	.w5(32'hb9ebf1b4),
	.w6(32'hba28c3a9),
	.w7(32'hb947b6db),
	.w8(32'hba1b3969),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6968cc),
	.w1(32'hba89cde3),
	.w2(32'hbb3eb9dd),
	.w3(32'hbb4550bb),
	.w4(32'hba179bb4),
	.w5(32'hbb227b95),
	.w6(32'hbaa05e52),
	.w7(32'h3a1fba67),
	.w8(32'hbaccbad9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ef07d),
	.w1(32'h39686bbd),
	.w2(32'hbac29516),
	.w3(32'h3a2d4d39),
	.w4(32'h395f04ca),
	.w5(32'hba6af85e),
	.w6(32'hba985428),
	.w7(32'hb9b20f94),
	.w8(32'hba863484),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eaf7f),
	.w1(32'hbb048043),
	.w2(32'hbb1bdd2b),
	.w3(32'hbac64dfa),
	.w4(32'hba7eedea),
	.w5(32'hba1ed050),
	.w6(32'hbaf64b02),
	.w7(32'h39163352),
	.w8(32'hba898f63),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62136a),
	.w1(32'h3ac50b68),
	.w2(32'hbb406c96),
	.w3(32'hba831bde),
	.w4(32'h3afa3088),
	.w5(32'hbb472af7),
	.w6(32'hba90030a),
	.w7(32'h3a89e92e),
	.w8(32'hbb6c4ba4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6aef5f),
	.w1(32'h3a33f48e),
	.w2(32'hbacff4b5),
	.w3(32'hbae8dc5f),
	.w4(32'h39215dcd),
	.w5(32'hba2025ed),
	.w6(32'hb98dc968),
	.w7(32'h3a3227e9),
	.w8(32'hba3db560),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b5464),
	.w1(32'h3a850313),
	.w2(32'h39db12e8),
	.w3(32'h3938dec5),
	.w4(32'h3a00902e),
	.w5(32'h39d5df93),
	.w6(32'h3989f55e),
	.w7(32'h39c19267),
	.w8(32'h39f69bce),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23948f),
	.w1(32'h3b41e678),
	.w2(32'h3a3886f1),
	.w3(32'h3a01787f),
	.w4(32'h3b4e0da4),
	.w5(32'h3959015a),
	.w6(32'h3a03c10b),
	.w7(32'h3ad9bfa3),
	.w8(32'hb9b0058c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d33d9),
	.w1(32'hb91851cc),
	.w2(32'hba5646fe),
	.w3(32'hbb05c096),
	.w4(32'h3ab75e4c),
	.w5(32'h3a2f805b),
	.w6(32'hbb21b5d4),
	.w7(32'h3acb7457),
	.w8(32'hba423d87),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b051ded),
	.w1(32'h3a7b4509),
	.w2(32'h3a0c8f9b),
	.w3(32'h3a866c20),
	.w4(32'h3a920fc5),
	.w5(32'h38e06b11),
	.w6(32'hba8a96a6),
	.w7(32'h3a45938d),
	.w8(32'h39aa79df),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79c525),
	.w1(32'hba0bce63),
	.w2(32'hb96bba9e),
	.w3(32'hba0f0801),
	.w4(32'hba5021c6),
	.w5(32'hb9eb9953),
	.w6(32'hba1522b0),
	.w7(32'hb986ea48),
	.w8(32'hba52e90e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319378),
	.w1(32'h393a3bea),
	.w2(32'hb75e72d5),
	.w3(32'hba2a7236),
	.w4(32'hb90faf71),
	.w5(32'h39466e5a),
	.w6(32'hb93d5417),
	.w7(32'hb8bb1c0e),
	.w8(32'hb9e3aca6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f43da),
	.w1(32'hbabb5754),
	.w2(32'hbba333e3),
	.w3(32'hbac0f9ab),
	.w4(32'hb852d091),
	.w5(32'hbb549535),
	.w6(32'hba7aea2d),
	.w7(32'hbac0d506),
	.w8(32'hbb04d38a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988725e),
	.w1(32'h3b86dbc0),
	.w2(32'h39cf7d58),
	.w3(32'h395335e5),
	.w4(32'h3aedb20b),
	.w5(32'h3a5d78de),
	.w6(32'h3b1fccf8),
	.w7(32'h3ad3f20e),
	.w8(32'h398251ac),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a903f28),
	.w1(32'h3ad78809),
	.w2(32'hba4b9375),
	.w3(32'h399927fb),
	.w4(32'h3a8f11ce),
	.w5(32'hba3087c5),
	.w6(32'hb9da3432),
	.w7(32'h3a08c48e),
	.w8(32'hbad530f7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c12bc),
	.w1(32'h3a482bda),
	.w2(32'h39d79f8e),
	.w3(32'hba39b7ff),
	.w4(32'h3a2155f8),
	.w5(32'h3a2eacca),
	.w6(32'h39cfd2cf),
	.w7(32'h3a0c4be7),
	.w8(32'h391e3fc4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e7f649),
	.w1(32'hb909eae6),
	.w2(32'hbb0ac6a2),
	.w3(32'h38d74dee),
	.w4(32'hb9993bdf),
	.w5(32'hbb3c7dc7),
	.w6(32'hba97f468),
	.w7(32'hbaf63ec6),
	.w8(32'hbb68f3bc),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fb2ea),
	.w1(32'h3914c8ed),
	.w2(32'h39739d02),
	.w3(32'hba4c34af),
	.w4(32'h3727d8f6),
	.w5(32'hb9783ee5),
	.w6(32'h39b69d68),
	.w7(32'hb7981056),
	.w8(32'hb8b9c194),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f02dc2),
	.w1(32'hb911e405),
	.w2(32'h39952415),
	.w3(32'hb9c38e50),
	.w4(32'hb99a9d71),
	.w5(32'h38a3526a),
	.w6(32'hb9c19d65),
	.w7(32'h377758aa),
	.w8(32'h37cf23ed),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397566d9),
	.w1(32'h3a41df6a),
	.w2(32'hbad41e90),
	.w3(32'hb921f1fe),
	.w4(32'h3ad15d7f),
	.w5(32'hba17f100),
	.w6(32'hb99f9245),
	.w7(32'h398e5d2f),
	.w8(32'hbab4e899),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a11f6),
	.w1(32'hbb02de62),
	.w2(32'hbb904bfb),
	.w3(32'hbb49ad97),
	.w4(32'hba500d64),
	.w5(32'hbbb142ad),
	.w6(32'hbb8b7574),
	.w7(32'h3985fdc9),
	.w8(32'hbb29be35),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96ce8e),
	.w1(32'h3b0a396b),
	.w2(32'h3ac7df94),
	.w3(32'h3a8280a6),
	.w4(32'h3b15ece0),
	.w5(32'h3a958ff9),
	.w6(32'hb917b1a7),
	.w7(32'h3a789d08),
	.w8(32'h39589b90),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a353ef4),
	.w1(32'h3b027d74),
	.w2(32'hbaea24ba),
	.w3(32'h3911958b),
	.w4(32'h3a991a91),
	.w5(32'hbade02f9),
	.w6(32'hba21ac90),
	.w7(32'h396b8100),
	.w8(32'hbb4e031f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a102d2f),
	.w1(32'hb8f8a422),
	.w2(32'hbab49997),
	.w3(32'hb91cbdbf),
	.w4(32'h3a86707a),
	.w5(32'hb9be5f8d),
	.w6(32'hb94f5ac2),
	.w7(32'h3a5c082f),
	.w8(32'hba9bbba7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9bddb),
	.w1(32'hbb20043f),
	.w2(32'hbbd897bb),
	.w3(32'hbb9dcb91),
	.w4(32'hba4ae057),
	.w5(32'hbb9a8616),
	.w6(32'hbb9d0239),
	.w7(32'h390d2631),
	.w8(32'hbb8c6aaf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c0510),
	.w1(32'hbaaa07ad),
	.w2(32'hbb91e568),
	.w3(32'hbb206039),
	.w4(32'h39766d7d),
	.w5(32'hbb07b7e4),
	.w6(32'hbb10aeb8),
	.w7(32'hba37a376),
	.w8(32'hbb407aa6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eaeb0),
	.w1(32'hbac53827),
	.w2(32'hbb224517),
	.w3(32'hbb2600e9),
	.w4(32'hbab48cd9),
	.w5(32'hbb00b5e4),
	.w6(32'hbb192c74),
	.w7(32'hba8c1fca),
	.w8(32'hbb1d5792),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65b718),
	.w1(32'h39513514),
	.w2(32'h3a0130ec),
	.w3(32'hb6e667ee),
	.w4(32'h380e1b91),
	.w5(32'h39df4531),
	.w6(32'h39bd0be8),
	.w7(32'h39e1cd73),
	.w8(32'h3a643d43),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1f0d),
	.w1(32'hb8aa8915),
	.w2(32'hbb0d6bd9),
	.w3(32'hbab39670),
	.w4(32'h39b71667),
	.w5(32'hb9b8153e),
	.w6(32'hb9ddeea1),
	.w7(32'h3a1a5ec1),
	.w8(32'hb961e485),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f71bf),
	.w1(32'hba2da66a),
	.w2(32'hb8c971ff),
	.w3(32'h393dfca0),
	.w4(32'hba76f31c),
	.w5(32'hb9fbfedc),
	.w6(32'hba34b35f),
	.w7(32'hb9d1c0c6),
	.w8(32'hb95bea3f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b7216),
	.w1(32'hb9983443),
	.w2(32'hba2cef57),
	.w3(32'hba16e0a5),
	.w4(32'hb9bcc3c0),
	.w5(32'hba2c06e0),
	.w6(32'hbaf5ee0a),
	.w7(32'hbad7e177),
	.w8(32'hbb01fc39),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf99a7c),
	.w1(32'hbabcb44e),
	.w2(32'h3ae4fc65),
	.w3(32'hbb10cb11),
	.w4(32'hb984cf4d),
	.w5(32'hb6866917),
	.w6(32'hbb04fc5d),
	.w7(32'hb9d438ea),
	.w8(32'hba80f563),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b9fbb),
	.w1(32'h395a3eb6),
	.w2(32'hbb0e6dd5),
	.w3(32'hbb4d7c5f),
	.w4(32'h3a0c457b),
	.w5(32'hb8e0f057),
	.w6(32'hbb2f9a23),
	.w7(32'hb9d0d2a3),
	.w8(32'hbae4aa64),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68bec4),
	.w1(32'h399f50ac),
	.w2(32'hba424c2a),
	.w3(32'h3a72d81e),
	.w4(32'h3a26cb31),
	.w5(32'h39d9590a),
	.w6(32'h35d6161b),
	.w7(32'h392c62af),
	.w8(32'h3a1b0e7c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76e6b0),
	.w1(32'h3aa4558a),
	.w2(32'h3a828b59),
	.w3(32'h3a084254),
	.w4(32'h3a8c6e9e),
	.w5(32'h3a6cd3e1),
	.w6(32'h3a9bda3f),
	.w7(32'h3a81c132),
	.w8(32'h3a16e047),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1886dc),
	.w1(32'hba160321),
	.w2(32'h394ac284),
	.w3(32'h398f3b17),
	.w4(32'h3a8c7677),
	.w5(32'hb8fe147e),
	.w6(32'hb9c45be7),
	.w7(32'hb7fb1279),
	.w8(32'h3a026a15),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9bc2c),
	.w1(32'hb862de3f),
	.w2(32'hbb1314b9),
	.w3(32'hbae3392b),
	.w4(32'h3a81f0fc),
	.w5(32'hba8ee99f),
	.w6(32'h398d35d9),
	.w7(32'h3a886b00),
	.w8(32'hba8216d9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9415cc),
	.w1(32'hbb68d8fe),
	.w2(32'hb9cdf53c),
	.w3(32'hbb5f0ebf),
	.w4(32'hbadeaa20),
	.w5(32'h3a95fab4),
	.w6(32'hbb026a2c),
	.w7(32'hb906c874),
	.w8(32'hb98335c8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362b0c),
	.w1(32'h39087329),
	.w2(32'h3a2b035b),
	.w3(32'hb9ea81b0),
	.w4(32'h39a78dc6),
	.w5(32'h387f92be),
	.w6(32'hba00c522),
	.w7(32'h39137c41),
	.w8(32'hb937db7b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b073),
	.w1(32'hbb25237d),
	.w2(32'hbbcea012),
	.w3(32'hbb8801ce),
	.w4(32'h3a33253b),
	.w5(32'hbb6a0b01),
	.w6(32'hb8384a6c),
	.w7(32'h3b550089),
	.w8(32'hba918f4d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9998c),
	.w1(32'h39c8e10a),
	.w2(32'hbbc35dcb),
	.w3(32'hbb08d28f),
	.w4(32'h3ba7000f),
	.w5(32'hba904799),
	.w6(32'hbaba00df),
	.w7(32'h3b828e6c),
	.w8(32'hbb324a08),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5577f),
	.w1(32'hbacc38c6),
	.w2(32'hba8a5130),
	.w3(32'hb9a797a3),
	.w4(32'hbae403e2),
	.w5(32'hbacccb98),
	.w6(32'hba021b70),
	.w7(32'hba346024),
	.w8(32'hba67d08a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972a21e),
	.w1(32'h3aabb08f),
	.w2(32'h3a4c9360),
	.w3(32'hb9669809),
	.w4(32'h3a69bbf8),
	.w5(32'h398e2b28),
	.w6(32'h3ae0f365),
	.w7(32'h3a226cf4),
	.w8(32'h3b29be6c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b303e55),
	.w1(32'hb8be3731),
	.w2(32'hb72a052d),
	.w3(32'h3b033c8d),
	.w4(32'h3a02caf8),
	.w5(32'h39ca31d3),
	.w6(32'h380d74fe),
	.w7(32'hb857ddda),
	.w8(32'hba0b9e04),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985b57c),
	.w1(32'h391a699c),
	.w2(32'hb9472916),
	.w3(32'hb949815d),
	.w4(32'h39671f14),
	.w5(32'hb94f70a1),
	.w6(32'hb8d773f0),
	.w7(32'hb9987dcc),
	.w8(32'h370f73fd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37abcab4),
	.w1(32'hbaa25f1a),
	.w2(32'hbafddf03),
	.w3(32'hb9c62445),
	.w4(32'hbacab2bb),
	.w5(32'hbb0d03c6),
	.w6(32'h395948ae),
	.w7(32'hba5a2cff),
	.w8(32'hbadf096c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34a4dc),
	.w1(32'hba69b3cc),
	.w2(32'hbabe5615),
	.w3(32'hbae7e089),
	.w4(32'hba01b12d),
	.w5(32'hbace580a),
	.w6(32'hbb1f81d3),
	.w7(32'hba5ec848),
	.w8(32'hbb34e8bf),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251b0a),
	.w1(32'hbb100dbc),
	.w2(32'hbb44bb10),
	.w3(32'hbb490046),
	.w4(32'hba81fdb5),
	.w5(32'hba9fcc94),
	.w6(32'hbba4c264),
	.w7(32'hbb09b78c),
	.w8(32'hbb2c571e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b4e5e),
	.w1(32'h3a375114),
	.w2(32'h39254b5d),
	.w3(32'h38d28db7),
	.w4(32'h39c58b5f),
	.w5(32'h399e8a9d),
	.w6(32'hba5bcfa0),
	.w7(32'hb74576b8),
	.w8(32'hb96347b7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fff4d),
	.w1(32'hbb256a93),
	.w2(32'hbbbba721),
	.w3(32'hba6b4f78),
	.w4(32'hba0525ae),
	.w5(32'hbb55c834),
	.w6(32'hbb6c5d58),
	.w7(32'hbb049d86),
	.w8(32'hbbb1f270),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aee36),
	.w1(32'hba781912),
	.w2(32'hba9b326c),
	.w3(32'hbb816bea),
	.w4(32'hba54a8a4),
	.w5(32'hbaac099c),
	.w6(32'hba9f6734),
	.w7(32'hba2ec45d),
	.w8(32'hbabb8206),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9365e2c),
	.w1(32'hb93a4a62),
	.w2(32'h3a108ec0),
	.w3(32'hb9e27af9),
	.w4(32'hb88c0a27),
	.w5(32'h39bb3de0),
	.w6(32'hb93c08d9),
	.w7(32'h3a07c110),
	.w8(32'h3a036ea8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc30b),
	.w1(32'hbb29ddbb),
	.w2(32'hbad9288e),
	.w3(32'hba938351),
	.w4(32'hbaa85a84),
	.w5(32'hb9a00f9c),
	.w6(32'hbab57aae),
	.w7(32'hb9b5932c),
	.w8(32'h3a036a5f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cae952),
	.w1(32'h3a54987b),
	.w2(32'h39aaefe9),
	.w3(32'h39bb65a6),
	.w4(32'h3a025a57),
	.w5(32'h3a1d97dc),
	.w6(32'h3a0db96b),
	.w7(32'h39dea484),
	.w8(32'h37877ec0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf998f7),
	.w1(32'hb880dad4),
	.w2(32'hbacfd3aa),
	.w3(32'hba6f6670),
	.w4(32'h3a07ce85),
	.w5(32'hbb0752b6),
	.w6(32'hbae87f52),
	.w7(32'hb9b02944),
	.w8(32'hbb53b602),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48d5b8),
	.w1(32'h3aa88094),
	.w2(32'hbb03212f),
	.w3(32'hbb1c9f8a),
	.w4(32'h3b41c85b),
	.w5(32'h3a1afb50),
	.w6(32'hbb3268e2),
	.w7(32'h39dfeeb4),
	.w8(32'hbb6a6d91),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed7173),
	.w1(32'h37f65df1),
	.w2(32'hbb18ca0a),
	.w3(32'h39cfc5b0),
	.w4(32'h39c8329b),
	.w5(32'hbacf6887),
	.w6(32'hbb1b2c5c),
	.w7(32'hba4ca942),
	.w8(32'hbb4e6c94),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8c2cd),
	.w1(32'h3a7f88b2),
	.w2(32'h3ab70d4b),
	.w3(32'hb9912616),
	.w4(32'h3a72b884),
	.w5(32'h39a82fed),
	.w6(32'h392b471e),
	.w7(32'h3a3dad30),
	.w8(32'h3aa9bb4f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac921e),
	.w1(32'h3b49f8f9),
	.w2(32'hbb393bf2),
	.w3(32'h366e50bd),
	.w4(32'h3b5f516e),
	.w5(32'hba963cd1),
	.w6(32'hb7db625a),
	.w7(32'h3a50d734),
	.w8(32'hbb731924),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3cd56),
	.w1(32'hba9c518e),
	.w2(32'hbb11c280),
	.w3(32'hba0d72c4),
	.w4(32'hb9d0ffaa),
	.w5(32'hba71a192),
	.w6(32'hbb0bf9e2),
	.w7(32'hb98f7005),
	.w8(32'hbaa629fd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88bf3b),
	.w1(32'hbb086697),
	.w2(32'hbb8523c0),
	.w3(32'hbb839be0),
	.w4(32'hbaa9a469),
	.w5(32'hbb3e76be),
	.w6(32'hbb969de7),
	.w7(32'hbb0fbc8b),
	.w8(32'hbb81f9f5),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e975),
	.w1(32'h38187588),
	.w2(32'hb9a95e27),
	.w3(32'h3a18f6ef),
	.w4(32'h39be7dc9),
	.w5(32'hb9c2aece),
	.w6(32'hb8a5fda1),
	.w7(32'hb9228a5a),
	.w8(32'hb95e5b63),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b0ad4),
	.w1(32'h38bf15d6),
	.w2(32'h3a06205a),
	.w3(32'hb9a0a794),
	.w4(32'h39418b50),
	.w5(32'h399b3c40),
	.w6(32'h397763f7),
	.w7(32'h39c59a28),
	.w8(32'h39d775da),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1af54b),
	.w1(32'hbab1ec10),
	.w2(32'hbb1b40f5),
	.w3(32'hbaa2dfff),
	.w4(32'h39306a44),
	.w5(32'hbae502f1),
	.w6(32'hbb5168f7),
	.w7(32'h38c15467),
	.w8(32'hbb107494),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34db5a),
	.w1(32'hb9d79244),
	.w2(32'hbb5c6c89),
	.w3(32'hbb0a4990),
	.w4(32'h385e695f),
	.w5(32'hbb81a3b6),
	.w6(32'hbafec2b2),
	.w7(32'hb8a85d12),
	.w8(32'hbb5d3b6e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b0d8c),
	.w1(32'hba189988),
	.w2(32'hbb3319a2),
	.w3(32'hbad59824),
	.w4(32'h3a816d51),
	.w5(32'hbab8c4a2),
	.w6(32'hbb551b89),
	.w7(32'h38c46e65),
	.w8(32'hbaa387ee),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba667b71),
	.w1(32'hbae94e3d),
	.w2(32'hba81a575),
	.w3(32'hbabf0e3e),
	.w4(32'hbb2549b5),
	.w5(32'hba9aa177),
	.w6(32'h3a86cd9b),
	.w7(32'hb9b5fe85),
	.w8(32'hba618f81),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b73c2),
	.w1(32'hba227b01),
	.w2(32'hb9c9de2b),
	.w3(32'h39b4c2f9),
	.w4(32'hb9c44ceb),
	.w5(32'hb8de567c),
	.w6(32'hba2de97d),
	.w7(32'hb9c9c80d),
	.w8(32'hb87028da),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9b530),
	.w1(32'hb9896f6f),
	.w2(32'h39e768f1),
	.w3(32'hba2ab1c3),
	.w4(32'h39a40747),
	.w5(32'h3a133836),
	.w6(32'h39aa03e2),
	.w7(32'h39cb2f95),
	.w8(32'h39500ef8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2da3ff),
	.w1(32'hba8e068b),
	.w2(32'hbaf4bac9),
	.w3(32'hbb08b66d),
	.w4(32'hbb868007),
	.w5(32'hbba05db1),
	.w6(32'hbb2ee8d4),
	.w7(32'h3a06b35f),
	.w8(32'hbaf7a8c9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf536ed),
	.w1(32'hbb66ff50),
	.w2(32'hbb9d9b73),
	.w3(32'hbba7f1cb),
	.w4(32'hbb0590ed),
	.w5(32'hbb6ad94d),
	.w6(32'hbb8e5a77),
	.w7(32'hb9d05e15),
	.w8(32'hbb52f8b1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88824e),
	.w1(32'hbb0c6a2c),
	.w2(32'hbb053521),
	.w3(32'hbb0ffed4),
	.w4(32'hbaba5daf),
	.w5(32'hbaca4791),
	.w6(32'hbb0129f6),
	.w7(32'h37c5eda1),
	.w8(32'hbaf0d33d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39240030),
	.w1(32'h3b2fb96f),
	.w2(32'h3a8aae34),
	.w3(32'hbac53a4d),
	.w4(32'h3aba547d),
	.w5(32'hb96e4ef4),
	.w6(32'hbb06329c),
	.w7(32'hb9c4d2f2),
	.w8(32'hbae2b9e7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29ae52),
	.w1(32'hba8a0a77),
	.w2(32'hbb54051f),
	.w3(32'hbb3d43af),
	.w4(32'h3a46e31c),
	.w5(32'hbac25202),
	.w6(32'hbb4b8d12),
	.w7(32'hba554c97),
	.w8(32'hbb31164d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa17659),
	.w1(32'h3901bc24),
	.w2(32'h3a32ba39),
	.w3(32'h3a73d662),
	.w4(32'h39e30e6f),
	.w5(32'h39c2ca8e),
	.w6(32'h3a09480f),
	.w7(32'h3a4f9efb),
	.w8(32'h3a18bb0e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9f81d),
	.w1(32'hb9d5a7d4),
	.w2(32'hb9e3fab7),
	.w3(32'h3971fc9d),
	.w4(32'hb9ae19ad),
	.w5(32'h39a64676),
	.w6(32'h39c91237),
	.w7(32'hb826382a),
	.w8(32'h39886bf5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924508),
	.w1(32'h395dcdec),
	.w2(32'h3aab0adb),
	.w3(32'h3ab5fc76),
	.w4(32'hba32681f),
	.w5(32'h393e9472),
	.w6(32'h38ca1d5e),
	.w7(32'h3abd188c),
	.w8(32'h3a99b148),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacfd40),
	.w1(32'h3a40b508),
	.w2(32'h3aa30809),
	.w3(32'h3abd7313),
	.w4(32'h3a41db76),
	.w5(32'h3a4bcb19),
	.w6(32'h398c05b2),
	.w7(32'h3a2e42eb),
	.w8(32'h39962447),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9ecd7),
	.w1(32'hba3ddd0a),
	.w2(32'hbae75e10),
	.w3(32'h391e1d86),
	.w4(32'hba6a9575),
	.w5(32'hbb12da7e),
	.w6(32'h39e5730f),
	.w7(32'hba23428b),
	.w8(32'hbaaf631e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62064e),
	.w1(32'hba7892df),
	.w2(32'hbb3f918a),
	.w3(32'hbae70620),
	.w4(32'h3a07d7fb),
	.w5(32'hbadd63e4),
	.w6(32'hbabe1aa3),
	.w7(32'h3965052c),
	.w8(32'hbb084379),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1cdd3),
	.w1(32'h3b571228),
	.w2(32'hba6f15b7),
	.w3(32'hba3f95b2),
	.w4(32'h3aff5e45),
	.w5(32'hb9a60b3d),
	.w6(32'h3a372fc8),
	.w7(32'h3a0ceb42),
	.w8(32'hba2394cf),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd0899),
	.w1(32'hba09776b),
	.w2(32'hb81c4c93),
	.w3(32'h3ad7cf59),
	.w4(32'hb9d2da20),
	.w5(32'h37b4112f),
	.w6(32'hba062179),
	.w7(32'h38ba9a8b),
	.w8(32'h3a075a38),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2d390),
	.w1(32'hbb921b5e),
	.w2(32'hbb852b62),
	.w3(32'hbb64c6a1),
	.w4(32'hbb766f9c),
	.w5(32'hbb0a0a21),
	.w6(32'hbb668b15),
	.w7(32'hb8e1a2c5),
	.w8(32'hbade1f67),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14d56a),
	.w1(32'hba997670),
	.w2(32'hba42f221),
	.w3(32'hba69b726),
	.w4(32'hba1331fd),
	.w5(32'hba2e99b4),
	.w6(32'hbaa71d29),
	.w7(32'h38467758),
	.w8(32'hba1fc0be),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe6dac),
	.w1(32'hb9c0fb5e),
	.w2(32'h388d573a),
	.w3(32'h3905d854),
	.w4(32'hba265da6),
	.w5(32'hb6c50de4),
	.w6(32'hb9b837a9),
	.w7(32'hb9b7a3cc),
	.w8(32'hb917bebd),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4208e),
	.w1(32'h39d4cbfe),
	.w2(32'hba98d677),
	.w3(32'hba473c50),
	.w4(32'h3a02793d),
	.w5(32'hb9c1b31f),
	.w6(32'hb8d557b5),
	.w7(32'h399a0402),
	.w8(32'hb9acd6f3),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b8bae),
	.w1(32'h39e15826),
	.w2(32'h3a716bbb),
	.w3(32'h38bd8ec2),
	.w4(32'h3a0a5a2f),
	.w5(32'h3a236af9),
	.w6(32'h3a1a84ea),
	.w7(32'h3a82f2f8),
	.w8(32'h3a89e699),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71fc72),
	.w1(32'hba04ca73),
	.w2(32'hb997621d),
	.w3(32'h3a244918),
	.w4(32'hb99183d9),
	.w5(32'hb9b93f47),
	.w6(32'hb9e3e141),
	.w7(32'hba021688),
	.w8(32'hba3a5f24),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eca65a),
	.w1(32'hb9693c78),
	.w2(32'h38068182),
	.w3(32'hb9b8bf08),
	.w4(32'hba004383),
	.w5(32'hb881ee1f),
	.w6(32'hb959037d),
	.w7(32'hb9408aa6),
	.w8(32'hb8d96c2b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a9edd),
	.w1(32'hb99f2996),
	.w2(32'h3a2f6287),
	.w3(32'hb8a44eb3),
	.w4(32'hb9fb4dd7),
	.w5(32'hb98e6c63),
	.w6(32'hb9263e58),
	.w7(32'h39bef241),
	.w8(32'hb8d1d63c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a422e),
	.w1(32'h3a2d1393),
	.w2(32'hb9b12cd8),
	.w3(32'hbaac8eab),
	.w4(32'hb98489cb),
	.w5(32'hba49fc10),
	.w6(32'hbaf11ed1),
	.w7(32'hba4b30ef),
	.w8(32'hba8b0ffd),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb392343),
	.w1(32'hbb5713ae),
	.w2(32'hbbfa387a),
	.w3(32'hbb490530),
	.w4(32'hbb137726),
	.w5(32'hbba6c029),
	.w6(32'hbb5d5533),
	.w7(32'hba4910f6),
	.w8(32'hbb3636c2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1dbba),
	.w1(32'hbaafb479),
	.w2(32'hbb5e3e3f),
	.w3(32'h3a27ed7f),
	.w4(32'hb93c249f),
	.w5(32'hba83a6b0),
	.w6(32'hba3aa097),
	.w7(32'h3a443a14),
	.w8(32'hba1ad97e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4860),
	.w1(32'hba88d92e),
	.w2(32'hbb41c9db),
	.w3(32'hbaf82004),
	.w4(32'h398d1300),
	.w5(32'hbab24245),
	.w6(32'hbab7a61b),
	.w7(32'h399947aa),
	.w8(32'hbadabc39),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00a8aa),
	.w1(32'h3a12fd66),
	.w2(32'hba60b61d),
	.w3(32'h392dd89b),
	.w4(32'hb904a093),
	.w5(32'hb9f9d647),
	.w6(32'hb9ca5f12),
	.w7(32'h38044701),
	.w8(32'hb905bf32),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba768bae),
	.w1(32'hba3d5f02),
	.w2(32'hb9811022),
	.w3(32'hba2e9e37),
	.w4(32'hba4ede6f),
	.w5(32'hb904e198),
	.w6(32'hb9ee1fe7),
	.w7(32'hb9ca2488),
	.w8(32'hb9bec817),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d17eae),
	.w1(32'h399a2db3),
	.w2(32'h3a1c0759),
	.w3(32'hb8f2cfd6),
	.w4(32'h397e0706),
	.w5(32'h39d72a3d),
	.w6(32'h39048e36),
	.w7(32'h39abc295),
	.w8(32'h39a9e869),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adeb07),
	.w1(32'h39e3e9ed),
	.w2(32'h3a2c854b),
	.w3(32'h39d44b7a),
	.w4(32'h39dab86d),
	.w5(32'h3a1beb18),
	.w6(32'h39a6813b),
	.w7(32'h39b7eb66),
	.w8(32'h39bde0d4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cebe3),
	.w1(32'hbb7328dc),
	.w2(32'hbb9a045a),
	.w3(32'hbb2b4c3b),
	.w4(32'hba94c3f0),
	.w5(32'hbb5304ca),
	.w6(32'hbb6c4fae),
	.w7(32'hb9d3c943),
	.w8(32'hbb173645),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a3214),
	.w1(32'h3aa9afba),
	.w2(32'h3a05220a),
	.w3(32'hba07d2d0),
	.w4(32'h3a8e65f3),
	.w5(32'h38c191ba),
	.w6(32'h3a95079e),
	.w7(32'hb97bb23e),
	.w8(32'h3845c5dd),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a40884),
	.w1(32'h3ab3c148),
	.w2(32'h3aa2ce0b),
	.w3(32'hb9c920a6),
	.w4(32'h3a9801a7),
	.w5(32'h3a6209fa),
	.w6(32'hb975a383),
	.w7(32'h3a049df4),
	.w8(32'h393cf3c0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ce6be),
	.w1(32'hb9a55293),
	.w2(32'hba309116),
	.w3(32'hbacb9390),
	.w4(32'h38b27964),
	.w5(32'hb8cb91aa),
	.w6(32'hb9b388b6),
	.w7(32'h399f5b1c),
	.w8(32'h3862d1ef),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396de84d),
	.w1(32'h378e2a7d),
	.w2(32'h399b8a6c),
	.w3(32'h38b3b6bc),
	.w4(32'hb98610ba),
	.w5(32'h385ca409),
	.w6(32'hb8df83d6),
	.w7(32'h3829bfb7),
	.w8(32'h38f36d6e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5968e),
	.w1(32'hbac5ba6a),
	.w2(32'hba4b5298),
	.w3(32'hba23a17c),
	.w4(32'hbadb58df),
	.w5(32'hbae32709),
	.w6(32'hba9657f4),
	.w7(32'h39ebd515),
	.w8(32'hb95251ee),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39629ffd),
	.w1(32'h3b0107a4),
	.w2(32'h3abc81e5),
	.w3(32'h39add870),
	.w4(32'h3ae92bba),
	.w5(32'h3acf1d73),
	.w6(32'h3a839be0),
	.w7(32'h3a93132a),
	.w8(32'h3a2be86c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966af5),
	.w1(32'hbb319cf5),
	.w2(32'hbbc858f0),
	.w3(32'hbb851472),
	.w4(32'h3abd014f),
	.w5(32'hb91976e1),
	.w6(32'hbb6fc6d0),
	.w7(32'h3b0fc7a9),
	.w8(32'hba5a7d47),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a91dab),
	.w1(32'hba2c005e),
	.w2(32'hba502505),
	.w3(32'hb7bfcfd9),
	.w4(32'hba2764ad),
	.w5(32'hba7437d8),
	.w6(32'hba080469),
	.w7(32'hba2f33bd),
	.w8(32'hba4ae5b8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d85e),
	.w1(32'h3aefdcd8),
	.w2(32'h3aca0012),
	.w3(32'hbab444c2),
	.w4(32'h3afdc108),
	.w5(32'h39e5725b),
	.w6(32'hbb8ef6fd),
	.w7(32'hb9cb7e5e),
	.w8(32'h3a08718e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule