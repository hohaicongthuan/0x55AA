module layer_10_featuremap_83(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58001e),
	.w1(32'h3b566ec9),
	.w2(32'h3b26df6f),
	.w3(32'hbb363698),
	.w4(32'hba226ec7),
	.w5(32'hbb1fbf39),
	.w6(32'hbbd93f2b),
	.w7(32'h3ad4b76f),
	.w8(32'hbb172b2b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01c103),
	.w1(32'h3c7bc001),
	.w2(32'hbb07a1ad),
	.w3(32'hba291919),
	.w4(32'hb8c05643),
	.w5(32'h3a4d5748),
	.w6(32'hba88ffa4),
	.w7(32'hbb4cd375),
	.w8(32'h3b95598f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d1fc),
	.w1(32'h3b2d23f2),
	.w2(32'h3be7deb9),
	.w3(32'h3cf30feb),
	.w4(32'hbc20a246),
	.w5(32'hbb3a76ee),
	.w6(32'h3c1964fd),
	.w7(32'hbafc2c7a),
	.w8(32'hbb82ea4a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9348c0),
	.w1(32'h3a24b099),
	.w2(32'h3913d63e),
	.w3(32'hbc15e289),
	.w4(32'hbb7844c9),
	.w5(32'hbbb02f5d),
	.w6(32'hbbde70a7),
	.w7(32'hbbaa11f0),
	.w8(32'hba87913c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa63e27),
	.w1(32'h3b20e050),
	.w2(32'hbb8e4115),
	.w3(32'h3b59741b),
	.w4(32'hbb6dd516),
	.w5(32'h3ab03e51),
	.w6(32'h3b0e1ec8),
	.w7(32'h3b994be7),
	.w8(32'h3ca8cdb6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4262d4),
	.w1(32'h3c1676ca),
	.w2(32'h3a08a1ba),
	.w3(32'h3bbf9c01),
	.w4(32'hba7bb5ee),
	.w5(32'hbc058a70),
	.w6(32'h3ac54621),
	.w7(32'hbb0965a0),
	.w8(32'hbc49308a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c1d60),
	.w1(32'hbb75cb69),
	.w2(32'hbb6a53ff),
	.w3(32'h3a0c51d7),
	.w4(32'h3a0a8fc1),
	.w5(32'hbc1d9508),
	.w6(32'h3b614db5),
	.w7(32'h3b7923a6),
	.w8(32'h39e27e13),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1a3ed),
	.w1(32'h3c62a10b),
	.w2(32'h3be9f4a1),
	.w3(32'hbb7afd56),
	.w4(32'hbb76efe2),
	.w5(32'h3a76d4f5),
	.w6(32'h3c663d05),
	.w7(32'h3bc22e33),
	.w8(32'hbc0a390c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ace10),
	.w1(32'h3ba64526),
	.w2(32'h3c1fdd66),
	.w3(32'h3b286412),
	.w4(32'hbc1fddc2),
	.w5(32'h3b1dfe5c),
	.w6(32'hb975e98e),
	.w7(32'hbb3f1de0),
	.w8(32'hb9f41754),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec2828),
	.w1(32'hbaacaf2b),
	.w2(32'hbbb3f32a),
	.w3(32'hbb12b3ee),
	.w4(32'hbb5b509f),
	.w5(32'hbc00c0fb),
	.w6(32'hbc15f60b),
	.w7(32'hbb2fe5e6),
	.w8(32'hba9e3d91),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92d23e),
	.w1(32'h3a32607d),
	.w2(32'hba2fe3a4),
	.w3(32'h3aebcaf5),
	.w4(32'h3bb92b49),
	.w5(32'hbb0c8a8f),
	.w6(32'h3a5db8b7),
	.w7(32'hbaa7f91c),
	.w8(32'h39a8ab2f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c24d3),
	.w1(32'h3baf700f),
	.w2(32'h3b86cae6),
	.w3(32'hbb084753),
	.w4(32'h3ac8c938),
	.w5(32'h3b04cdd3),
	.w6(32'h3abe945a),
	.w7(32'h3ae4bd21),
	.w8(32'hb8d9ff0d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849609),
	.w1(32'hba85befb),
	.w2(32'hbbb1c5be),
	.w3(32'hbbf3ea4b),
	.w4(32'h3915b9b6),
	.w5(32'hbac03c87),
	.w6(32'hbb8aab75),
	.w7(32'hbc0772c3),
	.w8(32'hbbad8d05),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ebb8f),
	.w1(32'h3c0c1c59),
	.w2(32'h3a44abbc),
	.w3(32'hbb04a8e9),
	.w4(32'h3b9c5cfb),
	.w5(32'hbb12dd73),
	.w6(32'h3b6c3e57),
	.w7(32'h3adebf27),
	.w8(32'h3c3a2712),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f34c),
	.w1(32'hb94b3e7f),
	.w2(32'hbacf04d2),
	.w3(32'h3b252b6f),
	.w4(32'hba014cc9),
	.w5(32'h3b8dced0),
	.w6(32'hbbb8168a),
	.w7(32'hbc15bccd),
	.w8(32'hba14917c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6a39e),
	.w1(32'h3a71b5f0),
	.w2(32'hbbbee089),
	.w3(32'hbbd18a67),
	.w4(32'hbaa60727),
	.w5(32'hbbe62b27),
	.w6(32'h3ad80bbc),
	.w7(32'hba80d90d),
	.w8(32'hbc2e6e52),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0600d4),
	.w1(32'hbb924e32),
	.w2(32'hba59f4ca),
	.w3(32'h3ba4d47a),
	.w4(32'hb81e2332),
	.w5(32'h3b08da0d),
	.w6(32'h3b19c690),
	.w7(32'h3a2232f3),
	.w8(32'h3a5daa58),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9eb92),
	.w1(32'h3b971714),
	.w2(32'hbc5308c0),
	.w3(32'hbb100c19),
	.w4(32'hbbde5a71),
	.w5(32'hbb5300b4),
	.w6(32'hbc697ee6),
	.w7(32'h3a063942),
	.w8(32'hbb9aedea),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced1637),
	.w1(32'hbbbb2708),
	.w2(32'hbbf490a9),
	.w3(32'hbaa51cdc),
	.w4(32'h3acdd1f0),
	.w5(32'hbae9eec6),
	.w6(32'h3a266b0f),
	.w7(32'hbba710cb),
	.w8(32'h38b66dd8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58d86),
	.w1(32'h3bb1aba0),
	.w2(32'h3ba037d8),
	.w3(32'hbb759181),
	.w4(32'hbaab48e7),
	.w5(32'h38206cf7),
	.w6(32'h3b5ddb15),
	.w7(32'h3a85d556),
	.w8(32'hbb33fd32),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb988c07),
	.w1(32'hbb4c398b),
	.w2(32'hb9b307f4),
	.w3(32'hbbbd5655),
	.w4(32'hbb2a382b),
	.w5(32'h3c801703),
	.w6(32'hbae1cfe4),
	.w7(32'hbb8ad82c),
	.w8(32'hb9727a44),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43303e),
	.w1(32'h39d35b06),
	.w2(32'hba62e711),
	.w3(32'hb920860d),
	.w4(32'h3baf57cf),
	.w5(32'hbb950843),
	.w6(32'h3b9343b9),
	.w7(32'h3aaa2c11),
	.w8(32'h3a19f64f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57edfd),
	.w1(32'h3b81a0b9),
	.w2(32'hbb3760f6),
	.w3(32'hbb49ee45),
	.w4(32'h3b6a035d),
	.w5(32'h3bf5e857),
	.w6(32'h3c7bca88),
	.w7(32'hbacd43af),
	.w8(32'h3b168b5a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0d3fd),
	.w1(32'hbb25a795),
	.w2(32'hbb312ee8),
	.w3(32'hbbb14701),
	.w4(32'h3ba34a55),
	.w5(32'hbbb8f468),
	.w6(32'hbba7feb7),
	.w7(32'h3c016059),
	.w8(32'hbbd5c5b8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89bfd2),
	.w1(32'h3b06e355),
	.w2(32'h3bc39f84),
	.w3(32'h3b66126d),
	.w4(32'h3b028540),
	.w5(32'hbb250904),
	.w6(32'hbad22ccb),
	.w7(32'hba66d80e),
	.w8(32'hbb8ff79b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24186c),
	.w1(32'h3a49c165),
	.w2(32'hbacbf218),
	.w3(32'hb95d034f),
	.w4(32'h3c9802ac),
	.w5(32'hb974aa74),
	.w6(32'h3ba5914f),
	.w7(32'h3cb95d29),
	.w8(32'hbb4b31f1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a363c5),
	.w1(32'h3a046562),
	.w2(32'h3b990ad5),
	.w3(32'h3a87cb7f),
	.w4(32'h3bcafb2e),
	.w5(32'h3b896869),
	.w6(32'h3ccb472a),
	.w7(32'h3be73a27),
	.w8(32'hbac3a73b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269f44),
	.w1(32'hbb1ee269),
	.w2(32'h3b19be1b),
	.w3(32'hbb09201b),
	.w4(32'hbb99aa4f),
	.w5(32'hbbf5e8c9),
	.w6(32'h3a6ad9df),
	.w7(32'h3cbbc745),
	.w8(32'hbb8ad7d5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a1830),
	.w1(32'h3a3ecc15),
	.w2(32'h3c82afb1),
	.w3(32'hbb3322f5),
	.w4(32'h3925fa5f),
	.w5(32'hbb88e495),
	.w6(32'hbb933193),
	.w7(32'h3a6f9b3f),
	.w8(32'h3b126501),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185240),
	.w1(32'hbb201934),
	.w2(32'hbbd5be25),
	.w3(32'hbb577d91),
	.w4(32'h3b24a241),
	.w5(32'hbbdc9ec2),
	.w6(32'hbb0f9e10),
	.w7(32'hbbc90699),
	.w8(32'hbbb9efa4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39916b1c),
	.w1(32'hbb868f94),
	.w2(32'h3996999c),
	.w3(32'h3aa694c6),
	.w4(32'h3ac274e7),
	.w5(32'hba3ac5a3),
	.w6(32'hbabedbf0),
	.w7(32'hbb1bc437),
	.w8(32'hbbcfa33e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce0a6),
	.w1(32'hb9da97e8),
	.w2(32'hbaeb1f36),
	.w3(32'h3aa5f1cd),
	.w4(32'hbaf96309),
	.w5(32'h3bcabf29),
	.w6(32'hbb463fbc),
	.w7(32'h3c9095fd),
	.w8(32'h3b247243),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6ad5),
	.w1(32'h3b9b3889),
	.w2(32'h3b88f47f),
	.w3(32'hbbd1f1f9),
	.w4(32'h3b961a72),
	.w5(32'h3af1f430),
	.w6(32'h3b0cb58f),
	.w7(32'hbb330e00),
	.w8(32'h396afd07),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c006),
	.w1(32'h3c265491),
	.w2(32'hbc8e09ac),
	.w3(32'h3ab01a52),
	.w4(32'hbb48c449),
	.w5(32'hbb290e03),
	.w6(32'hbb351ec0),
	.w7(32'hbbce07ab),
	.w8(32'h3b88bc81),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840d17),
	.w1(32'hbb8a8936),
	.w2(32'hbae1a893),
	.w3(32'h3a5814c8),
	.w4(32'h3b1f3499),
	.w5(32'hb7dd98d0),
	.w6(32'hbad5f3f9),
	.w7(32'hba714682),
	.w8(32'hbaf4c59a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8e987),
	.w1(32'h3b8c4275),
	.w2(32'hba9978a0),
	.w3(32'hbaf3cc04),
	.w4(32'hbb96691f),
	.w5(32'h3a5b727c),
	.w6(32'h3c2771d8),
	.w7(32'h3b2159e7),
	.w8(32'hbb7f9080),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8add8),
	.w1(32'h3bafea49),
	.w2(32'hbbc157da),
	.w3(32'hbbc6e20c),
	.w4(32'h3b2ef56e),
	.w5(32'h3b0b02e7),
	.w6(32'hbb6242eb),
	.w7(32'hba2f5114),
	.w8(32'hbb876a8b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a3fe),
	.w1(32'hba408668),
	.w2(32'hbb3616f8),
	.w3(32'hbbfd9d0e),
	.w4(32'h3ccb8807),
	.w5(32'h3b1e9ec4),
	.w6(32'h3b472671),
	.w7(32'h3bc9f64f),
	.w8(32'h3aa03c9c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3593f7),
	.w1(32'hbbdc06ca),
	.w2(32'hba13a45c),
	.w3(32'h3b9931db),
	.w4(32'hbb6973f2),
	.w5(32'h3a4444fb),
	.w6(32'hba58fc14),
	.w7(32'hba4d2e0c),
	.w8(32'h3ab30f61),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6d1fe),
	.w1(32'hbb264b83),
	.w2(32'hbaf31835),
	.w3(32'hbaa6ebe4),
	.w4(32'h3c5f307c),
	.w5(32'hbb648b7b),
	.w6(32'h3cb45120),
	.w7(32'hbb668404),
	.w8(32'h3cad9191),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962a3e7),
	.w1(32'hbaf6fc97),
	.w2(32'hbada1169),
	.w3(32'h3cf34596),
	.w4(32'hba8e4c32),
	.w5(32'hb9f7db9a),
	.w6(32'hb903183c),
	.w7(32'hbb5814aa),
	.w8(32'hba25ceac),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba258a5),
	.w1(32'hbb2e6ccc),
	.w2(32'h3b5ecf47),
	.w3(32'hbba7c6ec),
	.w4(32'h3ca9e711),
	.w5(32'h3bff6340),
	.w6(32'h3a20dd57),
	.w7(32'h3b2e1a92),
	.w8(32'hbb73341f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45da64),
	.w1(32'h3a4753be),
	.w2(32'hbbc48382),
	.w3(32'h39d31449),
	.w4(32'h3bd18f77),
	.w5(32'h3b96b215),
	.w6(32'h3b6403ed),
	.w7(32'h3c0d663e),
	.w8(32'h39451b71),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b260578),
	.w1(32'hba686da5),
	.w2(32'hbc06f163),
	.w3(32'hbbe7e75a),
	.w4(32'hbb76c6a9),
	.w5(32'hbbabbca7),
	.w6(32'hbc317ed7),
	.w7(32'h3c1ece68),
	.w8(32'hbbee91d9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163096),
	.w1(32'h3ba177b9),
	.w2(32'hbb9a276e),
	.w3(32'hbb88d391),
	.w4(32'hba8a39b3),
	.w5(32'h3b541029),
	.w6(32'hbbd001e7),
	.w7(32'hbb6860f2),
	.w8(32'hbb0eae87),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3178a9),
	.w1(32'hbbb9fb1a),
	.w2(32'hbac54b5e),
	.w3(32'hbb997f6c),
	.w4(32'hbb0e55fc),
	.w5(32'hbb464e1c),
	.w6(32'hbb4c6700),
	.w7(32'h3b29d36e),
	.w8(32'hbbc99ea7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85f73f),
	.w1(32'hba5838ff),
	.w2(32'hbb66457f),
	.w3(32'h3cb7f235),
	.w4(32'hbad44c8e),
	.w5(32'h3b53368c),
	.w6(32'hbb39c7ed),
	.w7(32'h3b77143c),
	.w8(32'hbbd62903),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8aa16),
	.w1(32'h3a868687),
	.w2(32'hbb85c617),
	.w3(32'hbaf12d90),
	.w4(32'h3c543f20),
	.w5(32'hb9de9533),
	.w6(32'h3b8a1553),
	.w7(32'hbb7ee64d),
	.w8(32'h3bf897e5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e0259),
	.w1(32'h3bb5b59e),
	.w2(32'h3c194450),
	.w3(32'hbb5518ca),
	.w4(32'hbaf357d9),
	.w5(32'h38631f5d),
	.w6(32'hba1a827f),
	.w7(32'hbb62833b),
	.w8(32'h3af3956f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c2d31),
	.w1(32'h3a80526c),
	.w2(32'h3b2d9387),
	.w3(32'h3b0ffb2b),
	.w4(32'h3b7ef3e5),
	.w5(32'h39fdb467),
	.w6(32'hbb8e06ae),
	.w7(32'h3a42f39c),
	.w8(32'hbb49e509),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47548c),
	.w1(32'h3b1163e1),
	.w2(32'hbaea8f88),
	.w3(32'h3aaf3697),
	.w4(32'h3b87ac7e),
	.w5(32'hb8835b4f),
	.w6(32'h3993e17a),
	.w7(32'h398c09cf),
	.w8(32'h39bd313d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831f23),
	.w1(32'h3b67c62a),
	.w2(32'hbbdfb742),
	.w3(32'hba769b5b),
	.w4(32'hbb97633a),
	.w5(32'h3b180cd0),
	.w6(32'hbc6e210c),
	.w7(32'h3a969ab6),
	.w8(32'hbb19b530),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04952),
	.w1(32'hba8c7dc8),
	.w2(32'hbb93b398),
	.w3(32'hbb8d3671),
	.w4(32'hbba0adf3),
	.w5(32'h3b492c84),
	.w6(32'h3b91c38e),
	.w7(32'hbb607c6f),
	.w8(32'h3c466d0b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed50f9),
	.w1(32'hbc03ea80),
	.w2(32'hbbac49d5),
	.w3(32'hbb2a4bd9),
	.w4(32'hbc29cf6c),
	.w5(32'hbb05b6af),
	.w6(32'hbbf22bcb),
	.w7(32'h3acd0b92),
	.w8(32'hbc28800c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7886b8),
	.w1(32'h3bbf038b),
	.w2(32'hbb8195d0),
	.w3(32'h3ad05083),
	.w4(32'h3bc76819),
	.w5(32'h3a2ca922),
	.w6(32'hbbb4653f),
	.w7(32'hbb8e95ea),
	.w8(32'hbc074932),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a93a9),
	.w1(32'hbaa24663),
	.w2(32'hbb22c226),
	.w3(32'h3ae5fae8),
	.w4(32'h398010f5),
	.w5(32'h3b773804),
	.w6(32'h3adc2d6f),
	.w7(32'h3bd193c0),
	.w8(32'hbb54d402),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f146f),
	.w1(32'hbb1b3b0e),
	.w2(32'hbb83554d),
	.w3(32'h3bc9b5d4),
	.w4(32'hba80b5f6),
	.w5(32'hb9139b98),
	.w6(32'h3cb23ed2),
	.w7(32'hba152ca6),
	.w8(32'hba8cc2b4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f8088),
	.w1(32'h3b5dd10b),
	.w2(32'hbb89363a),
	.w3(32'hbbb29fc8),
	.w4(32'h3b6771b1),
	.w5(32'hbb0e6293),
	.w6(32'hbaad23a5),
	.w7(32'hbaa3e0fb),
	.w8(32'hbb921cab),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e818d),
	.w1(32'hbbbd232f),
	.w2(32'h3b0fa86d),
	.w3(32'h3b10ac0e),
	.w4(32'h3b7e31ca),
	.w5(32'hba941a19),
	.w6(32'h3b2cd9c4),
	.w7(32'h3a89a12d),
	.w8(32'h39a1ef61),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e3626),
	.w1(32'hbb1ab56e),
	.w2(32'hbb60d324),
	.w3(32'h3b3352f1),
	.w4(32'h3a7fb867),
	.w5(32'h3ae6d314),
	.w6(32'hb9893aff),
	.w7(32'h3b2b5e1d),
	.w8(32'hbaf4eb7e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea6d4),
	.w1(32'h3c1ed228),
	.w2(32'h3b70dfe5),
	.w3(32'h39f9a5f2),
	.w4(32'h3b030b55),
	.w5(32'hbbf576a2),
	.w6(32'h3b81c1cb),
	.w7(32'h3a5b5e4c),
	.w8(32'h3adcf12b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8e82),
	.w1(32'h3af68d68),
	.w2(32'hba5856ac),
	.w3(32'hbaf2f6ad),
	.w4(32'h3b3f39c2),
	.w5(32'h3bf62a97),
	.w6(32'hb9a33634),
	.w7(32'h3b52ef01),
	.w8(32'hba83df37),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2417db),
	.w1(32'h3a5a1493),
	.w2(32'hbc298246),
	.w3(32'h3a6bab12),
	.w4(32'hb984d436),
	.w5(32'hbae46521),
	.w6(32'hba816a14),
	.w7(32'h3ad4a41e),
	.w8(32'h3bab5ed5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0d879),
	.w1(32'hbc369501),
	.w2(32'h3b555a5c),
	.w3(32'hbbb64345),
	.w4(32'hbac739f3),
	.w5(32'h3cd32f6c),
	.w6(32'hb931cc2f),
	.w7(32'h3ab75ee7),
	.w8(32'hbb419881),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4f2c),
	.w1(32'h3ab16155),
	.w2(32'h3af75e77),
	.w3(32'h3ad8b1d3),
	.w4(32'hba8bff97),
	.w5(32'h3be084cd),
	.w6(32'h3a753ffc),
	.w7(32'h3bde65c9),
	.w8(32'hbb08b1c1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa072b0),
	.w1(32'hbae0b11d),
	.w2(32'h3a299887),
	.w3(32'h3b109a32),
	.w4(32'hbadb2912),
	.w5(32'h38421bac),
	.w6(32'h3c3d9a80),
	.w7(32'h3c927175),
	.w8(32'hbc6061d1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c3836),
	.w1(32'h3b8a1962),
	.w2(32'h3aceea37),
	.w3(32'h3bd8ec61),
	.w4(32'hbb7dc908),
	.w5(32'hba92cf93),
	.w6(32'hb8916b67),
	.w7(32'hb8b1e3be),
	.w8(32'hbb0ec33a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d3cc),
	.w1(32'h3ca1e64b),
	.w2(32'hbc2b250b),
	.w3(32'h3aa07808),
	.w4(32'hbacc6a0a),
	.w5(32'hba3162f6),
	.w6(32'hb8f1de07),
	.w7(32'hbadb7edf),
	.w8(32'hbb9450f2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2823f),
	.w1(32'h39fddc79),
	.w2(32'hb9fcb55e),
	.w3(32'hbb1fe21c),
	.w4(32'h3ae6562e),
	.w5(32'h3b09a217),
	.w6(32'hbaac401b),
	.w7(32'hba31ddfb),
	.w8(32'hbac49b00),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba99dd),
	.w1(32'hbac80ddc),
	.w2(32'hbc02b243),
	.w3(32'hbc1ee740),
	.w4(32'h3ac5ec99),
	.w5(32'h3aacb5d4),
	.w6(32'hba2667b4),
	.w7(32'hbabaaad0),
	.w8(32'h3ca41a13),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b43b14),
	.w1(32'h3b802bb7),
	.w2(32'h3a488ced),
	.w3(32'hbbd31e53),
	.w4(32'h3b613e72),
	.w5(32'hbb20906d),
	.w6(32'hbb4a76aa),
	.w7(32'h3a22e3f4),
	.w8(32'h3b3897c8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fbcab),
	.w1(32'h3b8c4763),
	.w2(32'h3aae4b82),
	.w3(32'h3a0f6aa6),
	.w4(32'h3b768a94),
	.w5(32'hbb095d02),
	.w6(32'hbb3b87fc),
	.w7(32'hb9d803dd),
	.w8(32'hbbf65469),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c239ec6),
	.w1(32'hba1dec86),
	.w2(32'hbb112561),
	.w3(32'hbb063161),
	.w4(32'h3b567edb),
	.w5(32'h3bae33a6),
	.w6(32'hbb03332b),
	.w7(32'hbb179870),
	.w8(32'hba80e8e3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad918b2),
	.w1(32'hb90f5bff),
	.w2(32'hbb4a9ca4),
	.w3(32'hbb3c740c),
	.w4(32'hb842e005),
	.w5(32'hba0eae6a),
	.w6(32'h3c00262b),
	.w7(32'hba983f7c),
	.w8(32'hbb2a9be6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab31259),
	.w1(32'h3b5f3c26),
	.w2(32'h38dae590),
	.w3(32'h3b7e8c4b),
	.w4(32'hbb368518),
	.w5(32'h3a3704e2),
	.w6(32'h3b4eada0),
	.w7(32'hb783f2fb),
	.w8(32'h3b99cc63),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03bfc4),
	.w1(32'hbbd2e8f2),
	.w2(32'hba2f9313),
	.w3(32'hba9dbe67),
	.w4(32'h3af04991),
	.w5(32'h3b1eb03a),
	.w6(32'hbb0e175f),
	.w7(32'hbb4f7643),
	.w8(32'hba63f95b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0be58c),
	.w1(32'h39c55f16),
	.w2(32'hbb0ee561),
	.w3(32'hbb9ccd2c),
	.w4(32'hbb912a7e),
	.w5(32'hbb939ea0),
	.w6(32'h39180ea8),
	.w7(32'h3a86b73c),
	.w8(32'hb809c8b0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e47e6),
	.w1(32'hba66530c),
	.w2(32'h3ae14b6f),
	.w3(32'h3bb3b5b9),
	.w4(32'h3a427f97),
	.w5(32'h39fac763),
	.w6(32'hbb6a6ee7),
	.w7(32'hbb9427cf),
	.w8(32'h3a6fd740),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38655a97),
	.w1(32'hb93d4d88),
	.w2(32'h3ac9a8f3),
	.w3(32'h37e01c5b),
	.w4(32'hb9cd35e0),
	.w5(32'hbbb1563e),
	.w6(32'hbb820f3e),
	.w7(32'hbaf8c746),
	.w8(32'hba4e0e80),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab64527),
	.w1(32'hb8a4499b),
	.w2(32'hbc8bf844),
	.w3(32'h3880b67e),
	.w4(32'h3b6b1026),
	.w5(32'h3adcfcae),
	.w6(32'h375b468c),
	.w7(32'hbc1e44a7),
	.w8(32'h3b7b8178),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5442cc),
	.w1(32'hbae6c8ab),
	.w2(32'hbb31449c),
	.w3(32'hba98cacf),
	.w4(32'h3a137d16),
	.w5(32'hbb085bfe),
	.w6(32'hba6bf47f),
	.w7(32'h3b3afbe5),
	.w8(32'hba81f2ea),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949aa5c),
	.w1(32'h3afcc0a8),
	.w2(32'h3b119f57),
	.w3(32'h3b5061a3),
	.w4(32'h38881151),
	.w5(32'h3b74dd05),
	.w6(32'h3a33d51f),
	.w7(32'h3b32e171),
	.w8(32'h3c053fb9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089cd5),
	.w1(32'hba85beaa),
	.w2(32'h3b231ddf),
	.w3(32'hba8ff795),
	.w4(32'hba871216),
	.w5(32'hba50350a),
	.w6(32'hbb1efbd4),
	.w7(32'hbb00d81f),
	.w8(32'hbb32115e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391037b9),
	.w1(32'hbb4f0c1a),
	.w2(32'hbb1e11f8),
	.w3(32'h3988330e),
	.w4(32'h3ac79a94),
	.w5(32'hbb4ad5a3),
	.w6(32'h3adb9587),
	.w7(32'h3bcf8c4d),
	.w8(32'hbba05f90),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72fac8),
	.w1(32'h3b3bd198),
	.w2(32'hbd639af2),
	.w3(32'hbb96320e),
	.w4(32'h3cc059c1),
	.w5(32'hbac35506),
	.w6(32'hb98157d3),
	.w7(32'hbbe2abe3),
	.w8(32'hba4ff8da),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada1536),
	.w1(32'h3a308905),
	.w2(32'h3bcad125),
	.w3(32'hba89b015),
	.w4(32'hba373fd5),
	.w5(32'h3b69bc2c),
	.w6(32'h3beb06da),
	.w7(32'h3d23e274),
	.w8(32'h3a7ad3df),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e36a),
	.w1(32'h3d3ba557),
	.w2(32'h3c4c1a6a),
	.w3(32'h3bb6ffe3),
	.w4(32'h3bc08c1f),
	.w5(32'hba80f8c2),
	.w6(32'hbac60c3c),
	.w7(32'hbb374ee6),
	.w8(32'h3bd7054a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37f3f8),
	.w1(32'hbaa77080),
	.w2(32'hbb4165d6),
	.w3(32'h3850373f),
	.w4(32'h3b32fc82),
	.w5(32'h3ceeb3d2),
	.w6(32'h3b24cb90),
	.w7(32'h3b5ff74b),
	.w8(32'h39ab23cf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd440df),
	.w1(32'hbb1b7004),
	.w2(32'h3c124e64),
	.w3(32'h3b429a96),
	.w4(32'h3acf15d0),
	.w5(32'hbc1f8108),
	.w6(32'hbbe39a20),
	.w7(32'hbbaaff8a),
	.w8(32'hbaa35b40),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052728),
	.w1(32'h3b5e9110),
	.w2(32'h3b9e852c),
	.w3(32'hbb80f75a),
	.w4(32'hbbf2d652),
	.w5(32'hbb0d4aba),
	.w6(32'h3abdd9a9),
	.w7(32'h3b81013d),
	.w8(32'hbc06dae6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2395d),
	.w1(32'h3af1ae63),
	.w2(32'hbb43bd94),
	.w3(32'h3a4f5f00),
	.w4(32'hbb98c520),
	.w5(32'h3b5ba7d7),
	.w6(32'hba79e489),
	.w7(32'h3b8ff20e),
	.w8(32'h3978f051),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fa90e),
	.w1(32'h3af7df29),
	.w2(32'h3c610ed2),
	.w3(32'h3bcce23e),
	.w4(32'h3ba0f162),
	.w5(32'h3a5e3591),
	.w6(32'h3aa18653),
	.w7(32'h3b250c68),
	.w8(32'hb78509d1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba718822),
	.w1(32'h3bc68c4a),
	.w2(32'h3bdb9914),
	.w3(32'hbcfbecc2),
	.w4(32'hbb10d8d0),
	.w5(32'h3aad416c),
	.w6(32'hbc9047be),
	.w7(32'hbbe72fa4),
	.w8(32'hbb56b8b3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee0376),
	.w1(32'h3c5f7b4d),
	.w2(32'hbd48dc1b),
	.w3(32'hbafcde36),
	.w4(32'h3c0475f7),
	.w5(32'h3b915346),
	.w6(32'hba138914),
	.w7(32'hbbd4083b),
	.w8(32'hbb5bf628),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af69999),
	.w1(32'h3baa3d90),
	.w2(32'hb92b8bab),
	.w3(32'h3b3c9d2d),
	.w4(32'h3bec6533),
	.w5(32'h3c011367),
	.w6(32'hba4b5e01),
	.w7(32'h3c097bc4),
	.w8(32'h3cd97f0d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa392),
	.w1(32'hbb6d8351),
	.w2(32'hbaf46cde),
	.w3(32'h3aec7def),
	.w4(32'h3b1b0e5b),
	.w5(32'hbc85389d),
	.w6(32'hb96f7ecd),
	.w7(32'h3a1849f4),
	.w8(32'hbafaa072),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d51dc),
	.w1(32'h3cfc5d56),
	.w2(32'h3ae1444e),
	.w3(32'h3d50bb7a),
	.w4(32'h3b9eadea),
	.w5(32'hbac3ec58),
	.w6(32'h3a637814),
	.w7(32'h3b0241fd),
	.w8(32'hb77ae727),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14de0b),
	.w1(32'h3c0d8609),
	.w2(32'hbbf130b8),
	.w3(32'hb9ccc170),
	.w4(32'h3ba1c29f),
	.w5(32'hbb5ed428),
	.w6(32'hbadd774b),
	.w7(32'h3a34813d),
	.w8(32'h3be5d758),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f974),
	.w1(32'hbd8b01ed),
	.w2(32'hba881dff),
	.w3(32'h3b5d3412),
	.w4(32'h3b3c0bb4),
	.w5(32'h3c084cdf),
	.w6(32'hba3f869e),
	.w7(32'h3c4a0abe),
	.w8(32'hbd1fb939),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c5e0b),
	.w1(32'hbae70429),
	.w2(32'h3bcfe4b8),
	.w3(32'h3aa76155),
	.w4(32'hba1b5965),
	.w5(32'hba2a8527),
	.w6(32'h3b95f635),
	.w7(32'hb98a8d9a),
	.w8(32'h3b5aa3d4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359ff8),
	.w1(32'hbb2fe469),
	.w2(32'hbab432e6),
	.w3(32'h3b7cbbe0),
	.w4(32'hbc9cdacf),
	.w5(32'h3bcffc63),
	.w6(32'h3af352d3),
	.w7(32'h3c308453),
	.w8(32'hbb6e3e67),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998d268),
	.w1(32'hbaec79de),
	.w2(32'hbd6ce1e2),
	.w3(32'hbbfb2eab),
	.w4(32'h3bff8c3f),
	.w5(32'hbb822b28),
	.w6(32'hbd5d60e1),
	.w7(32'hbbaa11c2),
	.w8(32'hbb9aeb90),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fceef),
	.w1(32'h3afad80a),
	.w2(32'h3d272448),
	.w3(32'h3cdf23a6),
	.w4(32'hbb8e1af1),
	.w5(32'hbae951e6),
	.w6(32'h37985a81),
	.w7(32'hbb837853),
	.w8(32'hbc448fed),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c32bb),
	.w1(32'hbbc5913b),
	.w2(32'h3cd83d4d),
	.w3(32'h39cfce2b),
	.w4(32'hbb8a6376),
	.w5(32'hba370926),
	.w6(32'hba00fd19),
	.w7(32'hbb41759e),
	.w8(32'hbb07d82e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd0d14),
	.w1(32'h3cf6e99e),
	.w2(32'h3bb784ab),
	.w3(32'h3c1a78a4),
	.w4(32'hba7c334c),
	.w5(32'h3b831158),
	.w6(32'hba158d19),
	.w7(32'hbbcbf186),
	.w8(32'h3acc8a3c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a755),
	.w1(32'h3ae24f8e),
	.w2(32'h3b04cc10),
	.w3(32'h3bbe0aa5),
	.w4(32'hba1c775c),
	.w5(32'h3b924643),
	.w6(32'h3ba87054),
	.w7(32'hbc36e3cd),
	.w8(32'hb9a03906),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb417e99),
	.w1(32'h3b1b547a),
	.w2(32'hbb7331ec),
	.w3(32'hbb1a73bd),
	.w4(32'h387ee6d4),
	.w5(32'h3a1e814c),
	.w6(32'hbaea4ec7),
	.w7(32'h3b0a831e),
	.w8(32'h3a0e867e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9772b5),
	.w1(32'hbbca9044),
	.w2(32'hb9fa34d2),
	.w3(32'hba18fbeb),
	.w4(32'hbaa96a73),
	.w5(32'h39cbe3c1),
	.w6(32'hbb5b77d8),
	.w7(32'h398e4030),
	.w8(32'hbb68ea22),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ddca6),
	.w1(32'hbb35b4e2),
	.w2(32'hbbfe45f1),
	.w3(32'h3cf4f448),
	.w4(32'hbb0c77a2),
	.w5(32'hbb6371ee),
	.w6(32'hba5ad430),
	.w7(32'hbb022973),
	.w8(32'hbb2fb752),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717164),
	.w1(32'h3b1d3fb1),
	.w2(32'h3bc9fdb1),
	.w3(32'hbb27e204),
	.w4(32'h3b8ba02e),
	.w5(32'hbb91dee7),
	.w6(32'hbc5f4dfe),
	.w7(32'hbb3b9de5),
	.w8(32'h3b6a87ac),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649076),
	.w1(32'h3b540887),
	.w2(32'h3bcf5c8d),
	.w3(32'hbb998224),
	.w4(32'h39688dcd),
	.w5(32'h3b8f052f),
	.w6(32'hbc3b0c0c),
	.w7(32'hbb387974),
	.w8(32'h39dbff1c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c181a11),
	.w1(32'hbc11a40a),
	.w2(32'hbb85e5e4),
	.w3(32'hb9bdbdf5),
	.w4(32'hbb433466),
	.w5(32'hbb23ea08),
	.w6(32'hbb9e202f),
	.w7(32'hbb071252),
	.w8(32'h3b98de05),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe79980),
	.w1(32'hbb4918a4),
	.w2(32'hbc4cfbe0),
	.w3(32'hbb8d0172),
	.w4(32'h3ab4227e),
	.w5(32'hbaa5dc29),
	.w6(32'h3b9960bd),
	.w7(32'hb9ff0093),
	.w8(32'h3d8e557f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9797e),
	.w1(32'hbb1ccee1),
	.w2(32'h3a01e5b4),
	.w3(32'hbc8633e1),
	.w4(32'hbbb0d62c),
	.w5(32'hbbab340a),
	.w6(32'hbc109d5b),
	.w7(32'h39b243c7),
	.w8(32'hbb4316eb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa769bc),
	.w1(32'h3aa60e17),
	.w2(32'h3b16b125),
	.w3(32'hbb4392c0),
	.w4(32'hbb36ca21),
	.w5(32'h3a9b77c6),
	.w6(32'hbb34dbf3),
	.w7(32'h3bf173e5),
	.w8(32'hbb56adba),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a140f82),
	.w1(32'h3c289953),
	.w2(32'hb8c1dcba),
	.w3(32'hbc018ea1),
	.w4(32'hbbcc0fa8),
	.w5(32'hbbc6b7ca),
	.w6(32'hbc1bafaa),
	.w7(32'h3bb637e1),
	.w8(32'h3b4aa733),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5c9de),
	.w1(32'hbb827269),
	.w2(32'h3abb9c43),
	.w3(32'h3aefc3fe),
	.w4(32'h3a6108ab),
	.w5(32'h3a89dc16),
	.w6(32'h3b982a3a),
	.w7(32'h3b934b5f),
	.w8(32'hb9a87392),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb212ce),
	.w1(32'hbbf21d57),
	.w2(32'h394d28c8),
	.w3(32'hbb62ddf6),
	.w4(32'h3a83474c),
	.w5(32'h3c0261b1),
	.w6(32'h3b16656c),
	.w7(32'hbaa9580a),
	.w8(32'h3b36abd4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d6975),
	.w1(32'h3b2d1665),
	.w2(32'h3cb400a3),
	.w3(32'h39326d6f),
	.w4(32'h3be63b04),
	.w5(32'h3b459647),
	.w6(32'h3ae1e3f6),
	.w7(32'hbace113f),
	.w8(32'h3ac537d4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d1f11),
	.w1(32'hbc0b74dc),
	.w2(32'h3acbbb15),
	.w3(32'hbb60d36b),
	.w4(32'h3b08b1ad),
	.w5(32'h3a078413),
	.w6(32'hbc2a4afc),
	.w7(32'h3bf07053),
	.w8(32'h3bd3d665),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e25fd),
	.w1(32'h3a83b34e),
	.w2(32'h3c84d3fd),
	.w3(32'hbb9823cc),
	.w4(32'h3c5cf3ea),
	.w5(32'hbb8b6d7c),
	.w6(32'hbcfae40e),
	.w7(32'hbd896d67),
	.w8(32'h3abbdc2f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24bb7f),
	.w1(32'h3b3f9c92),
	.w2(32'hbb7eaeb8),
	.w3(32'hbba35076),
	.w4(32'hbb0fbf01),
	.w5(32'h3bf750b2),
	.w6(32'hbb27ed6c),
	.w7(32'h3acd42b1),
	.w8(32'hb9d550b4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f395),
	.w1(32'h376c3559),
	.w2(32'h398cddfe),
	.w3(32'hbd1dabc3),
	.w4(32'h3b7983d4),
	.w5(32'hbd1bf638),
	.w6(32'hba6c0f9f),
	.w7(32'hbc26c729),
	.w8(32'hbb6f8d43),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b89d0),
	.w1(32'h3cd7b0b9),
	.w2(32'h3a33ec26),
	.w3(32'hb5476de1),
	.w4(32'hbc040d01),
	.w5(32'h3c3ab41e),
	.w6(32'hbbace8ea),
	.w7(32'h3996991c),
	.w8(32'hbb80e91e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aae4f),
	.w1(32'hbb5a199a),
	.w2(32'hbaf3b7bc),
	.w3(32'hbc1502e9),
	.w4(32'h3aa6308d),
	.w5(32'hb9f85d8c),
	.w6(32'h3c785829),
	.w7(32'hbb9e12e2),
	.w8(32'h3bb89d62),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb1bb7),
	.w1(32'h350c5572),
	.w2(32'h3bdb7ba2),
	.w3(32'hbad11f4c),
	.w4(32'hbcf59769),
	.w5(32'h3bcd41f8),
	.w6(32'hbd031743),
	.w7(32'hb9ad082f),
	.w8(32'hba00965a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79236c),
	.w1(32'h3aab26d1),
	.w2(32'h3b47d31d),
	.w3(32'hbb7333ba),
	.w4(32'h3b646124),
	.w5(32'hbcd976e8),
	.w6(32'hbad6531f),
	.w7(32'hbc43d54c),
	.w8(32'hbb895982),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3573f5),
	.w1(32'h3b4cc277),
	.w2(32'h3b10aa2d),
	.w3(32'hbc2dc903),
	.w4(32'h3b0c2aed),
	.w5(32'hbb1fbb09),
	.w6(32'h3d0fd67a),
	.w7(32'hbab08554),
	.w8(32'hbac27682),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf02b8),
	.w1(32'hbb880b2f),
	.w2(32'hbc8aa108),
	.w3(32'hbb210310),
	.w4(32'hbc089512),
	.w5(32'hbbcac203),
	.w6(32'hbb186601),
	.w7(32'h3bad48b9),
	.w8(32'hbd821902),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90cfce),
	.w1(32'h3a6d421d),
	.w2(32'hbc1451ca),
	.w3(32'h3a3d236b),
	.w4(32'hba83a3cd),
	.w5(32'hb83bb9ea),
	.w6(32'hbab64061),
	.w7(32'h3a0a94c8),
	.w8(32'h3beea6f7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6b87b),
	.w1(32'hbb9924b4),
	.w2(32'h3b05de1c),
	.w3(32'hbcd1103b),
	.w4(32'h3b4fb450),
	.w5(32'h3a1ec1c9),
	.w6(32'hb8d41052),
	.w7(32'h3cf0b6c4),
	.w8(32'hbc342d54),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b7e02),
	.w1(32'h3c8a811f),
	.w2(32'hb782d8e7),
	.w3(32'hbc413dbd),
	.w4(32'h3b21a295),
	.w5(32'h3a8e1c13),
	.w6(32'hbb558e15),
	.w7(32'hba63f494),
	.w8(32'h3b4e1b13),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143885),
	.w1(32'h3b3f1161),
	.w2(32'hbb9ae0c4),
	.w3(32'hbcee6c29),
	.w4(32'hbabd474f),
	.w5(32'hbc4895f1),
	.w6(32'h3b79374a),
	.w7(32'hbcab53b8),
	.w8(32'h3b4ac9d9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e74b5),
	.w1(32'h3b344497),
	.w2(32'hbb2a89a0),
	.w3(32'hba868f57),
	.w4(32'hbac23853),
	.w5(32'hb9be0de4),
	.w6(32'hbccd197c),
	.w7(32'hba038a7d),
	.w8(32'h3bbca1e7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd22152c),
	.w1(32'hbc2641ff),
	.w2(32'hbbd5c9a2),
	.w3(32'hbb1e7fdf),
	.w4(32'hbc840f96),
	.w5(32'h3c950fe5),
	.w6(32'hbb472ab5),
	.w7(32'hba416b2f),
	.w8(32'hbb9198af),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c56d),
	.w1(32'h377a49d8),
	.w2(32'hbc1307dc),
	.w3(32'h3b895a4b),
	.w4(32'h3a6e9d59),
	.w5(32'hba8cc2e8),
	.w6(32'hbb7f147a),
	.w7(32'h3b039212),
	.w8(32'h3b230523),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3070c0),
	.w1(32'hbb20c105),
	.w2(32'hbc0929d6),
	.w3(32'hb8e829f3),
	.w4(32'h3d6e4fb3),
	.w5(32'hbb16cbe2),
	.w6(32'hbb4ded50),
	.w7(32'h3a9e9c5d),
	.w8(32'hbb9d0789),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6359f),
	.w1(32'hbc29a16e),
	.w2(32'h3b8502c4),
	.w3(32'hbb53f39c),
	.w4(32'h3b96c157),
	.w5(32'hbb191872),
	.w6(32'hbb38ba0a),
	.w7(32'hbb710e90),
	.w8(32'h3b01504d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bef13),
	.w1(32'h3a95fc17),
	.w2(32'h3b6dc2f5),
	.w3(32'h3a20717f),
	.w4(32'h3ae2e107),
	.w5(32'h3c83cf2e),
	.w6(32'hbb9319f3),
	.w7(32'hbb91d41d),
	.w8(32'hbb56d2c3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55cca1),
	.w1(32'h3a6dfc4a),
	.w2(32'hbae03604),
	.w3(32'h3aac2968),
	.w4(32'h3b5338cf),
	.w5(32'hbc104711),
	.w6(32'h3b65fdf3),
	.w7(32'h3b4b4174),
	.w8(32'hba10e27e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889cb6e),
	.w1(32'h3b06ee6e),
	.w2(32'h3bbdfd23),
	.w3(32'hbb1389cf),
	.w4(32'h3b2bef04),
	.w5(32'h3b4fbf28),
	.w6(32'h3a99c158),
	.w7(32'hbae87c8f),
	.w8(32'h39d23124),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b97dd),
	.w1(32'h3d3a3b0d),
	.w2(32'hbbf0b102),
	.w3(32'hbc40d6e6),
	.w4(32'h3ba6e5c4),
	.w5(32'hbb211caf),
	.w6(32'hbc014767),
	.w7(32'hbc76fcc7),
	.w8(32'hbbece3c7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d304c4),
	.w1(32'hbb890b63),
	.w2(32'h3b41319f),
	.w3(32'h3adf25c7),
	.w4(32'h3a7537f4),
	.w5(32'h3b40fba1),
	.w6(32'hb9a36bf7),
	.w7(32'hb7b7aa4a),
	.w8(32'h3b351876),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6565),
	.w1(32'h3ad1ba36),
	.w2(32'h3a998b8d),
	.w3(32'h3bff94fd),
	.w4(32'h3b77d4bb),
	.w5(32'h39ce96ba),
	.w6(32'h3cb8ea32),
	.w7(32'hbb42556f),
	.w8(32'hbb435f16),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d912b),
	.w1(32'hbabf486c),
	.w2(32'h3c11caaa),
	.w3(32'hbab960e6),
	.w4(32'h3c8f1a0e),
	.w5(32'h3bad058f),
	.w6(32'hb9f5bcd8),
	.w7(32'h3a07ee06),
	.w8(32'h3c7be0d0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e0a60),
	.w1(32'h3b65c2f8),
	.w2(32'h3c0595cb),
	.w3(32'h3a8d5614),
	.w4(32'hba9e2835),
	.w5(32'hbb9cc260),
	.w6(32'h3b46cd46),
	.w7(32'h3c114298),
	.w8(32'hbb212529),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e10eb),
	.w1(32'hbbd0b072),
	.w2(32'h3bb3c63b),
	.w3(32'h3b6c7c2d),
	.w4(32'h3bf44e60),
	.w5(32'hba3ae2f2),
	.w6(32'hba7af4df),
	.w7(32'hb9014066),
	.w8(32'hbb3df131),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b822c),
	.w1(32'hbaf919d8),
	.w2(32'hbb909402),
	.w3(32'hbc62168f),
	.w4(32'hbbc7e421),
	.w5(32'hbbd050e9),
	.w6(32'hbbf79ce3),
	.w7(32'hbbab1068),
	.w8(32'h3b7e7fb7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb884c93),
	.w1(32'h39ab4ad6),
	.w2(32'h3c7d3f00),
	.w3(32'h3b66cd9e),
	.w4(32'hbbb6dabb),
	.w5(32'h3a8af327),
	.w6(32'h3b06e225),
	.w7(32'hba93d543),
	.w8(32'hbbbfc1ed),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfcac8a),
	.w1(32'h3b91c623),
	.w2(32'hbbb0fa82),
	.w3(32'h3c827759),
	.w4(32'hb9122843),
	.w5(32'hbc210048),
	.w6(32'hbc26017c),
	.w7(32'hba661f98),
	.w8(32'hbb7aced8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b03f4),
	.w1(32'hb9fb510b),
	.w2(32'h3ab5b4ea),
	.w3(32'hbb34967a),
	.w4(32'h3b0e715c),
	.w5(32'hbacc9aaf),
	.w6(32'h3c143811),
	.w7(32'hbcd8fcdc),
	.w8(32'hbc5bf4f4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868e0a),
	.w1(32'hbb5b1b26),
	.w2(32'h39d91781),
	.w3(32'hba56fa6c),
	.w4(32'h3ba2505e),
	.w5(32'h3c3da930),
	.w6(32'hbd3ee240),
	.w7(32'hba7b5553),
	.w8(32'h3c12abd3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a7e87),
	.w1(32'hbbaddde0),
	.w2(32'h3c1bc421),
	.w3(32'hbadb4478),
	.w4(32'hbb0d4442),
	.w5(32'hbac0cbf8),
	.w6(32'hbbaea30c),
	.w7(32'hbb0b7546),
	.w8(32'h3afbab92),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb30b4),
	.w1(32'h39e2e067),
	.w2(32'hbc819c17),
	.w3(32'hbab7f194),
	.w4(32'hb80b833a),
	.w5(32'h3ae1bd67),
	.w6(32'h3c1b9599),
	.w7(32'hbab9ce92),
	.w8(32'hbc968d66),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8cd6d),
	.w1(32'hbaaa3e4a),
	.w2(32'h3a1e39f2),
	.w3(32'hbb8c41e1),
	.w4(32'hbb65b3f7),
	.w5(32'h3b8eeaaf),
	.w6(32'hbc245deb),
	.w7(32'h3ae694fe),
	.w8(32'h3b1b331f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb28e1a),
	.w1(32'hbad8b3e6),
	.w2(32'h3d13d870),
	.w3(32'hba0b05c1),
	.w4(32'h3c2aa74c),
	.w5(32'hbc187d6b),
	.w6(32'hbce08ec9),
	.w7(32'hbc1ed9e9),
	.w8(32'hbc01b67c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61e1d8),
	.w1(32'hbb08291e),
	.w2(32'h3bf1f56d),
	.w3(32'hbb567a5c),
	.w4(32'h3b18f65e),
	.w5(32'hbb1ee69e),
	.w6(32'h3b92fd7b),
	.w7(32'h3aca9b93),
	.w8(32'h3bea1e30),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bab45),
	.w1(32'hbc62023e),
	.w2(32'h3a260a05),
	.w3(32'hbb8f68c5),
	.w4(32'h3b21bed1),
	.w5(32'h393320a7),
	.w6(32'h3b4e51f8),
	.w7(32'hba2d20dd),
	.w8(32'h3adce977),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3f5d6),
	.w1(32'hb95c86b5),
	.w2(32'h38811adb),
	.w3(32'hbcdbefe5),
	.w4(32'hba72820a),
	.w5(32'hbb5d54bd),
	.w6(32'hbb892304),
	.w7(32'hbca24807),
	.w8(32'h3b9829bd),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62063c),
	.w1(32'hbb460f46),
	.w2(32'h3b2b2902),
	.w3(32'hbb7fcbe7),
	.w4(32'h3bf8881c),
	.w5(32'hbd11144a),
	.w6(32'hb9ea6338),
	.w7(32'h3c9c419d),
	.w8(32'h3c8145c6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99dfb7),
	.w1(32'h3bc0458d),
	.w2(32'hbbbc8244),
	.w3(32'hbabdff53),
	.w4(32'h3b33a2b4),
	.w5(32'h37e702f3),
	.w6(32'hbbc5f580),
	.w7(32'hbbd88b7e),
	.w8(32'h3ac99817),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1e0fd),
	.w1(32'h3808d656),
	.w2(32'h3c4ccf86),
	.w3(32'hba0bf9e0),
	.w4(32'hb9e9036c),
	.w5(32'h3ba2ef6f),
	.w6(32'hbb8715c7),
	.w7(32'h3b18c964),
	.w8(32'hbb37a9cd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13322d),
	.w1(32'h3addcadc),
	.w2(32'h3b37ec1d),
	.w3(32'hbacebebe),
	.w4(32'hbc186719),
	.w5(32'hbc04e501),
	.w6(32'hbbec9e0e),
	.w7(32'hbb980aa3),
	.w8(32'h3c5d9e50),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2c52),
	.w1(32'h39d586e0),
	.w2(32'hbb3c1a00),
	.w3(32'h3be3a0d1),
	.w4(32'hbb30f415),
	.w5(32'h39e799e4),
	.w6(32'h3a7c5fe6),
	.w7(32'h3ab5b63b),
	.w8(32'hb9bca72b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6af98e),
	.w1(32'hbb12988f),
	.w2(32'hbb59141e),
	.w3(32'h3b07636a),
	.w4(32'hbb0ae9e0),
	.w5(32'h3acb0760),
	.w6(32'hba35c130),
	.w7(32'h3a8eda3a),
	.w8(32'hbc376210),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aa0d6),
	.w1(32'h3aa1d16c),
	.w2(32'h3be1d990),
	.w3(32'hbc2efab9),
	.w4(32'hbac37b35),
	.w5(32'hbb4cb925),
	.w6(32'hbb0f71f7),
	.w7(32'h3ba07b58),
	.w8(32'h3b6e0f74),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1bcb),
	.w1(32'hbafc5716),
	.w2(32'hbbcfcb17),
	.w3(32'hba6bdd1d),
	.w4(32'h3bed6cb7),
	.w5(32'h3b55cc27),
	.w6(32'hba91d51d),
	.w7(32'hbbf9b4fd),
	.w8(32'hbb4eda49),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1043bb),
	.w1(32'h3af3e9ef),
	.w2(32'hbb69ef7b),
	.w3(32'h397ed0e7),
	.w4(32'h3b71c3a0),
	.w5(32'h3a3b3646),
	.w6(32'hbb9feec6),
	.w7(32'h3b41afb5),
	.w8(32'hb9ebb88f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef9440),
	.w1(32'h3b7390e2),
	.w2(32'h3b1e3ced),
	.w3(32'hbb5d8aca),
	.w4(32'h3af0ee8f),
	.w5(32'hb8aa2887),
	.w6(32'hbb1804bf),
	.w7(32'hbb6408bb),
	.w8(32'hbca02b12),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf731c),
	.w1(32'hbbb3f769),
	.w2(32'hbc8247af),
	.w3(32'hbc4e1f58),
	.w4(32'hbc098d72),
	.w5(32'hbc1558a0),
	.w6(32'h3c1ae32f),
	.w7(32'hbad85435),
	.w8(32'h3c10b8a6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8590e3),
	.w1(32'hbb5f350f),
	.w2(32'h3b6e7df1),
	.w3(32'hbbc3483f),
	.w4(32'h3b85583f),
	.w5(32'hbba0bc09),
	.w6(32'hbbef5f27),
	.w7(32'hb95e1592),
	.w8(32'h3b215a98),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf31f),
	.w1(32'h3c2315d7),
	.w2(32'h3c24c9c6),
	.w3(32'h3b9f4c82),
	.w4(32'h3c9d7b75),
	.w5(32'hbba7a108),
	.w6(32'hbb90378f),
	.w7(32'h3bc8f602),
	.w8(32'hbb9eef61),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e107),
	.w1(32'hba4e30b3),
	.w2(32'hbbab88aa),
	.w3(32'h3af86831),
	.w4(32'hba43acff),
	.w5(32'hb9f0fa4d),
	.w6(32'h3b217d52),
	.w7(32'hbbbc45ad),
	.w8(32'hbd81300e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40c7f6),
	.w1(32'h3c36b0ef),
	.w2(32'h3b43aae3),
	.w3(32'h3cae43cc),
	.w4(32'h3b7be090),
	.w5(32'hbd0af6ec),
	.w6(32'hbc287efd),
	.w7(32'hbc29afb0),
	.w8(32'hbbdf2767),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c9876),
	.w1(32'h3b8cbc65),
	.w2(32'hb97d846a),
	.w3(32'hbc20c608),
	.w4(32'hbb4f67a6),
	.w5(32'hbb49bdac),
	.w6(32'hbc2b2f88),
	.w7(32'hbba58b65),
	.w8(32'h3b2bfc64),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf039d),
	.w1(32'h3b364570),
	.w2(32'hba9ed9e0),
	.w3(32'h3a574d2f),
	.w4(32'h3a32f19f),
	.w5(32'h3ad8eac9),
	.w6(32'h3b89d710),
	.w7(32'hbcd403e8),
	.w8(32'hbb85244b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c6805),
	.w1(32'hbc384eb6),
	.w2(32'hbbded637),
	.w3(32'hbb66d6c3),
	.w4(32'h3c32919d),
	.w5(32'hbbd111e6),
	.w6(32'h3aee3fdc),
	.w7(32'hbb908962),
	.w8(32'hba8a0329),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb916b5b),
	.w1(32'hbae82b03),
	.w2(32'hbaa0fdde),
	.w3(32'h3bb174a5),
	.w4(32'h3902a453),
	.w5(32'hbb229b02),
	.w6(32'hbb4b9a52),
	.w7(32'h3b5e41b9),
	.w8(32'hbca8d97f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46e931),
	.w1(32'hbb8f1207),
	.w2(32'hbb3aa57d),
	.w3(32'hba4f3a9e),
	.w4(32'h3b38f04e),
	.w5(32'hbbb1c803),
	.w6(32'h3bb7affb),
	.w7(32'hbc237f7b),
	.w8(32'h37d84887),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea319a),
	.w1(32'hbc80a696),
	.w2(32'h3d51946c),
	.w3(32'hbad64646),
	.w4(32'hba5f1be2),
	.w5(32'h3bb6faee),
	.w6(32'hbb744e99),
	.w7(32'h38731784),
	.w8(32'hbc2150b3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9610e69),
	.w1(32'hbb934939),
	.w2(32'h3b6629fe),
	.w3(32'h3be8f73a),
	.w4(32'hbbe5fbe0),
	.w5(32'hbc7e0d9d),
	.w6(32'hbaca4d93),
	.w7(32'h3a88543e),
	.w8(32'h3b4c032d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1182e1),
	.w1(32'h3b39a7c8),
	.w2(32'hbb42ab57),
	.w3(32'hba426796),
	.w4(32'h39da7f9e),
	.w5(32'hbb6e3b4c),
	.w6(32'h3ae9aeb4),
	.w7(32'h3abd79ce),
	.w8(32'hbbbe2dca),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57b0d7),
	.w1(32'h3d171e01),
	.w2(32'hbb9ca98d),
	.w3(32'h3c4cbbaa),
	.w4(32'hb8951ade),
	.w5(32'hbc110fe5),
	.w6(32'hb8b39a90),
	.w7(32'h3b88436e),
	.w8(32'h3cb61fbe),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba755db),
	.w1(32'hbb44ea93),
	.w2(32'h3bdb546a),
	.w3(32'hbbc3320c),
	.w4(32'h3c31257b),
	.w5(32'hba468b4b),
	.w6(32'hbc13b9a9),
	.w7(32'hbc156026),
	.w8(32'h3bab71e7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd48083),
	.w1(32'hbb0346ca),
	.w2(32'hbcb2e19e),
	.w3(32'hbd6878a1),
	.w4(32'h3a9e4a3f),
	.w5(32'hb73b5f3c),
	.w6(32'h3bafafc3),
	.w7(32'hbc4e552c),
	.w8(32'hbc75ff05),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9799ee),
	.w1(32'h3a6faa9e),
	.w2(32'h3b955897),
	.w3(32'h3a1bb1bf),
	.w4(32'hba018e52),
	.w5(32'hbb9b6ce8),
	.w6(32'hbbd17d72),
	.w7(32'hbb558b6d),
	.w8(32'hbbc4f755),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f5690),
	.w1(32'hbb47fab4),
	.w2(32'hbb56220a),
	.w3(32'h3acc8bac),
	.w4(32'hbaab5ff6),
	.w5(32'h390c3bd3),
	.w6(32'hbb1b3c48),
	.w7(32'h3c54beab),
	.w8(32'hbbaa7250),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb48766),
	.w1(32'hbc04fdea),
	.w2(32'hbc436197),
	.w3(32'hbae01ed5),
	.w4(32'hbb71ce03),
	.w5(32'hbc4807a7),
	.w6(32'hbbf778cf),
	.w7(32'h3b2e60dc),
	.w8(32'hbc4aca8a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7548fb),
	.w1(32'hbc4d974e),
	.w2(32'hbb98b9b5),
	.w3(32'hbc18de76),
	.w4(32'h3a23f559),
	.w5(32'hbbbbfe3e),
	.w6(32'hbc7c22cf),
	.w7(32'hbb4f9b14),
	.w8(32'h3b747f7e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ee00a),
	.w1(32'h3b471c59),
	.w2(32'hbac44b99),
	.w3(32'hbb9e52c3),
	.w4(32'hbc5a3378),
	.w5(32'hbbce85e4),
	.w6(32'hbacff19b),
	.w7(32'hbaa8fdfe),
	.w8(32'hbbd01b5d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034218),
	.w1(32'hbb5f5b2c),
	.w2(32'h3b92b6d1),
	.w3(32'h3700075d),
	.w4(32'h3c097e3e),
	.w5(32'hbbb845d8),
	.w6(32'h3b030e46),
	.w7(32'hbb3cdfff),
	.w8(32'hbbe0d110),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb517363),
	.w1(32'hbbaa05cf),
	.w2(32'hbcaf3592),
	.w3(32'h3b7e2cac),
	.w4(32'hba02d771),
	.w5(32'h3b3eaa81),
	.w6(32'hbc8e996f),
	.w7(32'h3bb886ba),
	.w8(32'hbb4f7863),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06a801),
	.w1(32'h3a2f7519),
	.w2(32'hbbc56364),
	.w3(32'hbb3dca31),
	.w4(32'hbb2db731),
	.w5(32'h3a23a333),
	.w6(32'h39124fa2),
	.w7(32'hbbbf7e57),
	.w8(32'h3a5409a2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e30d0),
	.w1(32'h3c7a6857),
	.w2(32'hbbb06224),
	.w3(32'hbbe97365),
	.w4(32'h3c8f8df3),
	.w5(32'h3b349a18),
	.w6(32'hbba82a8c),
	.w7(32'hbc4076e4),
	.w8(32'h3bbfa445),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9f69),
	.w1(32'hbb04c6df),
	.w2(32'hbbf24e22),
	.w3(32'h3c48704b),
	.w4(32'h3bad184d),
	.w5(32'h3c06a0b1),
	.w6(32'hbbb5ba2e),
	.w7(32'hbaef1368),
	.w8(32'h3a08028a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c9b5),
	.w1(32'hbb7eac81),
	.w2(32'hbcafd4ce),
	.w3(32'hbb88b467),
	.w4(32'h3be68034),
	.w5(32'hbbd30cba),
	.w6(32'h3bd9627a),
	.w7(32'h3b95ca56),
	.w8(32'h3b0a32ab),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb478866),
	.w1(32'h3c5a980b),
	.w2(32'hbb842fc9),
	.w3(32'hbc8cff41),
	.w4(32'h3b84e1b1),
	.w5(32'h3b8b9f80),
	.w6(32'hbb1be34d),
	.w7(32'hbc122a7f),
	.w8(32'hbc3b0fe2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba457fdd),
	.w1(32'hbb5f64bb),
	.w2(32'h3b999c6c),
	.w3(32'hbbff1fc1),
	.w4(32'h3819aec6),
	.w5(32'hbbf16d31),
	.w6(32'h3b261670),
	.w7(32'h3a2d8069),
	.w8(32'hbbc11272),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76cda5),
	.w1(32'hbbd3210f),
	.w2(32'hbbd09c22),
	.w3(32'h3c100776),
	.w4(32'h3b87c1aa),
	.w5(32'h3c2e21d7),
	.w6(32'hbb70ca0a),
	.w7(32'hba665c9e),
	.w8(32'h3c17b5c6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38a8e6),
	.w1(32'h3bc262ad),
	.w2(32'hb9d288f3),
	.w3(32'hbb36d214),
	.w4(32'h3b520f07),
	.w5(32'hbbfe2b4b),
	.w6(32'hbb32d10d),
	.w7(32'hbbc0d298),
	.w8(32'hba407ee9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ca776),
	.w1(32'h3b231bff),
	.w2(32'h3b8c9e0c),
	.w3(32'hbbe4d08d),
	.w4(32'hbaa4ebe8),
	.w5(32'hba37728e),
	.w6(32'hbaacbc7f),
	.w7(32'h3bebf626),
	.w8(32'hbb931dea),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93fb45),
	.w1(32'hbba7c439),
	.w2(32'hbbb9650a),
	.w3(32'hbb0de2f7),
	.w4(32'h3bb4ab73),
	.w5(32'hbbfa08b1),
	.w6(32'h3c276258),
	.w7(32'h3a3245aa),
	.w8(32'h3b8677a1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8104fb),
	.w1(32'hbc04539c),
	.w2(32'hba9f018c),
	.w3(32'h3b23a958),
	.w4(32'hb89ef3e3),
	.w5(32'hbbd89a2b),
	.w6(32'h3ae1bcc5),
	.w7(32'hbc260973),
	.w8(32'hbba626cd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a570c38),
	.w1(32'hbb8923e7),
	.w2(32'h3bc374b6),
	.w3(32'h39cf4111),
	.w4(32'hbba691e0),
	.w5(32'hbc1eadcb),
	.w6(32'h3a0e3fa9),
	.w7(32'h3b237c2f),
	.w8(32'h3b227444),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe94a3),
	.w1(32'h3c0d97a8),
	.w2(32'hbb94a0d9),
	.w3(32'hbbe4d5e8),
	.w4(32'h3a5d1dbf),
	.w5(32'h3aa464fc),
	.w6(32'hbb99e1ad),
	.w7(32'hba02c710),
	.w8(32'hbb6c4f4c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3546c5),
	.w1(32'h3c382288),
	.w2(32'h3bb40c5a),
	.w3(32'h3b8c71d3),
	.w4(32'h3aa5b802),
	.w5(32'h3bc42863),
	.w6(32'hb8d731da),
	.w7(32'h3c05c273),
	.w8(32'h3b0293ca),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af35fcf),
	.w1(32'hbbe8e868),
	.w2(32'hbacd7fe7),
	.w3(32'h3c751105),
	.w4(32'hbc4d8f3a),
	.w5(32'h3cba7842),
	.w6(32'h3be91584),
	.w7(32'hbc08fdc8),
	.w8(32'hba8b32c9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc22ab),
	.w1(32'hbb59ae73),
	.w2(32'h3c196b9f),
	.w3(32'hbb05d7d6),
	.w4(32'h3bb3b180),
	.w5(32'h3bd1d325),
	.w6(32'h3a096660),
	.w7(32'h3bd539a3),
	.w8(32'h3814523d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4af6b),
	.w1(32'hbba349da),
	.w2(32'h3b83a0d8),
	.w3(32'hbb904951),
	.w4(32'hba92ccbb),
	.w5(32'hbb9cf070),
	.w6(32'h3b09a13b),
	.w7(32'h3afcee45),
	.w8(32'hbbae8525),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab5f37),
	.w1(32'hbbbf3861),
	.w2(32'hbb865d00),
	.w3(32'hbb98bd36),
	.w4(32'h39d8a8c2),
	.w5(32'hbc22d315),
	.w6(32'h3c97548f),
	.w7(32'h3bce6750),
	.w8(32'hba5d5f6a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74bd8a),
	.w1(32'h3c2cb823),
	.w2(32'h36e7368d),
	.w3(32'hba802eaf),
	.w4(32'h3b75349b),
	.w5(32'h3c1c4154),
	.w6(32'hbbd12f24),
	.w7(32'h3a680a8d),
	.w8(32'hb8c52325),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58839e),
	.w1(32'h3ab28169),
	.w2(32'hbb549807),
	.w3(32'hbbe0ee27),
	.w4(32'hba566e82),
	.w5(32'hbc2436c3),
	.w6(32'h3c6ac381),
	.w7(32'hbb8ce8d1),
	.w8(32'hbb986fae),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39881109),
	.w1(32'hbc07d89a),
	.w2(32'h39a73d44),
	.w3(32'hbb8cfb1e),
	.w4(32'h3bd6e6a7),
	.w5(32'h3c2134d2),
	.w6(32'hbb8b5e9c),
	.w7(32'hbaa23013),
	.w8(32'hbb12e2db),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64945),
	.w1(32'hbba9a760),
	.w2(32'hbbf31b82),
	.w3(32'hbb8e8a28),
	.w4(32'hbaabeb34),
	.w5(32'h3bdb8abc),
	.w6(32'hbc65eba0),
	.w7(32'hbab7ee06),
	.w8(32'hbc0ed153),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03bd19),
	.w1(32'h3b58edc8),
	.w2(32'h3a38eaca),
	.w3(32'hbb9bf1ef),
	.w4(32'hba87dcc7),
	.w5(32'hbaf4a777),
	.w6(32'hbb497417),
	.w7(32'h3be47680),
	.w8(32'hba02e281),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7cef6),
	.w1(32'h3984be9f),
	.w2(32'h3b63e90e),
	.w3(32'h3b9a19a2),
	.w4(32'h3b13c300),
	.w5(32'h3b8591ac),
	.w6(32'hbba0e8f1),
	.w7(32'h39246c5f),
	.w8(32'h3b49e6e8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dc4ff),
	.w1(32'hbc1b2e72),
	.w2(32'h3a8b40e3),
	.w3(32'hbb90b69b),
	.w4(32'h3b8e1332),
	.w5(32'h3b619101),
	.w6(32'h3bad7a33),
	.w7(32'h3b29d183),
	.w8(32'hba53f3d8),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cca25),
	.w1(32'h3b217e19),
	.w2(32'h3be7dad8),
	.w3(32'h3c8fcc08),
	.w4(32'h3be15059),
	.w5(32'h3c0339bd),
	.w6(32'hb8b569cb),
	.w7(32'h3cb4387b),
	.w8(32'hbbc9a0db),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3601ab),
	.w1(32'hbb79fded),
	.w2(32'hbc959058),
	.w3(32'h3acaa559),
	.w4(32'h3a9d4456),
	.w5(32'hbc443c7c),
	.w6(32'h3b10c536),
	.w7(32'hbc856f38),
	.w8(32'hbbfbebac),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69809b),
	.w1(32'h397d9def),
	.w2(32'hbb7c0413),
	.w3(32'h3b49551f),
	.w4(32'hbbd10359),
	.w5(32'hbaeea2ff),
	.w6(32'hba8c1e36),
	.w7(32'hbbc4f2b9),
	.w8(32'h3a432827),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5caa),
	.w1(32'hbb0015f5),
	.w2(32'h39572273),
	.w3(32'h3b8bffe3),
	.w4(32'hbaef37a0),
	.w5(32'hbbdd425b),
	.w6(32'hb91d4135),
	.w7(32'h3b64d38d),
	.w8(32'hbb678b36),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcee5b6),
	.w1(32'h3bff6870),
	.w2(32'hba032dae),
	.w3(32'h3a8ae457),
	.w4(32'h38c3013f),
	.w5(32'h3b764242),
	.w6(32'h3bcc737e),
	.w7(32'hbb275d7a),
	.w8(32'h3c559690),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc87c7b),
	.w1(32'hbc2f9620),
	.w2(32'h3c6f508c),
	.w3(32'h3c1edb50),
	.w4(32'h3c7896a0),
	.w5(32'hbc76c8d3),
	.w6(32'hbbbeeb88),
	.w7(32'hbbd0fe57),
	.w8(32'hbc161743),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59974c),
	.w1(32'hbbb53c59),
	.w2(32'hbbdff7ab),
	.w3(32'hbb7b3598),
	.w4(32'h39f99ce5),
	.w5(32'h3cbbdc0f),
	.w6(32'h3c278aa9),
	.w7(32'h389677ad),
	.w8(32'hbb635ce4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ece6c),
	.w1(32'h3a76c669),
	.w2(32'h3c388420),
	.w3(32'hbb8d60f6),
	.w4(32'hbc23f1d2),
	.w5(32'h3c1dd8c4),
	.w6(32'hbb228f8c),
	.w7(32'h3c0dd772),
	.w8(32'hbb6327cb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92daeb3),
	.w1(32'hbc2047b4),
	.w2(32'hbb088d22),
	.w3(32'h3c8bd161),
	.w4(32'h3c091129),
	.w5(32'h3936c90f),
	.w6(32'hba4c1ab7),
	.w7(32'h3a9d56eb),
	.w8(32'h3b226108),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5c17f),
	.w1(32'hbb076308),
	.w2(32'hba99aedd),
	.w3(32'h3a9bf815),
	.w4(32'h3af49653),
	.w5(32'h3b3b683d),
	.w6(32'h3bf19ae3),
	.w7(32'hbb17ed18),
	.w8(32'h3c974f4b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24f5f4),
	.w1(32'h3980c7fd),
	.w2(32'hbad83341),
	.w3(32'hbb354bd9),
	.w4(32'hba41faa1),
	.w5(32'hbbe91307),
	.w6(32'hbba68a9f),
	.w7(32'hbb2a1f89),
	.w8(32'h3a212714),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0fdd7),
	.w1(32'hbb33e886),
	.w2(32'h3ab9b493),
	.w3(32'h3bafc8c3),
	.w4(32'hba5d4037),
	.w5(32'hbac81486),
	.w6(32'hbb2be5e4),
	.w7(32'hbb9166a0),
	.w8(32'hbb25e369),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cd1ab),
	.w1(32'h3b5bd4b1),
	.w2(32'h3a4659a6),
	.w3(32'h3b3dd687),
	.w4(32'hb9c3b986),
	.w5(32'h3c0656db),
	.w6(32'h3a1c5df1),
	.w7(32'h3b29337c),
	.w8(32'hba4ca144),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa1549),
	.w1(32'hbab020b5),
	.w2(32'h3bb9f1dc),
	.w3(32'hbb02b3ec),
	.w4(32'h3b4bd97a),
	.w5(32'h3a41dd07),
	.w6(32'h3b5cf540),
	.w7(32'h39ad700e),
	.w8(32'h3b3148a5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb8ba3),
	.w1(32'h3b7b24ac),
	.w2(32'h3b6c17b6),
	.w3(32'h3aba62e6),
	.w4(32'h3b4ac89c),
	.w5(32'h3abe2ef1),
	.w6(32'hbb0c8a99),
	.w7(32'hbb05ea32),
	.w8(32'h3a49cbd8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bc215),
	.w1(32'h38d48dbe),
	.w2(32'hb9e61796),
	.w3(32'h3ab2a173),
	.w4(32'h3c698266),
	.w5(32'h3a43fcaf),
	.w6(32'h39a93e26),
	.w7(32'h3aafe516),
	.w8(32'hbaddd056),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f4108),
	.w1(32'hbc1d9f0c),
	.w2(32'hbb6492df),
	.w3(32'h39b355cf),
	.w4(32'hbab45c77),
	.w5(32'hbb27250a),
	.w6(32'hba860917),
	.w7(32'h3b84eadb),
	.w8(32'hbbabcfeb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00ad6d),
	.w1(32'h3c38ba95),
	.w2(32'hbb3eadb1),
	.w3(32'hbb39a940),
	.w4(32'h3c800355),
	.w5(32'hba544c7d),
	.w6(32'h3b3d2e0c),
	.w7(32'hbba3104b),
	.w8(32'hba6d4a09),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf4010),
	.w1(32'h3aabf688),
	.w2(32'hba519fa1),
	.w3(32'hbb8b6047),
	.w4(32'h3bba4bdc),
	.w5(32'h37c26082),
	.w6(32'h3babc474),
	.w7(32'hbaa903f3),
	.w8(32'h3c33acff),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fe4f4),
	.w1(32'h3b2a690e),
	.w2(32'hbb49836e),
	.w3(32'hba586acc),
	.w4(32'h382551e1),
	.w5(32'h3b3a4d09),
	.w6(32'h3c7f084c),
	.w7(32'hbc64c20e),
	.w8(32'h3900d8b0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1054e),
	.w1(32'h3b0e4d8d),
	.w2(32'hbafb11ea),
	.w3(32'hbb8f49b1),
	.w4(32'h3b1dc6c0),
	.w5(32'hb981f712),
	.w6(32'hbb7fc8f1),
	.w7(32'hba9c46c3),
	.w8(32'h3b339794),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beabc79),
	.w1(32'hbbbfee1d),
	.w2(32'h3b306965),
	.w3(32'hbb250383),
	.w4(32'h3a94067e),
	.w5(32'h39f439bd),
	.w6(32'h3aff7c49),
	.w7(32'hbae7ad13),
	.w8(32'hbaec00e2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45a867),
	.w1(32'h3a8f11c2),
	.w2(32'hbb9d26a1),
	.w3(32'hba84702b),
	.w4(32'hb99af703),
	.w5(32'hbc294e97),
	.w6(32'hbb100e41),
	.w7(32'hbb26fea2),
	.w8(32'hbb5d7d21),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09cb5f),
	.w1(32'hbc0ba3c2),
	.w2(32'hbb8ae89d),
	.w3(32'hbb125593),
	.w4(32'h3ac6a0db),
	.w5(32'hbc2c9627),
	.w6(32'hbb958b69),
	.w7(32'h3c99c70a),
	.w8(32'hbb42a632),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddaf92),
	.w1(32'hb8464f23),
	.w2(32'hbb251e18),
	.w3(32'hbacedaf7),
	.w4(32'hbb13d0dc),
	.w5(32'h3a35f9c6),
	.w6(32'hbb51c05b),
	.w7(32'h3b6e1f0c),
	.w8(32'hbb921d24),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e301e),
	.w1(32'h3b057155),
	.w2(32'h3c702fde),
	.w3(32'h3bb6e382),
	.w4(32'h399eb56a),
	.w5(32'hb87eec66),
	.w6(32'h3a81255d),
	.w7(32'hbb89cf79),
	.w8(32'hba49b02f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4663ba),
	.w1(32'hbb69131d),
	.w2(32'h3a33c040),
	.w3(32'h3ab5e3d2),
	.w4(32'h3b696a32),
	.w5(32'hb99fbcd5),
	.w6(32'h3757a285),
	.w7(32'hbab154ac),
	.w8(32'h3bd88e6c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7aa532a),
	.w1(32'hbbe77fe7),
	.w2(32'h3a762fb6),
	.w3(32'h3aea8624),
	.w4(32'hbb0c4b67),
	.w5(32'h3b8d7c98),
	.w6(32'h38f5f2f9),
	.w7(32'hbb2a912d),
	.w8(32'h3b9dda5d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f8cec),
	.w1(32'h399f54a9),
	.w2(32'h39ceead5),
	.w3(32'h3b87651c),
	.w4(32'h3abdc736),
	.w5(32'hb9d95e46),
	.w6(32'hba47ea80),
	.w7(32'h3b6ba37b),
	.w8(32'hba770327),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14745c),
	.w1(32'h3a2b76c4),
	.w2(32'h3b9e6582),
	.w3(32'hbb3a2a96),
	.w4(32'h3a5c5632),
	.w5(32'hba983954),
	.w6(32'hbb69125f),
	.w7(32'h3ad006e6),
	.w8(32'hb85a2e99),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cdd13),
	.w1(32'hbb1f265f),
	.w2(32'hbad13d8b),
	.w3(32'h3990252d),
	.w4(32'hba57dc47),
	.w5(32'h3c18c5f4),
	.w6(32'h3ab259d6),
	.w7(32'h3ad685ee),
	.w8(32'h39b4bd3c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bdbf3),
	.w1(32'h3aa98d0e),
	.w2(32'h3a846ae2),
	.w3(32'h3b47eccb),
	.w4(32'h3b1cc8e3),
	.w5(32'h3af90729),
	.w6(32'hbb2a2c98),
	.w7(32'h3b143b46),
	.w8(32'hba82ae63),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebd25e),
	.w1(32'h3b226152),
	.w2(32'h3b267806),
	.w3(32'h3a30f417),
	.w4(32'hbb11831a),
	.w5(32'h39393502),
	.w6(32'hba32b5ec),
	.w7(32'h39b4c41a),
	.w8(32'h3a71ec68),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8923b2),
	.w1(32'hbc83d212),
	.w2(32'h3b44af5b),
	.w3(32'h3b442166),
	.w4(32'h3b314b00),
	.w5(32'h399fa456),
	.w6(32'hbc17ba85),
	.w7(32'h3b1efc20),
	.w8(32'h3b7f9ad3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b459),
	.w1(32'h3a641fb5),
	.w2(32'hba8234f9),
	.w3(32'h3adf75d4),
	.w4(32'hba0c67c2),
	.w5(32'h3b466824),
	.w6(32'h3b743e1a),
	.w7(32'h3afedd69),
	.w8(32'hb918d896),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea868),
	.w1(32'h3b17f571),
	.w2(32'h3b3405ca),
	.w3(32'h3a0517c0),
	.w4(32'h3b3e3347),
	.w5(32'hbb902a9e),
	.w6(32'h3b69fe0e),
	.w7(32'h3c0c9e32),
	.w8(32'h3b1c3244),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3cb43),
	.w1(32'h3a50e381),
	.w2(32'hbb2ee26b),
	.w3(32'hbafcea27),
	.w4(32'h3a6f1d3b),
	.w5(32'hbaec05ba),
	.w6(32'hbc0ea3cf),
	.w7(32'h379abe41),
	.w8(32'h39295699),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a908f66),
	.w1(32'h39ef3863),
	.w2(32'h3b55c1f8),
	.w3(32'hb9dc9bf3),
	.w4(32'h3a855dc2),
	.w5(32'hb95220ae),
	.w6(32'h3a678c56),
	.w7(32'hbb12d8e5),
	.w8(32'hbc176b03),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5eecc9),
	.w1(32'h3cb20fb4),
	.w2(32'hbc012368),
	.w3(32'h3af40c43),
	.w4(32'hbb58234f),
	.w5(32'hba8c1534),
	.w6(32'hbb9d805e),
	.w7(32'hbb3b6523),
	.w8(32'h3b01195a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule